// This is the unpowered netlist.
module wrapped_6502 (clk,
    io_oeb,
    rst,
    io_in,
    io_out);
 input clk;
 output io_oeb;
 input rst;
 input [9:0] io_in;
 output [26:0] io_out;

 wire net12;
 wire net13;
 wire \MOS6502.ABH[0] ;
 wire \MOS6502.ABH[1] ;
 wire \MOS6502.ABH[2] ;
 wire \MOS6502.ABH[3] ;
 wire \MOS6502.ABH[4] ;
 wire \MOS6502.ABH[5] ;
 wire \MOS6502.ABH[6] ;
 wire \MOS6502.ABH[7] ;
 wire \MOS6502.ABL[0] ;
 wire \MOS6502.ABL[1] ;
 wire \MOS6502.ABL[2] ;
 wire \MOS6502.ABL[3] ;
 wire \MOS6502.ABL[4] ;
 wire \MOS6502.ABL[5] ;
 wire \MOS6502.ABL[6] ;
 wire \MOS6502.ABL[7] ;
 wire \MOS6502.ADD[0] ;
 wire \MOS6502.ADD[1] ;
 wire \MOS6502.ADD[2] ;
 wire \MOS6502.ADD[3] ;
 wire \MOS6502.ADD[4] ;
 wire \MOS6502.ADD[5] ;
 wire \MOS6502.ADD[6] ;
 wire \MOS6502.ADD[7] ;
 wire \MOS6502.AI[7] ;
 wire \MOS6502.ALU.AI7 ;
 wire \MOS6502.ALU.BI7 ;
 wire \MOS6502.ALU.CO ;
 wire \MOS6502.ALU.HC ;
 wire \MOS6502.ALU.temp[0] ;
 wire \MOS6502.ALU.temp[1] ;
 wire \MOS6502.ALU.temp[2] ;
 wire \MOS6502.ALU.temp[3] ;
 wire \MOS6502.ALU.temp[4] ;
 wire \MOS6502.ALU.temp[5] ;
 wire \MOS6502.ALU.temp[6] ;
 wire \MOS6502.ALU.temp[7] ;
 wire \MOS6502.ALU.temp_BI[7] ;
 wire \MOS6502.ALU.temp_HC ;
 wire \MOS6502.AXYS[0][0] ;
 wire \MOS6502.AXYS[0][1] ;
 wire \MOS6502.AXYS[0][2] ;
 wire \MOS6502.AXYS[0][3] ;
 wire \MOS6502.AXYS[0][4] ;
 wire \MOS6502.AXYS[0][5] ;
 wire \MOS6502.AXYS[0][6] ;
 wire \MOS6502.AXYS[0][7] ;
 wire \MOS6502.AXYS[1][0] ;
 wire \MOS6502.AXYS[1][1] ;
 wire \MOS6502.AXYS[1][2] ;
 wire \MOS6502.AXYS[1][3] ;
 wire \MOS6502.AXYS[1][4] ;
 wire \MOS6502.AXYS[1][5] ;
 wire \MOS6502.AXYS[1][6] ;
 wire \MOS6502.AXYS[1][7] ;
 wire \MOS6502.AXYS[2][0] ;
 wire \MOS6502.AXYS[2][1] ;
 wire \MOS6502.AXYS[2][2] ;
 wire \MOS6502.AXYS[2][3] ;
 wire \MOS6502.AXYS[2][4] ;
 wire \MOS6502.AXYS[2][5] ;
 wire \MOS6502.AXYS[2][6] ;
 wire \MOS6502.AXYS[2][7] ;
 wire \MOS6502.AXYS[3][0] ;
 wire \MOS6502.AXYS[3][1] ;
 wire \MOS6502.AXYS[3][2] ;
 wire \MOS6502.AXYS[3][3] ;
 wire \MOS6502.AXYS[3][4] ;
 wire \MOS6502.AXYS[3][5] ;
 wire \MOS6502.AXYS[3][6] ;
 wire \MOS6502.AXYS[3][7] ;
 wire \MOS6502.C ;
 wire \MOS6502.D ;
 wire \MOS6502.I ;
 wire \MOS6502.IRHOLD[0] ;
 wire \MOS6502.IRHOLD[1] ;
 wire \MOS6502.IRHOLD[2] ;
 wire \MOS6502.IRHOLD[3] ;
 wire \MOS6502.IRHOLD[4] ;
 wire \MOS6502.IRHOLD[5] ;
 wire \MOS6502.IRHOLD[6] ;
 wire \MOS6502.IRHOLD[7] ;
 wire \MOS6502.IRHOLD_valid ;
 wire \MOS6502.IR[5] ;
 wire \MOS6502.IR[6] ;
 wire \MOS6502.IR[7] ;
 wire \MOS6502.N ;
 wire \MOS6502.NMI_1 ;
 wire \MOS6502.NMI_edge ;
 wire \MOS6502.PC[0] ;
 wire \MOS6502.PC[10] ;
 wire \MOS6502.PC[11] ;
 wire \MOS6502.PC[12] ;
 wire \MOS6502.PC[13] ;
 wire \MOS6502.PC[14] ;
 wire \MOS6502.PC[15] ;
 wire \MOS6502.PC[1] ;
 wire \MOS6502.PC[2] ;
 wire \MOS6502.PC[3] ;
 wire \MOS6502.PC[4] ;
 wire \MOS6502.PC[5] ;
 wire \MOS6502.PC[6] ;
 wire \MOS6502.PC[7] ;
 wire \MOS6502.PC[8] ;
 wire \MOS6502.PC[9] ;
 wire \MOS6502.V ;
 wire \MOS6502.Z ;
 wire \MOS6502.adc_bcd ;
 wire \MOS6502.adc_sbc ;
 wire \MOS6502.adj_bcd ;
 wire \MOS6502.backwards ;
 wire \MOS6502.bit_ins ;
 wire \MOS6502.clc ;
 wire \MOS6502.cld ;
 wire \MOS6502.cli ;
 wire \MOS6502.clv ;
 wire \MOS6502.compare ;
 wire \MOS6502.cond_code[0] ;
 wire \MOS6502.cond_code[1] ;
 wire \MOS6502.cond_code[2] ;
 wire \MOS6502.dst_reg[0] ;
 wire \MOS6502.dst_reg[1] ;
 wire \MOS6502.inc ;
 wire \MOS6502.index_y ;
 wire \MOS6502.load_only ;
 wire \MOS6502.load_reg ;
 wire \MOS6502.op[0] ;
 wire \MOS6502.op[1] ;
 wire \MOS6502.op[2] ;
 wire \MOS6502.op[3] ;
 wire \MOS6502.php ;
 wire \MOS6502.plp ;
 wire \MOS6502.res ;
 wire \MOS6502.rotate ;
 wire \MOS6502.sec ;
 wire \MOS6502.sed ;
 wire \MOS6502.sei ;
 wire \MOS6502.shift ;
 wire \MOS6502.shift_right ;
 wire \MOS6502.src_reg[0] ;
 wire \MOS6502.src_reg[1] ;
 wire \MOS6502.state[0] ;
 wire \MOS6502.state[1] ;
 wire \MOS6502.state[2] ;
 wire \MOS6502.state[3] ;
 wire \MOS6502.state[4] ;
 wire \MOS6502.state[5] ;
 wire \MOS6502.store ;
 wire \MOS6502.write_back ;
 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire clknet_0_clk;
 wire clknet_4_0_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire net1;
 wire net10;
 wire net11;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;

 sky130_fd_sc_hd__diode_2 ANTENNA__0974__A (.DIODE(_0356_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0975__A0 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__0978__A0 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__0981__A0 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__1001__B (.DIODE(_0380_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1007__B (.DIODE(_0380_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1016__B (.DIODE(_0395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1032__A (.DIODE(_0410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1033__B1 (.DIODE(\MOS6502.store ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1049__B (.DIODE(_0426_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1057__A (.DIODE(_0380_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1071__B2 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__1074__A (.DIODE(_0426_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1084__C (.DIODE(_0461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1093__A1 (.DIODE(_0380_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1097__B2 (.DIODE(\MOS6502.load_only ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1097__C1 (.DIODE(_0474_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1106__D (.DIODE(_0461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1114__A2 (.DIODE(_0461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1117__A2 (.DIODE(_0461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1126__B (.DIODE(_0503_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1127__B2 (.DIODE(\MOS6502.ADD[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1128__A1 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__1139__B (.DIODE(_0516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1140__A1 (.DIODE(\MOS6502.ABH[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1140__B2 (.DIODE(\MOS6502.ADD[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1141__A1 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__1148__A1 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__1149__A1 (.DIODE(\MOS6502.ADD[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1150__A2 (.DIODE(_0525_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1151__B2 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__1163__A1 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__1164__A1 (.DIODE(\MOS6502.ADD[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1165__A2 (.DIODE(_0540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1167__B2 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__1177__A (.DIODE(_0426_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1179__B2 (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__1186__A1 (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__1187__A1 (.DIODE(\MOS6502.ADD[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1196__A1 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__1197__A1 (.DIODE(\MOS6502.ADD[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1200__A1 (.DIODE(_0426_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1201__A (.DIODE(\MOS6502.load_only ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1210__B1 (.DIODE(\MOS6502.ALU.CO ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1211__B1 (.DIODE(_0410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1219__B2 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__1231__A1 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__1232__A1 (.DIODE(\MOS6502.ADD[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1233__A2 (.DIODE(_0608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1238__B2 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__1247__A1 (.DIODE(_0426_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1257__A1 (.DIODE(_0426_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1260__A1 (.DIODE(_0426_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1265__B (.DIODE(_0640_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1266__A1 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__1267__A1 (.DIODE(\MOS6502.ADD[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1269__B2 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__1276__A (.DIODE(_0426_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1284__B2 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__1291__A1 (.DIODE(_0426_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1310__A (.DIODE(_0461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1318__A (.DIODE(_0356_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1318__B (.DIODE(_0461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1319__A1 (.DIODE(_0677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1319__A2 (.DIODE(_0678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1322__A (.DIODE(_0356_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1322__B (.DIODE(_0689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1323__A1 (.DIODE(\MOS6502.ADD[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1328__B (.DIODE(\MOS6502.ALU.CO ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1334__B (.DIODE(_0380_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1335__B2 (.DIODE(\MOS6502.ADD[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1341__B1 (.DIODE(_0677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1342__A1 (.DIODE(\MOS6502.ADD[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1346__A1 (.DIODE(_0678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1347__A1 (.DIODE(\MOS6502.ADD[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1347__C1 (.DIODE(_0677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1351__A1 (.DIODE(\MOS6502.ADD[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1351__C1 (.DIODE(_0677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1355__A1 (.DIODE(\MOS6502.ADD[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1355__C1 (.DIODE(_0677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1359__A1 (.DIODE(\MOS6502.ADD[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1359__C1 (.DIODE(_0677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1363__A (.DIODE(_0677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1364__A1 (.DIODE(\MOS6502.ADD[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1370__A (.DIODE(_0677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1370__B (.DIODE(_0678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1373__A1 (.DIODE(\MOS6502.ADD[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1374__A1 (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__1376__A1 (.DIODE(\MOS6502.ADD[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1377__A1 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__1381__A1 (.DIODE(\MOS6502.ADD[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1382__A1 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__1384__A1 (.DIODE(\MOS6502.ADD[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1385__A1 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__1385__B2 (.DIODE(\MOS6502.PC[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1389__A1 (.DIODE(\MOS6502.ADD[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1390__A1 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__1392__A1 (.DIODE(\MOS6502.ADD[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1393__A1 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__1397__A1 (.DIODE(\MOS6502.ADD[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1397__B2 (.DIODE(\MOS6502.ABH[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1398__A1 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__1398__B2 (.DIODE(\MOS6502.PC[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1403__A1 (.DIODE(\MOS6502.ADD[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1404__A1 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__1411__A1 (.DIODE(_0426_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1412__B2 (.DIODE(_0410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1414__A0 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__1415__A (.DIODE(_0356_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1416__A0 (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__1417__A (.DIODE(_0356_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1419__A0 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__1422__A0 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__1424__A0 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__1434__A1 (.DIODE(_0410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1435__B1 (.DIODE(_0689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1436__A1 (.DIODE(\MOS6502.ALU.CO ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1436__A2 (.DIODE(\MOS6502.store ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1437__A1 (.DIODE(\MOS6502.ALU.CO ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1437__A2 (.DIODE(\MOS6502.store ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1445__A (.DIODE(_0689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1450__A (.DIODE(_0678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1452__A (.DIODE(_0689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1462__A (.DIODE(_0689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1469__A (.DIODE(_0689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1470__A (.DIODE(_0689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1472__A (.DIODE(_0410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1473__A (.DIODE(_0689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1477__A (.DIODE(_0814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1488__A (.DIODE(_0689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1506__D1 (.DIODE(_0678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1512__A (.DIODE(_0410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1514__A (.DIODE(\MOS6502.ALU.CO ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1514__C (.DIODE(\MOS6502.store ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1515__B2 (.DIODE(_0678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1534__A1_N (.DIODE(_0410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1535__C (.DIODE(_0814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1539__A (.DIODE(_0883_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1543__B1 (.DIODE(_0883_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1547__A1 (.DIODE(_0380_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1552__A (.DIODE(_0395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1556__B (.DIODE(_0677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1557__A (.DIODE(_0410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1560__A1 (.DIODE(_0410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1562__A1 (.DIODE(\MOS6502.ADD[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1562__A2 (.DIODE(_0902_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1562__B2 (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__1566__B (.DIODE(_0902_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1569__B (.DIODE(_0902_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1572__B2 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__1572__C1 (.DIODE(_0913_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1573__B1 (.DIODE(_0902_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1573__B2 (.DIODE(\MOS6502.ADD[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1575__B2 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__1575__C1 (.DIODE(_0913_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1576__A1_N (.DIODE(_0608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1576__B1 (.DIODE(_0902_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1576__B2 (.DIODE(\MOS6502.ADD[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1578__B2 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__1579__A1_N (.DIODE(_0540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1579__B1 (.DIODE(_0902_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1579__B2 (.DIODE(\MOS6502.ADD[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1581__B2 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__1582__A1_N (.DIODE(_0525_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1582__B1 (.DIODE(_0902_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1582__B2 (.DIODE(\MOS6502.ADD[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1584__B2 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__1585__A1_N (.DIODE(_0503_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1585__B1 (.DIODE(_0902_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1585__B2 (.DIODE(\MOS6502.ADD[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1587__B2 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__1588__A1_N (.DIODE(_0516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1588__B1 (.DIODE(_0902_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1588__B2 (.DIODE(\MOS6502.ADD[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1590__B2 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__1591__A1_N (.DIODE(_0640_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1591__B1 (.DIODE(_0902_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1591__B2 (.DIODE(\MOS6502.ADD[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1593__A1 (.DIODE(\MOS6502.ADD[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1594__A (.DIODE(_0395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1596__A1 (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__1597__A2 (.DIODE(_0913_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1598__A1 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__1599__A1 (.DIODE(\MOS6502.ADD[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1599__B1 (.DIODE(_0913_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1601__A1 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__1601__B2 (.DIODE(\MOS6502.ADD[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1602__A2 (.DIODE(_0913_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1603__A1 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__1603__B2 (.DIODE(\MOS6502.ADD[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1604__A1 (.DIODE(\MOS6502.PC[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1604__A2 (.DIODE(_0913_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1605__A1 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__1605__B2 (.DIODE(\MOS6502.ADD[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1606__A2 (.DIODE(_0913_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1607__A1 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__1607__B2 (.DIODE(\MOS6502.ADD[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1608__A2 (.DIODE(_0913_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1609__A1 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__1609__B2 (.DIODE(\MOS6502.ADD[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1610__A1 (.DIODE(\MOS6502.PC[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1610__A2 (.DIODE(_0913_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1610__B2 (.DIODE(\MOS6502.ABH[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1611__A1 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__1611__B2 (.DIODE(\MOS6502.ADD[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1612__A2 (.DIODE(_0913_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1613__B (.DIODE(_0395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1614__A1 (.DIODE(\MOS6502.php ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1616__A1 (.DIODE(\MOS6502.php ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1616__B1_N (.DIODE(_0395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1617__B2 (.DIODE(\MOS6502.ADD[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1621__B2 (.DIODE(\MOS6502.ADD[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1624__B2 (.DIODE(\MOS6502.ADD[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1625__B (.DIODE(_0608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1627__B2 (.DIODE(\MOS6502.PC[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1628__B2 (.DIODE(\MOS6502.ADD[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1629__A2 (.DIODE(_0540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1630__A2 (.DIODE(_0395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1630__B1 (.DIODE(\MOS6502.ADD[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1632__A1 (.DIODE(\MOS6502.php ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1634__A2 (.DIODE(_0525_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1635__B (.DIODE(_0503_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1636__A2 (.DIODE(_0395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1636__B1 (.DIODE(\MOS6502.ADD[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1639__A (.DIODE(_0960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1641__A1 (.DIODE(\MOS6502.PC[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1641__B2 (.DIODE(\MOS6502.ADD[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1642__A2_N (.DIODE(_0516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1644__A2_N (.DIODE(_0640_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1644__B2 (.DIODE(\MOS6502.ADD[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1646__A (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__1647__A (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__1648__A (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__1649__A (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__1650__A (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__1651__A (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__1653__A0 (.DIODE(\MOS6502.ADD[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1653__A1 (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__1658__S (.DIODE(_0970_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1663__A (.DIODE(\MOS6502.ADD[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1664__B1 (.DIODE(\MOS6502.ADD[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1666__A1 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__1667__S (.DIODE(_0970_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1669__A (.DIODE(\MOS6502.ADD[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1670__A (.DIODE(\MOS6502.ADD[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1673__B1 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__1674__S (.DIODE(_0970_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1677__A (.DIODE(\MOS6502.ADD[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1679__A1 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__1680__S (.DIODE(_0970_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1682__A0 (.DIODE(\MOS6502.ADD[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1682__A1 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__1683__S (.DIODE(_0970_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1685__A (.DIODE(\MOS6502.ALU.CO ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1686__A (.DIODE(\MOS6502.ALU.CO ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1687__B1 (.DIODE(\MOS6502.ADD[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1688__A (.DIODE(\MOS6502.ADD[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1690__A1 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__1691__S (.DIODE(_0970_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1693__A (.DIODE(\MOS6502.ADD[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1694__A (.DIODE(\MOS6502.ADD[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1697__B1 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__1698__S (.DIODE(_0970_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1701__A (.DIODE(\MOS6502.ADD[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1704__A1 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__1704__A2 (.DIODE(_0410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1704__A3 (.DIODE(_0380_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1705__A1 (.DIODE(_0163_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1705__S (.DIODE(_0970_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1723__A1 (.DIODE(_0163_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1728__A (.DIODE(_0677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1729__B (.DIODE(_0678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1735__B (.DIODE(_0474_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1738__S (.DIODE(_0187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1740__S (.DIODE(_0187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1742__S (.DIODE(_0187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1744__S (.DIODE(_0187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1746__S (.DIODE(_0187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1748__S (.DIODE(_0187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1750__S (.DIODE(_0187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1752__S (.DIODE(_0187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1755__A1 (.DIODE(\MOS6502.ADD[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1757__A1 (.DIODE(\MOS6502.ALU.CO ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1758__A0 (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__1761__A2_N (.DIODE(_0883_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1761__B1 (.DIODE(_0395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1766__A (.DIODE(\MOS6502.ADD[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1766__B (.DIODE(\MOS6502.ADD[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1766__C (.DIODE(\MOS6502.ADD[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1766__D (.DIODE(\MOS6502.ADD[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1767__A (.DIODE(\MOS6502.ADD[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1767__B (.DIODE(\MOS6502.ADD[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1767__C (.DIODE(\MOS6502.ADD[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1767__D (.DIODE(\MOS6502.ADD[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1769__A0 (.DIODE(\MOS6502.ADD[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1769__A1 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__1770__B1_N (.DIODE(_0395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1777__A0 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__1777__A1 (.DIODE(\MOS6502.ADD[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1778__B1 (.DIODE(_0678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1779__A1 (.DIODE(_0395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1783__A1 (.DIODE(\MOS6502.ADD[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1784__A0 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__1785__A (.DIODE(_0678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1787__A1 (.DIODE(_0224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1791__A0 (.DIODE(\MOS6502.ADD[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1792__A0 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__1794__A2 (.DIODE(_0678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1796__A (.DIODE(_0814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1800__A (.DIODE(\MOS6502.ADD[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1800__B (.DIODE(\MOS6502.ALU.CO ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1802__A2 (.DIODE(\MOS6502.ADD[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1802__C1 (.DIODE(_0883_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1803__A1 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__1803__A2 (.DIODE(_0224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1804__A4 (.DIODE(_0883_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1807__A (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__1807__B (.DIODE(_0474_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1809__A0 (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__1811__A0 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__1813__A0 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__1815__A0 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__1817__A0 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__1819__A0 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__1821__A0 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__1823__A0 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__1825__A (.DIODE(_0883_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1827__A1 (.DIODE(_0474_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1827__B1 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__1845__A (.DIODE(_0224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1848__A (.DIODE(_0883_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1849__A2 (.DIODE(_0274_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1849__B1 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__1864__B1 (.DIODE(_0883_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1874__S (.DIODE(_0224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1877__A0 (.DIODE(\MOS6502.store ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1877__S (.DIODE(_0224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1879__B (.DIODE(_0883_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1881__A0 (.DIODE(\MOS6502.load_only ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1881__S (.DIODE(_0224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1885__A2 (.DIODE(_0274_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1889__B (.DIODE(_0224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1890__A2 (.DIODE(_0274_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1895__A2 (.DIODE(_0274_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1897__S (.DIODE(_0224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1899__A2 (.DIODE(_0274_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1900__C (.DIODE(_0883_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1910__S (.DIODE(_0224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1914__A2 (.DIODE(_0274_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1915__S (.DIODE(_0224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1918__B2 (.DIODE(_0274_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1921__A2 (.DIODE(_0274_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1923__A2 (.DIODE(_0274_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1924__A2 (.DIODE(_0274_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1928__A1 (.DIODE(\MOS6502.php ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1931__A2 (.DIODE(_0814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1932__S (.DIODE(_0187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1934__S (.DIODE(_0187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1944__A0 (.DIODE(\MOS6502.ABH[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1950__S (.DIODE(_0336_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1952__S (.DIODE(_0336_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1954__S (.DIODE(_0336_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1956__S (.DIODE(_0336_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1958__S (.DIODE(_0336_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1960__S (.DIODE(_0336_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1962__S (.DIODE(_0336_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1964__A1 (.DIODE(_0163_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1964__S (.DIODE(_0336_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1982__A1 (.DIODE(_0163_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1988__CLK (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1989__CLK (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__2018__CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__2022__CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__2025__CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__2041__CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__2042__CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__2044__CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__2044__D (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__2045__CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__2046__CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__2048__CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__2071__CLK (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__2075__CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__2090__CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__2093__CLK (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__2094__CLK (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__2095__CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__2096__CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_clk_A (.DIODE(clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_0_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_10_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_11_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_12_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_13_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_14_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_15_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_1_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_2_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_3_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_4_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_5_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_6_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_7_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_8_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_9_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_input10_A (.DIODE(io_in[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input11_A (.DIODE(rst));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_A (.DIODE(io_in[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_A (.DIODE(io_in[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input3_A (.DIODE(io_in[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input4_A (.DIODE(io_in[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input5_A (.DIODE(io_in[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input6_A (.DIODE(io_in[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input7_A (.DIODE(io_in[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input8_A (.DIODE(io_in[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input9_A (.DIODE(io_in[8]));
 sky130_fd_sc_hd__decap_3 FILLER_0_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_460 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_439 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_439 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_442 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_412 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_439 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_39 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_275 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_386 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_341 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_400 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_424 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_387 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_410 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_425 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_255 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_286 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_356 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_366 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_378 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_404 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_226 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_329 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_340 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_375 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_204 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_254 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_311 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_348 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_368 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_159 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_244 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_259 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_351 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_272 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_347 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_355 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_400 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_168 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_272 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_328 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_382 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_396 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_416 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_427 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_131 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_173 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_243 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_287 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_352 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_183 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_271 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_336 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_443 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_150 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_243 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_255 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_375 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_407 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_414 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_164 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_207 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_207 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_240 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_276 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_331 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_397 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_436 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_458 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_162 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_236 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_424 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_434 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_453 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_325 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_376 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_395 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_426 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_152 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_211 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_300 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_402 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_180 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_190 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_210 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_220 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_348 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_392 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_243 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_364 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_380 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_156 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_352 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_131 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_245 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_291 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_366 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_431 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_206 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_394 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_162 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_241 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_411 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_420 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_158 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_439 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_208 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_353 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_434 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_170 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_275 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_378 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_444 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_247 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_352 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_366 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_159 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_171 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_217 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_226 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_329 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_372 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_435 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_239 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_248 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_355 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_412 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_432 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_219 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_272 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_291 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_315 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_332 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_382 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_191 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_353 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_379 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_406 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_183 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_383 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_131 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_256 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_367 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_450 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_203 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_312 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_354 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_416 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_423 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_173 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_426 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_176 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_244 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_382 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_410 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_208 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_230 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_340 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_392 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_396 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_458 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_133 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_310 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_434 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_126 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_162 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_226 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_340 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_132 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_178 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_328 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_178 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_235 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_275 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_318 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_336 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_344 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_375 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_435 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_184 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_403 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_436 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_114 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_160 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_323 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_96 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_188 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_348 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_216 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_341 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_347 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_411 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_189 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_352 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_378 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_453 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_326 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_342 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_235 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_326 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_411 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_453 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_212 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_238 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_352 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_276 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_282 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_245 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_453 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_229 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_246 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_411 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_432 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_453 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_154 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_229 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_292 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_460 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_93 ();
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 ();
 sky130_fd_sc_hd__inv_2 _0972_ (.A(\MOS6502.I ),
    .Y(_0355_));
 sky130_fd_sc_hd__a21oi_4 _0973_ (.A1(_0355_),
    .A2(net9),
    .B1(\MOS6502.NMI_edge ),
    .Y(_0356_));
 sky130_fd_sc_hd__clkbuf_4 _0974_ (.A(_0356_),
    .X(_0357_));
 sky130_fd_sc_hd__mux2_2 _0975_ (.A0(net8),
    .A1(\MOS6502.IRHOLD[7] ),
    .S(\MOS6502.IRHOLD_valid ),
    .X(_0358_));
 sky130_fd_sc_hd__nand2_4 _0976_ (.A(_0357_),
    .B(_0358_),
    .Y(_0359_));
 sky130_fd_sc_hd__clkinv_2 _0977_ (.A(_0359_),
    .Y(\MOS6502.IR[7] ));
 sky130_fd_sc_hd__mux2_1 _0978_ (.A0(net6),
    .A1(\MOS6502.IRHOLD[5] ),
    .S(\MOS6502.IRHOLD_valid ),
    .X(_0360_));
 sky130_fd_sc_hd__nand2_1 _0979_ (.A(_0357_),
    .B(_0360_),
    .Y(_0361_));
 sky130_fd_sc_hd__clkinv_2 _0980_ (.A(_0361_),
    .Y(\MOS6502.IR[5] ));
 sky130_fd_sc_hd__mux2_1 _0981_ (.A0(net7),
    .A1(\MOS6502.IRHOLD[6] ),
    .S(\MOS6502.IRHOLD_valid ),
    .X(_0362_));
 sky130_fd_sc_hd__nand2_4 _0982_ (.A(_0357_),
    .B(_0362_),
    .Y(_0363_));
 sky130_fd_sc_hd__inv_2 _0983_ (.A(_0363_),
    .Y(\MOS6502.IR[6] ));
 sky130_fd_sc_hd__or2b_1 _0984_ (.A(\MOS6502.state[5] ),
    .B_N(\MOS6502.state[4] ),
    .X(_0364_));
 sky130_fd_sc_hd__clkbuf_4 _0985_ (.A(_0364_),
    .X(_0365_));
 sky130_fd_sc_hd__buf_2 _0986_ (.A(\MOS6502.state[2] ),
    .X(_0366_));
 sky130_fd_sc_hd__clkbuf_2 _0987_ (.A(_0366_),
    .X(_0367_));
 sky130_fd_sc_hd__inv_2 _0988_ (.A(\MOS6502.state[3] ),
    .Y(_0368_));
 sky130_fd_sc_hd__buf_2 _0989_ (.A(\MOS6502.state[1] ),
    .X(_0369_));
 sky130_fd_sc_hd__nand2_1 _0990_ (.A(_0369_),
    .B(\MOS6502.state[0] ),
    .Y(_0370_));
 sky130_fd_sc_hd__or3_2 _0991_ (.A(_0367_),
    .B(_0368_),
    .C(_0370_),
    .X(_0371_));
 sky130_fd_sc_hd__or2_2 _0992_ (.A(\MOS6502.state[4] ),
    .B(\MOS6502.state[5] ),
    .X(_0372_));
 sky130_fd_sc_hd__buf_2 _0993_ (.A(_0372_),
    .X(_0373_));
 sky130_fd_sc_hd__or2b_1 _0994_ (.A(\MOS6502.state[1] ),
    .B_N(\MOS6502.state[0] ),
    .X(_0374_));
 sky130_fd_sc_hd__or3_2 _0995_ (.A(_0366_),
    .B(_0368_),
    .C(_0374_),
    .X(_0375_));
 sky130_fd_sc_hd__or2_1 _0996_ (.A(_0373_),
    .B(_0375_),
    .X(_0376_));
 sky130_fd_sc_hd__o21ai_1 _0997_ (.A1(_0365_),
    .A2(_0371_),
    .B1(_0376_),
    .Y(_0377_));
 sky130_fd_sc_hd__clkbuf_2 _0998_ (.A(\MOS6502.state[0] ),
    .X(_0378_));
 sky130_fd_sc_hd__buf_2 _0999_ (.A(\MOS6502.state[3] ),
    .X(_0379_));
 sky130_fd_sc_hd__or4bb_4 _1000_ (.A(_0378_),
    .B(_0366_),
    .C_N(_0379_),
    .D_N(_0369_),
    .X(_0380_));
 sky130_fd_sc_hd__nor2_1 _1001_ (.A(_0373_),
    .B(_0380_),
    .Y(_0381_));
 sky130_fd_sc_hd__or2b_1 _1002_ (.A(\MOS6502.state[4] ),
    .B_N(\MOS6502.state[5] ),
    .X(_0382_));
 sky130_fd_sc_hd__buf_2 _1003_ (.A(_0382_),
    .X(_0383_));
 sky130_fd_sc_hd__or4b_1 _1004_ (.A(\MOS6502.state[0] ),
    .B(\MOS6502.state[2] ),
    .C(\MOS6502.state[3] ),
    .D_N(\MOS6502.state[1] ),
    .X(_0384_));
 sky130_fd_sc_hd__clkbuf_2 _1005_ (.A(_0384_),
    .X(_0385_));
 sky130_fd_sc_hd__nor2_2 _1006_ (.A(_0383_),
    .B(_0385_),
    .Y(_0386_));
 sky130_fd_sc_hd__nor2_2 _1007_ (.A(_0365_),
    .B(_0380_),
    .Y(_0387_));
 sky130_fd_sc_hd__or4b_2 _1008_ (.A(\MOS6502.state[1] ),
    .B(_0378_),
    .C(_0366_),
    .D_N(_0379_),
    .X(_0388_));
 sky130_fd_sc_hd__nor2_1 _1009_ (.A(_0373_),
    .B(_0388_),
    .Y(_0389_));
 sky130_fd_sc_hd__or2_1 _1010_ (.A(_0387_),
    .B(_0389_),
    .X(_0390_));
 sky130_fd_sc_hd__or4_2 _1011_ (.A(_0377_),
    .B(_0381_),
    .C(_0386_),
    .D(_0390_),
    .X(_0391_));
 sky130_fd_sc_hd__buf_2 _1012_ (.A(_0383_),
    .X(_0392_));
 sky130_fd_sc_hd__nand4b_4 _1013_ (.A_N(\MOS6502.state[0] ),
    .B(_0366_),
    .C(_0379_),
    .D(_0369_),
    .Y(_0393_));
 sky130_fd_sc_hd__nor2_1 _1014_ (.A(_0392_),
    .B(_0393_),
    .Y(_0394_));
 sky130_fd_sc_hd__buf_2 _1015_ (.A(_0394_),
    .X(_0395_));
 sky130_fd_sc_hd__or2_1 _1016_ (.A(_0391_),
    .B(_0395_),
    .X(_0396_));
 sky130_fd_sc_hd__clkbuf_4 _1017_ (.A(_0396_),
    .X(_0397_));
 sky130_fd_sc_hd__clkbuf_4 _1018_ (.A(_0373_),
    .X(_0398_));
 sky130_fd_sc_hd__or4b_1 _1019_ (.A(\MOS6502.state[1] ),
    .B(\MOS6502.state[0] ),
    .C(\MOS6502.state[3] ),
    .D_N(\MOS6502.state[2] ),
    .X(_0399_));
 sky130_fd_sc_hd__clkbuf_2 _1020_ (.A(_0399_),
    .X(_0400_));
 sky130_fd_sc_hd__nor2_1 _1021_ (.A(_0398_),
    .B(_0400_),
    .Y(_0401_));
 sky130_fd_sc_hd__or3_2 _1022_ (.A(_0367_),
    .B(_0379_),
    .C(_0374_),
    .X(_0402_));
 sky130_fd_sc_hd__nor2_1 _1023_ (.A(_0373_),
    .B(_0402_),
    .Y(_0403_));
 sky130_fd_sc_hd__buf_2 _1024_ (.A(\MOS6502.state[4] ),
    .X(_0404_));
 sky130_fd_sc_hd__nand2_1 _1025_ (.A(_0404_),
    .B(\MOS6502.state[5] ),
    .Y(_0405_));
 sky130_fd_sc_hd__nor2_1 _1026_ (.A(_0402_),
    .B(_0405_),
    .Y(_0406_));
 sky130_fd_sc_hd__nand2_2 _1027_ (.A(_0366_),
    .B(_0379_),
    .Y(_0407_));
 sky130_fd_sc_hd__nor3_1 _1028_ (.A(_0370_),
    .B(_0392_),
    .C(_0407_),
    .Y(_0408_));
 sky130_fd_sc_hd__or4_2 _1029_ (.A(_0401_),
    .B(_0403_),
    .C(_0406_),
    .D(_0408_),
    .X(_0409_));
 sky130_fd_sc_hd__buf_2 _1030_ (.A(_0365_),
    .X(_0410_));
 sky130_fd_sc_hd__or2_1 _1031_ (.A(_0379_),
    .B(_0374_),
    .X(_0411_));
 sky130_fd_sc_hd__nor2_1 _1032_ (.A(_0410_),
    .B(_0411_),
    .Y(_0412_));
 sky130_fd_sc_hd__o21a_1 _1033_ (.A1(_0409_),
    .A2(_0412_),
    .B1(\MOS6502.store ),
    .X(_0413_));
 sky130_fd_sc_hd__nor2_4 _1034_ (.A(_0397_),
    .B(_0413_),
    .Y(io_oeb));
 sky130_fd_sc_hd__inv_2 _1035_ (.A(io_oeb),
    .Y(io_out[26]));
 sky130_fd_sc_hd__or2_2 _1036_ (.A(_0374_),
    .B(_0407_),
    .X(_0414_));
 sky130_fd_sc_hd__nor2_2 _1037_ (.A(_0373_),
    .B(_0414_),
    .Y(_0415_));
 sky130_fd_sc_hd__or4bb_4 _1038_ (.A(_0366_),
    .B(\MOS6502.state[3] ),
    .C_N(_0369_),
    .D_N(_0378_),
    .X(_0416_));
 sky130_fd_sc_hd__nor2_1 _1039_ (.A(_0383_),
    .B(_0416_),
    .Y(_0417_));
 sky130_fd_sc_hd__nor2_1 _1040_ (.A(_0383_),
    .B(_0400_),
    .Y(_0418_));
 sky130_fd_sc_hd__or2_1 _1041_ (.A(_0417_),
    .B(_0418_),
    .X(_0419_));
 sky130_fd_sc_hd__or2_1 _1042_ (.A(_0415_),
    .B(_0419_),
    .X(_0420_));
 sky130_fd_sc_hd__clkbuf_4 _1043_ (.A(_0420_),
    .X(_0421_));
 sky130_fd_sc_hd__or4bb_4 _1044_ (.A(_0378_),
    .B(_0379_),
    .C_N(_0367_),
    .D_N(_0369_),
    .X(_0422_));
 sky130_fd_sc_hd__nor2_2 _1045_ (.A(_0373_),
    .B(_0422_),
    .Y(_0423_));
 sky130_fd_sc_hd__a221o_4 _1046_ (.A1(\MOS6502.op[2] ),
    .A2(_0421_),
    .B1(_0423_),
    .B2(\MOS6502.backwards ),
    .C1(_0391_),
    .X(_0424_));
 sky130_fd_sc_hd__and2_1 _1047_ (.A(\MOS6502.op[3] ),
    .B(_0421_),
    .X(_0425_));
 sky130_fd_sc_hd__clkbuf_4 _1048_ (.A(_0425_),
    .X(_0426_));
 sky130_fd_sc_hd__nor2_1 _1049_ (.A(_0424_),
    .B(_0426_),
    .Y(_0427_));
 sky130_fd_sc_hd__or4bb_4 _1050_ (.A(_0369_),
    .B(_0379_),
    .C_N(_0367_),
    .D_N(_0378_),
    .X(_0428_));
 sky130_fd_sc_hd__nor2_4 _1051_ (.A(_0372_),
    .B(_0428_),
    .Y(_0429_));
 sky130_fd_sc_hd__or3_1 _1052_ (.A(_0370_),
    .B(_0373_),
    .C(_0407_),
    .X(_0430_));
 sky130_fd_sc_hd__o21ai_1 _1053_ (.A1(_0404_),
    .A2(_0422_),
    .B1(_0430_),
    .Y(_0431_));
 sky130_fd_sc_hd__and4b_1 _1054_ (.A_N(_0366_),
    .B(\MOS6502.state[3] ),
    .C(\MOS6502.state[1] ),
    .D(\MOS6502.state[0] ),
    .X(_0432_));
 sky130_fd_sc_hd__xor2_1 _1055_ (.A(\MOS6502.state[4] ),
    .B(\MOS6502.state[5] ),
    .X(_0433_));
 sky130_fd_sc_hd__and2_1 _1056_ (.A(_0404_),
    .B(\MOS6502.state[5] ),
    .X(_0434_));
 sky130_fd_sc_hd__nor2_1 _1057_ (.A(_0380_),
    .B(_0434_),
    .Y(_0435_));
 sky130_fd_sc_hd__a21o_1 _1058_ (.A1(_0432_),
    .A2(_0433_),
    .B1(_0435_),
    .X(_0436_));
 sky130_fd_sc_hd__or2_1 _1059_ (.A(_0365_),
    .B(_0393_),
    .X(_0437_));
 sky130_fd_sc_hd__or3b_4 _1060_ (.A(_0379_),
    .B(_0370_),
    .C_N(_0367_),
    .X(_0438_));
 sky130_fd_sc_hd__or2_2 _1061_ (.A(_0392_),
    .B(_0438_),
    .X(_0439_));
 sky130_fd_sc_hd__or4bb_2 _1062_ (.A(_0431_),
    .B(_0436_),
    .C_N(_0437_),
    .D_N(_0439_),
    .X(_0440_));
 sky130_fd_sc_hd__or2_1 _1063_ (.A(_0417_),
    .B(_0429_),
    .X(_0441_));
 sky130_fd_sc_hd__buf_2 _1064_ (.A(_0441_),
    .X(_0442_));
 sky130_fd_sc_hd__or2_1 _1065_ (.A(_0383_),
    .B(_0411_),
    .X(_0443_));
 sky130_fd_sc_hd__nor3_1 _1066_ (.A(_0378_),
    .B(_0365_),
    .C(_0407_),
    .Y(_0444_));
 sky130_fd_sc_hd__and2b_1 _1067_ (.A_N(_0369_),
    .B(_0444_),
    .X(_0445_));
 sky130_fd_sc_hd__nor4_1 _1068_ (.A(_0386_),
    .B(_0389_),
    .C(_0418_),
    .D(_0445_),
    .Y(_0446_));
 sky130_fd_sc_hd__and4b_1 _1069_ (.A_N(_0442_),
    .B(_0443_),
    .C(_0376_),
    .D(_0446_),
    .X(_0447_));
 sky130_fd_sc_hd__nor2b_4 _1070_ (.A(_0440_),
    .B_N(_0447_),
    .Y(_0448_));
 sky130_fd_sc_hd__a22o_1 _1071_ (.A1(\MOS6502.PC[5] ),
    .A2(_0429_),
    .B1(_0448_),
    .B2(net6),
    .X(_0449_));
 sky130_fd_sc_hd__mux2_1 _1072_ (.A0(_0427_),
    .A1(_0424_),
    .S(_0449_),
    .X(_0450_));
 sky130_fd_sc_hd__inv_2 _1073_ (.A(_0424_),
    .Y(_0451_));
 sky130_fd_sc_hd__inv_2 _1074_ (.A(_0426_),
    .Y(_0452_));
 sky130_fd_sc_hd__nor2_1 _1075_ (.A(_0451_),
    .B(_0452_),
    .Y(_0453_));
 sky130_fd_sc_hd__or2_1 _1076_ (.A(_0450_),
    .B(_0453_),
    .X(_0454_));
 sky130_fd_sc_hd__nand2_1 _1077_ (.A(\MOS6502.shift_right ),
    .B(_0421_),
    .Y(_0455_));
 sky130_fd_sc_hd__buf_2 _1078_ (.A(_0455_),
    .X(_0456_));
 sky130_fd_sc_hd__nor2_1 _1079_ (.A(\MOS6502.state[4] ),
    .B(\MOS6502.state[5] ),
    .Y(_0457_));
 sky130_fd_sc_hd__nor2_1 _1080_ (.A(\MOS6502.state[1] ),
    .B(\MOS6502.state[0] ),
    .Y(_0458_));
 sky130_fd_sc_hd__and2_1 _1081_ (.A(_0366_),
    .B(\MOS6502.state[3] ),
    .X(_0459_));
 sky130_fd_sc_hd__and3_1 _1082_ (.A(_0457_),
    .B(_0458_),
    .C(_0459_),
    .X(_0460_));
 sky130_fd_sc_hd__buf_2 _1083_ (.A(_0460_),
    .X(_0461_));
 sky130_fd_sc_hd__nor3_2 _1084_ (.A(_0403_),
    .B(_0421_),
    .C(_0461_),
    .Y(_0462_));
 sky130_fd_sc_hd__a21oi_1 _1085_ (.A1(\MOS6502.op[0] ),
    .A2(_0421_),
    .B1(_0462_),
    .Y(_0463_));
 sky130_fd_sc_hd__buf_2 _1086_ (.A(_0463_),
    .X(_0464_));
 sky130_fd_sc_hd__buf_2 _1087_ (.A(_0423_),
    .X(_0465_));
 sky130_fd_sc_hd__buf_2 _1088_ (.A(_0377_),
    .X(_0466_));
 sky130_fd_sc_hd__a31o_1 _1089_ (.A1(_0371_),
    .A2(_0422_),
    .A3(_0438_),
    .B1(_0383_),
    .X(_0467_));
 sky130_fd_sc_hd__and2_1 _1090_ (.A(_0430_),
    .B(_0467_),
    .X(_0468_));
 sky130_fd_sc_hd__or3b_1 _1091_ (.A(_0466_),
    .B(_0381_),
    .C_N(_0468_),
    .X(_0469_));
 sky130_fd_sc_hd__clkbuf_2 _1092_ (.A(_0469_),
    .X(_0470_));
 sky130_fd_sc_hd__a21oi_2 _1093_ (.A1(_0380_),
    .A2(_0428_),
    .B1(_0383_),
    .Y(_0471_));
 sky130_fd_sc_hd__nor2_1 _1094_ (.A(_0387_),
    .B(_0471_),
    .Y(_0472_));
 sky130_fd_sc_hd__or2_1 _1095_ (.A(_0373_),
    .B(_0414_),
    .X(_0473_));
 sky130_fd_sc_hd__o21a_1 _1096_ (.A1(_0367_),
    .A2(_0443_),
    .B1(_0437_),
    .X(_0474_));
 sky130_fd_sc_hd__o221a_1 _1097_ (.A1(_0404_),
    .A2(_0385_),
    .B1(_0473_),
    .B2(\MOS6502.load_only ),
    .C1(_0474_),
    .X(_0475_));
 sky130_fd_sc_hd__o22ai_2 _1098_ (.A1(_0372_),
    .A2(_0393_),
    .B1(_0416_),
    .B2(_0365_),
    .Y(_0476_));
 sky130_fd_sc_hd__or4_2 _1099_ (.A(\MOS6502.state[1] ),
    .B(\MOS6502.state[0] ),
    .C(_0366_),
    .D(\MOS6502.state[3] ),
    .X(_0477_));
 sky130_fd_sc_hd__nor2_1 _1100_ (.A(_0405_),
    .B(_0477_),
    .Y(_0478_));
 sky130_fd_sc_hd__or2_1 _1101_ (.A(_0476_),
    .B(_0478_),
    .X(_0479_));
 sky130_fd_sc_hd__nor2_1 _1102_ (.A(_0389_),
    .B(_0479_),
    .Y(_0480_));
 sky130_fd_sc_hd__and4_1 _1103_ (.A(_0472_),
    .B(_0446_),
    .C(_0475_),
    .D(_0480_),
    .X(_0481_));
 sky130_fd_sc_hd__buf_2 _1104_ (.A(_0481_),
    .X(_0482_));
 sky130_fd_sc_hd__nor2_1 _1105_ (.A(_0372_),
    .B(_0385_),
    .Y(_0483_));
 sky130_fd_sc_hd__nor4_2 _1106_ (.A(_0476_),
    .B(_0478_),
    .C(_0483_),
    .D(_0461_),
    .Y(_0484_));
 sky130_fd_sc_hd__o22ai_1 _1107_ (.A1(_0404_),
    .A2(_0388_),
    .B1(_0393_),
    .B2(_0365_),
    .Y(_0485_));
 sky130_fd_sc_hd__a32o_1 _1108_ (.A1(_0458_),
    .A2(_0459_),
    .A3(_0433_),
    .B1(_0457_),
    .B2(_0432_),
    .X(_0486_));
 sky130_fd_sc_hd__or3_1 _1109_ (.A(_0365_),
    .B(_0370_),
    .C(_0407_),
    .X(_0487_));
 sky130_fd_sc_hd__or2_1 _1110_ (.A(_0383_),
    .B(_0385_),
    .X(_0488_));
 sky130_fd_sc_hd__and4bb_1 _1111_ (.A_N(_0485_),
    .B_N(_0486_),
    .C(_0487_),
    .D(_0488_),
    .X(_0489_));
 sky130_fd_sc_hd__nand4b_4 _1112_ (.A_N(\MOS6502.src_reg[0] ),
    .B(_0472_),
    .C(_0484_),
    .D(_0489_),
    .Y(_0490_));
 sky130_fd_sc_hd__o31a_1 _1113_ (.A1(_0476_),
    .A2(_0478_),
    .A3(_0483_),
    .B1(\MOS6502.index_y ),
    .X(_0491_));
 sky130_fd_sc_hd__a211o_2 _1114_ (.A1(\MOS6502.dst_reg[0] ),
    .A2(_0461_),
    .B1(_0484_),
    .C1(_0491_),
    .X(_0492_));
 sky130_fd_sc_hd__and2_2 _1115_ (.A(_0490_),
    .B(_0492_),
    .X(_0493_));
 sky130_fd_sc_hd__and4_1 _1116_ (.A(\MOS6502.src_reg[1] ),
    .B(_0472_),
    .C(_0484_),
    .D(_0489_),
    .X(_0494_));
 sky130_fd_sc_hd__a2111o_2 _1117_ (.A1(\MOS6502.dst_reg[1] ),
    .A2(_0461_),
    .B1(_0494_),
    .C1(_0479_),
    .D1(_0483_),
    .X(_0495_));
 sky130_fd_sc_hd__buf_4 _1118_ (.A(_0495_),
    .X(_0496_));
 sky130_fd_sc_hd__nor2_8 _1119_ (.A(_0493_),
    .B(_0496_),
    .Y(_0497_));
 sky130_fd_sc_hd__nand2_1 _1120_ (.A(_0490_),
    .B(_0492_),
    .Y(_0498_));
 sky130_fd_sc_hd__buf_4 _1121_ (.A(_0498_),
    .X(_0499_));
 sky130_fd_sc_hd__nor2_8 _1122_ (.A(_0499_),
    .B(_0496_),
    .Y(_0500_));
 sky130_fd_sc_hd__or2_1 _1123_ (.A(\MOS6502.AXYS[2][5] ),
    .B(_0493_),
    .X(_0501_));
 sky130_fd_sc_hd__o211a_1 _1124_ (.A1(\MOS6502.AXYS[3][5] ),
    .A2(_0499_),
    .B1(_0496_),
    .C1(_0501_),
    .X(_0502_));
 sky130_fd_sc_hd__a221oi_4 _1125_ (.A1(\MOS6502.AXYS[0][5] ),
    .A2(_0497_),
    .B1(_0500_),
    .B2(\MOS6502.AXYS[1][5] ),
    .C1(_0502_),
    .Y(_0503_));
 sky130_fd_sc_hd__nor2_1 _1126_ (.A(_0482_),
    .B(_0503_),
    .Y(_0504_));
 sky130_fd_sc_hd__a221o_1 _1127_ (.A1(\MOS6502.ABH[5] ),
    .A2(_0465_),
    .B1(_0470_),
    .B2(\MOS6502.ADD[5] ),
    .C1(_0504_),
    .X(_0505_));
 sky130_fd_sc_hd__a21oi_1 _1128_ (.A1(net6),
    .A2(_0442_),
    .B1(_0505_),
    .Y(_0506_));
 sky130_fd_sc_hd__a21bo_1 _1129_ (.A1(_0449_),
    .A2(_0464_),
    .B1_N(_0506_),
    .X(_0507_));
 sky130_fd_sc_hd__a21o_1 _1130_ (.A1(\MOS6502.op[1] ),
    .A2(_0421_),
    .B1(_0462_),
    .X(_0508_));
 sky130_fd_sc_hd__or2_1 _1131_ (.A(_0463_),
    .B(_0508_),
    .X(_0509_));
 sky130_fd_sc_hd__and2_1 _1132_ (.A(_0463_),
    .B(_0508_),
    .X(_0510_));
 sky130_fd_sc_hd__inv_2 _1133_ (.A(_0510_),
    .Y(_0511_));
 sky130_fd_sc_hd__and2b_1 _1134_ (.A_N(_0506_),
    .B(_0449_),
    .X(_0512_));
 sky130_fd_sc_hd__mux2_1 _1135_ (.A0(_0509_),
    .A1(_0511_),
    .S(_0512_),
    .X(_0513_));
 sky130_fd_sc_hd__or2_1 _1136_ (.A(\MOS6502.AXYS[2][6] ),
    .B(_0493_),
    .X(_0514_));
 sky130_fd_sc_hd__o211a_1 _1137_ (.A1(\MOS6502.AXYS[3][6] ),
    .A2(_0499_),
    .B1(_0496_),
    .C1(_0514_),
    .X(_0515_));
 sky130_fd_sc_hd__a221oi_4 _1138_ (.A1(\MOS6502.AXYS[0][6] ),
    .A2(_0497_),
    .B1(_0500_),
    .B2(\MOS6502.AXYS[1][6] ),
    .C1(_0515_),
    .Y(_0516_));
 sky130_fd_sc_hd__nor2_1 _1139_ (.A(_0482_),
    .B(_0516_),
    .Y(_0517_));
 sky130_fd_sc_hd__a221o_1 _1140_ (.A1(\MOS6502.ABH[6] ),
    .A2(_0465_),
    .B1(_0470_),
    .B2(\MOS6502.ADD[6] ),
    .C1(_0517_),
    .X(_0518_));
 sky130_fd_sc_hd__a21oi_1 _1141_ (.A1(net7),
    .A2(_0442_),
    .B1(_0518_),
    .Y(_0519_));
 sky130_fd_sc_hd__nor2_1 _1142_ (.A(_0456_),
    .B(_0519_),
    .Y(_0520_));
 sky130_fd_sc_hd__a31o_1 _1143_ (.A1(_0456_),
    .A2(_0507_),
    .A3(_0513_),
    .B1(_0520_),
    .X(_0521_));
 sky130_fd_sc_hd__or2b_1 _1144_ (.A(_0454_),
    .B_N(_0521_),
    .X(_0522_));
 sky130_fd_sc_hd__or2_1 _1145_ (.A(\MOS6502.AXYS[2][4] ),
    .B(_0493_),
    .X(_0523_));
 sky130_fd_sc_hd__o211a_1 _1146_ (.A1(\MOS6502.AXYS[3][4] ),
    .A2(_0499_),
    .B1(_0496_),
    .C1(_0523_),
    .X(_0524_));
 sky130_fd_sc_hd__a221oi_4 _1147_ (.A1(\MOS6502.AXYS[0][4] ),
    .A2(_0497_),
    .B1(_0500_),
    .B2(\MOS6502.AXYS[1][4] ),
    .C1(_0524_),
    .Y(_0525_));
 sky130_fd_sc_hd__a22o_1 _1148_ (.A1(net5),
    .A2(_0442_),
    .B1(_0465_),
    .B2(\MOS6502.ABH[4] ),
    .X(_0526_));
 sky130_fd_sc_hd__a21oi_1 _1149_ (.A1(\MOS6502.ADD[4] ),
    .A2(_0470_),
    .B1(_0526_),
    .Y(_0527_));
 sky130_fd_sc_hd__o21a_1 _1150_ (.A1(_0482_),
    .A2(_0525_),
    .B1(_0527_),
    .X(_0528_));
 sky130_fd_sc_hd__a22o_1 _1151_ (.A1(\MOS6502.PC[4] ),
    .A2(_0429_),
    .B1(_0448_),
    .B2(net5),
    .X(_0529_));
 sky130_fd_sc_hd__nand2_1 _1152_ (.A(_0464_),
    .B(_0529_),
    .Y(_0530_));
 sky130_fd_sc_hd__o21ai_1 _1153_ (.A1(_0528_),
    .A2(_0530_),
    .B1(_0509_),
    .Y(_0531_));
 sky130_fd_sc_hd__or3b_1 _1154_ (.A(_0508_),
    .B(_0528_),
    .C_N(_0529_),
    .X(_0532_));
 sky130_fd_sc_hd__a22o_1 _1155_ (.A1(_0528_),
    .A2(_0530_),
    .B1(_0531_),
    .B2(_0532_),
    .X(_0533_));
 sky130_fd_sc_hd__mux2_1 _1156_ (.A0(_0506_),
    .A1(_0533_),
    .S(_0456_),
    .X(_0534_));
 sky130_fd_sc_hd__or2_2 _1157_ (.A(_0427_),
    .B(_0453_),
    .X(_0535_));
 sky130_fd_sc_hd__mux2_1 _1158_ (.A0(_0535_),
    .A1(_0424_),
    .S(_0529_),
    .X(_0536_));
 sky130_fd_sc_hd__nor2_1 _1159_ (.A(_0534_),
    .B(_0536_),
    .Y(_0537_));
 sky130_fd_sc_hd__or2_1 _1160_ (.A(\MOS6502.AXYS[2][3] ),
    .B(_0493_),
    .X(_0538_));
 sky130_fd_sc_hd__o211a_1 _1161_ (.A1(\MOS6502.AXYS[3][3] ),
    .A2(_0499_),
    .B1(_0496_),
    .C1(_0538_),
    .X(_0539_));
 sky130_fd_sc_hd__a221oi_4 _1162_ (.A1(\MOS6502.AXYS[0][3] ),
    .A2(_0497_),
    .B1(_0500_),
    .B2(\MOS6502.AXYS[1][3] ),
    .C1(_0539_),
    .Y(_0540_));
 sky130_fd_sc_hd__a22o_1 _1163_ (.A1(net4),
    .A2(_0442_),
    .B1(_0465_),
    .B2(\MOS6502.ABH[3] ),
    .X(_0541_));
 sky130_fd_sc_hd__a21oi_1 _1164_ (.A1(\MOS6502.ADD[3] ),
    .A2(_0470_),
    .B1(_0541_),
    .Y(_0542_));
 sky130_fd_sc_hd__o21a_1 _1165_ (.A1(_0482_),
    .A2(_0540_),
    .B1(_0542_),
    .X(_0543_));
 sky130_fd_sc_hd__a21oi_2 _1166_ (.A1(\MOS6502.op[1] ),
    .A2(_0421_),
    .B1(_0462_),
    .Y(_0544_));
 sky130_fd_sc_hd__a22o_1 _1167_ (.A1(\MOS6502.PC[3] ),
    .A2(_0429_),
    .B1(_0448_),
    .B2(net4),
    .X(_0545_));
 sky130_fd_sc_hd__nand2_1 _1168_ (.A(_0544_),
    .B(_0545_),
    .Y(_0546_));
 sky130_fd_sc_hd__nand2_1 _1169_ (.A(_0464_),
    .B(_0545_),
    .Y(_0547_));
 sky130_fd_sc_hd__o21ai_1 _1170_ (.A1(_0543_),
    .A2(_0547_),
    .B1(_0509_),
    .Y(_0548_));
 sky130_fd_sc_hd__o21a_1 _1171_ (.A1(_0543_),
    .A2(_0546_),
    .B1(_0548_),
    .X(_0549_));
 sky130_fd_sc_hd__and2_1 _1172_ (.A(\MOS6502.shift_right ),
    .B(_0421_),
    .X(_0550_));
 sky130_fd_sc_hd__a21o_1 _1173_ (.A1(_0543_),
    .A2(_0547_),
    .B1(_0550_),
    .X(_0551_));
 sky130_fd_sc_hd__o22a_1 _1174_ (.A1(_0456_),
    .A2(_0528_),
    .B1(_0549_),
    .B2(_0551_),
    .X(_0552_));
 sky130_fd_sc_hd__mux2_1 _1175_ (.A0(_0535_),
    .A1(_0424_),
    .S(_0545_),
    .X(_0553_));
 sky130_fd_sc_hd__clkinv_2 _1176_ (.A(_0553_),
    .Y(_0554_));
 sky130_fd_sc_hd__or2_1 _1177_ (.A(_0426_),
    .B(_0553_),
    .X(_0555_));
 sky130_fd_sc_hd__mux2_1 _1178_ (.A0(_0554_),
    .A1(_0555_),
    .S(_0552_),
    .X(_0556_));
 sky130_fd_sc_hd__a22oi_4 _1179_ (.A1(\MOS6502.PC[0] ),
    .A2(_0429_),
    .B1(_0448_),
    .B2(net1),
    .Y(_0557_));
 sky130_fd_sc_hd__mux2_1 _1180_ (.A0(_0424_),
    .A1(_0535_),
    .S(_0557_),
    .X(_0558_));
 sky130_fd_sc_hd__and3_1 _1181_ (.A(\MOS6502.AXYS[1][0] ),
    .B(_0490_),
    .C(_0492_),
    .X(_0559_));
 sky130_fd_sc_hd__a21oi_1 _1182_ (.A1(\MOS6502.AXYS[0][0] ),
    .A2(_0498_),
    .B1(_0559_),
    .Y(_0560_));
 sky130_fd_sc_hd__a21o_1 _1183_ (.A1(_0490_),
    .A2(_0492_),
    .B1(\MOS6502.AXYS[2][0] ),
    .X(_0561_));
 sky130_fd_sc_hd__o21ai_1 _1184_ (.A1(\MOS6502.AXYS[3][0] ),
    .A2(_0498_),
    .B1(_0561_),
    .Y(_0562_));
 sky130_fd_sc_hd__mux2_1 _1185_ (.A0(_0560_),
    .A1(_0562_),
    .S(_0495_),
    .X(_0563_));
 sky130_fd_sc_hd__a22o_1 _1186_ (.A1(net1),
    .A2(_0442_),
    .B1(_0423_),
    .B2(\MOS6502.ABH[0] ),
    .X(_0564_));
 sky130_fd_sc_hd__a21oi_1 _1187_ (.A1(\MOS6502.ADD[0] ),
    .A2(_0470_),
    .B1(_0564_),
    .Y(_0565_));
 sky130_fd_sc_hd__o21a_1 _1188_ (.A1(_0482_),
    .A2(_0563_),
    .B1(_0565_),
    .X(_0566_));
 sky130_fd_sc_hd__o21ai_1 _1189_ (.A1(_0557_),
    .A2(_0566_),
    .B1(_0464_),
    .Y(_0567_));
 sky130_fd_sc_hd__a211o_1 _1190_ (.A1(_0544_),
    .A2(_0557_),
    .B1(_0566_),
    .C1(_0510_),
    .X(_0568_));
 sky130_fd_sc_hd__a221o_1 _1191_ (.A1(_0557_),
    .A2(_0566_),
    .B1(_0567_),
    .B2(_0568_),
    .C1(_0550_),
    .X(_0569_));
 sky130_fd_sc_hd__inv_2 _1192_ (.A(_0482_),
    .Y(_0570_));
 sky130_fd_sc_hd__mux2_1 _1193_ (.A0(\MOS6502.AXYS[1][1] ),
    .A1(\MOS6502.AXYS[0][1] ),
    .S(_0498_),
    .X(_0571_));
 sky130_fd_sc_hd__mux2_1 _1194_ (.A0(\MOS6502.AXYS[3][1] ),
    .A1(\MOS6502.AXYS[2][1] ),
    .S(_0498_),
    .X(_0572_));
 sky130_fd_sc_hd__mux2_1 _1195_ (.A0(_0571_),
    .A1(_0572_),
    .S(_0495_),
    .X(_0573_));
 sky130_fd_sc_hd__a22o_1 _1196_ (.A1(net2),
    .A2(_0442_),
    .B1(_0423_),
    .B2(\MOS6502.ABH[1] ),
    .X(_0574_));
 sky130_fd_sc_hd__a21o_1 _1197_ (.A1(\MOS6502.ADD[1] ),
    .A2(_0470_),
    .B1(_0574_),
    .X(_0575_));
 sky130_fd_sc_hd__a21oi_1 _1198_ (.A1(_0570_),
    .A2(_0573_),
    .B1(_0575_),
    .Y(_0576_));
 sky130_fd_sc_hd__or2_1 _1199_ (.A(_0455_),
    .B(_0576_),
    .X(_0577_));
 sky130_fd_sc_hd__o211ai_1 _1200_ (.A1(_0426_),
    .A2(_0558_),
    .B1(_0569_),
    .C1(_0577_),
    .Y(_0578_));
 sky130_fd_sc_hd__inv_2 _1201_ (.A(\MOS6502.load_only ),
    .Y(_0579_));
 sky130_fd_sc_hd__inv_2 _1202_ (.A(\MOS6502.shift ),
    .Y(_0580_));
 sky130_fd_sc_hd__a32o_1 _1203_ (.A1(_0579_),
    .A2(_0580_),
    .A3(_0415_),
    .B1(_0421_),
    .B2(\MOS6502.rotate ),
    .X(_0581_));
 sky130_fd_sc_hd__nand2_1 _1204_ (.A(\MOS6502.C ),
    .B(_0581_),
    .Y(_0582_));
 sky130_fd_sc_hd__inv_2 _1205_ (.A(\MOS6502.rotate ),
    .Y(_0583_));
 sky130_fd_sc_hd__a32o_1 _1206_ (.A1(_0580_),
    .A2(\MOS6502.inc ),
    .A3(_0419_),
    .B1(_0415_),
    .B2(\MOS6502.compare ),
    .X(_0584_));
 sky130_fd_sc_hd__nor2_1 _1207_ (.A(_0398_),
    .B(_0416_),
    .Y(_0585_));
 sky130_fd_sc_hd__nor2_1 _1208_ (.A(_0365_),
    .B(_0400_),
    .Y(_0586_));
 sky130_fd_sc_hd__or2_1 _1209_ (.A(_0585_),
    .B(_0586_),
    .X(_0587_));
 sky130_fd_sc_hd__o21a_1 _1210_ (.A1(_0465_),
    .A2(_0587_),
    .B1(\MOS6502.ALU.CO ),
    .X(_0588_));
 sky130_fd_sc_hd__a21oi_1 _1211_ (.A1(_0385_),
    .A2(_0393_),
    .B1(_0410_),
    .Y(_0589_));
 sky130_fd_sc_hd__or4b_1 _1212_ (.A(_0471_),
    .B(_0588_),
    .C(_0589_),
    .D_N(_0468_),
    .X(_0590_));
 sky130_fd_sc_hd__a21oi_1 _1213_ (.A1(_0583_),
    .A2(_0584_),
    .B1(_0590_),
    .Y(_0591_));
 sky130_fd_sc_hd__nand2_1 _1214_ (.A(_0582_),
    .B(_0591_),
    .Y(_0592_));
 sky130_fd_sc_hd__nor2_1 _1215_ (.A(_0550_),
    .B(_0453_),
    .Y(_0593_));
 sky130_fd_sc_hd__a21oi_1 _1216_ (.A1(_0577_),
    .A2(_0569_),
    .B1(_0558_),
    .Y(_0594_));
 sky130_fd_sc_hd__a31o_1 _1217_ (.A1(_0578_),
    .A2(_0592_),
    .A3(_0593_),
    .B1(_0594_),
    .X(_0595_));
 sky130_fd_sc_hd__clkinv_2 _1218_ (.A(_0535_),
    .Y(_0596_));
 sky130_fd_sc_hd__a22o_1 _1219_ (.A1(\MOS6502.PC[1] ),
    .A2(_0429_),
    .B1(_0448_),
    .B2(net2),
    .X(_0597_));
 sky130_fd_sc_hd__mux2_1 _1220_ (.A0(_0596_),
    .A1(_0451_),
    .S(_0597_),
    .X(_0598_));
 sky130_fd_sc_hd__nor2_1 _1221_ (.A(_0464_),
    .B(_0544_),
    .Y(_0599_));
 sky130_fd_sc_hd__and2b_1 _1222_ (.A_N(_0576_),
    .B(_0597_),
    .X(_0600_));
 sky130_fd_sc_hd__mux2_1 _1223_ (.A0(_0464_),
    .A1(_0544_),
    .S(_0600_),
    .X(_0601_));
 sky130_fd_sc_hd__a21bo_1 _1224_ (.A1(_0464_),
    .A2(_0597_),
    .B1_N(_0576_),
    .X(_0602_));
 sky130_fd_sc_hd__o211a_1 _1225_ (.A1(_0599_),
    .A2(_0601_),
    .B1(_0602_),
    .C1(_0455_),
    .X(_0603_));
 sky130_fd_sc_hd__and3_1 _1226_ (.A(\MOS6502.AXYS[1][2] ),
    .B(_0490_),
    .C(_0492_),
    .X(_0604_));
 sky130_fd_sc_hd__a21oi_1 _1227_ (.A1(\MOS6502.AXYS[0][2] ),
    .A2(_0499_),
    .B1(_0604_),
    .Y(_0605_));
 sky130_fd_sc_hd__a21o_1 _1228_ (.A1(_0490_),
    .A2(_0492_),
    .B1(\MOS6502.AXYS[2][2] ),
    .X(_0606_));
 sky130_fd_sc_hd__o21ai_1 _1229_ (.A1(\MOS6502.AXYS[3][2] ),
    .A2(_0499_),
    .B1(_0606_),
    .Y(_0607_));
 sky130_fd_sc_hd__mux2_1 _1230_ (.A0(_0605_),
    .A1(_0607_),
    .S(_0495_),
    .X(_0608_));
 sky130_fd_sc_hd__a22o_1 _1231_ (.A1(net3),
    .A2(_0442_),
    .B1(_0423_),
    .B2(\MOS6502.ABH[2] ),
    .X(_0609_));
 sky130_fd_sc_hd__a21oi_1 _1232_ (.A1(\MOS6502.ADD[2] ),
    .A2(_0470_),
    .B1(_0609_),
    .Y(_0610_));
 sky130_fd_sc_hd__o21a_1 _1233_ (.A1(_0482_),
    .A2(_0608_),
    .B1(_0610_),
    .X(_0611_));
 sky130_fd_sc_hd__nor2_1 _1234_ (.A(_0456_),
    .B(_0611_),
    .Y(_0612_));
 sky130_fd_sc_hd__a211o_1 _1235_ (.A1(_0452_),
    .A2(_0598_),
    .B1(_0603_),
    .C1(_0612_),
    .X(_0613_));
 sky130_fd_sc_hd__o21a_1 _1236_ (.A1(_0612_),
    .A2(_0603_),
    .B1(_0598_),
    .X(_0614_));
 sky130_fd_sc_hd__a21oi_1 _1237_ (.A1(_0595_),
    .A2(_0613_),
    .B1(_0614_),
    .Y(_0615_));
 sky130_fd_sc_hd__a22o_1 _1238_ (.A1(\MOS6502.PC[2] ),
    .A2(_0429_),
    .B1(_0448_),
    .B2(net3),
    .X(_0616_));
 sky130_fd_sc_hd__nor2_1 _1239_ (.A(_0508_),
    .B(_0611_),
    .Y(_0617_));
 sky130_fd_sc_hd__nand2_1 _1240_ (.A(_0463_),
    .B(_0616_),
    .Y(_0618_));
 sky130_fd_sc_hd__o21a_1 _1241_ (.A1(_0611_),
    .A2(_0618_),
    .B1(_0509_),
    .X(_0619_));
 sky130_fd_sc_hd__a21oi_1 _1242_ (.A1(_0616_),
    .A2(_0617_),
    .B1(_0619_),
    .Y(_0620_));
 sky130_fd_sc_hd__a21o_1 _1243_ (.A1(_0611_),
    .A2(_0618_),
    .B1(_0550_),
    .X(_0621_));
 sky130_fd_sc_hd__o22a_1 _1244_ (.A1(_0456_),
    .A2(_0543_),
    .B1(_0620_),
    .B2(_0621_),
    .X(_0622_));
 sky130_fd_sc_hd__mux2_1 _1245_ (.A0(_0535_),
    .A1(_0424_),
    .S(_0616_),
    .X(_0623_));
 sky130_fd_sc_hd__or2_1 _1246_ (.A(_0622_),
    .B(_0623_),
    .X(_0624_));
 sky130_fd_sc_hd__o21ai_1 _1247_ (.A1(_0426_),
    .A2(_0623_),
    .B1(_0622_),
    .Y(_0625_));
 sky130_fd_sc_hd__nand2_1 _1248_ (.A(_0624_),
    .B(_0625_),
    .Y(_0626_));
 sky130_fd_sc_hd__o21a_1 _1249_ (.A1(_0615_),
    .A2(_0626_),
    .B1(_0624_),
    .X(_0627_));
 sky130_fd_sc_hd__o22a_1 _1250_ (.A1(_0552_),
    .A2(_0553_),
    .B1(_0556_),
    .B2(_0627_),
    .X(_0628_));
 sky130_fd_sc_hd__xor2_1 _1251_ (.A(_0615_),
    .B(_0626_),
    .X(\MOS6502.ALU.temp[2] ));
 sky130_fd_sc_hd__or2b_1 _1252_ (.A(_0614_),
    .B_N(_0613_),
    .X(_0629_));
 sky130_fd_sc_hd__xnor2_1 _1253_ (.A(_0595_),
    .B(_0629_),
    .Y(\MOS6502.ALU.temp[1] ));
 sky130_fd_sc_hd__o211ai_1 _1254_ (.A1(_0615_),
    .A2(_0626_),
    .B1(_0556_),
    .C1(_0624_),
    .Y(_0630_));
 sky130_fd_sc_hd__and2_1 _1255_ (.A(\MOS6502.adc_bcd ),
    .B(_0415_),
    .X(_0631_));
 sky130_fd_sc_hd__o211ai_2 _1256_ (.A1(\MOS6502.ALU.temp[2] ),
    .A2(\MOS6502.ALU.temp[1] ),
    .B1(_0630_),
    .C1(_0631_),
    .Y(_0632_));
 sky130_fd_sc_hd__o21a_1 _1257_ (.A1(_0426_),
    .A2(_0536_),
    .B1(_0534_),
    .X(_0633_));
 sky130_fd_sc_hd__or2_1 _1258_ (.A(_0537_),
    .B(_0633_),
    .X(_0634_));
 sky130_fd_sc_hd__a21oi_1 _1259_ (.A1(_0628_),
    .A2(_0632_),
    .B1(_0634_),
    .Y(_0635_));
 sky130_fd_sc_hd__o21bai_1 _1260_ (.A1(_0426_),
    .A2(_0454_),
    .B1_N(_0521_),
    .Y(_0636_));
 sky130_fd_sc_hd__o211ai_1 _1261_ (.A1(_0537_),
    .A2(_0635_),
    .B1(_0636_),
    .C1(_0522_),
    .Y(_0637_));
 sky130_fd_sc_hd__or2_1 _1262_ (.A(\MOS6502.AXYS[2][7] ),
    .B(_0493_),
    .X(_0638_));
 sky130_fd_sc_hd__o211a_1 _1263_ (.A1(\MOS6502.AXYS[3][7] ),
    .A2(_0499_),
    .B1(_0496_),
    .C1(_0638_),
    .X(_0639_));
 sky130_fd_sc_hd__a221oi_4 _1264_ (.A1(\MOS6502.AXYS[0][7] ),
    .A2(_0497_),
    .B1(_0500_),
    .B2(\MOS6502.AXYS[1][7] ),
    .C1(_0639_),
    .Y(_0640_));
 sky130_fd_sc_hd__nor2_1 _1265_ (.A(_0482_),
    .B(_0640_),
    .Y(_0641_));
 sky130_fd_sc_hd__a22o_1 _1266_ (.A1(net8),
    .A2(_0442_),
    .B1(_0465_),
    .B2(\MOS6502.ABH[7] ),
    .X(_0642_));
 sky130_fd_sc_hd__a211o_1 _1267_ (.A1(\MOS6502.ADD[7] ),
    .A2(_0470_),
    .B1(_0641_),
    .C1(_0642_),
    .X(_0643_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _1268_ (.A(_0643_),
    .X(\MOS6502.AI[7] ));
 sky130_fd_sc_hd__a22o_1 _1269_ (.A1(\MOS6502.PC[6] ),
    .A2(_0429_),
    .B1(_0448_),
    .B2(net7),
    .X(_0644_));
 sky130_fd_sc_hd__and2b_1 _1270_ (.A_N(_0519_),
    .B(_0644_),
    .X(_0645_));
 sky130_fd_sc_hd__mux2_1 _1271_ (.A0(_0464_),
    .A1(_0544_),
    .S(_0645_),
    .X(_0646_));
 sky130_fd_sc_hd__a21bo_1 _1272_ (.A1(_0464_),
    .A2(_0644_),
    .B1_N(_0519_),
    .X(_0647_));
 sky130_fd_sc_hd__o211a_1 _1273_ (.A1(_0599_),
    .A2(_0646_),
    .B1(_0647_),
    .C1(_0456_),
    .X(_0648_));
 sky130_fd_sc_hd__a21oi_1 _1274_ (.A1(_0550_),
    .A2(\MOS6502.AI[7] ),
    .B1(_0648_),
    .Y(_0649_));
 sky130_fd_sc_hd__mux2_1 _1275_ (.A0(_0427_),
    .A1(_0424_),
    .S(_0644_),
    .X(_0650_));
 sky130_fd_sc_hd__or2_1 _1276_ (.A(_0426_),
    .B(_0650_),
    .X(_0651_));
 sky130_fd_sc_hd__or3_1 _1277_ (.A(_0453_),
    .B(_0649_),
    .C(_0650_),
    .X(_0652_));
 sky130_fd_sc_hd__a21bo_1 _1278_ (.A1(_0649_),
    .A2(_0651_),
    .B1_N(_0652_),
    .X(_0653_));
 sky130_fd_sc_hd__a21o_1 _1279_ (.A1(_0522_),
    .A2(_0637_),
    .B1(_0653_),
    .X(_0654_));
 sky130_fd_sc_hd__nand3_1 _1280_ (.A(_0522_),
    .B(_0637_),
    .C(_0653_),
    .Y(_0655_));
 sky130_fd_sc_hd__and2_1 _1281_ (.A(_0654_),
    .B(_0655_),
    .X(_0656_));
 sky130_fd_sc_hd__clkbuf_1 _1282_ (.A(_0656_),
    .X(\MOS6502.ALU.temp[6] ));
 sky130_fd_sc_hd__nand2_1 _1283_ (.A(_0628_),
    .B(_0632_),
    .Y(\MOS6502.ALU.temp_HC ));
 sky130_fd_sc_hd__a22o_1 _1284_ (.A1(\MOS6502.PC[7] ),
    .A2(_0429_),
    .B1(_0448_),
    .B2(net8),
    .X(_0657_));
 sky130_fd_sc_hd__a21oi_1 _1285_ (.A1(_0464_),
    .A2(_0657_),
    .B1(\MOS6502.AI[7] ),
    .Y(_0658_));
 sky130_fd_sc_hd__o21ai_1 _1286_ (.A1(_0509_),
    .A2(_0657_),
    .B1(_0456_),
    .Y(_0659_));
 sky130_fd_sc_hd__a31o_1 _1287_ (.A1(_0510_),
    .A2(\MOS6502.AI[7] ),
    .A3(_0657_),
    .B1(_0659_),
    .X(_0660_));
 sky130_fd_sc_hd__o2bb2a_1 _1288_ (.A1_N(_0550_),
    .A2_N(_0592_),
    .B1(_0658_),
    .B2(_0660_),
    .X(_0661_));
 sky130_fd_sc_hd__mux2_1 _1289_ (.A0(_0535_),
    .A1(_0424_),
    .S(_0657_),
    .X(_0662_));
 sky130_fd_sc_hd__or2_1 _1290_ (.A(_0661_),
    .B(_0662_),
    .X(_0663_));
 sky130_fd_sc_hd__o21ai_1 _1291_ (.A1(_0426_),
    .A2(_0662_),
    .B1(_0661_),
    .Y(_0664_));
 sky130_fd_sc_hd__nand2_1 _1292_ (.A(_0663_),
    .B(_0664_),
    .Y(_0665_));
 sky130_fd_sc_hd__a21o_1 _1293_ (.A1(_0652_),
    .A2(_0654_),
    .B1(_0665_),
    .X(_0666_));
 sky130_fd_sc_hd__nand3_1 _1294_ (.A(_0652_),
    .B(_0654_),
    .C(_0665_),
    .Y(_0667_));
 sky130_fd_sc_hd__and2_1 _1295_ (.A(_0666_),
    .B(_0667_),
    .X(_0668_));
 sky130_fd_sc_hd__clkbuf_1 _1296_ (.A(_0668_),
    .X(\MOS6502.ALU.temp[7] ));
 sky130_fd_sc_hd__a211o_1 _1297_ (.A1(_0663_),
    .A2(_0666_),
    .B1(_0456_),
    .C1(_0566_),
    .X(_0669_));
 sky130_fd_sc_hd__o211ai_1 _1298_ (.A1(_0456_),
    .A2(_0566_),
    .B1(_0663_),
    .C1(_0666_),
    .Y(_0670_));
 sky130_fd_sc_hd__a211o_1 _1299_ (.A1(_0522_),
    .A2(_0636_),
    .B1(_0635_),
    .C1(_0537_),
    .X(_0671_));
 sky130_fd_sc_hd__and2_1 _1300_ (.A(_0637_),
    .B(_0671_),
    .X(_0672_));
 sky130_fd_sc_hd__clkbuf_1 _1301_ (.A(_0672_),
    .X(\MOS6502.ALU.temp[5] ));
 sky130_fd_sc_hd__o2111a_1 _1302_ (.A1(\MOS6502.ALU.temp[6] ),
    .A2(\MOS6502.ALU.temp[5] ),
    .B1(_0666_),
    .C1(_0631_),
    .D1(_0667_),
    .X(_0673_));
 sky130_fd_sc_hd__a21o_1 _1303_ (.A1(_0669_),
    .A2(_0670_),
    .B1(_0673_),
    .X(_0001_));
 sky130_fd_sc_hd__and2_1 _1304_ (.A(\MOS6502.D ),
    .B(\MOS6502.adc_sbc ),
    .X(_0674_));
 sky130_fd_sc_hd__clkbuf_1 _1305_ (.A(_0674_),
    .X(_0000_));
 sky130_fd_sc_hd__and2b_1 _1306_ (.A_N(_0594_),
    .B(_0578_),
    .X(_0675_));
 sky130_fd_sc_hd__nand2_1 _1307_ (.A(_0592_),
    .B(_0593_),
    .Y(_0676_));
 sky130_fd_sc_hd__xnor2_1 _1308_ (.A(_0675_),
    .B(_0676_),
    .Y(\MOS6502.ALU.temp[0] ));
 sky130_fd_sc_hd__buf_2 _1309_ (.A(_0381_),
    .X(_0677_));
 sky130_fd_sc_hd__clkbuf_4 _1310_ (.A(_0461_),
    .X(_0678_));
 sky130_fd_sc_hd__nor2_1 _1311_ (.A(\MOS6502.state[5] ),
    .B(_0438_),
    .Y(_0679_));
 sky130_fd_sc_hd__and2_1 _1312_ (.A(_0365_),
    .B(_0383_),
    .X(_0680_));
 sky130_fd_sc_hd__nor2_1 _1313_ (.A(_0375_),
    .B(_0680_),
    .Y(_0681_));
 sky130_fd_sc_hd__nor2_1 _1314_ (.A(_0414_),
    .B(_0680_),
    .Y(_0682_));
 sky130_fd_sc_hd__a211o_2 _1315_ (.A1(_0404_),
    .A2(_0679_),
    .B1(_0681_),
    .C1(_0682_),
    .X(_0683_));
 sky130_fd_sc_hd__or2_1 _1316_ (.A(_0423_),
    .B(_0683_),
    .X(_0684_));
 sky130_fd_sc_hd__buf_2 _1317_ (.A(_0684_),
    .X(_0685_));
 sky130_fd_sc_hd__nand2_2 _1318_ (.A(_0356_),
    .B(_0461_),
    .Y(_0686_));
 sky130_fd_sc_hd__o31ai_2 _1319_ (.A1(_0677_),
    .A2(_0678_),
    .A3(_0685_),
    .B1(_0686_),
    .Y(_0687_));
 sky130_fd_sc_hd__or4_1 _1320_ (.A(_0369_),
    .B(_0378_),
    .C(_0373_),
    .D(_0407_),
    .X(_0688_));
 sky130_fd_sc_hd__clkbuf_4 _1321_ (.A(_0688_),
    .X(_0689_));
 sky130_fd_sc_hd__nor2_4 _1322_ (.A(_0356_),
    .B(_0689_),
    .Y(_0690_));
 sky130_fd_sc_hd__a22o_1 _1323_ (.A1(\MOS6502.ADD[0] ),
    .A2(_0684_),
    .B1(_0690_),
    .B2(\MOS6502.ABL[0] ),
    .X(_0691_));
 sky130_fd_sc_hd__a21oi_1 _1324_ (.A1(\MOS6502.PC[0] ),
    .A2(_0687_),
    .B1(_0691_),
    .Y(_0692_));
 sky130_fd_sc_hd__nor2_1 _1325_ (.A(_0681_),
    .B(_0679_),
    .Y(_0693_));
 sky130_fd_sc_hd__or3_1 _1326_ (.A(_0378_),
    .B(_0367_),
    .C(_0379_),
    .X(_0694_));
 sky130_fd_sc_hd__and3_1 _1327_ (.A(_0371_),
    .B(_0428_),
    .C(_0694_),
    .X(_0695_));
 sky130_fd_sc_hd__xnor2_1 _1328_ (.A(\MOS6502.backwards ),
    .B(\MOS6502.ALU.CO ),
    .Y(_0696_));
 sky130_fd_sc_hd__nand2_1 _1329_ (.A(_0423_),
    .B(_0696_),
    .Y(_0697_));
 sky130_fd_sc_hd__o211a_1 _1330_ (.A1(_0398_),
    .A2(_0695_),
    .B1(_0697_),
    .C1(_0686_),
    .X(_0698_));
 sky130_fd_sc_hd__o211a_1 _1331_ (.A1(_0404_),
    .A2(_0414_),
    .B1(_0693_),
    .C1(_0698_),
    .X(_0699_));
 sky130_fd_sc_hd__xor2_1 _1332_ (.A(_0692_),
    .B(_0699_),
    .X(_0002_));
 sky130_fd_sc_hd__or2_1 _1333_ (.A(_0692_),
    .B(_0699_),
    .X(_0700_));
 sky130_fd_sc_hd__or2_1 _1334_ (.A(_0398_),
    .B(_0380_),
    .X(_0701_));
 sky130_fd_sc_hd__a2bb2o_1 _1335_ (.A1_N(\MOS6502.res ),
    .A2_N(_0701_),
    .B1(_0685_),
    .B2(\MOS6502.ADD[1] ),
    .X(_0702_));
 sky130_fd_sc_hd__a221o_1 _1336_ (.A1(\MOS6502.PC[1] ),
    .A2(_0687_),
    .B1(_0690_),
    .B2(\MOS6502.ABL[1] ),
    .C1(_0702_),
    .X(_0703_));
 sky130_fd_sc_hd__and2b_1 _1337_ (.A_N(_0700_),
    .B(_0703_),
    .X(_0704_));
 sky130_fd_sc_hd__and2b_1 _1338_ (.A_N(_0703_),
    .B(_0700_),
    .X(_0705_));
 sky130_fd_sc_hd__nor2_1 _1339_ (.A(_0704_),
    .B(_0705_),
    .Y(_0009_));
 sky130_fd_sc_hd__inv_2 _1340_ (.A(\MOS6502.NMI_edge ),
    .Y(_0706_));
 sky130_fd_sc_hd__o21a_1 _1341_ (.A1(_0706_),
    .A2(\MOS6502.res ),
    .B1(_0677_),
    .X(_0707_));
 sky130_fd_sc_hd__a22o_1 _1342_ (.A1(\MOS6502.ADD[2] ),
    .A2(_0685_),
    .B1(_0687_),
    .B2(\MOS6502.PC[2] ),
    .X(_0708_));
 sky130_fd_sc_hd__a211oi_2 _1343_ (.A1(\MOS6502.ABL[2] ),
    .A2(_0690_),
    .B1(_0707_),
    .C1(_0708_),
    .Y(_0709_));
 sky130_fd_sc_hd__xnor2_1 _1344_ (.A(_0704_),
    .B(_0709_),
    .Y(_0010_));
 sky130_fd_sc_hd__or3b_1 _1345_ (.A(_0709_),
    .B(_0700_),
    .C_N(_0703_),
    .X(_0710_));
 sky130_fd_sc_hd__o21ai_2 _1346_ (.A1(_0678_),
    .A2(_0685_),
    .B1(_0686_),
    .Y(_0711_));
 sky130_fd_sc_hd__a221o_1 _1347_ (.A1(\MOS6502.ADD[3] ),
    .A2(_0685_),
    .B1(_0690_),
    .B2(\MOS6502.ABL[3] ),
    .C1(_0677_),
    .X(_0712_));
 sky130_fd_sc_hd__a21oi_1 _1348_ (.A1(\MOS6502.PC[3] ),
    .A2(_0711_),
    .B1(_0712_),
    .Y(_0713_));
 sky130_fd_sc_hd__xor2_1 _1349_ (.A(_0710_),
    .B(_0713_),
    .X(_0011_));
 sky130_fd_sc_hd__or2_1 _1350_ (.A(_0710_),
    .B(_0713_),
    .X(_0714_));
 sky130_fd_sc_hd__a221o_1 _1351_ (.A1(\MOS6502.ADD[4] ),
    .A2(_0685_),
    .B1(_0690_),
    .B2(\MOS6502.ABL[4] ),
    .C1(_0677_),
    .X(_0715_));
 sky130_fd_sc_hd__a21oi_1 _1352_ (.A1(\MOS6502.PC[4] ),
    .A2(_0711_),
    .B1(_0715_),
    .Y(_0716_));
 sky130_fd_sc_hd__xor2_1 _1353_ (.A(_0714_),
    .B(_0716_),
    .X(_0012_));
 sky130_fd_sc_hd__or2_1 _1354_ (.A(_0714_),
    .B(_0716_),
    .X(_0717_));
 sky130_fd_sc_hd__a221o_1 _1355_ (.A1(\MOS6502.ADD[5] ),
    .A2(_0685_),
    .B1(_0690_),
    .B2(\MOS6502.ABL[5] ),
    .C1(_0677_),
    .X(_0718_));
 sky130_fd_sc_hd__a21oi_1 _1356_ (.A1(\MOS6502.PC[5] ),
    .A2(_0711_),
    .B1(_0718_),
    .Y(_0719_));
 sky130_fd_sc_hd__xor2_1 _1357_ (.A(_0717_),
    .B(_0719_),
    .X(_0013_));
 sky130_fd_sc_hd__or2_1 _1358_ (.A(_0717_),
    .B(_0719_),
    .X(_0720_));
 sky130_fd_sc_hd__a221o_1 _1359_ (.A1(\MOS6502.ADD[6] ),
    .A2(_0685_),
    .B1(_0690_),
    .B2(\MOS6502.ABL[6] ),
    .C1(_0677_),
    .X(_0721_));
 sky130_fd_sc_hd__a21oi_1 _1360_ (.A1(\MOS6502.PC[6] ),
    .A2(_0711_),
    .B1(_0721_),
    .Y(_0722_));
 sky130_fd_sc_hd__xor2_1 _1361_ (.A(_0720_),
    .B(_0722_),
    .X(_0014_));
 sky130_fd_sc_hd__or2_1 _1362_ (.A(_0720_),
    .B(_0722_),
    .X(_0723_));
 sky130_fd_sc_hd__buf_2 _1363_ (.A(_0677_),
    .X(_0724_));
 sky130_fd_sc_hd__a221o_1 _1364_ (.A1(\MOS6502.ADD[7] ),
    .A2(_0685_),
    .B1(_0690_),
    .B2(\MOS6502.ABL[7] ),
    .C1(_0724_),
    .X(_0725_));
 sky130_fd_sc_hd__a21oi_1 _1365_ (.A1(\MOS6502.PC[7] ),
    .A2(_0711_),
    .B1(_0725_),
    .Y(_0726_));
 sky130_fd_sc_hd__nor2_1 _1366_ (.A(_0723_),
    .B(_0726_),
    .Y(_0727_));
 sky130_fd_sc_hd__and2_1 _1367_ (.A(_0723_),
    .B(_0726_),
    .X(_0728_));
 sky130_fd_sc_hd__nor2_1 _1368_ (.A(_0727_),
    .B(_0728_),
    .Y(_0015_));
 sky130_fd_sc_hd__nor2_4 _1369_ (.A(_0398_),
    .B(_0438_),
    .Y(_0729_));
 sky130_fd_sc_hd__or4_1 _1370_ (.A(_0677_),
    .B(_0678_),
    .C(_0685_),
    .D(_0729_),
    .X(_0730_));
 sky130_fd_sc_hd__nand2_2 _1371_ (.A(_0686_),
    .B(_0730_),
    .Y(_0731_));
 sky130_fd_sc_hd__or2_2 _1372_ (.A(_0465_),
    .B(_0690_),
    .X(_0732_));
 sky130_fd_sc_hd__a221o_1 _1373_ (.A1(\MOS6502.ADD[0] ),
    .A2(_0729_),
    .B1(_0732_),
    .B2(\MOS6502.ABH[0] ),
    .C1(_0724_),
    .X(_0733_));
 sky130_fd_sc_hd__a221o_1 _1374_ (.A1(net1),
    .A2(_0683_),
    .B1(_0731_),
    .B2(\MOS6502.PC[8] ),
    .C1(_0733_),
    .X(_0734_));
 sky130_fd_sc_hd__xor2_1 _1375_ (.A(_0727_),
    .B(_0734_),
    .X(_0016_));
 sky130_fd_sc_hd__a221o_1 _1376_ (.A1(\MOS6502.ADD[1] ),
    .A2(_0729_),
    .B1(_0732_),
    .B2(\MOS6502.ABH[1] ),
    .C1(_0724_),
    .X(_0735_));
 sky130_fd_sc_hd__a221o_1 _1377_ (.A1(net2),
    .A2(_0683_),
    .B1(_0731_),
    .B2(\MOS6502.PC[9] ),
    .C1(_0735_),
    .X(_0736_));
 sky130_fd_sc_hd__and3_1 _1378_ (.A(_0727_),
    .B(_0734_),
    .C(_0736_),
    .X(_0737_));
 sky130_fd_sc_hd__a21oi_1 _1379_ (.A1(_0727_),
    .A2(_0734_),
    .B1(_0736_),
    .Y(_0738_));
 sky130_fd_sc_hd__nor2_1 _1380_ (.A(_0737_),
    .B(_0738_),
    .Y(_0017_));
 sky130_fd_sc_hd__a221o_1 _1381_ (.A1(\MOS6502.ADD[2] ),
    .A2(_0729_),
    .B1(_0732_),
    .B2(\MOS6502.ABH[2] ),
    .C1(_0724_),
    .X(_0739_));
 sky130_fd_sc_hd__a221o_1 _1382_ (.A1(net3),
    .A2(_0683_),
    .B1(_0731_),
    .B2(\MOS6502.PC[10] ),
    .C1(_0739_),
    .X(_0740_));
 sky130_fd_sc_hd__xor2_1 _1383_ (.A(_0737_),
    .B(_0740_),
    .X(_0003_));
 sky130_fd_sc_hd__a221o_1 _1384_ (.A1(\MOS6502.ADD[3] ),
    .A2(_0729_),
    .B1(_0732_),
    .B2(\MOS6502.ABH[3] ),
    .C1(_0724_),
    .X(_0741_));
 sky130_fd_sc_hd__a221o_1 _1385_ (.A1(net4),
    .A2(_0683_),
    .B1(_0731_),
    .B2(\MOS6502.PC[11] ),
    .C1(_0741_),
    .X(_0742_));
 sky130_fd_sc_hd__and3_1 _1386_ (.A(_0737_),
    .B(_0740_),
    .C(_0742_),
    .X(_0743_));
 sky130_fd_sc_hd__a21oi_1 _1387_ (.A1(_0737_),
    .A2(_0740_),
    .B1(_0742_),
    .Y(_0744_));
 sky130_fd_sc_hd__nor2_1 _1388_ (.A(_0743_),
    .B(_0744_),
    .Y(_0004_));
 sky130_fd_sc_hd__a221o_1 _1389_ (.A1(\MOS6502.ADD[4] ),
    .A2(_0729_),
    .B1(_0732_),
    .B2(\MOS6502.ABH[4] ),
    .C1(_0724_),
    .X(_0745_));
 sky130_fd_sc_hd__a221o_1 _1390_ (.A1(net5),
    .A2(_0683_),
    .B1(_0731_),
    .B2(\MOS6502.PC[12] ),
    .C1(_0745_),
    .X(_0746_));
 sky130_fd_sc_hd__xor2_1 _1391_ (.A(_0743_),
    .B(_0746_),
    .X(_0005_));
 sky130_fd_sc_hd__a221o_1 _1392_ (.A1(\MOS6502.ADD[5] ),
    .A2(_0729_),
    .B1(_0732_),
    .B2(\MOS6502.ABH[5] ),
    .C1(_0724_),
    .X(_0747_));
 sky130_fd_sc_hd__a221o_1 _1393_ (.A1(net6),
    .A2(_0683_),
    .B1(_0731_),
    .B2(\MOS6502.PC[13] ),
    .C1(_0747_),
    .X(_0748_));
 sky130_fd_sc_hd__and3_1 _1394_ (.A(_0743_),
    .B(_0746_),
    .C(_0748_),
    .X(_0749_));
 sky130_fd_sc_hd__a21oi_1 _1395_ (.A1(_0743_),
    .A2(_0746_),
    .B1(_0748_),
    .Y(_0750_));
 sky130_fd_sc_hd__nor2_1 _1396_ (.A(_0749_),
    .B(_0750_),
    .Y(_0006_));
 sky130_fd_sc_hd__a221o_1 _1397_ (.A1(\MOS6502.ADD[6] ),
    .A2(_0729_),
    .B1(_0732_),
    .B2(\MOS6502.ABH[6] ),
    .C1(_0724_),
    .X(_0751_));
 sky130_fd_sc_hd__a221o_1 _1398_ (.A1(net7),
    .A2(_0683_),
    .B1(_0731_),
    .B2(\MOS6502.PC[14] ),
    .C1(_0751_),
    .X(_0752_));
 sky130_fd_sc_hd__nand2_1 _1399_ (.A(_0749_),
    .B(_0752_),
    .Y(_0753_));
 sky130_fd_sc_hd__or2_1 _1400_ (.A(_0749_),
    .B(_0752_),
    .X(_0754_));
 sky130_fd_sc_hd__and2_1 _1401_ (.A(_0753_),
    .B(_0754_),
    .X(_0755_));
 sky130_fd_sc_hd__clkbuf_1 _1402_ (.A(_0755_),
    .X(_0007_));
 sky130_fd_sc_hd__a221o_1 _1403_ (.A1(\MOS6502.ADD[7] ),
    .A2(_0729_),
    .B1(_0732_),
    .B2(\MOS6502.ABH[7] ),
    .C1(_0724_),
    .X(_0756_));
 sky130_fd_sc_hd__a221o_1 _1404_ (.A1(net8),
    .A2(_0683_),
    .B1(_0731_),
    .B2(\MOS6502.PC[15] ),
    .C1(_0756_),
    .X(_0757_));
 sky130_fd_sc_hd__xnor2_1 _1405_ (.A(_0753_),
    .B(_0757_),
    .Y(_0008_));
 sky130_fd_sc_hd__and3_1 _1406_ (.A(_0634_),
    .B(_0628_),
    .C(_0632_),
    .X(_0758_));
 sky130_fd_sc_hd__nor2_1 _1407_ (.A(_0635_),
    .B(_0758_),
    .Y(\MOS6502.ALU.temp[4] ));
 sky130_fd_sc_hd__nor2_1 _1408_ (.A(_0556_),
    .B(_0627_),
    .Y(_0759_));
 sky130_fd_sc_hd__and2b_1 _1409_ (.A_N(_0759_),
    .B(_0630_),
    .X(_0760_));
 sky130_fd_sc_hd__clkbuf_1 _1410_ (.A(_0760_),
    .X(\MOS6502.ALU.temp[3] ));
 sky130_fd_sc_hd__a21oi_1 _1411_ (.A1(_0426_),
    .A2(_0661_),
    .B1(_0662_),
    .Y(\MOS6502.ALU.temp_BI[7] ));
 sky130_fd_sc_hd__o32a_1 _1412_ (.A1(\MOS6502.write_back ),
    .A2(_0398_),
    .A3(_0416_),
    .B1(_0400_),
    .B2(_0410_),
    .X(_0761_));
 sky130_fd_sc_hd__inv_2 _1413_ (.A(_0409_),
    .Y(_0762_));
 sky130_fd_sc_hd__mux2_1 _1414_ (.A0(net5),
    .A1(\MOS6502.IRHOLD[4] ),
    .S(\MOS6502.IRHOLD_valid ),
    .X(_0763_));
 sky130_fd_sc_hd__and2_2 _1415_ (.A(_0356_),
    .B(_0763_),
    .X(_0764_));
 sky130_fd_sc_hd__mux2_1 _1416_ (.A0(net1),
    .A1(\MOS6502.IRHOLD[0] ),
    .S(\MOS6502.IRHOLD_valid ),
    .X(_0765_));
 sky130_fd_sc_hd__and2_1 _1417_ (.A(_0356_),
    .B(_0765_),
    .X(_0766_));
 sky130_fd_sc_hd__clkbuf_2 _1418_ (.A(_0766_),
    .X(_0767_));
 sky130_fd_sc_hd__mux2_1 _1419_ (.A0(net2),
    .A1(\MOS6502.IRHOLD[1] ),
    .S(\MOS6502.IRHOLD_valid ),
    .X(_0768_));
 sky130_fd_sc_hd__nand2_1 _1420_ (.A(_0357_),
    .B(_0768_),
    .Y(_0769_));
 sky130_fd_sc_hd__nand2_2 _1421_ (.A(_0767_),
    .B(_0769_),
    .Y(_0770_));
 sky130_fd_sc_hd__mux2_1 _1422_ (.A0(net4),
    .A1(\MOS6502.IRHOLD[3] ),
    .S(\MOS6502.IRHOLD_valid ),
    .X(_0771_));
 sky130_fd_sc_hd__nand2_1 _1423_ (.A(_0357_),
    .B(_0771_),
    .Y(_0772_));
 sky130_fd_sc_hd__mux2_1 _1424_ (.A0(net3),
    .A1(\MOS6502.IRHOLD[2] ),
    .S(\MOS6502.IRHOLD_valid ),
    .X(_0773_));
 sky130_fd_sc_hd__and2_1 _1425_ (.A(_0357_),
    .B(_0773_),
    .X(_0774_));
 sky130_fd_sc_hd__or2_2 _1426_ (.A(_0772_),
    .B(_0774_),
    .X(_0775_));
 sky130_fd_sc_hd__buf_2 _1427_ (.A(_0763_),
    .X(_0776_));
 sky130_fd_sc_hd__nand2_2 _1428_ (.A(_0357_),
    .B(_0773_),
    .Y(_0777_));
 sky130_fd_sc_hd__nand2_1 _1429_ (.A(_0772_),
    .B(_0777_),
    .Y(_0778_));
 sky130_fd_sc_hd__or4_1 _1430_ (.A(_0359_),
    .B(_0776_),
    .C(_0767_),
    .D(_0778_),
    .X(_0779_));
 sky130_fd_sc_hd__o31a_1 _1431_ (.A1(_0764_),
    .A2(_0770_),
    .A3(_0775_),
    .B1(_0779_),
    .X(_0780_));
 sky130_fd_sc_hd__or2_1 _1432_ (.A(_0414_),
    .B(_0680_),
    .X(_0781_));
 sky130_fd_sc_hd__or3_1 _1433_ (.A(_0378_),
    .B(_0392_),
    .C(_0407_),
    .X(_0782_));
 sky130_fd_sc_hd__o211a_1 _1434_ (.A1(_0410_),
    .A2(_0411_),
    .B1(_0781_),
    .C1(_0782_),
    .X(_0783_));
 sky130_fd_sc_hd__o221a_1 _1435_ (.A1(\MOS6502.write_back ),
    .A2(_0762_),
    .B1(_0689_),
    .B2(_0780_),
    .C1(_0783_),
    .X(_0784_));
 sky130_fd_sc_hd__o31ai_1 _1436_ (.A1(\MOS6502.ALU.CO ),
    .A2(\MOS6502.store ),
    .A3(_0761_),
    .B1(_0784_),
    .Y(_0785_));
 sky130_fd_sc_hd__o21a_1 _1437_ (.A1(\MOS6502.ALU.CO ),
    .A2(\MOS6502.store ),
    .B1(_0586_),
    .X(_0786_));
 sky130_fd_sc_hd__and2_1 _1438_ (.A(_0357_),
    .B(_0768_),
    .X(_0787_));
 sky130_fd_sc_hd__or2_1 _1439_ (.A(_0767_),
    .B(_0787_),
    .X(_0788_));
 sky130_fd_sc_hd__or2_2 _1440_ (.A(_0778_),
    .B(_0788_),
    .X(_0789_));
 sky130_fd_sc_hd__nand2_1 _1441_ (.A(_0357_),
    .B(_0776_),
    .Y(_0790_));
 sky130_fd_sc_hd__nand2_1 _1442_ (.A(_0361_),
    .B(_0790_),
    .Y(_0791_));
 sky130_fd_sc_hd__or2_2 _1443_ (.A(_0358_),
    .B(_0363_),
    .X(_0792_));
 sky130_fd_sc_hd__or3_1 _1444_ (.A(_0789_),
    .B(_0791_),
    .C(_0792_),
    .X(_0793_));
 sky130_fd_sc_hd__nor2_1 _1445_ (.A(_0689_),
    .B(_0793_),
    .Y(_0794_));
 sky130_fd_sc_hd__or3_1 _1446_ (.A(_0785_),
    .B(_0786_),
    .C(_0794_),
    .X(_0795_));
 sky130_fd_sc_hd__nor2_1 _1447_ (.A(\MOS6502.IR[7] ),
    .B(_0791_),
    .Y(_0796_));
 sky130_fd_sc_hd__buf_2 _1448_ (.A(_0788_),
    .X(_0797_));
 sky130_fd_sc_hd__nor2_2 _1449_ (.A(_0775_),
    .B(_0797_),
    .Y(_0798_));
 sky130_fd_sc_hd__and3_1 _1450_ (.A(_0678_),
    .B(_0796_),
    .C(_0798_),
    .X(_0799_));
 sky130_fd_sc_hd__and2_1 _1451_ (.A(\MOS6502.write_back ),
    .B(_0409_),
    .X(_0800_));
 sky130_fd_sc_hd__or4_1 _1452_ (.A(_0689_),
    .B(_0764_),
    .C(_0771_),
    .D(_0777_),
    .X(_0801_));
 sky130_fd_sc_hd__o21ai_1 _1453_ (.A1(_0398_),
    .A2(_0393_),
    .B1(_0801_),
    .Y(_0802_));
 sky130_fd_sc_hd__nor2_1 _1454_ (.A(_0680_),
    .B(_0422_),
    .Y(_0803_));
 sky130_fd_sc_hd__or2_1 _1455_ (.A(_0802_),
    .B(_0803_),
    .X(_0804_));
 sky130_fd_sc_hd__and2b_1 _1456_ (.A_N(_0696_),
    .B(_0465_),
    .X(_0805_));
 sky130_fd_sc_hd__or4_1 _1457_ (.A(_0483_),
    .B(_0435_),
    .C(_0589_),
    .D(_0805_),
    .X(_0806_));
 sky130_fd_sc_hd__or3_1 _1458_ (.A(_0800_),
    .B(_0804_),
    .C(_0806_),
    .X(_0807_));
 sky130_fd_sc_hd__inv_2 _1459_ (.A(_0477_),
    .Y(_0808_));
 sky130_fd_sc_hd__a2bb2o_1 _1460_ (.A1_N(_0388_),
    .A2_N(_0434_),
    .B1(_0808_),
    .B2(_0392_),
    .X(_0809_));
 sky130_fd_sc_hd__buf_2 _1461_ (.A(_0790_),
    .X(_0810_));
 sky130_fd_sc_hd__or3_1 _1462_ (.A(_0689_),
    .B(_0810_),
    .C(_0789_),
    .X(_0811_));
 sky130_fd_sc_hd__or4b_1 _1463_ (.A(_0445_),
    .B(_0807_),
    .C(_0809_),
    .D_N(_0811_),
    .X(_0812_));
 sky130_fd_sc_hd__or3_1 _1464_ (.A(_0795_),
    .B(_0799_),
    .C(_0812_),
    .X(_0813_));
 sky130_fd_sc_hd__clkbuf_1 _1465_ (.A(_0813_),
    .X(_0018_));
 sky130_fd_sc_hd__nor2_2 _1466_ (.A(_0371_),
    .B(_0398_),
    .Y(_0814_));
 sky130_fd_sc_hd__or2_1 _1467_ (.A(_0361_),
    .B(_0776_),
    .X(_0815_));
 sky130_fd_sc_hd__or4_1 _1468_ (.A(\MOS6502.IR[7] ),
    .B(_0775_),
    .C(_0797_),
    .D(_0815_),
    .X(_0816_));
 sky130_fd_sc_hd__nor2_1 _1469_ (.A(_0689_),
    .B(_0816_),
    .Y(_0817_));
 sky130_fd_sc_hd__or4_1 _1470_ (.A(_0689_),
    .B(_0764_),
    .C(_0770_),
    .D(_0778_),
    .X(_0818_));
 sky130_fd_sc_hd__or3b_1 _1471_ (.A(_0417_),
    .B(_0817_),
    .C_N(_0818_),
    .X(_0819_));
 sky130_fd_sc_hd__nor2_1 _1472_ (.A(_0410_),
    .B(_0375_),
    .Y(_0820_));
 sky130_fd_sc_hd__buf_2 _1473_ (.A(_0689_),
    .X(_0821_));
 sky130_fd_sc_hd__or2_1 _1474_ (.A(_0772_),
    .B(_0777_),
    .X(_0822_));
 sky130_fd_sc_hd__or4_1 _1475_ (.A(_0797_),
    .B(_0791_),
    .C(_0792_),
    .D(_0822_),
    .X(_0823_));
 sky130_fd_sc_hd__nor2_1 _1476_ (.A(_0821_),
    .B(_0823_),
    .Y(_0824_));
 sky130_fd_sc_hd__or4_1 _1477_ (.A(_0814_),
    .B(_0819_),
    .C(_0820_),
    .D(_0824_),
    .X(_0825_));
 sky130_fd_sc_hd__mux4_1 _1478_ (.A0(\MOS6502.N ),
    .A1(\MOS6502.V ),
    .A2(\MOS6502.C ),
    .A3(\MOS6502.Z ),
    .S0(\MOS6502.cond_code[1] ),
    .S1(\MOS6502.cond_code[2] ),
    .X(_0826_));
 sky130_fd_sc_hd__xnor2_1 _1479_ (.A(\MOS6502.cond_code[0] ),
    .B(_0826_),
    .Y(_0827_));
 sky130_fd_sc_hd__nor2_1 _1480_ (.A(_0392_),
    .B(_0428_),
    .Y(_0828_));
 sky130_fd_sc_hd__a21o_1 _1481_ (.A1(_0429_),
    .A2(_0827_),
    .B1(_0828_),
    .X(_0829_));
 sky130_fd_sc_hd__nand2_1 _1482_ (.A(_0359_),
    .B(_0363_),
    .Y(_0830_));
 sky130_fd_sc_hd__or2_1 _1483_ (.A(_0815_),
    .B(_0830_),
    .X(_0831_));
 sky130_fd_sc_hd__or2_1 _1484_ (.A(_0792_),
    .B(_0815_),
    .X(_0832_));
 sky130_fd_sc_hd__a211o_1 _1485_ (.A1(_0831_),
    .A2(_0832_),
    .B1(_0821_),
    .C1(_0789_),
    .X(_0833_));
 sky130_fd_sc_hd__nor3b_1 _1486_ (.A(_0825_),
    .B(_0829_),
    .C_N(_0833_),
    .Y(_0834_));
 sky130_fd_sc_hd__a21o_1 _1487_ (.A1(_0770_),
    .A2(_0777_),
    .B1(_0772_),
    .X(_0835_));
 sky130_fd_sc_hd__or4_1 _1488_ (.A(_0689_),
    .B(_0790_),
    .C(_0770_),
    .D(_0778_),
    .X(_0836_));
 sky130_fd_sc_hd__o211a_1 _1489_ (.A1(_0367_),
    .A2(_0443_),
    .B1(_0836_),
    .C1(_0376_),
    .X(_0837_));
 sky130_fd_sc_hd__o31a_1 _1490_ (.A1(_0821_),
    .A2(_0810_),
    .A3(_0835_),
    .B1(_0837_),
    .X(_0838_));
 sky130_fd_sc_hd__nand3b_1 _1491_ (.A_N(_0807_),
    .B(_0834_),
    .C(_0838_),
    .Y(_0019_));
 sky130_fd_sc_hd__o21a_1 _1492_ (.A1(_0359_),
    .A2(_0776_),
    .B1(_0831_),
    .X(_0839_));
 sky130_fd_sc_hd__or2_1 _1493_ (.A(_0767_),
    .B(_0769_),
    .X(_0840_));
 sky130_fd_sc_hd__a211o_1 _1494_ (.A1(_0770_),
    .A2(_0840_),
    .B1(_0822_),
    .C1(_0764_),
    .X(_0841_));
 sky130_fd_sc_hd__o31a_1 _1495_ (.A1(_0797_),
    .A2(_0822_),
    .A3(_0839_),
    .B1(_0841_),
    .X(_0842_));
 sky130_fd_sc_hd__nor2_1 _1496_ (.A(_0767_),
    .B(_0775_),
    .Y(_0843_));
 sky130_fd_sc_hd__o31a_1 _1497_ (.A1(\MOS6502.IR[7] ),
    .A2(_0776_),
    .A3(_0787_),
    .B1(_0843_),
    .X(_0844_));
 sky130_fd_sc_hd__nand2_1 _1498_ (.A(_0796_),
    .B(_0798_),
    .Y(_0845_));
 sky130_fd_sc_hd__and3b_1 _1499_ (.A_N(_0844_),
    .B(_0845_),
    .C(_0793_),
    .X(_0846_));
 sky130_fd_sc_hd__or3_1 _1500_ (.A(_0797_),
    .B(_0822_),
    .C(_0832_),
    .X(_0847_));
 sky130_fd_sc_hd__o2111a_1 _1501_ (.A1(_0789_),
    .A2(_0831_),
    .B1(_0847_),
    .C1(_0816_),
    .D1(_0823_),
    .X(_0848_));
 sky130_fd_sc_hd__o21a_1 _1502_ (.A1(_0791_),
    .A2(_0830_),
    .B1(_0832_),
    .X(_0849_));
 sky130_fd_sc_hd__and2_1 _1503_ (.A(_0767_),
    .B(_0769_),
    .X(_0850_));
 sky130_fd_sc_hd__clkbuf_2 _1504_ (.A(_0850_),
    .X(_0851_));
 sky130_fd_sc_hd__o21ai_1 _1505_ (.A1(_0851_),
    .A2(_0774_),
    .B1(_0772_),
    .Y(_0852_));
 sky130_fd_sc_hd__o2111a_1 _1506_ (.A1(_0810_),
    .A2(_0789_),
    .B1(_0852_),
    .C1(_0780_),
    .D1(_0678_),
    .X(_0853_));
 sky130_fd_sc_hd__o221a_1 _1507_ (.A1(_0810_),
    .A2(_0835_),
    .B1(_0849_),
    .B2(_0789_),
    .C1(_0853_),
    .X(_0854_));
 sky130_fd_sc_hd__and4_1 _1508_ (.A(_0842_),
    .B(_0846_),
    .C(_0848_),
    .D(_0854_),
    .X(_0855_));
 sky130_fd_sc_hd__a31o_1 _1509_ (.A1(_0375_),
    .A2(_0400_),
    .A3(_0694_),
    .B1(_0392_),
    .X(_0856_));
 sky130_fd_sc_hd__o311a_1 _1510_ (.A1(_0398_),
    .A2(_0428_),
    .A3(_0827_),
    .B1(_0697_),
    .C1(_0473_),
    .X(_0857_));
 sky130_fd_sc_hd__or4bb_1 _1511_ (.A(_0679_),
    .B(_0855_),
    .C_N(_0856_),
    .D_N(_0857_),
    .X(_0858_));
 sky130_fd_sc_hd__nor2_1 _1512_ (.A(_0410_),
    .B(_0416_),
    .Y(_0859_));
 sky130_fd_sc_hd__a211o_1 _1513_ (.A1(_0432_),
    .A2(_0433_),
    .B1(_0858_),
    .C1(_0859_),
    .X(_0860_));
 sky130_fd_sc_hd__or3_1 _1514_ (.A(\MOS6502.ALU.CO ),
    .B(\MOS6502.write_back ),
    .C(\MOS6502.store ),
    .X(_0861_));
 sky130_fd_sc_hd__a22o_1 _1515_ (.A1(_0585_),
    .A2(_0861_),
    .B1(_0844_),
    .B2(_0678_),
    .X(_0862_));
 sky130_fd_sc_hd__or4b_1 _1516_ (.A(_0444_),
    .B(_0805_),
    .C(_0804_),
    .D_N(_0811_),
    .X(_0863_));
 sky130_fd_sc_hd__or4_1 _1517_ (.A(_0795_),
    .B(_0829_),
    .C(_0862_),
    .D(_0863_),
    .X(_0864_));
 sky130_fd_sc_hd__or3_1 _1518_ (.A(_0825_),
    .B(_0860_),
    .C(_0864_),
    .X(_0865_));
 sky130_fd_sc_hd__clkbuf_1 _1519_ (.A(_0865_),
    .X(_0020_));
 sky130_fd_sc_hd__nor2_1 _1520_ (.A(_0821_),
    .B(_0842_),
    .Y(_0866_));
 sky130_fd_sc_hd__o21ai_1 _1521_ (.A1(_0821_),
    .A2(_0847_),
    .B1(_0439_),
    .Y(_0867_));
 sky130_fd_sc_hd__or4_1 _1522_ (.A(_0821_),
    .B(_0810_),
    .C(_0771_),
    .D(_0777_),
    .X(_0868_));
 sky130_fd_sc_hd__nand2_1 _1523_ (.A(_0430_),
    .B(_0868_),
    .Y(_0869_));
 sky130_fd_sc_hd__nand2_1 _1524_ (.A(_0487_),
    .B(_0838_),
    .Y(_0870_));
 sky130_fd_sc_hd__or4_1 _1525_ (.A(_0862_),
    .B(_0867_),
    .C(_0869_),
    .D(_0870_),
    .X(_0871_));
 sky130_fd_sc_hd__or4b_1 _1526_ (.A(_0018_),
    .B(_0866_),
    .C(_0871_),
    .D_N(_0834_),
    .X(_0872_));
 sky130_fd_sc_hd__nor2_1 _1527_ (.A(_0860_),
    .B(_0872_),
    .Y(_0873_));
 sky130_fd_sc_hd__o21ai_1 _1528_ (.A1(_0388_),
    .A2(_0434_),
    .B1(_0376_),
    .Y(_0874_));
 sky130_fd_sc_hd__or4_1 _1529_ (.A(_0444_),
    .B(_0436_),
    .C(_0802_),
    .D(_0874_),
    .X(_0875_));
 sky130_fd_sc_hd__or4_1 _1530_ (.A(_0785_),
    .B(_0819_),
    .C(_0867_),
    .D(_0875_),
    .X(_0876_));
 sky130_fd_sc_hd__or4b_1 _1531_ (.A(_0858_),
    .B(_0873_),
    .C(_0876_),
    .D_N(_0833_),
    .X(_0877_));
 sky130_fd_sc_hd__clkbuf_1 _1532_ (.A(_0877_),
    .X(_0021_));
 sky130_fd_sc_hd__o211a_1 _1533_ (.A1(_0367_),
    .A2(_0370_),
    .B1(_0388_),
    .C1(_0422_),
    .X(_0878_));
 sky130_fd_sc_hd__a2bb2o_1 _1534_ (.A1_N(_0410_),
    .A2_N(_0878_),
    .B1(_0808_),
    .B2(_0404_),
    .X(_0879_));
 sky130_fd_sc_hd__nor3_1 _1535_ (.A(_0387_),
    .B(_0445_),
    .C(_0814_),
    .Y(_0880_));
 sky130_fd_sc_hd__nand2_1 _1536_ (.A(_0836_),
    .B(_0880_),
    .Y(_0881_));
 sky130_fd_sc_hd__or4_1 _1537_ (.A(_0589_),
    .B(_0786_),
    .C(_0820_),
    .D(_0881_),
    .X(_0882_));
 sky130_fd_sc_hd__buf_2 _1538_ (.A(_0821_),
    .X(_0883_));
 sky130_fd_sc_hd__nor2_1 _1539_ (.A(_0883_),
    .B(_0848_),
    .Y(_0884_));
 sky130_fd_sc_hd__or4_1 _1540_ (.A(_0869_),
    .B(_0879_),
    .C(_0882_),
    .D(_0884_),
    .X(_0885_));
 sky130_fd_sc_hd__clkbuf_1 _1541_ (.A(_0885_),
    .X(_0022_));
 sky130_fd_sc_hd__or2_1 _1542_ (.A(_0789_),
    .B(_0832_),
    .X(_0886_));
 sky130_fd_sc_hd__a21oi_1 _1543_ (.A1(_0886_),
    .A2(_0846_),
    .B1(_0883_),
    .Y(_0887_));
 sky130_fd_sc_hd__o41a_1 _1544_ (.A1(_0369_),
    .A2(_0378_),
    .A3(_0368_),
    .A4(_0392_),
    .B1(_0487_),
    .X(_0888_));
 sky130_fd_sc_hd__nand2_1 _1545_ (.A(_0467_),
    .B(_0888_),
    .Y(_0889_));
 sky130_fd_sc_hd__nand2_1 _1546_ (.A(_0801_),
    .B(_0868_),
    .Y(_0890_));
 sky130_fd_sc_hd__a31o_1 _1547_ (.A1(_0380_),
    .A2(_0411_),
    .A3(_0416_),
    .B1(_0392_),
    .X(_0891_));
 sky130_fd_sc_hd__or4b_1 _1548_ (.A(_0478_),
    .B(_0800_),
    .C(_0890_),
    .D_N(_0891_),
    .X(_0892_));
 sky130_fd_sc_hd__or3_1 _1549_ (.A(_0887_),
    .B(_0889_),
    .C(_0892_),
    .X(_0893_));
 sky130_fd_sc_hd__clkbuf_1 _1550_ (.A(_0893_),
    .X(_0023_));
 sky130_fd_sc_hd__a211o_2 _1551_ (.A1(_0367_),
    .A2(_0412_),
    .B1(_0729_),
    .C1(_0401_),
    .X(_0894_));
 sky130_fd_sc_hd__or3_1 _1552_ (.A(_0395_),
    .B(_0419_),
    .C(_0894_),
    .X(_0895_));
 sky130_fd_sc_hd__clkbuf_4 _1553_ (.A(_0895_),
    .X(_0896_));
 sky130_fd_sc_hd__a211oi_2 _1554_ (.A1(_0404_),
    .A2(_0679_),
    .B1(_0681_),
    .C1(_0587_),
    .Y(_0897_));
 sky130_fd_sc_hd__o21ai_4 _1555_ (.A1(\MOS6502.state[5] ),
    .A2(_0402_),
    .B1(_0897_),
    .Y(_0898_));
 sky130_fd_sc_hd__or3_1 _1556_ (.A(_0466_),
    .B(_0677_),
    .C(_0889_),
    .X(_0899_));
 sky130_fd_sc_hd__nor2_1 _1557_ (.A(_0410_),
    .B(_0477_),
    .Y(_0900_));
 sky130_fd_sc_hd__or4b_1 _1558_ (.A(_0406_),
    .B(_0859_),
    .C(_0465_),
    .D_N(_0430_),
    .X(_0901_));
 sky130_fd_sc_hd__or4_4 _1559_ (.A(_0898_),
    .B(_0899_),
    .C(_0900_),
    .D(_0901_),
    .X(_0902_));
 sky130_fd_sc_hd__o21bai_1 _1560_ (.A1(_0410_),
    .A2(_0385_),
    .B1_N(_0408_),
    .Y(_0903_));
 sky130_fd_sc_hd__clkbuf_4 _1561_ (.A(_0903_),
    .X(_0904_));
 sky130_fd_sc_hd__a22o_1 _1562_ (.A1(\MOS6502.ADD[0] ),
    .A2(_0902_),
    .B1(_0904_),
    .B2(net1),
    .X(_0905_));
 sky130_fd_sc_hd__buf_2 _1563_ (.A(_0390_),
    .X(_0906_));
 sky130_fd_sc_hd__nor3_2 _1564_ (.A(_0386_),
    .B(_0906_),
    .C(_0471_),
    .Y(_0907_));
 sky130_fd_sc_hd__or3_2 _1565_ (.A(_0386_),
    .B(_0906_),
    .C(_0471_),
    .X(_0908_));
 sky130_fd_sc_hd__nor4_4 _1566_ (.A(_0908_),
    .B(_0902_),
    .C(_0896_),
    .D(_0904_),
    .Y(_0909_));
 sky130_fd_sc_hd__a2bb2o_1 _1567_ (.A1_N(_0563_),
    .A2_N(_0907_),
    .B1(_0909_),
    .B2(\MOS6502.PC[0] ),
    .X(_0910_));
 sky130_fd_sc_hd__a211o_4 _1568_ (.A1(\MOS6502.ABL[0] ),
    .A2(_0896_),
    .B1(_0905_),
    .C1(_0910_),
    .X(io_out[10]));
 sky130_fd_sc_hd__or4_1 _1569_ (.A(_0908_),
    .B(_0902_),
    .C(_0896_),
    .D(_0904_),
    .X(_0911_));
 sky130_fd_sc_hd__clkbuf_4 _1570_ (.A(_0911_),
    .X(_0912_));
 sky130_fd_sc_hd__buf_4 _1571_ (.A(_0909_),
    .X(_0913_));
 sky130_fd_sc_hd__a221o_1 _1572_ (.A1(\MOS6502.ABL[1] ),
    .A2(_0896_),
    .B1(_0904_),
    .B2(net2),
    .C1(_0913_),
    .X(_0914_));
 sky130_fd_sc_hd__a22o_1 _1573_ (.A1(_0573_),
    .A2(_0908_),
    .B1(_0902_),
    .B2(\MOS6502.ADD[1] ),
    .X(_0915_));
 sky130_fd_sc_hd__o22a_4 _1574_ (.A1(\MOS6502.PC[1] ),
    .A2(_0912_),
    .B1(_0914_),
    .B2(_0915_),
    .X(io_out[11]));
 sky130_fd_sc_hd__a221o_1 _1575_ (.A1(\MOS6502.ABL[2] ),
    .A2(_0896_),
    .B1(_0904_),
    .B2(net3),
    .C1(_0913_),
    .X(_0916_));
 sky130_fd_sc_hd__a2bb2o_1 _1576_ (.A1_N(_0608_),
    .A2_N(_0907_),
    .B1(_0902_),
    .B2(\MOS6502.ADD[2] ),
    .X(_0917_));
 sky130_fd_sc_hd__o22a_4 _1577_ (.A1(\MOS6502.PC[2] ),
    .A2(_0912_),
    .B1(_0916_),
    .B2(_0917_),
    .X(io_out[12]));
 sky130_fd_sc_hd__a221o_1 _1578_ (.A1(\MOS6502.ABL[3] ),
    .A2(_0896_),
    .B1(_0904_),
    .B2(net4),
    .C1(_0909_),
    .X(_0918_));
 sky130_fd_sc_hd__a2bb2o_1 _1579_ (.A1_N(_0540_),
    .A2_N(_0907_),
    .B1(_0902_),
    .B2(\MOS6502.ADD[3] ),
    .X(_0919_));
 sky130_fd_sc_hd__o22a_4 _1580_ (.A1(\MOS6502.PC[3] ),
    .A2(_0912_),
    .B1(_0918_),
    .B2(_0919_),
    .X(io_out[13]));
 sky130_fd_sc_hd__a221o_1 _1581_ (.A1(\MOS6502.ABL[4] ),
    .A2(_0896_),
    .B1(_0904_),
    .B2(net5),
    .C1(_0909_),
    .X(_0920_));
 sky130_fd_sc_hd__a2bb2o_1 _1582_ (.A1_N(_0525_),
    .A2_N(_0907_),
    .B1(_0902_),
    .B2(\MOS6502.ADD[4] ),
    .X(_0921_));
 sky130_fd_sc_hd__o22a_4 _1583_ (.A1(\MOS6502.PC[4] ),
    .A2(_0912_),
    .B1(_0920_),
    .B2(_0921_),
    .X(io_out[14]));
 sky130_fd_sc_hd__a221o_1 _1584_ (.A1(\MOS6502.ABL[5] ),
    .A2(_0896_),
    .B1(_0904_),
    .B2(net6),
    .C1(_0909_),
    .X(_0922_));
 sky130_fd_sc_hd__a2bb2o_1 _1585_ (.A1_N(_0503_),
    .A2_N(_0907_),
    .B1(_0902_),
    .B2(\MOS6502.ADD[5] ),
    .X(_0923_));
 sky130_fd_sc_hd__o22a_4 _1586_ (.A1(\MOS6502.PC[5] ),
    .A2(_0912_),
    .B1(_0922_),
    .B2(_0923_),
    .X(io_out[15]));
 sky130_fd_sc_hd__a221o_1 _1587_ (.A1(\MOS6502.ABL[6] ),
    .A2(_0896_),
    .B1(_0904_),
    .B2(net7),
    .C1(_0909_),
    .X(_0924_));
 sky130_fd_sc_hd__a2bb2o_1 _1588_ (.A1_N(_0516_),
    .A2_N(_0907_),
    .B1(_0902_),
    .B2(\MOS6502.ADD[6] ),
    .X(_0925_));
 sky130_fd_sc_hd__o22a_4 _1589_ (.A1(\MOS6502.PC[6] ),
    .A2(_0912_),
    .B1(_0924_),
    .B2(_0925_),
    .X(io_out[16]));
 sky130_fd_sc_hd__a221o_1 _1590_ (.A1(\MOS6502.ABL[7] ),
    .A2(_0896_),
    .B1(_0904_),
    .B2(net8),
    .C1(_0909_),
    .X(_0926_));
 sky130_fd_sc_hd__a2bb2o_1 _1591_ (.A1_N(_0640_),
    .A2_N(_0907_),
    .B1(_0902_),
    .B2(\MOS6502.ADD[7] ),
    .X(_0927_));
 sky130_fd_sc_hd__o22a_4 _1592_ (.A1(\MOS6502.PC[7] ),
    .A2(_0912_),
    .B1(_0926_),
    .B2(_0927_),
    .X(io_out[17]));
 sky130_fd_sc_hd__a211o_1 _1593_ (.A1(\MOS6502.ADD[0] ),
    .A2(_0894_),
    .B1(_0899_),
    .C1(_0908_),
    .X(_0928_));
 sky130_fd_sc_hd__or3_1 _1594_ (.A(_0395_),
    .B(_0419_),
    .C(_0465_),
    .X(_0929_));
 sky130_fd_sc_hd__clkbuf_4 _1595_ (.A(_0929_),
    .X(_0930_));
 sky130_fd_sc_hd__a22o_1 _1596_ (.A1(net1),
    .A2(_0898_),
    .B1(_0930_),
    .B2(\MOS6502.ABH[0] ),
    .X(_0931_));
 sky130_fd_sc_hd__a211o_4 _1597_ (.A1(\MOS6502.PC[8] ),
    .A2(_0913_),
    .B1(_0928_),
    .C1(_0931_),
    .X(io_out[18]));
 sky130_fd_sc_hd__a22o_1 _1598_ (.A1(net2),
    .A2(_0898_),
    .B1(_0930_),
    .B2(\MOS6502.ABH[1] ),
    .X(_0932_));
 sky130_fd_sc_hd__a211o_1 _1599_ (.A1(\MOS6502.ADD[1] ),
    .A2(_0894_),
    .B1(_0913_),
    .C1(_0932_),
    .X(_0933_));
 sky130_fd_sc_hd__o21a_2 _1600_ (.A1(\MOS6502.PC[9] ),
    .A2(_0912_),
    .B1(_0933_),
    .X(io_out[19]));
 sky130_fd_sc_hd__a22o_1 _1601_ (.A1(net3),
    .A2(_0898_),
    .B1(_0894_),
    .B2(\MOS6502.ADD[2] ),
    .X(_0934_));
 sky130_fd_sc_hd__a221o_4 _1602_ (.A1(\MOS6502.PC[10] ),
    .A2(_0913_),
    .B1(_0930_),
    .B2(\MOS6502.ABH[2] ),
    .C1(_0934_),
    .X(io_out[20]));
 sky130_fd_sc_hd__a22o_1 _1603_ (.A1(net4),
    .A2(_0898_),
    .B1(_0894_),
    .B2(\MOS6502.ADD[3] ),
    .X(_0935_));
 sky130_fd_sc_hd__a221o_4 _1604_ (.A1(\MOS6502.PC[11] ),
    .A2(_0913_),
    .B1(_0930_),
    .B2(\MOS6502.ABH[3] ),
    .C1(_0935_),
    .X(io_out[21]));
 sky130_fd_sc_hd__a22o_1 _1605_ (.A1(net5),
    .A2(_0898_),
    .B1(_0894_),
    .B2(\MOS6502.ADD[4] ),
    .X(_0936_));
 sky130_fd_sc_hd__a221o_4 _1606_ (.A1(\MOS6502.PC[12] ),
    .A2(_0913_),
    .B1(_0930_),
    .B2(\MOS6502.ABH[4] ),
    .C1(_0936_),
    .X(io_out[22]));
 sky130_fd_sc_hd__a22o_1 _1607_ (.A1(net6),
    .A2(_0898_),
    .B1(_0894_),
    .B2(\MOS6502.ADD[5] ),
    .X(_0937_));
 sky130_fd_sc_hd__a221o_4 _1608_ (.A1(\MOS6502.PC[13] ),
    .A2(_0913_),
    .B1(_0930_),
    .B2(\MOS6502.ABH[5] ),
    .C1(_0937_),
    .X(io_out[23]));
 sky130_fd_sc_hd__a22o_1 _1609_ (.A1(net7),
    .A2(_0898_),
    .B1(_0894_),
    .B2(\MOS6502.ADD[6] ),
    .X(_0938_));
 sky130_fd_sc_hd__a221o_4 _1610_ (.A1(\MOS6502.PC[14] ),
    .A2(_0913_),
    .B1(_0930_),
    .B2(\MOS6502.ABH[6] ),
    .C1(_0938_),
    .X(io_out[24]));
 sky130_fd_sc_hd__a22o_1 _1611_ (.A1(net8),
    .A2(_0898_),
    .B1(_0894_),
    .B2(\MOS6502.ADD[7] ),
    .X(_0939_));
 sky130_fd_sc_hd__a221o_4 _1612_ (.A1(\MOS6502.PC[15] ),
    .A2(_0913_),
    .B1(_0930_),
    .B2(\MOS6502.ABH[7] ),
    .C1(_0939_),
    .X(io_out[25]));
 sky130_fd_sc_hd__nor2_2 _1613_ (.A(_0391_),
    .B(_0395_),
    .Y(_0940_));
 sky130_fd_sc_hd__a21o_2 _1614_ (.A1(\MOS6502.php ),
    .A2(_0386_),
    .B1(_0724_),
    .X(_0941_));
 sky130_fd_sc_hd__a22o_1 _1615_ (.A1(\MOS6502.PC[8] ),
    .A2(_0906_),
    .B1(_0941_),
    .B2(\MOS6502.C ),
    .X(_0942_));
 sky130_fd_sc_hd__o21bai_4 _1616_ (.A1(\MOS6502.php ),
    .A2(_0488_),
    .B1_N(_0395_),
    .Y(_0943_));
 sky130_fd_sc_hd__a22o_1 _1617_ (.A1(\MOS6502.PC[0] ),
    .A2(_0466_),
    .B1(_0943_),
    .B2(\MOS6502.ADD[0] ),
    .X(_0944_));
 sky130_fd_sc_hd__nand2_1 _1618_ (.A(_0940_),
    .B(_0563_),
    .Y(_0945_));
 sky130_fd_sc_hd__o31a_4 _1619_ (.A1(_0940_),
    .A2(_0942_),
    .A3(_0944_),
    .B1(_0945_),
    .X(io_out[0]));
 sky130_fd_sc_hd__a22o_1 _1620_ (.A1(\MOS6502.PC[1] ),
    .A2(_0466_),
    .B1(_0941_),
    .B2(\MOS6502.Z ),
    .X(_0946_));
 sky130_fd_sc_hd__a221o_1 _1621_ (.A1(\MOS6502.PC[9] ),
    .A2(_0906_),
    .B1(_0943_),
    .B2(\MOS6502.ADD[1] ),
    .C1(_0940_),
    .X(_0947_));
 sky130_fd_sc_hd__o22a_2 _1622_ (.A1(_0397_),
    .A2(_0573_),
    .B1(_0946_),
    .B2(_0947_),
    .X(io_out[1]));
 sky130_fd_sc_hd__a22o_1 _1623_ (.A1(\MOS6502.PC[2] ),
    .A2(_0466_),
    .B1(_0941_),
    .B2(\MOS6502.I ),
    .X(_0948_));
 sky130_fd_sc_hd__a22o_1 _1624_ (.A1(\MOS6502.PC[10] ),
    .A2(_0906_),
    .B1(_0943_),
    .B2(\MOS6502.ADD[2] ),
    .X(_0949_));
 sky130_fd_sc_hd__nand2_1 _1625_ (.A(_0940_),
    .B(_0608_),
    .Y(_0950_));
 sky130_fd_sc_hd__o31a_4 _1626_ (.A1(_0940_),
    .A2(_0948_),
    .A3(_0949_),
    .B1(_0950_),
    .X(io_out[2]));
 sky130_fd_sc_hd__a22o_1 _1627_ (.A1(\MOS6502.PC[3] ),
    .A2(_0466_),
    .B1(_0906_),
    .B2(\MOS6502.PC[11] ),
    .X(_0951_));
 sky130_fd_sc_hd__a221o_1 _1628_ (.A1(\MOS6502.D ),
    .A2(_0941_),
    .B1(_0943_),
    .B2(\MOS6502.ADD[3] ),
    .C1(_0951_),
    .X(_0952_));
 sky130_fd_sc_hd__o21bai_4 _1629_ (.A1(_0397_),
    .A2(_0540_),
    .B1_N(_0952_),
    .Y(io_out[3]));
 sky130_fd_sc_hd__o21a_1 _1630_ (.A1(_0386_),
    .A2(_0395_),
    .B1(\MOS6502.ADD[4] ),
    .X(_0953_));
 sky130_fd_sc_hd__a221o_1 _1631_ (.A1(\MOS6502.PC[4] ),
    .A2(_0466_),
    .B1(_0906_),
    .B2(\MOS6502.PC[12] ),
    .C1(_0953_),
    .X(_0954_));
 sky130_fd_sc_hd__a21oi_1 _1632_ (.A1(\MOS6502.php ),
    .A2(_0386_),
    .B1(_0954_),
    .Y(_0955_));
 sky130_fd_sc_hd__o31a_1 _1633_ (.A1(\MOS6502.NMI_edge ),
    .A2(net9),
    .A3(_0701_),
    .B1(_0955_),
    .X(_0956_));
 sky130_fd_sc_hd__o21ai_4 _1634_ (.A1(_0397_),
    .A2(_0525_),
    .B1(_0956_),
    .Y(io_out[4]));
 sky130_fd_sc_hd__nor2_1 _1635_ (.A(_0397_),
    .B(_0503_),
    .Y(_0957_));
 sky130_fd_sc_hd__o21a_1 _1636_ (.A1(_0386_),
    .A2(_0395_),
    .B1(\MOS6502.ADD[5] ),
    .X(_0958_));
 sky130_fd_sc_hd__a221o_1 _1637_ (.A1(\MOS6502.PC[5] ),
    .A2(_0466_),
    .B1(_0906_),
    .B2(\MOS6502.PC[13] ),
    .C1(_0941_),
    .X(_0959_));
 sky130_fd_sc_hd__or3_1 _1638_ (.A(_0957_),
    .B(_0958_),
    .C(_0959_),
    .X(_0960_));
 sky130_fd_sc_hd__buf_2 _1639_ (.A(_0960_),
    .X(io_out[5]));
 sky130_fd_sc_hd__a22o_1 _1640_ (.A1(\MOS6502.PC[6] ),
    .A2(_0466_),
    .B1(_0941_),
    .B2(\MOS6502.V ),
    .X(_0961_));
 sky130_fd_sc_hd__a221o_1 _1641_ (.A1(\MOS6502.PC[14] ),
    .A2(_0906_),
    .B1(_0943_),
    .B2(\MOS6502.ADD[6] ),
    .C1(_0940_),
    .X(_0962_));
 sky130_fd_sc_hd__o2bb2a_2 _1642_ (.A1_N(_0940_),
    .A2_N(_0516_),
    .B1(_0961_),
    .B2(_0962_),
    .X(io_out[6]));
 sky130_fd_sc_hd__a22o_1 _1643_ (.A1(\MOS6502.PC[7] ),
    .A2(_0466_),
    .B1(_0906_),
    .B2(\MOS6502.PC[15] ),
    .X(_0963_));
 sky130_fd_sc_hd__a2bb2o_1 _1644_ (.A1_N(_0397_),
    .A2_N(_0640_),
    .B1(_0943_),
    .B2(\MOS6502.ADD[7] ),
    .X(_0964_));
 sky130_fd_sc_hd__a211o_4 _1645_ (.A1(\MOS6502.N ),
    .A2(_0941_),
    .B1(_0963_),
    .C1(_0964_),
    .X(io_out[7]));
 sky130_fd_sc_hd__inv_2 _1646_ (.A(net11),
    .Y(_0024_));
 sky130_fd_sc_hd__inv_2 _1647_ (.A(net11),
    .Y(_0025_));
 sky130_fd_sc_hd__inv_2 _1648_ (.A(net11),
    .Y(_0026_));
 sky130_fd_sc_hd__inv_2 _1649_ (.A(net11),
    .Y(_0027_));
 sky130_fd_sc_hd__inv_2 _1650_ (.A(net11),
    .Y(_0028_));
 sky130_fd_sc_hd__inv_2 _1651_ (.A(net11),
    .Y(_0029_));
 sky130_fd_sc_hd__buf_2 _1652_ (.A(_0387_),
    .X(_0965_));
 sky130_fd_sc_hd__mux2_1 _1653_ (.A0(\MOS6502.ADD[0] ),
    .A1(net1),
    .S(_0965_),
    .X(_0966_));
 sky130_fd_sc_hd__or3b_1 _1654_ (.A(_0821_),
    .B(\MOS6502.plp ),
    .C_N(\MOS6502.load_reg ),
    .X(_0967_));
 sky130_fd_sc_hd__nand3_1 _1655_ (.A(_0880_),
    .B(_0888_),
    .C(_0967_),
    .Y(_0968_));
 sky130_fd_sc_hd__and3_1 _1656_ (.A(_0499_),
    .B(_0496_),
    .C(_0968_),
    .X(_0969_));
 sky130_fd_sc_hd__clkbuf_4 _1657_ (.A(_0969_),
    .X(_0970_));
 sky130_fd_sc_hd__mux2_1 _1658_ (.A0(\MOS6502.AXYS[2][0] ),
    .A1(_0966_),
    .S(_0970_),
    .X(_0971_));
 sky130_fd_sc_hd__clkbuf_1 _1659_ (.A(_0971_),
    .X(_0030_));
 sky130_fd_sc_hd__and3_1 _1660_ (.A(\MOS6502.adc_bcd ),
    .B(\MOS6502.adj_bcd ),
    .C(\MOS6502.ALU.HC ),
    .X(_0125_));
 sky130_fd_sc_hd__or2b_1 _1661_ (.A(\MOS6502.adc_bcd ),
    .B_N(\MOS6502.adj_bcd ),
    .X(_0126_));
 sky130_fd_sc_hd__nor2_1 _1662_ (.A(\MOS6502.ALU.HC ),
    .B(_0126_),
    .Y(_0127_));
 sky130_fd_sc_hd__or3_1 _1663_ (.A(\MOS6502.ADD[1] ),
    .B(_0125_),
    .C(_0127_),
    .X(_0128_));
 sky130_fd_sc_hd__o21a_1 _1664_ (.A1(_0125_),
    .A2(_0127_),
    .B1(\MOS6502.ADD[1] ),
    .X(_0129_));
 sky130_fd_sc_hd__nor2_1 _1665_ (.A(_0965_),
    .B(_0129_),
    .Y(_0130_));
 sky130_fd_sc_hd__a22o_1 _1666_ (.A1(net2),
    .A2(_0965_),
    .B1(_0128_),
    .B2(_0130_),
    .X(_0131_));
 sky130_fd_sc_hd__mux2_1 _1667_ (.A0(\MOS6502.AXYS[2][1] ),
    .A1(_0131_),
    .S(_0970_),
    .X(_0132_));
 sky130_fd_sc_hd__clkbuf_1 _1668_ (.A(_0132_),
    .X(_0031_));
 sky130_fd_sc_hd__or2_1 _1669_ (.A(\MOS6502.ADD[2] ),
    .B(_0125_),
    .X(_0133_));
 sky130_fd_sc_hd__nand2_1 _1670_ (.A(\MOS6502.ADD[2] ),
    .B(_0125_),
    .Y(_0134_));
 sky130_fd_sc_hd__a21oi_1 _1671_ (.A1(_0133_),
    .A2(_0134_),
    .B1(_0129_),
    .Y(_0135_));
 sky130_fd_sc_hd__a31o_1 _1672_ (.A1(_0129_),
    .A2(_0133_),
    .A3(_0134_),
    .B1(_0965_),
    .X(_0136_));
 sky130_fd_sc_hd__a2bb2o_1 _1673_ (.A1_N(_0135_),
    .A2_N(_0136_),
    .B1(net3),
    .B2(_0965_),
    .X(_0137_));
 sky130_fd_sc_hd__mux2_1 _1674_ (.A0(\MOS6502.AXYS[2][2] ),
    .A1(_0137_),
    .S(_0970_),
    .X(_0138_));
 sky130_fd_sc_hd__clkbuf_1 _1675_ (.A(_0138_),
    .X(_0032_));
 sky130_fd_sc_hd__a21bo_1 _1676_ (.A1(_0129_),
    .A2(_0133_),
    .B1_N(_0134_),
    .X(_0139_));
 sky130_fd_sc_hd__xnor2_1 _1677_ (.A(\MOS6502.ADD[3] ),
    .B(_0127_),
    .Y(_0140_));
 sky130_fd_sc_hd__xnor2_1 _1678_ (.A(_0139_),
    .B(_0140_),
    .Y(_0141_));
 sky130_fd_sc_hd__mux2_1 _1679_ (.A0(_0141_),
    .A1(net4),
    .S(_0965_),
    .X(_0142_));
 sky130_fd_sc_hd__mux2_1 _1680_ (.A0(\MOS6502.AXYS[2][3] ),
    .A1(_0142_),
    .S(_0970_),
    .X(_0143_));
 sky130_fd_sc_hd__clkbuf_1 _1681_ (.A(_0143_),
    .X(_0033_));
 sky130_fd_sc_hd__mux2_1 _1682_ (.A0(\MOS6502.ADD[4] ),
    .A1(net5),
    .S(_0965_),
    .X(_0144_));
 sky130_fd_sc_hd__mux2_1 _1683_ (.A0(\MOS6502.AXYS[2][4] ),
    .A1(_0144_),
    .S(_0970_),
    .X(_0145_));
 sky130_fd_sc_hd__clkbuf_1 _1684_ (.A(_0145_),
    .X(_0034_));
 sky130_fd_sc_hd__and3_1 _1685_ (.A(\MOS6502.ALU.CO ),
    .B(\MOS6502.adc_bcd ),
    .C(\MOS6502.adj_bcd ),
    .X(_0146_));
 sky130_fd_sc_hd__nor2_1 _1686_ (.A(\MOS6502.ALU.CO ),
    .B(_0126_),
    .Y(_0147_));
 sky130_fd_sc_hd__o21a_1 _1687_ (.A1(_0146_),
    .A2(_0147_),
    .B1(\MOS6502.ADD[5] ),
    .X(_0148_));
 sky130_fd_sc_hd__or3_1 _1688_ (.A(\MOS6502.ADD[5] ),
    .B(_0146_),
    .C(_0147_),
    .X(_0149_));
 sky130_fd_sc_hd__or3b_1 _1689_ (.A(_0387_),
    .B(_0148_),
    .C_N(_0149_),
    .X(_0150_));
 sky130_fd_sc_hd__a21bo_1 _1690_ (.A1(net6),
    .A2(_0965_),
    .B1_N(_0150_),
    .X(_0151_));
 sky130_fd_sc_hd__mux2_1 _1691_ (.A0(\MOS6502.AXYS[2][5] ),
    .A1(_0151_),
    .S(_0970_),
    .X(_0152_));
 sky130_fd_sc_hd__clkbuf_1 _1692_ (.A(_0152_),
    .X(_0035_));
 sky130_fd_sc_hd__or2_1 _1693_ (.A(\MOS6502.ADD[6] ),
    .B(_0146_),
    .X(_0153_));
 sky130_fd_sc_hd__nand2_1 _1694_ (.A(\MOS6502.ADD[6] ),
    .B(_0146_),
    .Y(_0154_));
 sky130_fd_sc_hd__a21oi_1 _1695_ (.A1(_0153_),
    .A2(_0154_),
    .B1(_0148_),
    .Y(_0155_));
 sky130_fd_sc_hd__a31o_1 _1696_ (.A1(_0148_),
    .A2(_0153_),
    .A3(_0154_),
    .B1(_0387_),
    .X(_0156_));
 sky130_fd_sc_hd__a2bb2o_1 _1697_ (.A1_N(_0155_),
    .A2_N(_0156_),
    .B1(net7),
    .B2(_0965_),
    .X(_0157_));
 sky130_fd_sc_hd__mux2_1 _1698_ (.A0(\MOS6502.AXYS[2][6] ),
    .A1(_0157_),
    .S(_0970_),
    .X(_0158_));
 sky130_fd_sc_hd__clkbuf_1 _1699_ (.A(_0158_),
    .X(_0036_));
 sky130_fd_sc_hd__a21bo_1 _1700_ (.A1(_0148_),
    .A2(_0153_),
    .B1_N(_0154_),
    .X(_0159_));
 sky130_fd_sc_hd__xnor2_1 _1701_ (.A(\MOS6502.ADD[7] ),
    .B(_0147_),
    .Y(_0160_));
 sky130_fd_sc_hd__nor2_1 _1702_ (.A(_0159_),
    .B(_0160_),
    .Y(_0161_));
 sky130_fd_sc_hd__a21o_1 _1703_ (.A1(_0159_),
    .A2(_0160_),
    .B1(_0965_),
    .X(_0162_));
 sky130_fd_sc_hd__o32a_2 _1704_ (.A1(net8),
    .A2(_0410_),
    .A3(_0380_),
    .B1(_0161_),
    .B2(_0162_),
    .X(_0163_));
 sky130_fd_sc_hd__mux2_1 _1705_ (.A0(\MOS6502.AXYS[2][7] ),
    .A1(_0163_),
    .S(_0970_),
    .X(_0164_));
 sky130_fd_sc_hd__clkbuf_1 _1706_ (.A(_0164_),
    .X(_0037_));
 sky130_fd_sc_hd__and2_1 _1707_ (.A(_0500_),
    .B(_0968_),
    .X(_0165_));
 sky130_fd_sc_hd__clkbuf_4 _1708_ (.A(_0165_),
    .X(_0166_));
 sky130_fd_sc_hd__mux2_1 _1709_ (.A0(\MOS6502.AXYS[1][0] ),
    .A1(_0966_),
    .S(_0166_),
    .X(_0167_));
 sky130_fd_sc_hd__clkbuf_1 _1710_ (.A(_0167_),
    .X(_0038_));
 sky130_fd_sc_hd__mux2_1 _1711_ (.A0(\MOS6502.AXYS[1][1] ),
    .A1(_0131_),
    .S(_0166_),
    .X(_0168_));
 sky130_fd_sc_hd__clkbuf_1 _1712_ (.A(_0168_),
    .X(_0039_));
 sky130_fd_sc_hd__mux2_1 _1713_ (.A0(\MOS6502.AXYS[1][2] ),
    .A1(_0137_),
    .S(_0166_),
    .X(_0169_));
 sky130_fd_sc_hd__clkbuf_1 _1714_ (.A(_0169_),
    .X(_0040_));
 sky130_fd_sc_hd__mux2_1 _1715_ (.A0(\MOS6502.AXYS[1][3] ),
    .A1(_0142_),
    .S(_0166_),
    .X(_0170_));
 sky130_fd_sc_hd__clkbuf_1 _1716_ (.A(_0170_),
    .X(_0041_));
 sky130_fd_sc_hd__mux2_1 _1717_ (.A0(\MOS6502.AXYS[1][4] ),
    .A1(_0144_),
    .S(_0166_),
    .X(_0171_));
 sky130_fd_sc_hd__clkbuf_1 _1718_ (.A(_0171_),
    .X(_0042_));
 sky130_fd_sc_hd__mux2_1 _1719_ (.A0(\MOS6502.AXYS[1][5] ),
    .A1(_0151_),
    .S(_0166_),
    .X(_0172_));
 sky130_fd_sc_hd__clkbuf_1 _1720_ (.A(_0172_),
    .X(_0043_));
 sky130_fd_sc_hd__mux2_1 _1721_ (.A0(\MOS6502.AXYS[1][6] ),
    .A1(_0157_),
    .S(_0166_),
    .X(_0173_));
 sky130_fd_sc_hd__clkbuf_1 _1722_ (.A(_0173_),
    .X(_0044_));
 sky130_fd_sc_hd__mux2_1 _1723_ (.A0(\MOS6502.AXYS[1][7] ),
    .A1(_0163_),
    .S(_0166_),
    .X(_0174_));
 sky130_fd_sc_hd__clkbuf_1 _1724_ (.A(_0174_),
    .X(_0045_));
 sky130_fd_sc_hd__a21oi_1 _1725_ (.A1(_0428_),
    .A2(_0477_),
    .B1(\MOS6502.state[5] ),
    .Y(_0175_));
 sky130_fd_sc_hd__nand2_1 _1726_ (.A(_0402_),
    .B(_0781_),
    .Y(_0176_));
 sky130_fd_sc_hd__or4_1 _1727_ (.A(_0389_),
    .B(_0828_),
    .C(_0479_),
    .D(_0803_),
    .X(_0177_));
 sky130_fd_sc_hd__or4_1 _1728_ (.A(_0677_),
    .B(_0401_),
    .C(_0421_),
    .D(_0177_),
    .X(_0178_));
 sky130_fd_sc_hd__or2_1 _1729_ (.A(_0394_),
    .B(_0678_),
    .X(_0179_));
 sky130_fd_sc_hd__or3_1 _1730_ (.A(_0874_),
    .B(_0903_),
    .C(_0179_),
    .X(_0180_));
 sky130_fd_sc_hd__nor2_1 _1731_ (.A(_0404_),
    .B(_0385_),
    .Y(_0181_));
 sky130_fd_sc_hd__or3_1 _1732_ (.A(_0181_),
    .B(_0486_),
    .C(_0587_),
    .X(_0182_));
 sky130_fd_sc_hd__or4_1 _1733_ (.A(_0440_),
    .B(_0178_),
    .C(_0180_),
    .D(_0182_),
    .X(_0183_));
 sky130_fd_sc_hd__or4b_1 _1734_ (.A(_0175_),
    .B(_0176_),
    .C(_0183_),
    .D_N(_0693_),
    .X(_0184_));
 sky130_fd_sc_hd__and3_1 _1735_ (.A(_0488_),
    .B(_0474_),
    .C(_0184_),
    .X(_0185_));
 sky130_fd_sc_hd__buf_2 _1736_ (.A(_0185_),
    .X(_0186_));
 sky130_fd_sc_hd__clkbuf_4 _1737_ (.A(_0186_),
    .X(_0187_));
 sky130_fd_sc_hd__mux2_1 _1738_ (.A0(\MOS6502.ABL[0] ),
    .A1(io_out[10]),
    .S(_0187_),
    .X(_0188_));
 sky130_fd_sc_hd__clkbuf_1 _1739_ (.A(_0188_),
    .X(_0046_));
 sky130_fd_sc_hd__mux2_1 _1740_ (.A0(\MOS6502.ABL[1] ),
    .A1(io_out[11]),
    .S(_0187_),
    .X(_0189_));
 sky130_fd_sc_hd__clkbuf_1 _1741_ (.A(_0189_),
    .X(_0047_));
 sky130_fd_sc_hd__mux2_1 _1742_ (.A0(\MOS6502.ABL[2] ),
    .A1(io_out[12]),
    .S(_0187_),
    .X(_0190_));
 sky130_fd_sc_hd__clkbuf_1 _1743_ (.A(_0190_),
    .X(_0048_));
 sky130_fd_sc_hd__mux2_1 _1744_ (.A0(\MOS6502.ABL[3] ),
    .A1(io_out[13]),
    .S(_0187_),
    .X(_0191_));
 sky130_fd_sc_hd__clkbuf_1 _1745_ (.A(_0191_),
    .X(_0049_));
 sky130_fd_sc_hd__mux2_1 _1746_ (.A0(\MOS6502.ABL[4] ),
    .A1(io_out[14]),
    .S(_0187_),
    .X(_0192_));
 sky130_fd_sc_hd__clkbuf_1 _1747_ (.A(_0192_),
    .X(_0050_));
 sky130_fd_sc_hd__mux2_1 _1748_ (.A0(\MOS6502.ABL[5] ),
    .A1(io_out[15]),
    .S(_0187_),
    .X(_0193_));
 sky130_fd_sc_hd__clkbuf_1 _1749_ (.A(_0193_),
    .X(_0051_));
 sky130_fd_sc_hd__mux2_1 _1750_ (.A0(\MOS6502.ABL[6] ),
    .A1(io_out[16]),
    .S(_0187_),
    .X(_0194_));
 sky130_fd_sc_hd__clkbuf_1 _1751_ (.A(_0194_),
    .X(_0052_));
 sky130_fd_sc_hd__mux2_1 _1752_ (.A0(\MOS6502.ABL[7] ),
    .A1(io_out[17]),
    .S(_0187_),
    .X(_0195_));
 sky130_fd_sc_hd__clkbuf_1 _1753_ (.A(_0195_),
    .X(_0053_));
 sky130_fd_sc_hd__clkinv_2 _1754_ (.A(\MOS6502.clc ),
    .Y(_0196_));
 sky130_fd_sc_hd__mux2_1 _1755_ (.A0(_0196_),
    .A1(\MOS6502.ADD[0] ),
    .S(\MOS6502.plp ),
    .X(_0197_));
 sky130_fd_sc_hd__or3_1 _1756_ (.A(\MOS6502.adc_sbc ),
    .B(\MOS6502.compare ),
    .C(\MOS6502.shift ),
    .X(_0198_));
 sky130_fd_sc_hd__mux2_1 _1757_ (.A0(_0197_),
    .A1(\MOS6502.ALU.CO ),
    .S(_0198_),
    .X(_0199_));
 sky130_fd_sc_hd__mux2_1 _1758_ (.A0(net1),
    .A1(_0199_),
    .S(_0439_),
    .X(_0200_));
 sky130_fd_sc_hd__buf_2 _1759_ (.A(\MOS6502.plp ),
    .X(_0201_));
 sky130_fd_sc_hd__or4_1 _1760_ (.A(_0201_),
    .B(_0369_),
    .C(\MOS6502.clc ),
    .D(\MOS6502.sec ),
    .X(_0202_));
 sky130_fd_sc_hd__a2bb2o_1 _1761_ (.A1_N(\MOS6502.write_back ),
    .A2_N(_0883_),
    .B1(_0395_),
    .B2(\MOS6502.shift ),
    .X(_0203_));
 sky130_fd_sc_hd__nor2_2 _1762_ (.A(_0392_),
    .B(_0438_),
    .Y(_0204_));
 sky130_fd_sc_hd__o22a_1 _1763_ (.A1(_0198_),
    .A2(_0202_),
    .B1(_0203_),
    .B2(_0204_),
    .X(_0205_));
 sky130_fd_sc_hd__mux2_1 _1764_ (.A0(\MOS6502.C ),
    .A1(_0200_),
    .S(_0205_),
    .X(_0206_));
 sky130_fd_sc_hd__clkbuf_1 _1765_ (.A(_0206_),
    .X(_0054_));
 sky130_fd_sc_hd__or4_1 _1766_ (.A(\MOS6502.ADD[4] ),
    .B(\MOS6502.ADD[5] ),
    .C(\MOS6502.ADD[6] ),
    .D(\MOS6502.ADD[7] ),
    .X(_0207_));
 sky130_fd_sc_hd__or4_1 _1767_ (.A(\MOS6502.ADD[0] ),
    .B(\MOS6502.ADD[1] ),
    .C(\MOS6502.ADD[2] ),
    .D(\MOS6502.ADD[3] ),
    .X(_0208_));
 sky130_fd_sc_hd__nor2_1 _1768_ (.A(_0207_),
    .B(_0208_),
    .Y(_0209_));
 sky130_fd_sc_hd__mux2_1 _1769_ (.A0(\MOS6502.ADD[1] ),
    .A1(net2),
    .S(_0204_),
    .X(_0210_));
 sky130_fd_sc_hd__o21ba_1 _1770_ (.A1(_0201_),
    .A2(_0204_),
    .B1_N(_0395_),
    .X(_0211_));
 sky130_fd_sc_hd__mux2_1 _1771_ (.A0(_0209_),
    .A1(_0210_),
    .S(_0211_),
    .X(_0212_));
 sky130_fd_sc_hd__o21a_1 _1772_ (.A1(_0499_),
    .A2(_0496_),
    .B1(\MOS6502.load_reg ),
    .X(_0213_));
 sky130_fd_sc_hd__or4_1 _1773_ (.A(_0201_),
    .B(\MOS6502.compare ),
    .C(_0821_),
    .D(_0213_),
    .X(_0214_));
 sky130_fd_sc_hd__o22a_1 _1774_ (.A1(_0204_),
    .A2(_0179_),
    .B1(_0214_),
    .B2(\MOS6502.bit_ins ),
    .X(_0215_));
 sky130_fd_sc_hd__mux2_1 _1775_ (.A0(\MOS6502.Z ),
    .A1(_0212_),
    .S(_0215_),
    .X(_0216_));
 sky130_fd_sc_hd__clkbuf_1 _1776_ (.A(_0216_),
    .X(_0055_));
 sky130_fd_sc_hd__mux2_1 _1777_ (.A0(net8),
    .A1(\MOS6502.ADD[7] ),
    .S(_0179_),
    .X(_0217_));
 sky130_fd_sc_hd__a211o_1 _1778_ (.A1(\MOS6502.bit_ins ),
    .A2(_0415_),
    .B1(_0678_),
    .C1(_0204_),
    .X(_0218_));
 sky130_fd_sc_hd__o21a_1 _1779_ (.A1(_0395_),
    .A2(_0218_),
    .B1(_0214_),
    .X(_0219_));
 sky130_fd_sc_hd__mux2_1 _1780_ (.A0(\MOS6502.N ),
    .A1(_0217_),
    .S(_0219_),
    .X(_0220_));
 sky130_fd_sc_hd__clkbuf_1 _1781_ (.A(_0220_),
    .X(_0056_));
 sky130_fd_sc_hd__clkinv_2 _1782_ (.A(\MOS6502.cld ),
    .Y(_0221_));
 sky130_fd_sc_hd__mux2_1 _1783_ (.A0(_0221_),
    .A1(\MOS6502.ADD[3] ),
    .S(_0201_),
    .X(_0222_));
 sky130_fd_sc_hd__mux2_1 _1784_ (.A0(net4),
    .A1(_0222_),
    .S(_0439_),
    .X(_0223_));
 sky130_fd_sc_hd__clkbuf_4 _1785_ (.A(_0678_),
    .X(_0224_));
 sky130_fd_sc_hd__or4_1 _1786_ (.A(_0201_),
    .B(\MOS6502.cld ),
    .C(\MOS6502.sed ),
    .D(_0821_),
    .X(_0225_));
 sky130_fd_sc_hd__o21a_1 _1787_ (.A1(_0224_),
    .A2(_0204_),
    .B1(_0225_),
    .X(_0226_));
 sky130_fd_sc_hd__mux2_1 _1788_ (.A0(\MOS6502.D ),
    .A1(_0223_),
    .S(_0226_),
    .X(_0227_));
 sky130_fd_sc_hd__clkbuf_1 _1789_ (.A(_0227_),
    .X(_0057_));
 sky130_fd_sc_hd__inv_2 _1790_ (.A(\MOS6502.cli ),
    .Y(_0228_));
 sky130_fd_sc_hd__mux2_1 _1791_ (.A0(\MOS6502.ADD[2] ),
    .A1(_0228_),
    .S(_0418_),
    .X(_0229_));
 sky130_fd_sc_hd__mux2_1 _1792_ (.A0(net3),
    .A1(_0229_),
    .S(_0439_),
    .X(_0230_));
 sky130_fd_sc_hd__o32a_1 _1793_ (.A1(\MOS6502.cli ),
    .A2(\MOS6502.sei ),
    .A3(_0400_),
    .B1(_0368_),
    .B2(_0201_),
    .X(_0231_));
 sky130_fd_sc_hd__o31a_1 _1794_ (.A1(_0418_),
    .A2(_0678_),
    .A3(_0204_),
    .B1(_0231_),
    .X(_0232_));
 sky130_fd_sc_hd__mux2_1 _1795_ (.A0(\MOS6502.I ),
    .A1(_0230_),
    .S(_0232_),
    .X(_0233_));
 sky130_fd_sc_hd__or2_1 _1796_ (.A(_0814_),
    .B(_0233_),
    .X(_0234_));
 sky130_fd_sc_hd__clkbuf_1 _1797_ (.A(_0234_),
    .X(_0058_));
 sky130_fd_sc_hd__nor2_1 _1798_ (.A(_0201_),
    .B(\MOS6502.clv ),
    .Y(_0235_));
 sky130_fd_sc_hd__xor2_1 _1799_ (.A(\MOS6502.ALU.BI7 ),
    .B(\MOS6502.ALU.AI7 ),
    .X(_0236_));
 sky130_fd_sc_hd__xnor2_1 _1800_ (.A(\MOS6502.ADD[7] ),
    .B(\MOS6502.ALU.CO ),
    .Y(_0237_));
 sky130_fd_sc_hd__xnor2_1 _1801_ (.A(_0236_),
    .B(_0237_),
    .Y(_0238_));
 sky130_fd_sc_hd__a221o_1 _1802_ (.A1(_0201_),
    .A2(\MOS6502.ADD[6] ),
    .B1(_0235_),
    .B2(_0238_),
    .C1(_0883_),
    .X(_0239_));
 sky130_fd_sc_hd__o21a_1 _1803_ (.A1(net7),
    .A2(_0224_),
    .B1(_0239_),
    .X(_0240_));
 sky130_fd_sc_hd__o41a_1 _1804_ (.A1(_0201_),
    .A2(\MOS6502.adc_sbc ),
    .A3(\MOS6502.clv ),
    .A4(_0883_),
    .B1(_0218_),
    .X(_0241_));
 sky130_fd_sc_hd__mux2_1 _1805_ (.A0(\MOS6502.V ),
    .A1(_0240_),
    .S(_0241_),
    .X(_0242_));
 sky130_fd_sc_hd__clkbuf_1 _1806_ (.A(_0242_),
    .X(_0059_));
 sky130_fd_sc_hd__or2_1 _1807_ (.A(net11),
    .B(_0474_),
    .X(_0243_));
 sky130_fd_sc_hd__buf_2 _1808_ (.A(_0243_),
    .X(_0244_));
 sky130_fd_sc_hd__mux2_1 _1809_ (.A0(net1),
    .A1(\MOS6502.IRHOLD[0] ),
    .S(_0244_),
    .X(_0245_));
 sky130_fd_sc_hd__clkbuf_1 _1810_ (.A(_0245_),
    .X(_0060_));
 sky130_fd_sc_hd__mux2_1 _1811_ (.A0(net2),
    .A1(\MOS6502.IRHOLD[1] ),
    .S(_0244_),
    .X(_0246_));
 sky130_fd_sc_hd__clkbuf_1 _1812_ (.A(_0246_),
    .X(_0061_));
 sky130_fd_sc_hd__mux2_1 _1813_ (.A0(net3),
    .A1(\MOS6502.IRHOLD[2] ),
    .S(_0244_),
    .X(_0247_));
 sky130_fd_sc_hd__clkbuf_1 _1814_ (.A(_0247_),
    .X(_0062_));
 sky130_fd_sc_hd__mux2_1 _1815_ (.A0(net4),
    .A1(\MOS6502.IRHOLD[3] ),
    .S(_0244_),
    .X(_0248_));
 sky130_fd_sc_hd__clkbuf_1 _1816_ (.A(_0248_),
    .X(_0063_));
 sky130_fd_sc_hd__mux2_1 _1817_ (.A0(net5),
    .A1(\MOS6502.IRHOLD[4] ),
    .S(_0244_),
    .X(_0249_));
 sky130_fd_sc_hd__clkbuf_1 _1818_ (.A(_0249_),
    .X(_0064_));
 sky130_fd_sc_hd__mux2_1 _1819_ (.A0(net6),
    .A1(\MOS6502.IRHOLD[5] ),
    .S(_0244_),
    .X(_0250_));
 sky130_fd_sc_hd__clkbuf_1 _1820_ (.A(_0250_),
    .X(_0065_));
 sky130_fd_sc_hd__mux2_1 _1821_ (.A0(net7),
    .A1(\MOS6502.IRHOLD[6] ),
    .S(_0244_),
    .X(_0251_));
 sky130_fd_sc_hd__clkbuf_1 _1822_ (.A(_0251_),
    .X(_0066_));
 sky130_fd_sc_hd__mux2_1 _1823_ (.A0(net8),
    .A1(\MOS6502.IRHOLD[7] ),
    .S(_0244_),
    .X(_0252_));
 sky130_fd_sc_hd__clkbuf_1 _1824_ (.A(_0252_),
    .X(_0067_));
 sky130_fd_sc_hd__buf_2 _1825_ (.A(_0883_),
    .X(_0253_));
 sky130_fd_sc_hd__nand2_1 _1826_ (.A(\MOS6502.IRHOLD_valid ),
    .B(_0253_),
    .Y(_0254_));
 sky130_fd_sc_hd__a21oi_1 _1827_ (.A1(_0474_),
    .A2(_0254_),
    .B1(net11),
    .Y(_0068_));
 sky130_fd_sc_hd__and3_1 _1828_ (.A(_0357_),
    .B(_0358_),
    .C(_0362_),
    .X(_0255_));
 sky130_fd_sc_hd__or2_1 _1829_ (.A(_0775_),
    .B(_0840_),
    .X(_0256_));
 sky130_fd_sc_hd__nor2_1 _1830_ (.A(_0791_),
    .B(_0256_),
    .Y(_0257_));
 sky130_fd_sc_hd__nand2_2 _1831_ (.A(\MOS6502.IR[7] ),
    .B(_0363_),
    .Y(_0258_));
 sky130_fd_sc_hd__nor2_1 _1832_ (.A(_0360_),
    .B(_0258_),
    .Y(_0259_));
 sky130_fd_sc_hd__a22o_1 _1833_ (.A1(_0255_),
    .A2(_0257_),
    .B1(_0259_),
    .B2(_0843_),
    .X(_0260_));
 sky130_fd_sc_hd__nand2_1 _1834_ (.A(_0359_),
    .B(_0810_),
    .Y(_0261_));
 sky130_fd_sc_hd__and3_1 _1835_ (.A(\MOS6502.IR[7] ),
    .B(_0363_),
    .C(_0776_),
    .X(_0262_));
 sky130_fd_sc_hd__nand2_1 _1836_ (.A(\MOS6502.IR[5] ),
    .B(_0262_),
    .Y(_0263_));
 sky130_fd_sc_hd__a21oi_1 _1837_ (.A1(_0261_),
    .A2(_0263_),
    .B1(_0256_),
    .Y(_0264_));
 sky130_fd_sc_hd__and2_1 _1838_ (.A(_0810_),
    .B(_0798_),
    .X(_0265_));
 sky130_fd_sc_hd__nor2_1 _1839_ (.A(_0359_),
    .B(\MOS6502.IR[5] ),
    .Y(_0266_));
 sky130_fd_sc_hd__or2_1 _1840_ (.A(_0767_),
    .B(_0777_),
    .X(_0267_));
 sky130_fd_sc_hd__buf_2 _1841_ (.A(_0361_),
    .X(_0268_));
 sky130_fd_sc_hd__or4_1 _1842_ (.A(_0268_),
    .B(_0764_),
    .C(_0767_),
    .D(_0258_),
    .X(_0269_));
 sky130_fd_sc_hd__o221a_1 _1843_ (.A1(_0770_),
    .A2(_0266_),
    .B1(_0263_),
    .B2(_0267_),
    .C1(_0269_),
    .X(_0270_));
 sky130_fd_sc_hd__or4b_1 _1844_ (.A(_0260_),
    .B(_0264_),
    .C(_0265_),
    .D_N(_0270_),
    .X(_0271_));
 sky130_fd_sc_hd__clkbuf_4 _1845_ (.A(_0224_),
    .X(_0272_));
 sky130_fd_sc_hd__mux2_1 _1846_ (.A0(\MOS6502.load_reg ),
    .A1(_0271_),
    .S(_0272_),
    .X(_0273_));
 sky130_fd_sc_hd__clkbuf_1 _1847_ (.A(_0273_),
    .X(_0069_));
 sky130_fd_sc_hd__clkbuf_4 _1848_ (.A(_0883_),
    .X(_0274_));
 sky130_fd_sc_hd__a21o_1 _1849_ (.A1(\MOS6502.res ),
    .A2(_0274_),
    .B1(net11),
    .X(_0070_));
 sky130_fd_sc_hd__nor2_1 _1850_ (.A(_0256_),
    .B(_0258_),
    .Y(_0275_));
 sky130_fd_sc_hd__a2111o_1 _1851_ (.A1(_0776_),
    .A2(_0777_),
    .B1(_0797_),
    .C1(_0258_),
    .D1(_0268_),
    .X(_0276_));
 sky130_fd_sc_hd__a21bo_1 _1852_ (.A1(_0266_),
    .A2(_0265_),
    .B1_N(_0276_),
    .X(_0277_));
 sky130_fd_sc_hd__a31o_1 _1853_ (.A1(_0268_),
    .A2(_0764_),
    .A3(_0275_),
    .B1(_0277_),
    .X(_0278_));
 sky130_fd_sc_hd__a21o_1 _1854_ (.A1(\MOS6502.dst_reg[0] ),
    .A2(_0253_),
    .B1(_0799_),
    .X(_0279_));
 sky130_fd_sc_hd__a21o_1 _1855_ (.A1(_0272_),
    .A2(_0278_),
    .B1(_0279_),
    .X(_0071_));
 sky130_fd_sc_hd__nor2_1 _1856_ (.A(_0767_),
    .B(_0769_),
    .Y(_0280_));
 sky130_fd_sc_hd__nor2_1 _1857_ (.A(_0268_),
    .B(_0258_),
    .Y(_0281_));
 sky130_fd_sc_hd__o21a_1 _1858_ (.A1(_0257_),
    .A2(_0265_),
    .B1(_0255_),
    .X(_0282_));
 sky130_fd_sc_hd__a211o_1 _1859_ (.A1(_0280_),
    .A2(_0281_),
    .B1(_0277_),
    .C1(_0282_),
    .X(_0283_));
 sky130_fd_sc_hd__mux2_1 _1860_ (.A0(\MOS6502.dst_reg[1] ),
    .A1(_0283_),
    .S(_0272_),
    .X(_0284_));
 sky130_fd_sc_hd__clkbuf_1 _1861_ (.A(_0284_),
    .X(_0072_));
 sky130_fd_sc_hd__or2_1 _1862_ (.A(\MOS6502.IR[6] ),
    .B(_0778_),
    .X(_0285_));
 sky130_fd_sc_hd__a21oi_1 _1863_ (.A1(\MOS6502.IR[6] ),
    .A2(_0776_),
    .B1(_0797_),
    .Y(_0286_));
 sky130_fd_sc_hd__a31o_1 _1864_ (.A1(_0266_),
    .A2(_0285_),
    .A3(_0286_),
    .B1(_0883_),
    .X(_0287_));
 sky130_fd_sc_hd__a31o_1 _1865_ (.A1(\MOS6502.IR[5] ),
    .A2(_0776_),
    .A3(_0275_),
    .B1(_0287_),
    .X(_0288_));
 sky130_fd_sc_hd__o21a_1 _1866_ (.A1(\MOS6502.src_reg[0] ),
    .A2(_0272_),
    .B1(_0288_),
    .X(_0073_));
 sky130_fd_sc_hd__inv_2 _1867_ (.A(_0267_),
    .Y(_0289_));
 sky130_fd_sc_hd__nor2_1 _1868_ (.A(_0797_),
    .B(_0815_),
    .Y(_0290_));
 sky130_fd_sc_hd__a22o_1 _1869_ (.A1(_0289_),
    .A2(_0259_),
    .B1(_0290_),
    .B2(_0255_),
    .X(_0291_));
 sky130_fd_sc_hd__o32a_1 _1870_ (.A1(_0260_),
    .A2(_0287_),
    .A3(_0291_),
    .B1(_0272_),
    .B2(\MOS6502.src_reg[1] ),
    .X(_0074_));
 sky130_fd_sc_hd__nand2_1 _1871_ (.A(_0810_),
    .B(_0772_),
    .Y(_0292_));
 sky130_fd_sc_hd__nor2_1 _1872_ (.A(_0777_),
    .B(_0840_),
    .Y(_0293_));
 sky130_fd_sc_hd__a32o_1 _1873_ (.A1(_0851_),
    .A2(_0777_),
    .A3(_0292_),
    .B1(_0293_),
    .B2(_0262_),
    .X(_0294_));
 sky130_fd_sc_hd__mux2_1 _1874_ (.A0(\MOS6502.index_y ),
    .A1(_0294_),
    .S(_0224_),
    .X(_0295_));
 sky130_fd_sc_hd__clkbuf_1 _1875_ (.A(_0295_),
    .X(_0075_));
 sky130_fd_sc_hd__o21a_1 _1876_ (.A1(_0851_),
    .A2(_0289_),
    .B1(_0259_),
    .X(_0296_));
 sky130_fd_sc_hd__mux2_1 _1877_ (.A0(\MOS6502.store ),
    .A1(_0296_),
    .S(_0224_),
    .X(_0297_));
 sky130_fd_sc_hd__clkbuf_1 _1878_ (.A(_0297_),
    .X(_0076_));
 sky130_fd_sc_hd__and2_1 _1879_ (.A(\MOS6502.write_back ),
    .B(_0883_),
    .X(_0298_));
 sky130_fd_sc_hd__a31o_1 _1880_ (.A1(_0272_),
    .A2(_0258_),
    .A3(_0293_),
    .B1(_0298_),
    .X(_0077_));
 sky130_fd_sc_hd__mux2_1 _1881_ (.A0(\MOS6502.load_only ),
    .A1(_0281_),
    .S(_0224_),
    .X(_0299_));
 sky130_fd_sc_hd__clkbuf_1 _1882_ (.A(_0299_),
    .X(_0078_));
 sky130_fd_sc_hd__and2_1 _1883_ (.A(_0272_),
    .B(_0255_),
    .X(_0300_));
 sky130_fd_sc_hd__a21o_1 _1884_ (.A1(\MOS6502.IR[5] ),
    .A2(_0293_),
    .B1(_0265_),
    .X(_0301_));
 sky130_fd_sc_hd__a22o_1 _1885_ (.A1(\MOS6502.inc ),
    .A2(_0274_),
    .B1(_0300_),
    .B2(_0301_),
    .X(_0079_));
 sky130_fd_sc_hd__or3b_2 _1886_ (.A(_0368_),
    .B(_0398_),
    .C_N(_0458_),
    .X(_0302_));
 sky130_fd_sc_hd__nor3_1 _1887_ (.A(_0268_),
    .B(_0363_),
    .C(_0302_),
    .Y(_0303_));
 sky130_fd_sc_hd__a22o_1 _1888_ (.A1(\MOS6502.adc_sbc ),
    .A2(_0302_),
    .B1(_0851_),
    .B2(_0303_),
    .X(_0080_));
 sky130_fd_sc_hd__and4_1 _1889_ (.A(_0359_),
    .B(_0224_),
    .C(_0778_),
    .D(_0280_),
    .X(_0304_));
 sky130_fd_sc_hd__a21o_1 _1890_ (.A1(\MOS6502.shift ),
    .A2(_0274_),
    .B1(_0304_),
    .X(_0081_));
 sky130_fd_sc_hd__and3_1 _1891_ (.A(_0359_),
    .B(_0851_),
    .C(_0303_),
    .X(_0305_));
 sky130_fd_sc_hd__a22o_1 _1892_ (.A1(\MOS6502.adc_bcd ),
    .A2(_0302_),
    .B1(_0305_),
    .B2(\MOS6502.D ),
    .X(_0082_));
 sky130_fd_sc_hd__and3b_1 _1893_ (.A_N(_0797_),
    .B(_0775_),
    .C(_0810_),
    .X(_0306_));
 sky130_fd_sc_hd__a21o_1 _1894_ (.A1(_0268_),
    .A2(_0851_),
    .B1(_0306_),
    .X(_0307_));
 sky130_fd_sc_hd__a22o_1 _1895_ (.A1(\MOS6502.compare ),
    .A2(_0274_),
    .B1(_0300_),
    .B2(_0307_),
    .X(_0083_));
 sky130_fd_sc_hd__nor2_1 _1896_ (.A(_0792_),
    .B(_0840_),
    .Y(_0308_));
 sky130_fd_sc_hd__mux2_1 _1897_ (.A0(\MOS6502.shift_right ),
    .A1(_0308_),
    .S(_0224_),
    .X(_0309_));
 sky130_fd_sc_hd__clkbuf_1 _1898_ (.A(_0309_),
    .X(_0084_));
 sky130_fd_sc_hd__a22o_1 _1899_ (.A1(\MOS6502.rotate ),
    .A2(_0274_),
    .B1(_0304_),
    .B2(\MOS6502.IR[5] ),
    .X(_0085_));
 sky130_fd_sc_hd__or4_1 _1900_ (.A(\MOS6502.IR[7] ),
    .B(\MOS6502.IR[5] ),
    .C(_0883_),
    .D(_0770_),
    .X(_0310_));
 sky130_fd_sc_hd__o21a_1 _1901_ (.A1(\MOS6502.op[0] ),
    .A2(_0272_),
    .B1(_0310_),
    .X(_0086_));
 sky130_fd_sc_hd__o211a_1 _1902_ (.A1(_0268_),
    .A2(_0363_),
    .B1(_0851_),
    .C1(_0359_),
    .X(_0311_));
 sky130_fd_sc_hd__a21o_1 _1903_ (.A1(_0268_),
    .A2(_0293_),
    .B1(_0306_),
    .X(_0312_));
 sky130_fd_sc_hd__o31a_1 _1904_ (.A1(_0851_),
    .A2(_0257_),
    .A3(_0312_),
    .B1(_0255_),
    .X(_0313_));
 sky130_fd_sc_hd__nor4_1 _1905_ (.A(_0268_),
    .B(_0777_),
    .C(_0797_),
    .D(_0831_),
    .Y(_0314_));
 sky130_fd_sc_hd__a31o_1 _1906_ (.A1(_0810_),
    .A2(_0798_),
    .A3(_0259_),
    .B1(_0308_),
    .X(_0315_));
 sky130_fd_sc_hd__or4_1 _1907_ (.A(_0311_),
    .B(_0313_),
    .C(_0314_),
    .D(_0315_),
    .X(_0316_));
 sky130_fd_sc_hd__nor2_1 _1908_ (.A(_0253_),
    .B(_0830_),
    .Y(_0317_));
 sky130_fd_sc_hd__o2bb2a_1 _1909_ (.A1_N(_0316_),
    .A2_N(_0317_),
    .B1(\MOS6502.op[1] ),
    .B2(_0272_),
    .X(_0087_));
 sky130_fd_sc_hd__mux2_1 _1910_ (.A0(\MOS6502.op[2] ),
    .A1(_0316_),
    .S(_0224_),
    .X(_0318_));
 sky130_fd_sc_hd__clkbuf_1 _1911_ (.A(_0318_),
    .X(_0088_));
 sky130_fd_sc_hd__a31o_1 _1912_ (.A1(_0359_),
    .A2(_0363_),
    .A3(_0280_),
    .B1(_0316_),
    .X(_0319_));
 sky130_fd_sc_hd__nor2_1 _1913_ (.A(_0358_),
    .B(_0253_),
    .Y(_0320_));
 sky130_fd_sc_hd__a22o_1 _1914_ (.A1(\MOS6502.op[3] ),
    .A2(_0274_),
    .B1(_0319_),
    .B2(_0320_),
    .X(_0089_));
 sky130_fd_sc_hd__mux2_1 _1915_ (.A0(\MOS6502.bit_ins ),
    .A1(_0314_),
    .S(_0224_),
    .X(_0321_));
 sky130_fd_sc_hd__clkbuf_1 _1916_ (.A(_0321_),
    .X(_0090_));
 sky130_fd_sc_hd__nand2_1 _1917_ (.A(_0272_),
    .B(_0798_),
    .Y(_0322_));
 sky130_fd_sc_hd__a2bb2o_1 _1918_ (.A1_N(_0322_),
    .A2_N(_0263_),
    .B1(\MOS6502.clv ),
    .B2(_0274_),
    .X(_0091_));
 sky130_fd_sc_hd__and3_1 _1919_ (.A(\MOS6502.IR[5] ),
    .B(_0776_),
    .C(_0798_),
    .X(_0323_));
 sky130_fd_sc_hd__nor2_1 _1920_ (.A(_0253_),
    .B(_0792_),
    .Y(_0324_));
 sky130_fd_sc_hd__a22o_1 _1921_ (.A1(\MOS6502.sei ),
    .A2(_0274_),
    .B1(_0323_),
    .B2(_0324_),
    .X(_0092_));
 sky130_fd_sc_hd__and3_1 _1922_ (.A(_0268_),
    .B(_0764_),
    .C(_0798_),
    .X(_0325_));
 sky130_fd_sc_hd__a22o_1 _1923_ (.A1(\MOS6502.cli ),
    .A2(_0274_),
    .B1(_0324_),
    .B2(_0325_),
    .X(_0093_));
 sky130_fd_sc_hd__a22o_1 _1924_ (.A1(\MOS6502.sed ),
    .A2(_0274_),
    .B1(_0300_),
    .B2(_0323_),
    .X(_0094_));
 sky130_fd_sc_hd__a22o_1 _1925_ (.A1(\MOS6502.cld ),
    .A2(_0253_),
    .B1(_0300_),
    .B2(_0325_),
    .X(_0095_));
 sky130_fd_sc_hd__a22o_1 _1926_ (.A1(\MOS6502.sec ),
    .A2(_0253_),
    .B1(_0317_),
    .B2(_0323_),
    .X(_0096_));
 sky130_fd_sc_hd__a22o_1 _1927_ (.A1(\MOS6502.clc ),
    .A2(_0253_),
    .B1(_0317_),
    .B2(_0325_),
    .X(_0097_));
 sky130_fd_sc_hd__a22o_1 _1928_ (.A1(\MOS6502.php ),
    .A2(_0253_),
    .B1(_0799_),
    .B2(_0363_),
    .X(_0098_));
 sky130_fd_sc_hd__a22o_1 _1929_ (.A1(_0201_),
    .A2(_0253_),
    .B1(_0817_),
    .B2(_0363_),
    .X(_0099_));
 sky130_fd_sc_hd__or3b_1 _1930_ (.A(\MOS6502.NMI_edge ),
    .B(\MOS6502.NMI_1 ),
    .C_N(net10),
    .X(_0326_));
 sky130_fd_sc_hd__o21ai_1 _1931_ (.A1(_0706_),
    .A2(_0814_),
    .B1(_0326_),
    .Y(_0100_));
 sky130_fd_sc_hd__mux2_1 _1932_ (.A0(\MOS6502.ABH[0] ),
    .A1(io_out[18]),
    .S(_0187_),
    .X(_0327_));
 sky130_fd_sc_hd__clkbuf_1 _1933_ (.A(_0327_),
    .X(_0101_));
 sky130_fd_sc_hd__mux2_1 _1934_ (.A0(\MOS6502.ABH[1] ),
    .A1(io_out[19]),
    .S(_0187_),
    .X(_0328_));
 sky130_fd_sc_hd__clkbuf_1 _1935_ (.A(_0328_),
    .X(_0102_));
 sky130_fd_sc_hd__mux2_1 _1936_ (.A0(\MOS6502.ABH[2] ),
    .A1(io_out[20]),
    .S(_0186_),
    .X(_0329_));
 sky130_fd_sc_hd__clkbuf_1 _1937_ (.A(_0329_),
    .X(_0103_));
 sky130_fd_sc_hd__mux2_1 _1938_ (.A0(\MOS6502.ABH[3] ),
    .A1(io_out[21]),
    .S(_0186_),
    .X(_0330_));
 sky130_fd_sc_hd__clkbuf_1 _1939_ (.A(_0330_),
    .X(_0104_));
 sky130_fd_sc_hd__mux2_1 _1940_ (.A0(\MOS6502.ABH[4] ),
    .A1(io_out[22]),
    .S(_0186_),
    .X(_0331_));
 sky130_fd_sc_hd__clkbuf_1 _1941_ (.A(_0331_),
    .X(_0105_));
 sky130_fd_sc_hd__mux2_1 _1942_ (.A0(\MOS6502.ABH[5] ),
    .A1(io_out[23]),
    .S(_0186_),
    .X(_0332_));
 sky130_fd_sc_hd__clkbuf_1 _1943_ (.A(_0332_),
    .X(_0106_));
 sky130_fd_sc_hd__mux2_1 _1944_ (.A0(\MOS6502.ABH[6] ),
    .A1(io_out[24]),
    .S(_0186_),
    .X(_0333_));
 sky130_fd_sc_hd__clkbuf_1 _1945_ (.A(_0333_),
    .X(_0107_));
 sky130_fd_sc_hd__mux2_1 _1946_ (.A0(\MOS6502.ABH[7] ),
    .A1(io_out[25]),
    .S(_0186_),
    .X(_0334_));
 sky130_fd_sc_hd__clkbuf_1 _1947_ (.A(_0334_),
    .X(_0108_));
 sky130_fd_sc_hd__and3_1 _1948_ (.A(_0493_),
    .B(_0496_),
    .C(_0968_),
    .X(_0335_));
 sky130_fd_sc_hd__clkbuf_4 _1949_ (.A(_0335_),
    .X(_0336_));
 sky130_fd_sc_hd__mux2_1 _1950_ (.A0(\MOS6502.AXYS[3][0] ),
    .A1(_0966_),
    .S(_0336_),
    .X(_0337_));
 sky130_fd_sc_hd__clkbuf_1 _1951_ (.A(_0337_),
    .X(_0109_));
 sky130_fd_sc_hd__mux2_1 _1952_ (.A0(\MOS6502.AXYS[3][1] ),
    .A1(_0131_),
    .S(_0336_),
    .X(_0338_));
 sky130_fd_sc_hd__clkbuf_1 _1953_ (.A(_0338_),
    .X(_0110_));
 sky130_fd_sc_hd__mux2_1 _1954_ (.A0(\MOS6502.AXYS[3][2] ),
    .A1(_0137_),
    .S(_0336_),
    .X(_0339_));
 sky130_fd_sc_hd__clkbuf_1 _1955_ (.A(_0339_),
    .X(_0111_));
 sky130_fd_sc_hd__mux2_1 _1956_ (.A0(\MOS6502.AXYS[3][3] ),
    .A1(_0142_),
    .S(_0336_),
    .X(_0340_));
 sky130_fd_sc_hd__clkbuf_1 _1957_ (.A(_0340_),
    .X(_0112_));
 sky130_fd_sc_hd__mux2_1 _1958_ (.A0(\MOS6502.AXYS[3][4] ),
    .A1(_0144_),
    .S(_0336_),
    .X(_0341_));
 sky130_fd_sc_hd__clkbuf_1 _1959_ (.A(_0341_),
    .X(_0113_));
 sky130_fd_sc_hd__mux2_1 _1960_ (.A0(\MOS6502.AXYS[3][5] ),
    .A1(_0151_),
    .S(_0336_),
    .X(_0342_));
 sky130_fd_sc_hd__clkbuf_1 _1961_ (.A(_0342_),
    .X(_0114_));
 sky130_fd_sc_hd__mux2_1 _1962_ (.A0(\MOS6502.AXYS[3][6] ),
    .A1(_0157_),
    .S(_0336_),
    .X(_0343_));
 sky130_fd_sc_hd__clkbuf_1 _1963_ (.A(_0343_),
    .X(_0115_));
 sky130_fd_sc_hd__mux2_1 _1964_ (.A0(\MOS6502.AXYS[3][7] ),
    .A1(_0163_),
    .S(_0336_),
    .X(_0344_));
 sky130_fd_sc_hd__clkbuf_1 _1965_ (.A(_0344_),
    .X(_0116_));
 sky130_fd_sc_hd__and2_1 _1966_ (.A(_0497_),
    .B(_0968_),
    .X(_0345_));
 sky130_fd_sc_hd__clkbuf_4 _1967_ (.A(_0345_),
    .X(_0346_));
 sky130_fd_sc_hd__mux2_1 _1968_ (.A0(\MOS6502.AXYS[0][0] ),
    .A1(_0966_),
    .S(_0346_),
    .X(_0347_));
 sky130_fd_sc_hd__clkbuf_1 _1969_ (.A(_0347_),
    .X(_0117_));
 sky130_fd_sc_hd__mux2_1 _1970_ (.A0(\MOS6502.AXYS[0][1] ),
    .A1(_0131_),
    .S(_0346_),
    .X(_0348_));
 sky130_fd_sc_hd__clkbuf_1 _1971_ (.A(_0348_),
    .X(_0118_));
 sky130_fd_sc_hd__mux2_1 _1972_ (.A0(\MOS6502.AXYS[0][2] ),
    .A1(_0137_),
    .S(_0346_),
    .X(_0349_));
 sky130_fd_sc_hd__clkbuf_1 _1973_ (.A(_0349_),
    .X(_0119_));
 sky130_fd_sc_hd__mux2_1 _1974_ (.A0(\MOS6502.AXYS[0][3] ),
    .A1(_0142_),
    .S(_0346_),
    .X(_0350_));
 sky130_fd_sc_hd__clkbuf_1 _1975_ (.A(_0350_),
    .X(_0120_));
 sky130_fd_sc_hd__mux2_1 _1976_ (.A0(\MOS6502.AXYS[0][4] ),
    .A1(_0144_),
    .S(_0346_),
    .X(_0351_));
 sky130_fd_sc_hd__clkbuf_1 _1977_ (.A(_0351_),
    .X(_0121_));
 sky130_fd_sc_hd__mux2_1 _1978_ (.A0(\MOS6502.AXYS[0][5] ),
    .A1(_0151_),
    .S(_0346_),
    .X(_0352_));
 sky130_fd_sc_hd__clkbuf_1 _1979_ (.A(_0352_),
    .X(_0122_));
 sky130_fd_sc_hd__mux2_1 _1980_ (.A0(\MOS6502.AXYS[0][6] ),
    .A1(_0157_),
    .S(_0346_),
    .X(_0353_));
 sky130_fd_sc_hd__clkbuf_1 _1981_ (.A(_0353_),
    .X(_0123_));
 sky130_fd_sc_hd__mux2_1 _1982_ (.A0(\MOS6502.AXYS[0][7] ),
    .A1(_0163_),
    .S(_0346_),
    .X(_0354_));
 sky130_fd_sc_hd__clkbuf_1 _1983_ (.A(_0354_),
    .X(_0124_));
 sky130_fd_sc_hd__dfrtp_2 _1984_ (.CLK(clknet_4_6_0_clk),
    .D(_0018_),
    .RESET_B(_0024_),
    .Q(\MOS6502.state[0] ));
 sky130_fd_sc_hd__dfrtp_2 _1985_ (.CLK(clknet_4_6_0_clk),
    .D(_0019_),
    .RESET_B(_0025_),
    .Q(\MOS6502.state[1] ));
 sky130_fd_sc_hd__dfrtp_1 _1986_ (.CLK(clknet_4_6_0_clk),
    .D(_0020_),
    .RESET_B(_0026_),
    .Q(\MOS6502.state[2] ));
 sky130_fd_sc_hd__dfstp_1 _1987_ (.CLK(clknet_4_6_0_clk),
    .D(_0021_),
    .SET_B(_0027_),
    .Q(\MOS6502.state[3] ));
 sky130_fd_sc_hd__dfrtp_1 _1988_ (.CLK(clknet_4_12_0_clk),
    .D(_0022_),
    .RESET_B(_0028_),
    .Q(\MOS6502.state[4] ));
 sky130_fd_sc_hd__dfrtp_4 _1989_ (.CLK(clknet_4_12_0_clk),
    .D(_0023_),
    .RESET_B(_0029_),
    .Q(\MOS6502.state[5] ));
 sky130_fd_sc_hd__dfxtp_1 _1990_ (.CLK(clknet_4_1_0_clk),
    .D(_0030_),
    .Q(\MOS6502.AXYS[2][0] ));
 sky130_fd_sc_hd__dfxtp_1 _1991_ (.CLK(clknet_4_1_0_clk),
    .D(_0031_),
    .Q(\MOS6502.AXYS[2][1] ));
 sky130_fd_sc_hd__dfxtp_1 _1992_ (.CLK(clknet_4_0_0_clk),
    .D(_0032_),
    .Q(\MOS6502.AXYS[2][2] ));
 sky130_fd_sc_hd__dfxtp_1 _1993_ (.CLK(clknet_4_0_0_clk),
    .D(_0033_),
    .Q(\MOS6502.AXYS[2][3] ));
 sky130_fd_sc_hd__dfxtp_1 _1994_ (.CLK(clknet_4_2_0_clk),
    .D(_0034_),
    .Q(\MOS6502.AXYS[2][4] ));
 sky130_fd_sc_hd__dfxtp_1 _1995_ (.CLK(clknet_4_0_0_clk),
    .D(_0035_),
    .Q(\MOS6502.AXYS[2][5] ));
 sky130_fd_sc_hd__dfxtp_1 _1996_ (.CLK(clknet_4_2_0_clk),
    .D(_0036_),
    .Q(\MOS6502.AXYS[2][6] ));
 sky130_fd_sc_hd__dfxtp_1 _1997_ (.CLK(clknet_4_0_0_clk),
    .D(_0037_),
    .Q(\MOS6502.AXYS[2][7] ));
 sky130_fd_sc_hd__dfxtp_1 _1998_ (.CLK(clknet_4_1_0_clk),
    .D(_0038_),
    .Q(\MOS6502.AXYS[1][0] ));
 sky130_fd_sc_hd__dfxtp_1 _1999_ (.CLK(clknet_4_3_0_clk),
    .D(_0039_),
    .Q(\MOS6502.AXYS[1][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2000_ (.CLK(clknet_4_0_0_clk),
    .D(_0040_),
    .Q(\MOS6502.AXYS[1][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2001_ (.CLK(clknet_4_2_0_clk),
    .D(_0041_),
    .Q(\MOS6502.AXYS[1][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2002_ (.CLK(clknet_4_2_0_clk),
    .D(_0042_),
    .Q(\MOS6502.AXYS[1][4] ));
 sky130_fd_sc_hd__dfxtp_1 _2003_ (.CLK(clknet_4_0_0_clk),
    .D(_0043_),
    .Q(\MOS6502.AXYS[1][5] ));
 sky130_fd_sc_hd__dfxtp_1 _2004_ (.CLK(clknet_4_3_0_clk),
    .D(_0044_),
    .Q(\MOS6502.AXYS[1][6] ));
 sky130_fd_sc_hd__dfxtp_1 _2005_ (.CLK(clknet_4_0_0_clk),
    .D(_0045_),
    .Q(\MOS6502.AXYS[1][7] ));
 sky130_fd_sc_hd__dfxtp_4 _2006_ (.CLK(clknet_4_8_0_clk),
    .D(_0001_),
    .Q(\MOS6502.ALU.CO ));
 sky130_fd_sc_hd__dfxtp_4 _2007_ (.CLK(clknet_4_8_0_clk),
    .D(\MOS6502.ALU.temp[7] ),
    .Q(\MOS6502.ADD[7] ));
 sky130_fd_sc_hd__dfxtp_1 _2008_ (.CLK(clknet_4_2_0_clk),
    .D(\MOS6502.ALU.temp_HC ),
    .Q(\MOS6502.ALU.HC ));
 sky130_fd_sc_hd__dfxtp_2 _2009_ (.CLK(clknet_4_8_0_clk),
    .D(\MOS6502.ALU.temp[0] ),
    .Q(\MOS6502.ADD[0] ));
 sky130_fd_sc_hd__dfxtp_4 _2010_ (.CLK(clknet_4_2_0_clk),
    .D(\MOS6502.ALU.temp[1] ),
    .Q(\MOS6502.ADD[1] ));
 sky130_fd_sc_hd__dfxtp_4 _2011_ (.CLK(clknet_4_8_0_clk),
    .D(\MOS6502.ALU.temp[2] ),
    .Q(\MOS6502.ADD[2] ));
 sky130_fd_sc_hd__dfxtp_4 _2012_ (.CLK(clknet_4_8_0_clk),
    .D(\MOS6502.ALU.temp[3] ),
    .Q(\MOS6502.ADD[3] ));
 sky130_fd_sc_hd__dfxtp_2 _2013_ (.CLK(clknet_4_10_0_clk),
    .D(\MOS6502.ALU.temp[4] ),
    .Q(\MOS6502.ADD[4] ));
 sky130_fd_sc_hd__dfxtp_2 _2014_ (.CLK(clknet_4_10_0_clk),
    .D(\MOS6502.ALU.temp[5] ),
    .Q(\MOS6502.ADD[5] ));
 sky130_fd_sc_hd__dfxtp_4 _2015_ (.CLK(clknet_4_10_0_clk),
    .D(\MOS6502.ALU.temp[6] ),
    .Q(\MOS6502.ADD[6] ));
 sky130_fd_sc_hd__dfxtp_1 _2016_ (.CLK(clknet_4_2_0_clk),
    .D(\MOS6502.AI[7] ),
    .Q(\MOS6502.ALU.AI7 ));
 sky130_fd_sc_hd__dfxtp_1 _2017_ (.CLK(clknet_4_2_0_clk),
    .D(\MOS6502.ALU.temp_BI[7] ),
    .Q(\MOS6502.ALU.BI7 ));
 sky130_fd_sc_hd__dfxtp_1 _2018_ (.CLK(clknet_4_14_0_clk),
    .D(_0002_),
    .Q(\MOS6502.PC[0] ));
 sky130_fd_sc_hd__dfxtp_1 _2019_ (.CLK(clknet_4_10_0_clk),
    .D(_0009_),
    .Q(\MOS6502.PC[1] ));
 sky130_fd_sc_hd__dfxtp_1 _2020_ (.CLK(clknet_4_10_0_clk),
    .D(_0010_),
    .Q(\MOS6502.PC[2] ));
 sky130_fd_sc_hd__dfxtp_1 _2021_ (.CLK(clknet_4_11_0_clk),
    .D(_0011_),
    .Q(\MOS6502.PC[3] ));
 sky130_fd_sc_hd__dfxtp_1 _2022_ (.CLK(clknet_4_9_0_clk),
    .D(_0012_),
    .Q(\MOS6502.PC[4] ));
 sky130_fd_sc_hd__dfxtp_1 _2023_ (.CLK(clknet_4_11_0_clk),
    .D(_0013_),
    .Q(\MOS6502.PC[5] ));
 sky130_fd_sc_hd__dfxtp_1 _2024_ (.CLK(clknet_4_11_0_clk),
    .D(_0014_),
    .Q(\MOS6502.PC[6] ));
 sky130_fd_sc_hd__dfxtp_1 _2025_ (.CLK(clknet_4_14_0_clk),
    .D(_0015_),
    .Q(\MOS6502.PC[7] ));
 sky130_fd_sc_hd__dfxtp_1 _2026_ (.CLK(clknet_4_13_0_clk),
    .D(_0016_),
    .Q(\MOS6502.PC[8] ));
 sky130_fd_sc_hd__dfxtp_1 _2027_ (.CLK(clknet_4_13_0_clk),
    .D(_0017_),
    .Q(\MOS6502.PC[9] ));
 sky130_fd_sc_hd__dfxtp_1 _2028_ (.CLK(clknet_4_13_0_clk),
    .D(_0003_),
    .Q(\MOS6502.PC[10] ));
 sky130_fd_sc_hd__dfxtp_1 _2029_ (.CLK(clknet_4_15_0_clk),
    .D(_0004_),
    .Q(\MOS6502.PC[11] ));
 sky130_fd_sc_hd__dfxtp_1 _2030_ (.CLK(clknet_4_15_0_clk),
    .D(_0005_),
    .Q(\MOS6502.PC[12] ));
 sky130_fd_sc_hd__dfxtp_1 _2031_ (.CLK(clknet_4_15_0_clk),
    .D(_0006_),
    .Q(\MOS6502.PC[13] ));
 sky130_fd_sc_hd__dfxtp_1 _2032_ (.CLK(clknet_4_15_0_clk),
    .D(_0007_),
    .Q(\MOS6502.PC[14] ));
 sky130_fd_sc_hd__dfxtp_1 _2033_ (.CLK(clknet_4_15_0_clk),
    .D(_0008_),
    .Q(\MOS6502.PC[15] ));
 sky130_fd_sc_hd__dfxtp_1 _2034_ (.CLK(clknet_4_10_0_clk),
    .D(_0046_),
    .Q(\MOS6502.ABL[0] ));
 sky130_fd_sc_hd__dfxtp_1 _2035_ (.CLK(clknet_4_10_0_clk),
    .D(_0047_),
    .Q(\MOS6502.ABL[1] ));
 sky130_fd_sc_hd__dfxtp_1 _2036_ (.CLK(clknet_4_10_0_clk),
    .D(_0048_),
    .Q(\MOS6502.ABL[2] ));
 sky130_fd_sc_hd__dfxtp_1 _2037_ (.CLK(clknet_4_10_0_clk),
    .D(_0049_),
    .Q(\MOS6502.ABL[3] ));
 sky130_fd_sc_hd__dfxtp_1 _2038_ (.CLK(clknet_4_10_0_clk),
    .D(_0050_),
    .Q(\MOS6502.ABL[4] ));
 sky130_fd_sc_hd__dfxtp_1 _2039_ (.CLK(clknet_4_11_0_clk),
    .D(_0051_),
    .Q(\MOS6502.ABL[5] ));
 sky130_fd_sc_hd__dfxtp_1 _2040_ (.CLK(clknet_4_11_0_clk),
    .D(_0052_),
    .Q(\MOS6502.ABL[6] ));
 sky130_fd_sc_hd__dfxtp_1 _2041_ (.CLK(clknet_4_14_0_clk),
    .D(_0053_),
    .Q(\MOS6502.ABL[7] ));
 sky130_fd_sc_hd__dfxtp_1 _2042_ (.CLK(clknet_4_14_0_clk),
    .D(_0054_),
    .Q(\MOS6502.C ));
 sky130_fd_sc_hd__dfxtp_1 _2043_ (.CLK(clknet_4_3_0_clk),
    .D(_0000_),
    .Q(\MOS6502.adj_bcd ));
 sky130_fd_sc_hd__dfxtp_1 _2044_ (.CLK(clknet_4_9_0_clk),
    .D(net8),
    .Q(\MOS6502.backwards ));
 sky130_fd_sc_hd__dfxtp_1 _2045_ (.CLK(clknet_4_9_0_clk),
    .D(_0055_),
    .Q(\MOS6502.Z ));
 sky130_fd_sc_hd__dfxtp_1 _2046_ (.CLK(clknet_4_9_0_clk),
    .D(_0056_),
    .Q(\MOS6502.N ));
 sky130_fd_sc_hd__dfxtp_1 _2047_ (.CLK(clknet_4_3_0_clk),
    .D(_0057_),
    .Q(\MOS6502.D ));
 sky130_fd_sc_hd__dfxtp_1 _2048_ (.CLK(clknet_4_14_0_clk),
    .D(_0058_),
    .Q(\MOS6502.I ));
 sky130_fd_sc_hd__dfxtp_1 _2049_ (.CLK(clknet_4_3_0_clk),
    .D(_0059_),
    .Q(\MOS6502.V ));
 sky130_fd_sc_hd__dfxtp_1 _2050_ (.CLK(clknet_4_7_0_clk),
    .D(_0060_),
    .Q(\MOS6502.IRHOLD[0] ));
 sky130_fd_sc_hd__dfxtp_1 _2051_ (.CLK(clknet_4_7_0_clk),
    .D(_0061_),
    .Q(\MOS6502.IRHOLD[1] ));
 sky130_fd_sc_hd__dfxtp_1 _2052_ (.CLK(clknet_4_7_0_clk),
    .D(_0062_),
    .Q(\MOS6502.IRHOLD[2] ));
 sky130_fd_sc_hd__dfxtp_1 _2053_ (.CLK(clknet_4_7_0_clk),
    .D(_0063_),
    .Q(\MOS6502.IRHOLD[3] ));
 sky130_fd_sc_hd__dfxtp_1 _2054_ (.CLK(clknet_4_7_0_clk),
    .D(_0064_),
    .Q(\MOS6502.IRHOLD[4] ));
 sky130_fd_sc_hd__dfxtp_1 _2055_ (.CLK(clknet_4_7_0_clk),
    .D(_0065_),
    .Q(\MOS6502.IRHOLD[5] ));
 sky130_fd_sc_hd__dfxtp_1 _2056_ (.CLK(clknet_4_7_0_clk),
    .D(_0066_),
    .Q(\MOS6502.IRHOLD[6] ));
 sky130_fd_sc_hd__dfxtp_1 _2057_ (.CLK(clknet_4_7_0_clk),
    .D(_0067_),
    .Q(\MOS6502.IRHOLD[7] ));
 sky130_fd_sc_hd__dfxtp_2 _2058_ (.CLK(clknet_4_7_0_clk),
    .D(_0068_),
    .Q(\MOS6502.IRHOLD_valid ));
 sky130_fd_sc_hd__dfxtp_1 _2059_ (.CLK(clknet_4_1_0_clk),
    .D(_0069_),
    .Q(\MOS6502.load_reg ));
 sky130_fd_sc_hd__dfxtp_1 _2060_ (.CLK(clknet_4_13_0_clk),
    .D(_0070_),
    .Q(\MOS6502.res ));
 sky130_fd_sc_hd__dfxtp_1 _2061_ (.CLK(clknet_4_5_0_clk),
    .D(_0071_),
    .Q(\MOS6502.dst_reg[0] ));
 sky130_fd_sc_hd__dfxtp_1 _2062_ (.CLK(clknet_4_5_0_clk),
    .D(_0072_),
    .Q(\MOS6502.dst_reg[1] ));
 sky130_fd_sc_hd__dfxtp_1 _2063_ (.CLK(clknet_4_5_0_clk),
    .D(_0073_),
    .Q(\MOS6502.src_reg[0] ));
 sky130_fd_sc_hd__dfxtp_1 _2064_ (.CLK(clknet_4_7_0_clk),
    .D(_0074_),
    .Q(\MOS6502.src_reg[1] ));
 sky130_fd_sc_hd__dfxtp_1 _2065_ (.CLK(clknet_4_6_0_clk),
    .D(_0075_),
    .Q(\MOS6502.index_y ));
 sky130_fd_sc_hd__dfxtp_1 _2066_ (.CLK(clknet_4_7_0_clk),
    .D(_0076_),
    .Q(\MOS6502.store ));
 sky130_fd_sc_hd__dfxtp_1 _2067_ (.CLK(clknet_4_5_0_clk),
    .D(_0077_),
    .Q(\MOS6502.write_back ));
 sky130_fd_sc_hd__dfxtp_1 _2068_ (.CLK(clknet_4_4_0_clk),
    .D(_0078_),
    .Q(\MOS6502.load_only ));
 sky130_fd_sc_hd__dfxtp_1 _2069_ (.CLK(clknet_4_5_0_clk),
    .D(_0079_),
    .Q(\MOS6502.inc ));
 sky130_fd_sc_hd__dfxtp_1 _2070_ (.CLK(clknet_4_4_0_clk),
    .D(_0080_),
    .Q(\MOS6502.adc_sbc ));
 sky130_fd_sc_hd__dfxtp_1 _2071_ (.CLK(clknet_4_12_0_clk),
    .D(_0081_),
    .Q(\MOS6502.shift ));
 sky130_fd_sc_hd__dfxtp_1 _2072_ (.CLK(clknet_4_3_0_clk),
    .D(_0082_),
    .Q(\MOS6502.adc_bcd ));
 sky130_fd_sc_hd__dfxtp_1 _2073_ (.CLK(clknet_4_5_0_clk),
    .D(_0083_),
    .Q(\MOS6502.compare ));
 sky130_fd_sc_hd__dfxtp_1 _2074_ (.CLK(clknet_4_1_0_clk),
    .D(_0084_),
    .Q(\MOS6502.shift_right ));
 sky130_fd_sc_hd__dfxtp_1 _2075_ (.CLK(clknet_4_9_0_clk),
    .D(_0085_),
    .Q(\MOS6502.rotate ));
 sky130_fd_sc_hd__dfxtp_1 _2076_ (.CLK(clknet_4_1_0_clk),
    .D(_0086_),
    .Q(\MOS6502.op[0] ));
 sky130_fd_sc_hd__dfxtp_1 _2077_ (.CLK(clknet_4_1_0_clk),
    .D(_0087_),
    .Q(\MOS6502.op[1] ));
 sky130_fd_sc_hd__dfxtp_1 _2078_ (.CLK(clknet_4_1_0_clk),
    .D(_0088_),
    .Q(\MOS6502.op[2] ));
 sky130_fd_sc_hd__dfxtp_1 _2079_ (.CLK(clknet_4_4_0_clk),
    .D(_0089_),
    .Q(\MOS6502.op[3] ));
 sky130_fd_sc_hd__dfxtp_1 _2080_ (.CLK(clknet_4_4_0_clk),
    .D(_0090_),
    .Q(\MOS6502.bit_ins ));
 sky130_fd_sc_hd__dfxtp_1 _2081_ (.CLK(clknet_4_1_0_clk),
    .D(_0091_),
    .Q(\MOS6502.clv ));
 sky130_fd_sc_hd__dfxtp_1 _2082_ (.CLK(clknet_4_7_0_clk),
    .D(_0092_),
    .Q(\MOS6502.sei ));
 sky130_fd_sc_hd__dfxtp_1 _2083_ (.CLK(clknet_4_6_0_clk),
    .D(_0093_),
    .Q(\MOS6502.cli ));
 sky130_fd_sc_hd__dfxtp_1 _2084_ (.CLK(clknet_4_4_0_clk),
    .D(_0094_),
    .Q(\MOS6502.sed ));
 sky130_fd_sc_hd__dfxtp_1 _2085_ (.CLK(clknet_4_4_0_clk),
    .D(_0095_),
    .Q(\MOS6502.cld ));
 sky130_fd_sc_hd__dfxtp_1 _2086_ (.CLK(clknet_4_5_0_clk),
    .D(_0096_),
    .Q(\MOS6502.sec ));
 sky130_fd_sc_hd__dfxtp_1 _2087_ (.CLK(clknet_4_5_0_clk),
    .D(_0097_),
    .Q(\MOS6502.clc ));
 sky130_fd_sc_hd__dfxtp_2 _2088_ (.CLK(clknet_4_6_0_clk),
    .D(_0098_),
    .Q(\MOS6502.php ));
 sky130_fd_sc_hd__dfxtp_1 _2089_ (.CLK(clknet_4_6_0_clk),
    .D(_0099_),
    .Q(\MOS6502.plp ));
 sky130_fd_sc_hd__dfxtp_1 _2090_ (.CLK(clknet_4_9_0_clk),
    .D(\MOS6502.IR[5] ),
    .Q(\MOS6502.cond_code[0] ));
 sky130_fd_sc_hd__dfxtp_1 _2091_ (.CLK(clknet_4_1_0_clk),
    .D(\MOS6502.IR[6] ),
    .Q(\MOS6502.cond_code[1] ));
 sky130_fd_sc_hd__dfxtp_1 _2092_ (.CLK(clknet_4_1_0_clk),
    .D(\MOS6502.IR[7] ),
    .Q(\MOS6502.cond_code[2] ));
 sky130_fd_sc_hd__dfxtp_1 _2093_ (.CLK(clknet_4_12_0_clk),
    .D(net10),
    .Q(\MOS6502.NMI_1 ));
 sky130_fd_sc_hd__dfxtp_1 _2094_ (.CLK(clknet_4_12_0_clk),
    .D(_0100_),
    .Q(\MOS6502.NMI_edge ));
 sky130_fd_sc_hd__dfxtp_1 _2095_ (.CLK(clknet_4_14_0_clk),
    .D(_0101_),
    .Q(\MOS6502.ABH[0] ));
 sky130_fd_sc_hd__dfxtp_1 _2096_ (.CLK(clknet_4_14_0_clk),
    .D(_0102_),
    .Q(\MOS6502.ABH[1] ));
 sky130_fd_sc_hd__dfxtp_1 _2097_ (.CLK(clknet_4_15_0_clk),
    .D(_0103_),
    .Q(\MOS6502.ABH[2] ));
 sky130_fd_sc_hd__dfxtp_1 _2098_ (.CLK(clknet_4_13_0_clk),
    .D(_0104_),
    .Q(\MOS6502.ABH[3] ));
 sky130_fd_sc_hd__dfxtp_1 _2099_ (.CLK(clknet_4_15_0_clk),
    .D(_0105_),
    .Q(\MOS6502.ABH[4] ));
 sky130_fd_sc_hd__dfxtp_1 _2100_ (.CLK(clknet_4_15_0_clk),
    .D(_0106_),
    .Q(\MOS6502.ABH[5] ));
 sky130_fd_sc_hd__dfxtp_1 _2101_ (.CLK(clknet_4_13_0_clk),
    .D(_0107_),
    .Q(\MOS6502.ABH[6] ));
 sky130_fd_sc_hd__dfxtp_1 _2102_ (.CLK(clknet_4_15_0_clk),
    .D(_0108_),
    .Q(\MOS6502.ABH[7] ));
 sky130_fd_sc_hd__dfxtp_1 _2103_ (.CLK(clknet_4_1_0_clk),
    .D(_0109_),
    .Q(\MOS6502.AXYS[3][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2104_ (.CLK(clknet_4_0_0_clk),
    .D(_0110_),
    .Q(\MOS6502.AXYS[3][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2105_ (.CLK(clknet_4_0_0_clk),
    .D(_0111_),
    .Q(\MOS6502.AXYS[3][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2106_ (.CLK(clknet_4_0_0_clk),
    .D(_0112_),
    .Q(\MOS6502.AXYS[3][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2107_ (.CLK(clknet_4_2_0_clk),
    .D(_0113_),
    .Q(\MOS6502.AXYS[3][4] ));
 sky130_fd_sc_hd__dfxtp_1 _2108_ (.CLK(clknet_4_0_0_clk),
    .D(_0114_),
    .Q(\MOS6502.AXYS[3][5] ));
 sky130_fd_sc_hd__dfxtp_1 _2109_ (.CLK(clknet_4_2_0_clk),
    .D(_0115_),
    .Q(\MOS6502.AXYS[3][6] ));
 sky130_fd_sc_hd__dfxtp_1 _2110_ (.CLK(clknet_4_0_0_clk),
    .D(_0116_),
    .Q(\MOS6502.AXYS[3][7] ));
 sky130_fd_sc_hd__dfxtp_1 _2111_ (.CLK(clknet_4_0_0_clk),
    .D(_0117_),
    .Q(\MOS6502.AXYS[0][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2112_ (.CLK(clknet_4_3_0_clk),
    .D(_0118_),
    .Q(\MOS6502.AXYS[0][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2113_ (.CLK(clknet_4_0_0_clk),
    .D(_0119_),
    .Q(\MOS6502.AXYS[0][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2114_ (.CLK(clknet_4_2_0_clk),
    .D(_0120_),
    .Q(\MOS6502.AXYS[0][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2115_ (.CLK(clknet_4_2_0_clk),
    .D(_0121_),
    .Q(\MOS6502.AXYS[0][4] ));
 sky130_fd_sc_hd__dfxtp_1 _2116_ (.CLK(clknet_4_0_0_clk),
    .D(_0122_),
    .Q(\MOS6502.AXYS[0][5] ));
 sky130_fd_sc_hd__dfxtp_1 _2117_ (.CLK(clknet_4_3_0_clk),
    .D(_0123_),
    .Q(\MOS6502.AXYS[0][6] ));
 sky130_fd_sc_hd__dfxtp_1 _2118_ (.CLK(clknet_4_0_0_clk),
    .D(_0124_),
    .Q(\MOS6502.AXYS[0][7] ));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sky130_fd_sc_hd__buf_4 input1 (.A(io_in[0]),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 input10 (.A(io_in[9]),
    .X(net10));
 sky130_fd_sc_hd__buf_4 input11 (.A(rst),
    .X(net11));
 sky130_fd_sc_hd__buf_4 input2 (.A(io_in[1]),
    .X(net2));
 sky130_fd_sc_hd__buf_4 input3 (.A(io_in[2]),
    .X(net3));
 sky130_fd_sc_hd__buf_4 input4 (.A(io_in[3]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_4 input5 (.A(io_in[4]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_4 input6 (.A(io_in[5]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_4 input7 (.A(io_in[6]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_4 input8 (.A(io_in[7]),
    .X(net8));
 sky130_fd_sc_hd__dlymetal6s2s_1 input9 (.A(io_in[8]),
    .X(net9));
 sky130_fd_sc_hd__conb_1 wrapped_6502_12 (.LO(net12));
 sky130_fd_sc_hd__conb_1 wrapped_6502_13 (.LO(net13));
 assign io_out[8] = net12;
 assign io_out[9] = net13;
endmodule

