// This is the unpowered netlist.
module multiplexer (design_clk_o,
    dso_tune,
    oeb_6502,
    oeb_as1802,
    oeb_as2650,
    oeb_as512512512,
    oeb_as5401,
    oeb_mc14500,
    rst_6502,
    rst_LCD,
    rst_as1802,
    rst_as2650,
    rst_as512512512,
    rst_as5401,
    rst_counter,
    rst_diceroll,
    rst_mc14500,
    rst_posit,
    rst_tbb1143,
    rst_tune,
    wb_clk_i,
    wb_rst_i,
    wbs_ack_o,
    wbs_cyc_i,
    wbs_stb_i,
    wbs_we_i,
    dsi_all,
    dso_6502,
    dso_LCD,
    dso_as1802,
    dso_as2650,
    dso_as512512512,
    dso_as5401,
    dso_counter,
    dso_diceroll,
    dso_mc14500,
    dso_multiplier,
    dso_posit,
    dso_tbb1143,
    io_in,
    io_oeb,
    io_out,
    wbs_adr_i,
    wbs_dat_i,
    wbs_dat_o);
 output design_clk_o;
 input dso_tune;
 input oeb_6502;
 input oeb_as1802;
 input oeb_as2650;
 input oeb_as512512512;
 input oeb_as5401;
 input oeb_mc14500;
 output rst_6502;
 output rst_LCD;
 output rst_as1802;
 output rst_as2650;
 output rst_as512512512;
 output rst_as5401;
 output rst_counter;
 output rst_diceroll;
 output rst_mc14500;
 output rst_posit;
 output rst_tbb1143;
 output rst_tune;
 input wb_clk_i;
 input wb_rst_i;
 output wbs_ack_o;
 input wbs_cyc_i;
 input wbs_stb_i;
 input wbs_we_i;
 output [27:0] dsi_all;
 input [26:0] dso_6502;
 input [7:0] dso_LCD;
 input [26:0] dso_as1802;
 input [26:0] dso_as2650;
 input [27:0] dso_as512512512;
 input [26:0] dso_as5401;
 input [11:0] dso_counter;
 input [7:0] dso_diceroll;
 input [8:0] dso_mc14500;
 input [7:0] dso_multiplier;
 input [3:0] dso_posit;
 input [7:0] dso_tbb1143;
 input [37:0] io_in;
 output [37:0] io_oeb;
 output [37:0] io_out;
 input [31:0] wbs_adr_i;
 input [31:0] wbs_dat_i;
 output [31:0] wbs_dat_o;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire \design_addr[0] ;
 wire \design_addr[1] ;
 wire \design_addr[2] ;
 wire \design_addr[3] ;
 wire clknet_0_wb_clk_i;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net487;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire wb_clk_override;
 wire \wb_counter[0] ;
 wire \wb_counter[10] ;
 wire \wb_counter[11] ;
 wire \wb_counter[12] ;
 wire \wb_counter[13] ;
 wire \wb_counter[14] ;
 wire \wb_counter[15] ;
 wire \wb_counter[16] ;
 wire \wb_counter[17] ;
 wire \wb_counter[18] ;
 wire \wb_counter[19] ;
 wire \wb_counter[20] ;
 wire \wb_counter[21] ;
 wire \wb_counter[22] ;
 wire \wb_counter[23] ;
 wire \wb_counter[5] ;
 wire \wb_counter[6] ;
 wire \wb_counter[7] ;
 wire \wb_counter[8] ;
 wire \wb_counter[9] ;
 wire \wb_design_addr_override[0] ;
 wire \wb_design_addr_override[1] ;
 wire \wb_design_addr_override[2] ;
 wire \wb_design_addr_override[3] ;
 wire wb_feedback_delay;
 wire \wb_io_override[0] ;
 wire \wb_io_override[10] ;
 wire \wb_io_override[11] ;
 wire \wb_io_override[12] ;
 wire \wb_io_override[13] ;
 wire \wb_io_override[14] ;
 wire \wb_io_override[15] ;
 wire \wb_io_override[16] ;
 wire \wb_io_override[17] ;
 wire \wb_io_override[18] ;
 wire \wb_io_override[19] ;
 wire \wb_io_override[1] ;
 wire \wb_io_override[20] ;
 wire \wb_io_override[21] ;
 wire \wb_io_override[22] ;
 wire \wb_io_override[23] ;
 wire \wb_io_override[24] ;
 wire \wb_io_override[25] ;
 wire \wb_io_override[26] ;
 wire \wb_io_override[27] ;
 wire \wb_io_override[2] ;
 wire \wb_io_override[3] ;
 wire \wb_io_override[4] ;
 wire \wb_io_override[5] ;
 wire \wb_io_override[6] ;
 wire \wb_io_override[7] ;
 wire \wb_io_override[8] ;
 wire \wb_io_override[9] ;
 wire wb_override;
 wire wb_rst_override;
 wire wb_single_step;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire clknet_3_0__leaf_wb_clk_i;
 wire clknet_3_1__leaf_wb_clk_i;
 wire clknet_3_2__leaf_wb_clk_i;
 wire clknet_3_3__leaf_wb_clk_i;
 wire clknet_3_4__leaf_wb_clk_i;
 wire clknet_3_5__leaf_wb_clk_i;
 wire clknet_3_6__leaf_wb_clk_i;
 wire clknet_3_7__leaf_wb_clk_i;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;

 sky130_fd_sc_hd__inv_2 _0446_ (.A(net516),
    .Y(_0172_));
 sky130_fd_sc_hd__inv_2 _0447_ (.A(net519),
    .Y(_0173_));
 sky130_fd_sc_hd__inv_2 _0448_ (.A(net525),
    .Y(_0174_));
 sky130_fd_sc_hd__clkinv_2 _0449_ (.A(net513),
    .Y(_0175_));
 sky130_fd_sc_hd__inv_2 _0450_ (.A(net358),
    .Y(_0176_));
 sky130_fd_sc_hd__inv_2 _0451_ (.A(\wb_design_addr_override[3] ),
    .Y(_0177_));
 sky130_fd_sc_hd__inv_2 _0452_ (.A(\wb_design_addr_override[2] ),
    .Y(_0178_));
 sky130_fd_sc_hd__inv_2 _0453_ (.A(net470),
    .Y(_0179_));
 sky130_fd_sc_hd__inv_2 _0454_ (.A(net269),
    .Y(_0180_));
 sky130_fd_sc_hd__clkinv_2 _0455_ (.A(net471),
    .Y(_0181_));
 sky130_fd_sc_hd__inv_2 _0456_ (.A(net474),
    .Y(_0182_));
 sky130_fd_sc_hd__inv_2 _0457_ (.A(net460),
    .Y(_0183_));
 sky130_fd_sc_hd__nor3_2 _0458_ (.A(net457),
    .B(net451),
    .C(net454),
    .Y(_0184_));
 sky130_fd_sc_hd__nor4b_2 _0459_ (.A(net456),
    .B(net449),
    .C(net452),
    .D_N(net458),
    .Y(_0185_));
 sky130_fd_sc_hd__mux2_4 _0460_ (.A0(net228),
    .A1(wb_rst_override),
    .S(net442),
    .X(_0186_));
 sky130_fd_sc_hd__nand2b_1 _0461_ (.A_N(net436),
    .B(net440),
    .Y(net364));
 sky130_fd_sc_hd__nor4b_4 _0462_ (.A(net458),
    .B(net449),
    .C(net453),
    .D_N(net455),
    .Y(_0187_));
 sky130_fd_sc_hd__nand2b_1 _0463_ (.A_N(net436),
    .B(net435),
    .Y(net366));
 sky130_fd_sc_hd__nand2_2 _0464_ (.A(net457),
    .B(net460),
    .Y(_0188_));
 sky130_fd_sc_hd__and3b_2 _0465_ (.A_N(net454),
    .B(net460),
    .C(net457),
    .X(_0189_));
 sky130_fd_sc_hd__and4bb_4 _0466_ (.A_N(net451),
    .B_N(net454),
    .C(net455),
    .D(net458),
    .X(_0190_));
 sky130_fd_sc_hd__nand2b_1 _0467_ (.A_N(_0186_),
    .B(_0190_),
    .Y(net360));
 sky130_fd_sc_hd__and2b_2 _0468_ (.A_N(net451),
    .B(net454),
    .X(_0191_));
 sky130_fd_sc_hd__nand2b_1 _0469_ (.A_N(net451),
    .B(net454),
    .Y(_0192_));
 sky130_fd_sc_hd__nor4b_4 _0470_ (.A(net455),
    .B(net458),
    .C(net450),
    .D_N(net453),
    .Y(_0193_));
 sky130_fd_sc_hd__nand2b_1 _0471_ (.A_N(net436),
    .B(net434),
    .Y(net367));
 sky130_fd_sc_hd__and4bb_4 _0472_ (.A_N(net455),
    .B_N(net451),
    .C(net454),
    .D(net458),
    .X(_0194_));
 sky130_fd_sc_hd__nand2b_1 _0473_ (.A_N(net436),
    .B(net433),
    .Y(net365));
 sky130_fd_sc_hd__and4bb_4 _0474_ (.A_N(net458),
    .B_N(net449),
    .C(net452),
    .D(net455),
    .X(_0195_));
 sky130_fd_sc_hd__nand2b_1 _0475_ (.A_N(net436),
    .B(_0195_),
    .Y(net369));
 sky130_fd_sc_hd__and4b_4 _0476_ (.A_N(net449),
    .B(net452),
    .C(net455),
    .D(net459),
    .X(_0196_));
 sky130_fd_sc_hd__or3_2 _0477_ (.A(_0186_),
    .B(_0188_),
    .C(_0192_),
    .X(net362));
 sky130_fd_sc_hd__nor3b_2 _0478_ (.A(net457),
    .B(net454),
    .C_N(net451),
    .Y(_0197_));
 sky130_fd_sc_hd__nor4b_4 _0479_ (.A(net455),
    .B(net458),
    .C(net452),
    .D_N(net450),
    .Y(_0198_));
 sky130_fd_sc_hd__nand2b_1 _0480_ (.A_N(net436),
    .B(net426),
    .Y(net359));
 sky130_fd_sc_hd__and4bb_4 _0481_ (.A_N(net455),
    .B_N(net452),
    .C(net449),
    .D(net458),
    .X(_0199_));
 sky130_fd_sc_hd__nand2b_1 _0482_ (.A_N(net436),
    .B(net423),
    .Y(net361));
 sky130_fd_sc_hd__and4bb_4 _0483_ (.A_N(net459),
    .B_N(net452),
    .C(net449),
    .D(net456),
    .X(_0200_));
 sky130_fd_sc_hd__nand2b_1 _0484_ (.A_N(net436),
    .B(_0200_),
    .Y(net370));
 sky130_fd_sc_hd__and4b_4 _0485_ (.A_N(net453),
    .B(net451),
    .C(net458),
    .D(net455),
    .X(_0201_));
 sky130_fd_sc_hd__nand2b_1 _0486_ (.A_N(net436),
    .B(_0201_),
    .Y(net368));
 sky130_fd_sc_hd__and4bb_2 _0487_ (.A_N(net455),
    .B_N(net458),
    .C(net450),
    .D(net453),
    .X(_0202_));
 sky130_fd_sc_hd__nand2b_1 _0488_ (.A_N(net436),
    .B(net420),
    .Y(net363));
 sky130_fd_sc_hd__and2_1 _0489_ (.A(net232),
    .B(net420),
    .X(_0203_));
 sky130_fd_sc_hd__a22o_2 _0490_ (.A1(net229),
    .A2(net425),
    .B1(net421),
    .B2(net230),
    .X(_0204_));
 sky130_fd_sc_hd__a22o_1 _0491_ (.A1(_0183_),
    .A2(_0191_),
    .B1(net429),
    .B2(net231),
    .X(_0205_));
 sky130_fd_sc_hd__o21a_1 _0492_ (.A1(_0183_),
    .A2(net233),
    .B1(_0184_),
    .X(_0206_));
 sky130_fd_sc_hd__or4_4 _0493_ (.A(_0203_),
    .B(_0204_),
    .C(_0205_),
    .D(_0206_),
    .X(net303));
 sky130_fd_sc_hd__nor2_2 _0494_ (.A(_0201_),
    .B(net303),
    .Y(_0207_));
 sky130_fd_sc_hd__inv_2 _0495_ (.A(_0207_),
    .Y(net302));
 sky130_fd_sc_hd__or2_1 _0496_ (.A(net435),
    .B(net302),
    .X(net300));
 sky130_fd_sc_hd__a211o_1 _0497_ (.A1(net231),
    .A2(net429),
    .B1(_0201_),
    .C1(_0184_),
    .X(_0208_));
 sky130_fd_sc_hd__or3_4 _0498_ (.A(_0203_),
    .B(_0204_),
    .C(_0208_),
    .X(net307));
 sky130_fd_sc_hd__or2_2 _0499_ (.A(net432),
    .B(net307),
    .X(net305));
 sky130_fd_sc_hd__a211o_4 _0500_ (.A1(net234),
    .A2(net434),
    .B1(net432),
    .C1(net307),
    .X(net304));
 sky130_fd_sc_hd__a21o_1 _0501_ (.A1(net232),
    .A2(net420),
    .B1(_0189_),
    .X(_0209_));
 sky130_fd_sc_hd__or3_4 _0502_ (.A(net440),
    .B(_0197_),
    .C(_0209_),
    .X(net309));
 sky130_fd_sc_hd__or2_4 _0503_ (.A(net422),
    .B(_0209_),
    .X(net311));
 sky130_fd_sc_hd__or2_4 _0504_ (.A(net433),
    .B(net311),
    .X(net312));
 sky130_fd_sc_hd__o21ba_2 _0505_ (.A1(net457),
    .A2(_0192_),
    .B1_N(_0209_),
    .X(_0210_));
 sky130_fd_sc_hd__inv_2 _0506_ (.A(_0210_),
    .Y(net313));
 sky130_fd_sc_hd__a21o_4 _0507_ (.A1(_0188_),
    .A2(_0191_),
    .B1(_0209_),
    .X(net315));
 sky130_fd_sc_hd__nor4_4 _0508_ (.A(net456),
    .B(net459),
    .C(net449),
    .D(net452),
    .Y(_0211_));
 sky130_fd_sc_hd__a211o_2 _0509_ (.A1(_0188_),
    .A2(_0191_),
    .B1(_0211_),
    .C1(_0189_),
    .X(net325));
 sky130_fd_sc_hd__or2_4 _0510_ (.A(net420),
    .B(net415),
    .X(net326));
 sky130_fd_sc_hd__or3_4 _0511_ (.A(_0184_),
    .B(_0189_),
    .C(_0191_),
    .X(net299));
 sky130_fd_sc_hd__and2_4 _0512_ (.A(net194),
    .B(_0200_),
    .X(_0212_));
 sky130_fd_sc_hd__a22o_1 _0513_ (.A1(net118),
    .A2(net437),
    .B1(_0201_),
    .B2(net182),
    .X(_0213_));
 sky130_fd_sc_hd__a221o_1 _0514_ (.A1(net36),
    .A2(net422),
    .B1(net420),
    .B2(net90),
    .C1(net414),
    .X(_0214_));
 sky130_fd_sc_hd__a22o_4 _0515_ (.A1(net28),
    .A2(_0190_),
    .B1(_0194_),
    .B2(net145),
    .X(_0215_));
 sky130_fd_sc_hd__a221o_1 _0516_ (.A1(net63),
    .A2(net430),
    .B1(net426),
    .B2(net1),
    .C1(_0213_),
    .X(_0216_));
 sky130_fd_sc_hd__or3_4 _0517_ (.A(_0214_),
    .B(_0215_),
    .C(_0216_),
    .X(net328));
 sky130_fd_sc_hd__a22o_1 _0518_ (.A1(net129),
    .A2(net437),
    .B1(_0201_),
    .B2(net183),
    .X(_0217_));
 sky130_fd_sc_hd__a22o_4 _0519_ (.A1(net29),
    .A2(_0190_),
    .B1(_0194_),
    .B2(net148),
    .X(_0218_));
 sky130_fd_sc_hd__a22o_1 _0520_ (.A1(net12),
    .A2(net428),
    .B1(net420),
    .B2(net101),
    .X(_0219_));
 sky130_fd_sc_hd__a221o_1 _0521_ (.A1(net157),
    .A2(_0187_),
    .B1(net423),
    .B2(net47),
    .C1(_0217_),
    .X(_0220_));
 sky130_fd_sc_hd__a211o_1 _0522_ (.A1(net74),
    .A2(net429),
    .B1(_0212_),
    .C1(_0219_),
    .X(_0221_));
 sky130_fd_sc_hd__or3_4 _0523_ (.A(_0218_),
    .B(_0220_),
    .C(_0221_),
    .X(net329));
 sky130_fd_sc_hd__o211a_2 _0524_ (.A1(net456),
    .A2(net459),
    .B1(net449),
    .C1(net452),
    .X(_0222_));
 sky130_fd_sc_hd__a21o_4 _0525_ (.A1(net194),
    .A2(_0200_),
    .B1(_0222_),
    .X(_0223_));
 sky130_fd_sc_hd__a22o_1 _0526_ (.A1(net158),
    .A2(net435),
    .B1(net425),
    .B2(net20),
    .X(_0224_));
 sky130_fd_sc_hd__a21o_1 _0527_ (.A1(net55),
    .A2(net421),
    .B1(_0224_),
    .X(_0225_));
 sky130_fd_sc_hd__a221o_4 _0528_ (.A1(net30),
    .A2(_0190_),
    .B1(_0194_),
    .B2(net149),
    .C1(_0223_),
    .X(_0226_));
 sky130_fd_sc_hd__a22o_4 _0529_ (.A1(net82),
    .A2(net431),
    .B1(net418),
    .B2(net110),
    .X(_0227_));
 sky130_fd_sc_hd__a221o_1 _0530_ (.A1(net137),
    .A2(net437),
    .B1(_0201_),
    .B2(net184),
    .C1(_0227_),
    .X(_0228_));
 sky130_fd_sc_hd__or3_4 _0531_ (.A(_0225_),
    .B(_0226_),
    .C(_0228_),
    .X(net330));
 sky130_fd_sc_hd__a22o_1 _0532_ (.A1(net138),
    .A2(net437),
    .B1(net421),
    .B2(net56),
    .X(_0229_));
 sky130_fd_sc_hd__a22o_2 _0533_ (.A1(net31),
    .A2(_0190_),
    .B1(_0194_),
    .B2(net150),
    .X(_0230_));
 sky130_fd_sc_hd__a22o_1 _0534_ (.A1(net159),
    .A2(net435),
    .B1(net428),
    .B2(net21),
    .X(_0231_));
 sky130_fd_sc_hd__a22o_1 _0535_ (.A1(net83),
    .A2(net431),
    .B1(net418),
    .B2(net111),
    .X(_0232_));
 sky130_fd_sc_hd__or4_4 _0536_ (.A(_0223_),
    .B(_0230_),
    .C(_0231_),
    .D(_0232_),
    .X(_0233_));
 sky130_fd_sc_hd__a211o_2 _0537_ (.A1(net185),
    .A2(_0201_),
    .B1(_0229_),
    .C1(_0233_),
    .X(net331));
 sky130_fd_sc_hd__a22o_1 _0538_ (.A1(net139),
    .A2(net439),
    .B1(net424),
    .B2(net57),
    .X(_0234_));
 sky130_fd_sc_hd__a21o_2 _0539_ (.A1(net151),
    .A2(net433),
    .B1(_0234_),
    .X(_0235_));
 sky130_fd_sc_hd__a221o_2 _0540_ (.A1(net22),
    .A2(net427),
    .B1(net419),
    .B2(net112),
    .C1(_0212_),
    .X(_0236_));
 sky130_fd_sc_hd__a22o_2 _0541_ (.A1(net160),
    .A2(net435),
    .B1(_0190_),
    .B2(net32),
    .X(_0237_));
 sky130_fd_sc_hd__a221o_4 _0542_ (.A1(net165),
    .A2(net434),
    .B1(net429),
    .B2(net84),
    .C1(_0237_),
    .X(_0238_));
 sky130_fd_sc_hd__or3_4 _0543_ (.A(_0235_),
    .B(_0236_),
    .C(_0238_),
    .X(net332));
 sky130_fd_sc_hd__a22o_1 _0544_ (.A1(net140),
    .A2(net438),
    .B1(net427),
    .B2(net23),
    .X(_0239_));
 sky130_fd_sc_hd__a21o_2 _0545_ (.A1(net152),
    .A2(net433),
    .B1(_0239_),
    .X(_0240_));
 sky130_fd_sc_hd__a22o_1 _0546_ (.A1(net33),
    .A2(_0190_),
    .B1(net419),
    .B2(net113),
    .X(_0241_));
 sky130_fd_sc_hd__a22o_2 _0547_ (.A1(net161),
    .A2(net435),
    .B1(net431),
    .B2(net85),
    .X(_0242_));
 sky130_fd_sc_hd__and2_1 _0548_ (.A(net58),
    .B(net423),
    .X(_0243_));
 sky130_fd_sc_hd__a22o_1 _0549_ (.A1(net166),
    .A2(_0193_),
    .B1(_0200_),
    .B2(net194),
    .X(_0244_));
 sky130_fd_sc_hd__or4_1 _0550_ (.A(_0241_),
    .B(_0242_),
    .C(_0243_),
    .D(_0244_),
    .X(_0245_));
 sky130_fd_sc_hd__or2_4 _0551_ (.A(_0240_),
    .B(_0245_),
    .X(net333));
 sky130_fd_sc_hd__a22o_1 _0552_ (.A1(net59),
    .A2(net423),
    .B1(net418),
    .B2(net114),
    .X(_0246_));
 sky130_fd_sc_hd__a22o_1 _0553_ (.A1(net34),
    .A2(_0190_),
    .B1(net432),
    .B2(net186),
    .X(_0247_));
 sky130_fd_sc_hd__a221o_1 _0554_ (.A1(net167),
    .A2(net434),
    .B1(net433),
    .B2(net153),
    .C1(_0247_),
    .X(_0248_));
 sky130_fd_sc_hd__a221o_1 _0555_ (.A1(net162),
    .A2(net435),
    .B1(net427),
    .B2(net24),
    .C1(_0246_),
    .X(_0249_));
 sky130_fd_sc_hd__a221o_2 _0556_ (.A1(net141),
    .A2(net438),
    .B1(net431),
    .B2(net86),
    .C1(_0223_),
    .X(_0250_));
 sky130_fd_sc_hd__or3_4 _0557_ (.A(_0248_),
    .B(_0249_),
    .C(_0250_),
    .X(net334));
 sky130_fd_sc_hd__a22o_2 _0558_ (.A1(net142),
    .A2(net439),
    .B1(net433),
    .B2(net154),
    .X(_0251_));
 sky130_fd_sc_hd__a221o_2 _0559_ (.A1(net25),
    .A2(net428),
    .B1(net424),
    .B2(net60),
    .C1(_0251_),
    .X(_0252_));
 sky130_fd_sc_hd__a22o_1 _0560_ (.A1(net163),
    .A2(net435),
    .B1(net432),
    .B2(net187),
    .X(_0253_));
 sky130_fd_sc_hd__a211o_1 _0561_ (.A1(net87),
    .A2(net429),
    .B1(_0212_),
    .C1(_0253_),
    .X(_0254_));
 sky130_fd_sc_hd__a22o_2 _0562_ (.A1(net168),
    .A2(net434),
    .B1(net418),
    .B2(net115),
    .X(_0255_));
 sky130_fd_sc_hd__a21o_1 _0563_ (.A1(net35),
    .A2(_0190_),
    .B1(_0255_),
    .X(_0256_));
 sky130_fd_sc_hd__or3_4 _0564_ (.A(_0252_),
    .B(_0254_),
    .C(_0256_),
    .X(net335));
 sky130_fd_sc_hd__a22o_1 _0565_ (.A1(net88),
    .A2(net431),
    .B1(net427),
    .B2(net26),
    .X(_0257_));
 sky130_fd_sc_hd__a221o_4 _0566_ (.A1(net143),
    .A2(net438),
    .B1(net435),
    .B2(net164),
    .C1(_0257_),
    .X(_0258_));
 sky130_fd_sc_hd__a22o_1 _0567_ (.A1(net169),
    .A2(net434),
    .B1(net433),
    .B2(net155),
    .X(_0259_));
 sky130_fd_sc_hd__a221o_4 _0568_ (.A1(net188),
    .A2(net432),
    .B1(net417),
    .B2(net174),
    .C1(_0259_),
    .X(_0260_));
 sky130_fd_sc_hd__a22o_1 _0569_ (.A1(net61),
    .A2(net423),
    .B1(net418),
    .B2(net116),
    .X(_0261_));
 sky130_fd_sc_hd__nor4_4 _0570_ (.A(_0223_),
    .B(_0258_),
    .C(_0260_),
    .D(_0261_),
    .Y(_0262_));
 sky130_fd_sc_hd__inv_2 _0571_ (.A(_0262_),
    .Y(net336));
 sky130_fd_sc_hd__a22o_2 _0572_ (.A1(net170),
    .A2(net434),
    .B1(net417),
    .B2(net175),
    .X(_0263_));
 sky130_fd_sc_hd__a22o_2 _0573_ (.A1(net144),
    .A2(net438),
    .B1(net432),
    .B2(net189),
    .X(_0264_));
 sky130_fd_sc_hd__a22o_1 _0574_ (.A1(net89),
    .A2(net431),
    .B1(net418),
    .B2(net117),
    .X(_0265_));
 sky130_fd_sc_hd__a221o_2 _0575_ (.A1(net27),
    .A2(net427),
    .B1(net423),
    .B2(net62),
    .C1(_0265_),
    .X(_0266_));
 sky130_fd_sc_hd__a21oi_1 _0576_ (.A1(net156),
    .A2(net433),
    .B1(_0263_),
    .Y(_0267_));
 sky130_fd_sc_hd__nor4b_4 _0577_ (.A(net414),
    .B(_0264_),
    .C(_0266_),
    .D_N(_0267_),
    .Y(_0268_));
 sky130_fd_sc_hd__inv_2 _0578_ (.A(_0268_),
    .Y(net338));
 sky130_fd_sc_hd__and2_1 _0579_ (.A(net37),
    .B(net423),
    .X(_0269_));
 sky130_fd_sc_hd__a21o_4 _0580_ (.A1(net194),
    .A2(_0200_),
    .B1(net435),
    .X(_0270_));
 sky130_fd_sc_hd__a22o_2 _0581_ (.A1(net190),
    .A2(net432),
    .B1(net417),
    .B2(net176),
    .X(_0271_));
 sky130_fd_sc_hd__a221o_1 _0582_ (.A1(net171),
    .A2(net434),
    .B1(net433),
    .B2(net146),
    .C1(_0270_),
    .X(_0272_));
 sky130_fd_sc_hd__a22o_1 _0583_ (.A1(net2),
    .A2(net427),
    .B1(net418),
    .B2(net91),
    .X(_0273_));
 sky130_fd_sc_hd__a221o_2 _0584_ (.A1(net119),
    .A2(net438),
    .B1(net431),
    .B2(net64),
    .C1(_0273_),
    .X(_0274_));
 sky130_fd_sc_hd__or4_4 _0585_ (.A(_0269_),
    .B(_0271_),
    .C(_0272_),
    .D(_0274_),
    .X(net339));
 sky130_fd_sc_hd__a22o_1 _0586_ (.A1(net120),
    .A2(net438),
    .B1(net432),
    .B2(net191),
    .X(_0275_));
 sky130_fd_sc_hd__a22o_1 _0587_ (.A1(net65),
    .A2(net431),
    .B1(net418),
    .B2(net92),
    .X(_0276_));
 sky130_fd_sc_hd__a211o_1 _0588_ (.A1(net38),
    .A2(net423),
    .B1(net414),
    .C1(_0275_),
    .X(_0277_));
 sky130_fd_sc_hd__a22o_1 _0589_ (.A1(net172),
    .A2(net434),
    .B1(net433),
    .B2(net147),
    .X(_0278_));
 sky130_fd_sc_hd__a221o_1 _0590_ (.A1(net3),
    .A2(net427),
    .B1(_0211_),
    .B2(net177),
    .C1(_0276_),
    .X(_0279_));
 sky130_fd_sc_hd__or3_4 _0591_ (.A(_0277_),
    .B(_0278_),
    .C(_0279_),
    .X(net340));
 sky130_fd_sc_hd__a22o_4 _0592_ (.A1(net4),
    .A2(net425),
    .B1(net422),
    .B2(net39),
    .X(_0280_));
 sky130_fd_sc_hd__a22o_2 _0593_ (.A1(net192),
    .A2(net432),
    .B1(net417),
    .B2(net178),
    .X(_0281_));
 sky130_fd_sc_hd__or3_1 _0594_ (.A(net456),
    .B(net459),
    .C(net93),
    .X(_0282_));
 sky130_fd_sc_hd__a32o_1 _0595_ (.A1(net449),
    .A2(net452),
    .A3(_0282_),
    .B1(net434),
    .B2(net173),
    .X(_0283_));
 sky130_fd_sc_hd__a2111o_4 _0596_ (.A1(net66),
    .A2(net429),
    .B1(_0270_),
    .C1(_0281_),
    .D1(_0283_),
    .X(_0284_));
 sky130_fd_sc_hd__a211oi_4 _0597_ (.A1(net121),
    .A2(net437),
    .B1(_0280_),
    .C1(_0284_),
    .Y(_0285_));
 sky130_fd_sc_hd__inv_2 _0598_ (.A(_0285_),
    .Y(net341));
 sky130_fd_sc_hd__a22o_1 _0599_ (.A1(net193),
    .A2(net432),
    .B1(net417),
    .B2(net179),
    .X(_0286_));
 sky130_fd_sc_hd__a221o_1 _0600_ (.A1(net122),
    .A2(net438),
    .B1(net418),
    .B2(net94),
    .C1(_0223_),
    .X(_0287_));
 sky130_fd_sc_hd__a22o_4 _0601_ (.A1(net5),
    .A2(net425),
    .B1(net421),
    .B2(net40),
    .X(_0288_));
 sky130_fd_sc_hd__a211o_1 _0602_ (.A1(net67),
    .A2(net431),
    .B1(_0286_),
    .C1(_0288_),
    .X(_0289_));
 sky130_fd_sc_hd__or2_4 _0603_ (.A(_0287_),
    .B(_0289_),
    .X(net342));
 sky130_fd_sc_hd__a221o_2 _0604_ (.A1(net123),
    .A2(net440),
    .B1(net423),
    .B2(net41),
    .C1(_0270_),
    .X(_0290_));
 sky130_fd_sc_hd__a22o_2 _0605_ (.A1(net95),
    .A2(net418),
    .B1(net417),
    .B2(net180),
    .X(_0291_));
 sky130_fd_sc_hd__a221o_1 _0606_ (.A1(net68),
    .A2(net429),
    .B1(net427),
    .B2(net6),
    .C1(_0291_),
    .X(_0292_));
 sky130_fd_sc_hd__or2_4 _0607_ (.A(_0290_),
    .B(_0292_),
    .X(net343));
 sky130_fd_sc_hd__a22o_1 _0608_ (.A1(net7),
    .A2(net427),
    .B1(net420),
    .B2(net96),
    .X(_0293_));
 sky130_fd_sc_hd__a22o_2 _0609_ (.A1(net124),
    .A2(net438),
    .B1(_0211_),
    .B2(net181),
    .X(_0294_));
 sky130_fd_sc_hd__a211o_1 _0610_ (.A1(net42),
    .A2(net423),
    .B1(net414),
    .C1(_0294_),
    .X(_0295_));
 sky130_fd_sc_hd__a211o_4 _0611_ (.A1(net69),
    .A2(net429),
    .B1(_0293_),
    .C1(_0295_),
    .X(net344));
 sky130_fd_sc_hd__a22o_2 _0612_ (.A1(net125),
    .A2(net437),
    .B1(net424),
    .B2(net43),
    .X(_0296_));
 sky130_fd_sc_hd__a311o_1 _0613_ (.A1(net450),
    .A2(net453),
    .A3(net97),
    .B1(_0222_),
    .C1(_0296_),
    .X(_0297_));
 sky130_fd_sc_hd__a221o_1 _0614_ (.A1(net70),
    .A2(net429),
    .B1(net427),
    .B2(net8),
    .C1(_0270_),
    .X(_0298_));
 sky130_fd_sc_hd__or2_4 _0615_ (.A(_0297_),
    .B(_0298_),
    .X(net345));
 sky130_fd_sc_hd__a22o_4 _0616_ (.A1(net126),
    .A2(net439),
    .B1(net420),
    .B2(net98),
    .X(_0299_));
 sky130_fd_sc_hd__a221o_2 _0617_ (.A1(net9),
    .A2(net425),
    .B1(net421),
    .B2(net44),
    .C1(_0299_),
    .X(_0300_));
 sky130_fd_sc_hd__a211o_2 _0618_ (.A1(net71),
    .A2(net430),
    .B1(net414),
    .C1(_0300_),
    .X(net346));
 sky130_fd_sc_hd__a31o_2 _0619_ (.A1(net450),
    .A2(net453),
    .A3(net99),
    .B1(_0222_),
    .X(_0301_));
 sky130_fd_sc_hd__a221o_1 _0620_ (.A1(net127),
    .A2(net437),
    .B1(net424),
    .B2(net45),
    .C1(_0301_),
    .X(_0302_));
 sky130_fd_sc_hd__a221o_1 _0621_ (.A1(net72),
    .A2(net430),
    .B1(net428),
    .B2(net10),
    .C1(_0270_),
    .X(_0303_));
 sky130_fd_sc_hd__or2_4 _0622_ (.A(_0302_),
    .B(_0303_),
    .X(net347));
 sky130_fd_sc_hd__a22o_4 _0623_ (.A1(net128),
    .A2(net439),
    .B1(net419),
    .B2(net100),
    .X(_0304_));
 sky130_fd_sc_hd__a221o_2 _0624_ (.A1(net11),
    .A2(net425),
    .B1(net421),
    .B2(net46),
    .C1(_0304_),
    .X(_0305_));
 sky130_fd_sc_hd__a211o_2 _0625_ (.A1(net73),
    .A2(net430),
    .B1(net414),
    .C1(_0305_),
    .X(net349));
 sky130_fd_sc_hd__a22o_2 _0626_ (.A1(net130),
    .A2(net438),
    .B1(net419),
    .B2(net102),
    .X(_0306_));
 sky130_fd_sc_hd__a221o_2 _0627_ (.A1(net13),
    .A2(net426),
    .B1(net424),
    .B2(net48),
    .C1(_0270_),
    .X(_0307_));
 sky130_fd_sc_hd__a211o_4 _0628_ (.A1(net75),
    .A2(net429),
    .B1(_0306_),
    .C1(_0307_),
    .X(net350));
 sky130_fd_sc_hd__a22o_4 _0629_ (.A1(net131),
    .A2(net439),
    .B1(net419),
    .B2(net103),
    .X(_0308_));
 sky130_fd_sc_hd__a221o_4 _0630_ (.A1(net14),
    .A2(net425),
    .B1(net421),
    .B2(net49),
    .C1(_0308_),
    .X(_0309_));
 sky130_fd_sc_hd__a211o_4 _0631_ (.A1(net76),
    .A2(net430),
    .B1(net414),
    .C1(_0309_),
    .X(net351));
 sky130_fd_sc_hd__a31o_2 _0632_ (.A1(net449),
    .A2(net452),
    .A3(net104),
    .B1(_0222_),
    .X(_0310_));
 sky130_fd_sc_hd__a221o_1 _0633_ (.A1(net132),
    .A2(net437),
    .B1(net424),
    .B2(net50),
    .C1(_0310_),
    .X(_0311_));
 sky130_fd_sc_hd__a221o_1 _0634_ (.A1(net77),
    .A2(net430),
    .B1(net428),
    .B2(net15),
    .C1(_0270_),
    .X(_0312_));
 sky130_fd_sc_hd__or2_4 _0635_ (.A(_0311_),
    .B(_0312_),
    .X(net352));
 sky130_fd_sc_hd__a22o_4 _0636_ (.A1(net133),
    .A2(net439),
    .B1(net419),
    .B2(net105),
    .X(_0313_));
 sky130_fd_sc_hd__a221o_4 _0637_ (.A1(net16),
    .A2(net425),
    .B1(net421),
    .B2(net51),
    .C1(_0313_),
    .X(_0314_));
 sky130_fd_sc_hd__a211o_2 _0638_ (.A1(net78),
    .A2(net430),
    .B1(net414),
    .C1(_0314_),
    .X(net353));
 sky130_fd_sc_hd__a221o_4 _0639_ (.A1(net79),
    .A2(net431),
    .B1(net419),
    .B2(net106),
    .C1(_0270_),
    .X(_0315_));
 sky130_fd_sc_hd__a22o_2 _0640_ (.A1(net17),
    .A2(net425),
    .B1(net421),
    .B2(net52),
    .X(_0316_));
 sky130_fd_sc_hd__a211o_4 _0641_ (.A1(net134),
    .A2(net437),
    .B1(_0315_),
    .C1(_0316_),
    .X(net354));
 sky130_fd_sc_hd__a221o_4 _0642_ (.A1(net80),
    .A2(_0196_),
    .B1(net419),
    .B2(net107),
    .C1(_0270_),
    .X(_0317_));
 sky130_fd_sc_hd__a22o_1 _0643_ (.A1(net135),
    .A2(net437),
    .B1(net426),
    .B2(net18),
    .X(_0318_));
 sky130_fd_sc_hd__a211o_4 _0644_ (.A1(net53),
    .A2(net422),
    .B1(_0317_),
    .C1(_0318_),
    .X(net355));
 sky130_fd_sc_hd__a22o_4 _0645_ (.A1(net136),
    .A2(net438),
    .B1(net419),
    .B2(net108),
    .X(_0319_));
 sky130_fd_sc_hd__a221o_4 _0646_ (.A1(net19),
    .A2(net425),
    .B1(net421),
    .B2(net54),
    .C1(_0319_),
    .X(_0320_));
 sky130_fd_sc_hd__a211o_2 _0647_ (.A1(net81),
    .A2(net430),
    .B1(net414),
    .C1(_0320_),
    .X(net356));
 sky130_fd_sc_hd__a211o_4 _0648_ (.A1(net109),
    .A2(net420),
    .B1(net414),
    .C1(_0197_),
    .X(net327));
 sky130_fd_sc_hd__mux2_2 _0649_ (.A0(clknet_3_0__leaf_wb_clk_i),
    .A1(wb_clk_override),
    .S(wb_single_step),
    .X(_0321_));
 sky130_fd_sc_hd__mux2_2 _0650_ (.A0(net196),
    .A1(_0321_),
    .S(net446),
    .X(net270));
 sky130_fd_sc_hd__and2b_1 _0651_ (.A_N(net442),
    .B(net197),
    .X(_0322_));
 sky130_fd_sc_hd__a31o_2 _0652_ (.A1(net448),
    .A2(\wb_io_override[0] ),
    .A3(net300),
    .B1(_0322_),
    .X(net271));
 sky130_fd_sc_hd__and2b_1 _0653_ (.A_N(net441),
    .B(net198),
    .X(_0323_));
 sky130_fd_sc_hd__a31o_1 _0654_ (.A1(net441),
    .A2(\wb_io_override[1] ),
    .A3(net302),
    .B1(_0323_),
    .X(net282));
 sky130_fd_sc_hd__and2b_1 _0655_ (.A_N(net441),
    .B(net199),
    .X(_0324_));
 sky130_fd_sc_hd__a31o_1 _0656_ (.A1(net441),
    .A2(\wb_io_override[2] ),
    .A3(net302),
    .B1(_0324_),
    .X(net291));
 sky130_fd_sc_hd__and2b_1 _0657_ (.A_N(net443),
    .B(net200),
    .X(_0325_));
 sky130_fd_sc_hd__a31o_1 _0658_ (.A1(net445),
    .A2(\wb_io_override[3] ),
    .A3(net303),
    .B1(_0325_),
    .X(net292));
 sky130_fd_sc_hd__and2b_1 _0659_ (.A_N(net441),
    .B(net201),
    .X(_0326_));
 sky130_fd_sc_hd__a31o_1 _0660_ (.A1(net441),
    .A2(\wb_io_override[4] ),
    .A3(net304),
    .B1(_0326_),
    .X(net293));
 sky130_fd_sc_hd__and2b_1 _0661_ (.A_N(net441),
    .B(net202),
    .X(_0327_));
 sky130_fd_sc_hd__a31o_1 _0662_ (.A1(net441),
    .A2(\wb_io_override[5] ),
    .A3(net305),
    .B1(_0327_),
    .X(net294));
 sky130_fd_sc_hd__and2b_1 _0663_ (.A_N(net441),
    .B(net203),
    .X(_0328_));
 sky130_fd_sc_hd__a31o_1 _0664_ (.A1(net441),
    .A2(\wb_io_override[6] ),
    .A3(net307),
    .B1(_0328_),
    .X(net295));
 sky130_fd_sc_hd__and2b_1 _0665_ (.A_N(net442),
    .B(net204),
    .X(_0329_));
 sky130_fd_sc_hd__a31o_1 _0666_ (.A1(net442),
    .A2(\wb_io_override[7] ),
    .A3(net307),
    .B1(_0329_),
    .X(net296));
 sky130_fd_sc_hd__and2b_1 _0667_ (.A_N(net442),
    .B(net205),
    .X(_0330_));
 sky130_fd_sc_hd__a31o_1 _0668_ (.A1(net443),
    .A2(\wb_io_override[8] ),
    .A3(net309),
    .B1(_0330_),
    .X(net297));
 sky130_fd_sc_hd__and2b_1 _0669_ (.A_N(net444),
    .B(net206),
    .X(_0331_));
 sky130_fd_sc_hd__a31o_1 _0670_ (.A1(net444),
    .A2(\wb_io_override[9] ),
    .A3(net309),
    .B1(_0331_),
    .X(net298));
 sky130_fd_sc_hd__and2b_1 _0671_ (.A_N(net443),
    .B(net207),
    .X(_0332_));
 sky130_fd_sc_hd__a31o_1 _0672_ (.A1(net444),
    .A2(\wb_io_override[10] ),
    .A3(net311),
    .B1(_0332_),
    .X(net272));
 sky130_fd_sc_hd__and2b_1 _0673_ (.A_N(net444),
    .B(net208),
    .X(_0333_));
 sky130_fd_sc_hd__a31o_1 _0674_ (.A1(net444),
    .A2(\wb_io_override[11] ),
    .A3(net311),
    .B1(_0333_),
    .X(net273));
 sky130_fd_sc_hd__and2b_1 _0675_ (.A_N(net444),
    .B(net209),
    .X(_0334_));
 sky130_fd_sc_hd__a31o_2 _0676_ (.A1(net448),
    .A2(\wb_io_override[12] ),
    .A3(net312),
    .B1(_0334_),
    .X(net274));
 sky130_fd_sc_hd__and2b_1 _0677_ (.A_N(net444),
    .B(net210),
    .X(_0335_));
 sky130_fd_sc_hd__a31o_1 _0678_ (.A1(net445),
    .A2(\wb_io_override[13] ),
    .A3(net313),
    .B1(_0335_),
    .X(net275));
 sky130_fd_sc_hd__and2b_1 _0679_ (.A_N(net444),
    .B(net211),
    .X(_0336_));
 sky130_fd_sc_hd__a31o_1 _0680_ (.A1(net446),
    .A2(\wb_io_override[14] ),
    .A3(net315),
    .B1(_0336_),
    .X(net276));
 sky130_fd_sc_hd__and2b_1 _0681_ (.A_N(wb_override),
    .B(net212),
    .X(_0337_));
 sky130_fd_sc_hd__a31o_1 _0682_ (.A1(net446),
    .A2(\wb_io_override[15] ),
    .A3(net315),
    .B1(_0337_),
    .X(net277));
 sky130_fd_sc_hd__and2b_1 _0683_ (.A_N(net445),
    .B(net213),
    .X(_0338_));
 sky130_fd_sc_hd__a31o_2 _0684_ (.A1(net447),
    .A2(\wb_io_override[16] ),
    .A3(net415),
    .B1(_0338_),
    .X(net278));
 sky130_fd_sc_hd__and2b_1 _0685_ (.A_N(net443),
    .B(net214),
    .X(_0339_));
 sky130_fd_sc_hd__a31o_2 _0686_ (.A1(net447),
    .A2(\wb_io_override[17] ),
    .A3(net415),
    .B1(_0339_),
    .X(net279));
 sky130_fd_sc_hd__and2b_1 _0687_ (.A_N(net443),
    .B(net215),
    .X(_0340_));
 sky130_fd_sc_hd__a31o_2 _0688_ (.A1(net447),
    .A2(\wb_io_override[18] ),
    .A3(net415),
    .B1(_0340_),
    .X(net280));
 sky130_fd_sc_hd__and2b_1 _0689_ (.A_N(net443),
    .B(net216),
    .X(_0341_));
 sky130_fd_sc_hd__a31o_2 _0690_ (.A1(net447),
    .A2(\wb_io_override[19] ),
    .A3(net415),
    .B1(_0341_),
    .X(net281));
 sky130_fd_sc_hd__and2b_1 _0691_ (.A_N(net443),
    .B(net217),
    .X(_0342_));
 sky130_fd_sc_hd__a31o_2 _0692_ (.A1(net447),
    .A2(\wb_io_override[20] ),
    .A3(net415),
    .B1(_0342_),
    .X(net283));
 sky130_fd_sc_hd__and2b_1 _0693_ (.A_N(net446),
    .B(net218),
    .X(_0343_));
 sky130_fd_sc_hd__a31o_1 _0694_ (.A1(net446),
    .A2(\wb_io_override[21] ),
    .A3(net326),
    .B1(_0343_),
    .X(net284));
 sky130_fd_sc_hd__and2b_1 _0695_ (.A_N(net445),
    .B(net219),
    .X(_0344_));
 sky130_fd_sc_hd__a31o_2 _0696_ (.A1(net447),
    .A2(\wb_io_override[22] ),
    .A3(net415),
    .B1(_0344_),
    .X(net285));
 sky130_fd_sc_hd__and2b_1 _0697_ (.A_N(net443),
    .B(net220),
    .X(_0345_));
 sky130_fd_sc_hd__a31o_1 _0698_ (.A1(net446),
    .A2(\wb_io_override[23] ),
    .A3(net326),
    .B1(_0345_),
    .X(net286));
 sky130_fd_sc_hd__and2b_1 _0699_ (.A_N(net447),
    .B(net221),
    .X(_0346_));
 sky130_fd_sc_hd__a31o_2 _0700_ (.A1(net447),
    .A2(\wb_io_override[24] ),
    .A3(net415),
    .B1(_0346_),
    .X(net287));
 sky130_fd_sc_hd__and2b_1 _0701_ (.A_N(net447),
    .B(net222),
    .X(_0347_));
 sky130_fd_sc_hd__a31o_2 _0702_ (.A1(net447),
    .A2(\wb_io_override[25] ),
    .A3(net415),
    .B1(_0347_),
    .X(net288));
 sky130_fd_sc_hd__and2b_1 _0703_ (.A_N(net445),
    .B(net223),
    .X(_0348_));
 sky130_fd_sc_hd__a31o_1 _0704_ (.A1(net446),
    .A2(\wb_io_override[26] ),
    .A3(net326),
    .B1(_0348_),
    .X(net289));
 sky130_fd_sc_hd__and2b_1 _0705_ (.A_N(net446),
    .B(net195),
    .X(_0349_));
 sky130_fd_sc_hd__a31o_1 _0706_ (.A1(net446),
    .A2(\wb_io_override[27] ),
    .A3(net299),
    .B1(_0349_),
    .X(net290));
 sky130_fd_sc_hd__and2_2 _0707_ (.A(net268),
    .B(net239),
    .X(_0350_));
 sky130_fd_sc_hd__nand2_2 _0708_ (.A(net268),
    .B(net239),
    .Y(_0351_));
 sky130_fd_sc_hd__and3_4 _0709_ (.A(net470),
    .B(net269),
    .C(_0350_),
    .X(_0352_));
 sky130_fd_sc_hd__mux2_1 _0710_ (.A0(\wb_design_addr_override[0] ),
    .A1(net262),
    .S(_0352_),
    .X(_0353_));
 sky130_fd_sc_hd__and2_1 _0711_ (.A(net461),
    .B(_0353_),
    .X(_0000_));
 sky130_fd_sc_hd__mux2_1 _0712_ (.A0(\wb_design_addr_override[1] ),
    .A1(net263),
    .S(_0352_),
    .X(_0354_));
 sky130_fd_sc_hd__and2_1 _0713_ (.A(net461),
    .B(_0354_),
    .X(_0001_));
 sky130_fd_sc_hd__mux2_1 _0714_ (.A0(\wb_design_addr_override[2] ),
    .A1(net264),
    .S(_0352_),
    .X(_0355_));
 sky130_fd_sc_hd__and2_1 _0715_ (.A(net462),
    .B(_0355_),
    .X(_0002_));
 sky130_fd_sc_hd__mux2_1 _0716_ (.A0(\wb_design_addr_override[3] ),
    .A1(net265),
    .S(_0352_),
    .X(_0356_));
 sky130_fd_sc_hd__and2_1 _0717_ (.A(net461),
    .B(_0356_),
    .X(_0003_));
 sky130_fd_sc_hd__nor2_1 _0718_ (.A(net474),
    .B(_0351_),
    .Y(_0005_));
 sky130_fd_sc_hd__and2_1 _0719_ (.A(net462),
    .B(_0352_),
    .X(_0357_));
 sky130_fd_sc_hd__mux2_1 _0720_ (.A0(wb_single_step),
    .A1(net260),
    .S(_0357_),
    .X(_0004_));
 sky130_fd_sc_hd__nand2_1 _0721_ (.A(_0179_),
    .B(net269),
    .Y(_0358_));
 sky130_fd_sc_hd__nor2_1 _0722_ (.A(net471),
    .B(_0358_),
    .Y(_0359_));
 sky130_fd_sc_hd__and3_1 _0723_ (.A(net236),
    .B(_0350_),
    .C(_0359_),
    .X(_0360_));
 sky130_fd_sc_hd__or4b_4 _0724_ (.A(net471),
    .B(_0351_),
    .C(_0358_),
    .D_N(net236),
    .X(_0361_));
 sky130_fd_sc_hd__or2_1 _0725_ (.A(\wb_counter[0] ),
    .B(net402),
    .X(_0362_));
 sky130_fd_sc_hd__o211a_1 _0726_ (.A1(net240),
    .A2(net413),
    .B1(_0362_),
    .C1(net461),
    .X(_0006_));
 sky130_fd_sc_hd__or2_1 _0727_ (.A(net337),
    .B(net402),
    .X(_0363_));
 sky130_fd_sc_hd__o211a_1 _0728_ (.A1(net251),
    .A2(net413),
    .B1(_0363_),
    .C1(net461),
    .X(_0007_));
 sky130_fd_sc_hd__or2_1 _0729_ (.A(net348),
    .B(net402),
    .X(_0364_));
 sky130_fd_sc_hd__o211a_1 _0730_ (.A1(net260),
    .A2(net413),
    .B1(_0364_),
    .C1(net461),
    .X(_0008_));
 sky130_fd_sc_hd__or2_1 _0731_ (.A(net357),
    .B(net402),
    .X(_0365_));
 sky130_fd_sc_hd__o211a_1 _0732_ (.A1(net261),
    .A2(net413),
    .B1(_0365_),
    .C1(net461),
    .X(_0009_));
 sky130_fd_sc_hd__nand2_1 _0733_ (.A(_0176_),
    .B(net413),
    .Y(_0366_));
 sky130_fd_sc_hd__o211a_1 _0734_ (.A1(net262),
    .A2(net413),
    .B1(_0366_),
    .C1(net462),
    .X(_0010_));
 sky130_fd_sc_hd__or2_1 _0735_ (.A(\wb_counter[5] ),
    .B(net402),
    .X(_0367_));
 sky130_fd_sc_hd__o211a_1 _0736_ (.A1(net263),
    .A2(net413),
    .B1(_0367_),
    .C1(net461),
    .X(_0011_));
 sky130_fd_sc_hd__or2_1 _0737_ (.A(\wb_counter[6] ),
    .B(net402),
    .X(_0368_));
 sky130_fd_sc_hd__o211a_1 _0738_ (.A1(net264),
    .A2(net413),
    .B1(_0368_),
    .C1(net464),
    .X(_0012_));
 sky130_fd_sc_hd__or2_1 _0739_ (.A(\wb_counter[7] ),
    .B(net401),
    .X(_0369_));
 sky130_fd_sc_hd__o211a_1 _0740_ (.A1(net265),
    .A2(net411),
    .B1(_0369_),
    .C1(net464),
    .X(_0013_));
 sky130_fd_sc_hd__nand2_1 _0741_ (.A(_0175_),
    .B(net413),
    .Y(_0370_));
 sky130_fd_sc_hd__o211a_1 _0742_ (.A1(net266),
    .A2(net413),
    .B1(_0370_),
    .C1(net467),
    .X(_0014_));
 sky130_fd_sc_hd__nand2_1 _0743_ (.A(_0174_),
    .B(net411),
    .Y(_0371_));
 sky130_fd_sc_hd__o211a_1 _0744_ (.A1(net267),
    .A2(net411),
    .B1(_0371_),
    .C1(net467),
    .X(_0015_));
 sky130_fd_sc_hd__or2_1 _0745_ (.A(\wb_counter[10] ),
    .B(net401),
    .X(_0372_));
 sky130_fd_sc_hd__o211a_1 _0746_ (.A1(net241),
    .A2(net411),
    .B1(_0372_),
    .C1(net464),
    .X(_0016_));
 sky130_fd_sc_hd__or2_1 _0747_ (.A(\wb_counter[11] ),
    .B(net401),
    .X(_0373_));
 sky130_fd_sc_hd__o211a_1 _0748_ (.A1(net242),
    .A2(net412),
    .B1(_0373_),
    .C1(net463),
    .X(_0017_));
 sky130_fd_sc_hd__or2_1 _0749_ (.A(\wb_counter[12] ),
    .B(net402),
    .X(_0374_));
 sky130_fd_sc_hd__o211a_1 _0750_ (.A1(net243),
    .A2(net412),
    .B1(_0374_),
    .C1(net463),
    .X(_0018_));
 sky130_fd_sc_hd__or2_1 _0751_ (.A(\wb_counter[13] ),
    .B(net402),
    .X(_0375_));
 sky130_fd_sc_hd__o211a_1 _0752_ (.A1(net244),
    .A2(net412),
    .B1(_0375_),
    .C1(net463),
    .X(_0019_));
 sky130_fd_sc_hd__nand2_1 _0753_ (.A(_0173_),
    .B(net411),
    .Y(_0376_));
 sky130_fd_sc_hd__o211a_1 _0754_ (.A1(net245),
    .A2(net411),
    .B1(_0376_),
    .C1(net463),
    .X(_0020_));
 sky130_fd_sc_hd__or2_1 _0755_ (.A(\wb_counter[15] ),
    .B(net401),
    .X(_0377_));
 sky130_fd_sc_hd__o211a_1 _0756_ (.A1(net246),
    .A2(net411),
    .B1(_0377_),
    .C1(net463),
    .X(_0021_));
 sky130_fd_sc_hd__or2_1 _0757_ (.A(\wb_counter[16] ),
    .B(net401),
    .X(_0378_));
 sky130_fd_sc_hd__o211a_1 _0758_ (.A1(net247),
    .A2(net412),
    .B1(_0378_),
    .C1(net463),
    .X(_0022_));
 sky130_fd_sc_hd__or2_1 _0759_ (.A(\wb_counter[17] ),
    .B(net402),
    .X(_0379_));
 sky130_fd_sc_hd__o211a_1 _0760_ (.A1(net248),
    .A2(net412),
    .B1(_0379_),
    .C1(net463),
    .X(_0023_));
 sky130_fd_sc_hd__or2_1 _0761_ (.A(\wb_counter[18] ),
    .B(net401),
    .X(_0380_));
 sky130_fd_sc_hd__o211a_1 _0762_ (.A1(net249),
    .A2(net412),
    .B1(_0380_),
    .C1(net464),
    .X(_0024_));
 sky130_fd_sc_hd__or2_1 _0763_ (.A(\wb_counter[19] ),
    .B(net401),
    .X(_0381_));
 sky130_fd_sc_hd__o211a_1 _0764_ (.A1(net250),
    .A2(net412),
    .B1(_0381_),
    .C1(net465),
    .X(_0025_));
 sky130_fd_sc_hd__or2_1 _0765_ (.A(\wb_counter[20] ),
    .B(net401),
    .X(_0382_));
 sky130_fd_sc_hd__o211a_1 _0766_ (.A1(net252),
    .A2(net411),
    .B1(_0382_),
    .C1(net463),
    .X(_0026_));
 sky130_fd_sc_hd__or2_1 _0767_ (.A(\wb_counter[21] ),
    .B(net401),
    .X(_0383_));
 sky130_fd_sc_hd__o211a_1 _0768_ (.A1(net253),
    .A2(net412),
    .B1(_0383_),
    .C1(net465),
    .X(_0027_));
 sky130_fd_sc_hd__or2_1 _0769_ (.A(\wb_counter[22] ),
    .B(net401),
    .X(_0384_));
 sky130_fd_sc_hd__o211a_1 _0770_ (.A1(net254),
    .A2(net412),
    .B1(_0384_),
    .C1(net463),
    .X(_0028_));
 sky130_fd_sc_hd__nand2_1 _0771_ (.A(_0172_),
    .B(net411),
    .Y(_0385_));
 sky130_fd_sc_hd__o211a_1 _0772_ (.A1(net255),
    .A2(net411),
    .B1(_0385_),
    .C1(net463),
    .X(_0029_));
 sky130_fd_sc_hd__and2_1 _0773_ (.A(net466),
    .B(wb_feedback_delay),
    .X(_0030_));
 sky130_fd_sc_hd__or4_1 _0774_ (.A(net469),
    .B(net476),
    .C(_0351_),
    .D(_0358_),
    .X(_0386_));
 sky130_fd_sc_hd__mux2_1 _0775_ (.A0(net240),
    .A1(\wb_io_override[0] ),
    .S(net409),
    .X(_0031_));
 sky130_fd_sc_hd__mux2_1 _0776_ (.A0(net251),
    .A1(\wb_io_override[1] ),
    .S(net407),
    .X(_0032_));
 sky130_fd_sc_hd__mux2_1 _0777_ (.A0(net260),
    .A1(\wb_io_override[2] ),
    .S(net407),
    .X(_0033_));
 sky130_fd_sc_hd__mux2_1 _0778_ (.A0(net261),
    .A1(\wb_io_override[3] ),
    .S(net407),
    .X(_0034_));
 sky130_fd_sc_hd__mux2_1 _0779_ (.A0(net262),
    .A1(\wb_io_override[4] ),
    .S(net407),
    .X(_0035_));
 sky130_fd_sc_hd__mux2_1 _0780_ (.A0(net263),
    .A1(\wb_io_override[5] ),
    .S(net407),
    .X(_0036_));
 sky130_fd_sc_hd__mux2_1 _0781_ (.A0(net264),
    .A1(\wb_io_override[6] ),
    .S(net407),
    .X(_0037_));
 sky130_fd_sc_hd__mux2_1 _0782_ (.A0(net265),
    .A1(\wb_io_override[7] ),
    .S(net408),
    .X(_0038_));
 sky130_fd_sc_hd__mux2_1 _0783_ (.A0(net266),
    .A1(\wb_io_override[8] ),
    .S(net407),
    .X(_0039_));
 sky130_fd_sc_hd__mux2_1 _0784_ (.A0(net267),
    .A1(\wb_io_override[9] ),
    .S(net407),
    .X(_0040_));
 sky130_fd_sc_hd__mux2_1 _0785_ (.A0(net241),
    .A1(\wb_io_override[10] ),
    .S(net407),
    .X(_0041_));
 sky130_fd_sc_hd__mux2_1 _0786_ (.A0(net242),
    .A1(\wb_io_override[11] ),
    .S(net408),
    .X(_0042_));
 sky130_fd_sc_hd__mux2_1 _0787_ (.A0(net243),
    .A1(\wb_io_override[12] ),
    .S(net410),
    .X(_0043_));
 sky130_fd_sc_hd__mux2_1 _0788_ (.A0(net244),
    .A1(\wb_io_override[13] ),
    .S(net410),
    .X(_0044_));
 sky130_fd_sc_hd__mux2_1 _0789_ (.A0(net245),
    .A1(\wb_io_override[14] ),
    .S(net408),
    .X(_0045_));
 sky130_fd_sc_hd__mux2_1 _0790_ (.A0(net246),
    .A1(\wb_io_override[15] ),
    .S(net409),
    .X(_0046_));
 sky130_fd_sc_hd__mux2_1 _0791_ (.A0(net247),
    .A1(\wb_io_override[16] ),
    .S(net408),
    .X(_0047_));
 sky130_fd_sc_hd__mux2_1 _0792_ (.A0(net248),
    .A1(\wb_io_override[17] ),
    .S(net409),
    .X(_0048_));
 sky130_fd_sc_hd__mux2_1 _0793_ (.A0(net249),
    .A1(\wb_io_override[18] ),
    .S(net410),
    .X(_0049_));
 sky130_fd_sc_hd__mux2_1 _0794_ (.A0(net250),
    .A1(\wb_io_override[19] ),
    .S(net409),
    .X(_0050_));
 sky130_fd_sc_hd__mux2_1 _0795_ (.A0(net252),
    .A1(\wb_io_override[20] ),
    .S(net407),
    .X(_0051_));
 sky130_fd_sc_hd__mux2_1 _0796_ (.A0(net253),
    .A1(\wb_io_override[21] ),
    .S(net410),
    .X(_0052_));
 sky130_fd_sc_hd__mux2_1 _0797_ (.A0(net254),
    .A1(\wb_io_override[22] ),
    .S(net409),
    .X(_0053_));
 sky130_fd_sc_hd__mux2_1 _0798_ (.A0(net255),
    .A1(\wb_io_override[23] ),
    .S(net410),
    .X(_0054_));
 sky130_fd_sc_hd__mux2_1 _0799_ (.A0(net256),
    .A1(\wb_io_override[24] ),
    .S(net410),
    .X(_0055_));
 sky130_fd_sc_hd__mux2_1 _0800_ (.A0(net257),
    .A1(\wb_io_override[25] ),
    .S(net410),
    .X(_0056_));
 sky130_fd_sc_hd__mux2_1 _0801_ (.A0(net258),
    .A1(\wb_io_override[26] ),
    .S(net410),
    .X(_0057_));
 sky130_fd_sc_hd__mux2_1 _0802_ (.A0(net259),
    .A1(\wb_io_override[27] ),
    .S(net410),
    .X(_0058_));
 sky130_fd_sc_hd__mux2_1 _0803_ (.A0(net224),
    .A1(\wb_design_addr_override[0] ),
    .S(net445),
    .X(_0387_));
 sky130_fd_sc_hd__mux2_1 _0804_ (.A0(net460),
    .A1(_0387_),
    .S(net462),
    .X(_0059_));
 sky130_fd_sc_hd__mux2_1 _0805_ (.A0(net225),
    .A1(\wb_design_addr_override[1] ),
    .S(net445),
    .X(_0388_));
 sky130_fd_sc_hd__mux2_1 _0806_ (.A0(net457),
    .A1(_0388_),
    .S(net462),
    .X(_0060_));
 sky130_fd_sc_hd__mux2_1 _0807_ (.A0(net226),
    .A1(\wb_design_addr_override[2] ),
    .S(net445),
    .X(_0389_));
 sky130_fd_sc_hd__mux2_1 _0808_ (.A0(net454),
    .A1(_0389_),
    .S(net462),
    .X(_0061_));
 sky130_fd_sc_hd__mux2_1 _0809_ (.A0(net227),
    .A1(\wb_design_addr_override[3] ),
    .S(net445),
    .X(_0390_));
 sky130_fd_sc_hd__mux2_1 _0810_ (.A0(net451),
    .A1(_0390_),
    .S(net462),
    .X(_0062_));
 sky130_fd_sc_hd__a211o_1 _0811_ (.A1(_0180_),
    .A2(net236),
    .B1(net472),
    .C1(net470),
    .X(_0391_));
 sky130_fd_sc_hd__nand2_2 _0812_ (.A(_0350_),
    .B(_0391_),
    .Y(_0392_));
 sky130_fd_sc_hd__nand2_1 _0813_ (.A(net372),
    .B(net406),
    .Y(_0393_));
 sky130_fd_sc_hd__nor2_1 _0814_ (.A(net469),
    .B(net303),
    .Y(_0394_));
 sky130_fd_sc_hd__a21o_1 _0815_ (.A1(\wb_counter[0] ),
    .A2(net469),
    .B1(net470),
    .X(_0395_));
 sky130_fd_sc_hd__a31o_1 _0816_ (.A1(net471),
    .A2(_0207_),
    .A3(net328),
    .B1(_0395_),
    .X(_0396_));
 sky130_fd_sc_hd__nor2_1 _0817_ (.A(net448),
    .B(_0179_),
    .Y(_0397_));
 sky130_fd_sc_hd__or3b_4 _0818_ (.A(_0397_),
    .B(net404),
    .C_N(_0396_),
    .X(_0398_));
 sky130_fd_sc_hd__a21oi_1 _0819_ (.A1(_0393_),
    .A2(_0398_),
    .B1(net474),
    .Y(_0063_));
 sky130_fd_sc_hd__nand2_1 _0820_ (.A(net383),
    .B(net406),
    .Y(_0399_));
 sky130_fd_sc_hd__a21o_1 _0821_ (.A1(net337),
    .A2(net469),
    .B1(net470),
    .X(_0400_));
 sky130_fd_sc_hd__a31o_1 _0822_ (.A1(net471),
    .A2(_0207_),
    .A3(net329),
    .B1(_0400_),
    .X(_0401_));
 sky130_fd_sc_hd__nor2_1 _0823_ (.A(wb_rst_override),
    .B(_0179_),
    .Y(_0402_));
 sky130_fd_sc_hd__or3b_4 _0824_ (.A(_0402_),
    .B(net404),
    .C_N(_0401_),
    .X(_0403_));
 sky130_fd_sc_hd__a21oi_1 _0825_ (.A1(_0399_),
    .A2(_0403_),
    .B1(net474),
    .Y(_0064_));
 sky130_fd_sc_hd__nand2_1 _0826_ (.A(net392),
    .B(net406),
    .Y(_0404_));
 sky130_fd_sc_hd__a21o_1 _0827_ (.A1(net348),
    .A2(net469),
    .B1(net470),
    .X(_0405_));
 sky130_fd_sc_hd__a31o_1 _0828_ (.A1(net471),
    .A2(_0207_),
    .A3(net330),
    .B1(_0405_),
    .X(_0406_));
 sky130_fd_sc_hd__nor2_1 _0829_ (.A(\wb_design_addr_override[0] ),
    .B(_0179_),
    .Y(_0407_));
 sky130_fd_sc_hd__or3b_4 _0830_ (.A(_0407_),
    .B(net404),
    .C_N(_0406_),
    .X(_0408_));
 sky130_fd_sc_hd__a21oi_1 _0831_ (.A1(_0404_),
    .A2(_0408_),
    .B1(net474),
    .Y(_0065_));
 sky130_fd_sc_hd__a221o_1 _0832_ (.A1(net357),
    .A2(net469),
    .B1(net331),
    .B2(_0394_),
    .C1(net470),
    .X(_0409_));
 sky130_fd_sc_hd__o211a_1 _0833_ (.A1(\wb_design_addr_override[1] ),
    .A2(_0179_),
    .B1(_0350_),
    .C1(_0391_),
    .X(_0410_));
 sky130_fd_sc_hd__a22o_1 _0834_ (.A1(net393),
    .A2(net404),
    .B1(_0409_),
    .B2(_0410_),
    .X(_0411_));
 sky130_fd_sc_hd__and2_1 _0835_ (.A(net466),
    .B(_0411_),
    .X(_0066_));
 sky130_fd_sc_hd__nand2_1 _0836_ (.A(net394),
    .B(net406),
    .Y(_0412_));
 sky130_fd_sc_hd__o31ai_4 _0837_ (.A1(_0235_),
    .A2(_0236_),
    .A3(_0238_),
    .B1(net472),
    .Y(_0413_));
 sky130_fd_sc_hd__o221a_1 _0838_ (.A1(_0176_),
    .A2(net471),
    .B1(net304),
    .B2(_0413_),
    .C1(_0179_),
    .X(_0414_));
 sky130_fd_sc_hd__a211o_2 _0839_ (.A1(_0178_),
    .A2(net470),
    .B1(net404),
    .C1(_0414_),
    .X(_0415_));
 sky130_fd_sc_hd__a21oi_1 _0840_ (.A1(_0412_),
    .A2(_0415_),
    .B1(net474),
    .Y(_0067_));
 sky130_fd_sc_hd__nand2_1 _0841_ (.A(net395),
    .B(net406),
    .Y(_0416_));
 sky130_fd_sc_hd__nor2_2 _0842_ (.A(net469),
    .B(net307),
    .Y(_0417_));
 sky130_fd_sc_hd__a221oi_2 _0843_ (.A1(\wb_counter[5] ),
    .A2(net469),
    .B1(net333),
    .B2(_0417_),
    .C1(net470),
    .Y(_0418_));
 sky130_fd_sc_hd__a211o_2 _0844_ (.A1(_0177_),
    .A2(net470),
    .B1(net404),
    .C1(_0418_),
    .X(_0419_));
 sky130_fd_sc_hd__a21oi_1 _0845_ (.A1(_0416_),
    .A2(_0419_),
    .B1(net474),
    .Y(_0068_));
 sky130_fd_sc_hd__a22oi_2 _0846_ (.A1(\wb_counter[6] ),
    .A2(net468),
    .B1(net334),
    .B2(_0417_),
    .Y(_0420_));
 sky130_fd_sc_hd__nor2_4 _0847_ (.A(net238),
    .B(net403),
    .Y(_0421_));
 sky130_fd_sc_hd__or2_4 _0848_ (.A(net238),
    .B(net403),
    .X(_0422_));
 sky130_fd_sc_hd__a2bb2o_1 _0849_ (.A1_N(_0420_),
    .A2_N(_0422_),
    .B1(net396),
    .B2(net403),
    .X(_0423_));
 sky130_fd_sc_hd__and2_1 _0850_ (.A(net465),
    .B(_0423_),
    .X(_0069_));
 sky130_fd_sc_hd__a22o_2 _0851_ (.A1(\wb_counter[7] ),
    .A2(net468),
    .B1(net335),
    .B2(_0417_),
    .X(_0424_));
 sky130_fd_sc_hd__a22o_1 _0852_ (.A1(net397),
    .A2(net405),
    .B1(net400),
    .B2(_0424_),
    .X(_0425_));
 sky130_fd_sc_hd__and2_1 _0853_ (.A(net465),
    .B(_0425_),
    .X(_0070_));
 sky130_fd_sc_hd__or2_1 _0854_ (.A(net468),
    .B(net309),
    .X(_0426_));
 sky130_fd_sc_hd__o22a_1 _0855_ (.A1(_0175_),
    .A2(net471),
    .B1(_0262_),
    .B2(_0426_),
    .X(_0427_));
 sky130_fd_sc_hd__o2bb2a_1 _0856_ (.A1_N(net398),
    .A2_N(net403),
    .B1(_0422_),
    .B2(_0427_),
    .X(_0428_));
 sky130_fd_sc_hd__nor2_1 _0857_ (.A(net474),
    .B(_0428_),
    .Y(_0071_));
 sky130_fd_sc_hd__o22a_1 _0858_ (.A1(_0174_),
    .A2(net471),
    .B1(_0268_),
    .B2(_0426_),
    .X(_0429_));
 sky130_fd_sc_hd__o2bb2a_1 _0859_ (.A1_N(net399),
    .A2_N(net403),
    .B1(_0422_),
    .B2(_0429_),
    .X(_0430_));
 sky130_fd_sc_hd__nor2_1 _0860_ (.A(net474),
    .B(_0430_),
    .Y(_0072_));
 sky130_fd_sc_hd__nor2_2 _0861_ (.A(net468),
    .B(net311),
    .Y(_0431_));
 sky130_fd_sc_hd__a22o_2 _0862_ (.A1(\wb_counter[10] ),
    .A2(net468),
    .B1(net339),
    .B2(_0431_),
    .X(_0432_));
 sky130_fd_sc_hd__a22o_1 _0863_ (.A1(net373),
    .A2(net405),
    .B1(_0421_),
    .B2(_0432_),
    .X(_0433_));
 sky130_fd_sc_hd__and2_1 _0864_ (.A(net465),
    .B(_0433_),
    .X(_0073_));
 sky130_fd_sc_hd__a22oi_4 _0865_ (.A1(\wb_counter[11] ),
    .A2(net468),
    .B1(net340),
    .B2(_0431_),
    .Y(_0434_));
 sky130_fd_sc_hd__o2bb2a_1 _0866_ (.A1_N(net374),
    .A2_N(net403),
    .B1(_0422_),
    .B2(_0434_),
    .X(_0435_));
 sky130_fd_sc_hd__nor2_1 _0867_ (.A(net474),
    .B(_0435_),
    .Y(_0074_));
 sky130_fd_sc_hd__o21ai_1 _0868_ (.A1(net312),
    .A2(_0285_),
    .B1(net472),
    .Y(_0436_));
 sky130_fd_sc_hd__or2_1 _0869_ (.A(\wb_counter[12] ),
    .B(net472),
    .X(_0437_));
 sky130_fd_sc_hd__a32o_1 _0870_ (.A1(net400),
    .A2(_0436_),
    .A3(_0437_),
    .B1(net403),
    .B2(net375),
    .X(_0438_));
 sky130_fd_sc_hd__and2_1 _0871_ (.A(net465),
    .B(_0438_),
    .X(_0075_));
 sky130_fd_sc_hd__a21o_1 _0872_ (.A1(_0210_),
    .A2(net342),
    .B1(net468),
    .X(_0439_));
 sky130_fd_sc_hd__or2_1 _0873_ (.A(\wb_counter[13] ),
    .B(net472),
    .X(_0440_));
 sky130_fd_sc_hd__a32o_1 _0874_ (.A1(net400),
    .A2(_0439_),
    .A3(_0440_),
    .B1(net403),
    .B2(net376),
    .X(_0441_));
 sky130_fd_sc_hd__and2_1 _0875_ (.A(net465),
    .B(_0441_),
    .X(_0076_));
 sky130_fd_sc_hd__nor2_2 _0876_ (.A(net468),
    .B(net315),
    .Y(_0442_));
 sky130_fd_sc_hd__o2bb2a_1 _0877_ (.A1_N(net343),
    .A2_N(_0442_),
    .B1(_0173_),
    .B2(net472),
    .X(_0443_));
 sky130_fd_sc_hd__o2bb2a_1 _0878_ (.A1_N(net377),
    .A2_N(net404),
    .B1(_0422_),
    .B2(_0443_),
    .X(_0444_));
 sky130_fd_sc_hd__nor2_1 _0879_ (.A(net475),
    .B(_0444_),
    .Y(_0077_));
 sky130_fd_sc_hd__a22oi_4 _0880_ (.A1(\wb_counter[15] ),
    .A2(net468),
    .B1(net344),
    .B2(_0442_),
    .Y(_0445_));
 sky130_fd_sc_hd__o2bb2a_1 _0881_ (.A1_N(net378),
    .A2_N(net404),
    .B1(_0422_),
    .B2(_0445_),
    .X(_0118_));
 sky130_fd_sc_hd__nor2_1 _0882_ (.A(net475),
    .B(_0118_),
    .Y(_0078_));
 sky130_fd_sc_hd__mux2_2 _0883_ (.A0(\wb_counter[16] ),
    .A1(net345),
    .S(net472),
    .X(_0119_));
 sky130_fd_sc_hd__a22o_1 _0884_ (.A1(net379),
    .A2(net405),
    .B1(net400),
    .B2(_0119_),
    .X(_0120_));
 sky130_fd_sc_hd__and2_1 _0885_ (.A(net466),
    .B(_0120_),
    .X(_0079_));
 sky130_fd_sc_hd__mux2_2 _0886_ (.A0(\wb_counter[17] ),
    .A1(net346),
    .S(net472),
    .X(_0121_));
 sky130_fd_sc_hd__a22oi_1 _0887_ (.A1(net380),
    .A2(net405),
    .B1(net400),
    .B2(_0121_),
    .Y(_0122_));
 sky130_fd_sc_hd__nor2_1 _0888_ (.A(net475),
    .B(_0122_),
    .Y(_0080_));
 sky130_fd_sc_hd__mux2_2 _0889_ (.A0(\wb_counter[18] ),
    .A1(net347),
    .S(net473),
    .X(_0123_));
 sky130_fd_sc_hd__a22o_1 _0890_ (.A1(net381),
    .A2(net405),
    .B1(_0421_),
    .B2(_0123_),
    .X(_0124_));
 sky130_fd_sc_hd__and2_1 _0891_ (.A(net466),
    .B(_0124_),
    .X(_0081_));
 sky130_fd_sc_hd__mux2_2 _0892_ (.A0(\wb_counter[19] ),
    .A1(net349),
    .S(net472),
    .X(_0125_));
 sky130_fd_sc_hd__a22oi_1 _0893_ (.A1(net382),
    .A2(net406),
    .B1(net400),
    .B2(_0125_),
    .Y(_0126_));
 sky130_fd_sc_hd__nor2_1 _0894_ (.A(net475),
    .B(_0126_),
    .Y(_0082_));
 sky130_fd_sc_hd__mux2_2 _0895_ (.A0(\wb_counter[20] ),
    .A1(net350),
    .S(net473),
    .X(_0127_));
 sky130_fd_sc_hd__a22o_1 _0896_ (.A1(net384),
    .A2(net405),
    .B1(net400),
    .B2(_0127_),
    .X(_0128_));
 sky130_fd_sc_hd__and2_1 _0897_ (.A(net466),
    .B(_0128_),
    .X(_0083_));
 sky130_fd_sc_hd__nor2_2 _0898_ (.A(net469),
    .B(net326),
    .Y(_0129_));
 sky130_fd_sc_hd__a22oi_4 _0899_ (.A1(\wb_counter[21] ),
    .A2(net468),
    .B1(net351),
    .B2(_0129_),
    .Y(_0130_));
 sky130_fd_sc_hd__o2bb2a_1 _0900_ (.A1_N(net385),
    .A2_N(net403),
    .B1(_0422_),
    .B2(_0130_),
    .X(_0131_));
 sky130_fd_sc_hd__nor2_1 _0901_ (.A(net475),
    .B(_0131_),
    .Y(_0084_));
 sky130_fd_sc_hd__mux2_1 _0902_ (.A0(\wb_counter[22] ),
    .A1(net352),
    .S(net473),
    .X(_0132_));
 sky130_fd_sc_hd__a22o_1 _0903_ (.A1(net386),
    .A2(net405),
    .B1(net400),
    .B2(_0132_),
    .X(_0133_));
 sky130_fd_sc_hd__and2_1 _0904_ (.A(net465),
    .B(_0133_),
    .X(_0085_));
 sky130_fd_sc_hd__o2bb2a_1 _0905_ (.A1_N(net353),
    .A2_N(_0129_),
    .B1(_0172_),
    .B2(net471),
    .X(_0134_));
 sky130_fd_sc_hd__o2bb2a_1 _0906_ (.A1_N(net387),
    .A2_N(net403),
    .B1(_0422_),
    .B2(_0134_),
    .X(_0135_));
 sky130_fd_sc_hd__nor2_1 _0907_ (.A(net475),
    .B(_0135_),
    .Y(_0086_));
 sky130_fd_sc_hd__a32o_1 _0908_ (.A1(net473),
    .A2(net354),
    .A3(net400),
    .B1(net405),
    .B2(net388),
    .X(_0136_));
 sky130_fd_sc_hd__and2_1 _0909_ (.A(net465),
    .B(_0136_),
    .X(_0087_));
 sky130_fd_sc_hd__a32o_1 _0910_ (.A1(net473),
    .A2(net355),
    .A3(_0421_),
    .B1(net405),
    .B2(net389),
    .X(_0137_));
 sky130_fd_sc_hd__and2_1 _0911_ (.A(net465),
    .B(_0137_),
    .X(_0088_));
 sky130_fd_sc_hd__nand2_1 _0912_ (.A(net390),
    .B(net405),
    .Y(_0138_));
 sky130_fd_sc_hd__or4b_2 _0913_ (.A(net469),
    .B(net326),
    .C(_0422_),
    .D_N(net356),
    .X(_0139_));
 sky130_fd_sc_hd__a21oi_1 _0914_ (.A1(_0138_),
    .A2(_0139_),
    .B1(net475),
    .Y(_0089_));
 sky130_fd_sc_hd__a32o_1 _0915_ (.A1(net473),
    .A2(net327),
    .A3(net400),
    .B1(net406),
    .B2(net391),
    .X(_0140_));
 sky130_fd_sc_hd__and2_1 _0916_ (.A(net466),
    .B(_0140_),
    .X(_0090_));
 sky130_fd_sc_hd__nand2_1 _0917_ (.A(net509),
    .B(net462),
    .Y(_0141_));
 sky130_fd_sc_hd__xnor2_1 _0918_ (.A(net509),
    .B(net476),
    .Y(_0091_));
 sky130_fd_sc_hd__xnor2_1 _0919_ (.A(net511),
    .B(_0141_),
    .Y(_0092_));
 sky130_fd_sc_hd__and4b_2 _0920_ (.A_N(net476),
    .B(net509),
    .C(net511),
    .D(net553),
    .X(_0142_));
 sky130_fd_sc_hd__a31o_1 _0921_ (.A1(net511),
    .A2(net509),
    .A3(net462),
    .B1(net553),
    .X(_0143_));
 sky130_fd_sc_hd__and2b_1 _0922_ (.A_N(_0142_),
    .B(net554),
    .X(_0093_));
 sky130_fd_sc_hd__nand2_1 _0923_ (.A(net556),
    .B(_0142_),
    .Y(_0144_));
 sky130_fd_sc_hd__or2_1 _0924_ (.A(net556),
    .B(_0142_),
    .X(_0145_));
 sky130_fd_sc_hd__and2_1 _0925_ (.A(net557),
    .B(_0145_),
    .X(_0094_));
 sky130_fd_sc_hd__xnor2_1 _0926_ (.A(net528),
    .B(net557),
    .Y(_0095_));
 sky130_fd_sc_hd__and4_2 _0927_ (.A(net544),
    .B(net528),
    .C(net556),
    .D(_0142_),
    .X(_0146_));
 sky130_fd_sc_hd__a31o_1 _0928_ (.A1(net528),
    .A2(net357),
    .A3(_0142_),
    .B1(net544),
    .X(_0147_));
 sky130_fd_sc_hd__and2b_1 _0929_ (.A_N(_0146_),
    .B(net545),
    .X(_0096_));
 sky130_fd_sc_hd__xor2_1 _0930_ (.A(net497),
    .B(_0146_),
    .X(_0097_));
 sky130_fd_sc_hd__and2_1 _0931_ (.A(net533),
    .B(net497),
    .X(_0148_));
 sky130_fd_sc_hd__and2_1 _0932_ (.A(_0146_),
    .B(_0148_),
    .X(_0149_));
 sky130_fd_sc_hd__a21oi_1 _0933_ (.A1(net497),
    .A2(_0146_),
    .B1(net533),
    .Y(_0150_));
 sky130_fd_sc_hd__nor2_1 _0934_ (.A(_0149_),
    .B(net534),
    .Y(_0098_));
 sky130_fd_sc_hd__xnor2_1 _0935_ (.A(net514),
    .B(_0149_),
    .Y(_0099_));
 sky130_fd_sc_hd__nor2_1 _0936_ (.A(_0174_),
    .B(net514),
    .Y(_0151_));
 sky130_fd_sc_hd__and3_1 _0937_ (.A(_0146_),
    .B(_0148_),
    .C(_0151_),
    .X(_0152_));
 sky130_fd_sc_hd__a21oi_1 _0938_ (.A1(net513),
    .A2(_0149_),
    .B1(net525),
    .Y(_0153_));
 sky130_fd_sc_hd__nor2_1 _0939_ (.A(_0152_),
    .B(net526),
    .Y(_0100_));
 sky130_fd_sc_hd__and4_2 _0940_ (.A(net522),
    .B(_0146_),
    .C(_0148_),
    .D(_0151_),
    .X(_0154_));
 sky130_fd_sc_hd__nor2_1 _0941_ (.A(net522),
    .B(_0152_),
    .Y(_0155_));
 sky130_fd_sc_hd__nor2_1 _0942_ (.A(_0154_),
    .B(net523),
    .Y(_0101_));
 sky130_fd_sc_hd__and2_2 _0943_ (.A(net530),
    .B(_0154_),
    .X(_0156_));
 sky130_fd_sc_hd__nor2_1 _0944_ (.A(net530),
    .B(_0154_),
    .Y(_0157_));
 sky130_fd_sc_hd__nor2_1 _0945_ (.A(_0156_),
    .B(net531),
    .Y(_0102_));
 sky130_fd_sc_hd__xor2_1 _0946_ (.A(net503),
    .B(_0156_),
    .X(_0103_));
 sky130_fd_sc_hd__and3_1 _0947_ (.A(net538),
    .B(net503),
    .C(_0156_),
    .X(_0158_));
 sky130_fd_sc_hd__a21oi_1 _0948_ (.A1(net503),
    .A2(_0156_),
    .B1(net538),
    .Y(_0159_));
 sky130_fd_sc_hd__nor2_1 _0949_ (.A(_0158_),
    .B(net539),
    .Y(_0104_));
 sky130_fd_sc_hd__and2_1 _0950_ (.A(net519),
    .B(_0158_),
    .X(_0160_));
 sky130_fd_sc_hd__xnor2_1 _0951_ (.A(net520),
    .B(_0158_),
    .Y(_0105_));
 sky130_fd_sc_hd__and4_1 _0952_ (.A(net536),
    .B(net519),
    .C(net538),
    .D(net503),
    .X(_0161_));
 sky130_fd_sc_hd__o2bb2a_1 _0953_ (.A1_N(_0156_),
    .A2_N(_0161_),
    .B1(_0160_),
    .B2(net536),
    .X(_0106_));
 sky130_fd_sc_hd__and4_2 _0954_ (.A(net541),
    .B(net530),
    .C(_0154_),
    .D(_0161_),
    .X(_0162_));
 sky130_fd_sc_hd__a21oi_1 _0955_ (.A1(_0156_),
    .A2(_0161_),
    .B1(net541),
    .Y(_0163_));
 sky130_fd_sc_hd__nor2_1 _0956_ (.A(_0162_),
    .B(net542),
    .Y(_0107_));
 sky130_fd_sc_hd__nand2_1 _0957_ (.A(net505),
    .B(_0162_),
    .Y(_0164_));
 sky130_fd_sc_hd__xor2_1 _0958_ (.A(net505),
    .B(_0162_),
    .X(_0108_));
 sky130_fd_sc_hd__xnor2_1 _0959_ (.A(net501),
    .B(_0164_),
    .Y(_0109_));
 sky130_fd_sc_hd__and4_2 _0960_ (.A(net547),
    .B(net501),
    .C(net505),
    .D(_0162_),
    .X(_0165_));
 sky130_fd_sc_hd__a31o_1 _0961_ (.A1(net501),
    .A2(net505),
    .A3(_0162_),
    .B1(net547),
    .X(_0166_));
 sky130_fd_sc_hd__and2b_1 _0962_ (.A_N(_0165_),
    .B(net548),
    .X(_0110_));
 sky130_fd_sc_hd__nand2_1 _0963_ (.A(net499),
    .B(_0165_),
    .Y(_0167_));
 sky130_fd_sc_hd__xor2_1 _0964_ (.A(net499),
    .B(_0165_),
    .X(_0111_));
 sky130_fd_sc_hd__xnor2_1 _0965_ (.A(net507),
    .B(_0167_),
    .Y(_0112_));
 sky130_fd_sc_hd__and4_1 _0966_ (.A(net550),
    .B(net507),
    .C(net499),
    .D(_0165_),
    .X(_0168_));
 sky130_fd_sc_hd__a31o_1 _0967_ (.A1(net507),
    .A2(net499),
    .A3(_0165_),
    .B1(net550),
    .X(_0169_));
 sky130_fd_sc_hd__and2b_1 _0968_ (.A_N(_0168_),
    .B(net551),
    .X(_0113_));
 sky130_fd_sc_hd__xnor2_1 _0969_ (.A(net517),
    .B(_0168_),
    .Y(_0114_));
 sky130_fd_sc_hd__mux2_1 _0970_ (.A0(wb_rst_override),
    .A1(net251),
    .S(_0352_),
    .X(_0170_));
 sky130_fd_sc_hd__and2_1 _0971_ (.A(net461),
    .B(_0170_),
    .X(_0115_));
 sky130_fd_sc_hd__mux2_1 _0972_ (.A0(wb_clk_override),
    .A1(net261),
    .S(_0357_),
    .X(_0116_));
 sky130_fd_sc_hd__mux2_1 _0973_ (.A0(net448),
    .A1(net240),
    .S(_0352_),
    .X(_0171_));
 sky130_fd_sc_hd__and2_1 _0974_ (.A(net461),
    .B(_0171_),
    .X(_0117_));
 sky130_fd_sc_hd__dfxtp_1 _0975_ (.CLK(clknet_3_1__leaf_wb_clk_i),
    .D(_0000_),
    .Q(\wb_design_addr_override[0] ));
 sky130_fd_sc_hd__dfxtp_2 _0976_ (.CLK(clknet_3_1__leaf_wb_clk_i),
    .D(_0001_),
    .Q(\wb_design_addr_override[1] ));
 sky130_fd_sc_hd__dfxtp_2 _0977_ (.CLK(clknet_3_0__leaf_wb_clk_i),
    .D(_0002_),
    .Q(\wb_design_addr_override[2] ));
 sky130_fd_sc_hd__dfxtp_1 _0978_ (.CLK(clknet_3_1__leaf_wb_clk_i),
    .D(_0003_),
    .Q(\wb_design_addr_override[3] ));
 sky130_fd_sc_hd__dfxtp_1 _0979_ (.CLK(clknet_3_0__leaf_wb_clk_i),
    .D(_0004_),
    .Q(wb_single_step));
 sky130_fd_sc_hd__dfxtp_1 _0980_ (.CLK(clknet_3_5__leaf_wb_clk_i),
    .D(_0005_),
    .Q(wb_feedback_delay));
 sky130_fd_sc_hd__dfxtp_4 _0981_ (.CLK(clknet_3_1__leaf_wb_clk_i),
    .D(_0006_),
    .Q(\wb_counter[0] ));
 sky130_fd_sc_hd__dfxtp_4 _0982_ (.CLK(clknet_3_1__leaf_wb_clk_i),
    .D(_0007_),
    .Q(net337));
 sky130_fd_sc_hd__dfxtp_4 _0983_ (.CLK(clknet_3_1__leaf_wb_clk_i),
    .D(_0008_),
    .Q(net348));
 sky130_fd_sc_hd__dfxtp_4 _0984_ (.CLK(clknet_3_1__leaf_wb_clk_i),
    .D(_0009_),
    .Q(net357));
 sky130_fd_sc_hd__dfxtp_4 _0985_ (.CLK(clknet_3_0__leaf_wb_clk_i),
    .D(_0010_),
    .Q(net358));
 sky130_fd_sc_hd__dfxtp_2 _0986_ (.CLK(clknet_3_3__leaf_wb_clk_i),
    .D(_0011_),
    .Q(\wb_counter[5] ));
 sky130_fd_sc_hd__dfxtp_2 _0987_ (.CLK(clknet_3_3__leaf_wb_clk_i),
    .D(_0012_),
    .Q(\wb_counter[6] ));
 sky130_fd_sc_hd__dfxtp_1 _0988_ (.CLK(clknet_3_3__leaf_wb_clk_i),
    .D(_0013_),
    .Q(\wb_counter[7] ));
 sky130_fd_sc_hd__dfxtp_1 _0989_ (.CLK(clknet_3_2__leaf_wb_clk_i),
    .D(_0014_),
    .Q(\wb_counter[8] ));
 sky130_fd_sc_hd__dfxtp_1 _0990_ (.CLK(clknet_3_2__leaf_wb_clk_i),
    .D(_0015_),
    .Q(\wb_counter[9] ));
 sky130_fd_sc_hd__dfxtp_1 _0991_ (.CLK(clknet_3_2__leaf_wb_clk_i),
    .D(_0016_),
    .Q(\wb_counter[10] ));
 sky130_fd_sc_hd__dfxtp_2 _0992_ (.CLK(clknet_3_2__leaf_wb_clk_i),
    .D(_0017_),
    .Q(\wb_counter[11] ));
 sky130_fd_sc_hd__dfxtp_2 _0993_ (.CLK(clknet_3_3__leaf_wb_clk_i),
    .D(_0018_),
    .Q(\wb_counter[12] ));
 sky130_fd_sc_hd__dfxtp_2 _0994_ (.CLK(clknet_3_6__leaf_wb_clk_i),
    .D(_0019_),
    .Q(\wb_counter[13] ));
 sky130_fd_sc_hd__dfxtp_1 _0995_ (.CLK(clknet_3_2__leaf_wb_clk_i),
    .D(_0020_),
    .Q(\wb_counter[14] ));
 sky130_fd_sc_hd__dfxtp_2 _0996_ (.CLK(clknet_3_3__leaf_wb_clk_i),
    .D(_0021_),
    .Q(\wb_counter[15] ));
 sky130_fd_sc_hd__dfxtp_1 _0997_ (.CLK(clknet_3_2__leaf_wb_clk_i),
    .D(_0022_),
    .Q(\wb_counter[16] ));
 sky130_fd_sc_hd__dfxtp_4 _0998_ (.CLK(clknet_3_6__leaf_wb_clk_i),
    .D(_0023_),
    .Q(\wb_counter[17] ));
 sky130_fd_sc_hd__dfxtp_2 _0999_ (.CLK(clknet_3_3__leaf_wb_clk_i),
    .D(_0024_),
    .Q(\wb_counter[18] ));
 sky130_fd_sc_hd__dfxtp_2 _1000_ (.CLK(clknet_3_6__leaf_wb_clk_i),
    .D(_0025_),
    .Q(\wb_counter[19] ));
 sky130_fd_sc_hd__dfxtp_2 _1001_ (.CLK(clknet_3_3__leaf_wb_clk_i),
    .D(_0026_),
    .Q(\wb_counter[20] ));
 sky130_fd_sc_hd__dfxtp_4 _1002_ (.CLK(clknet_3_6__leaf_wb_clk_i),
    .D(_0027_),
    .Q(\wb_counter[21] ));
 sky130_fd_sc_hd__dfxtp_1 _1003_ (.CLK(clknet_3_6__leaf_wb_clk_i),
    .D(_0028_),
    .Q(\wb_counter[22] ));
 sky130_fd_sc_hd__dfxtp_1 _1004_ (.CLK(clknet_3_2__leaf_wb_clk_i),
    .D(_0029_),
    .Q(\wb_counter[23] ));
 sky130_fd_sc_hd__dfxtp_1 _1005_ (.CLK(clknet_3_5__leaf_wb_clk_i),
    .D(_0030_),
    .Q(net371));
 sky130_fd_sc_hd__dfxtp_1 _1006_ (.CLK(clknet_3_1__leaf_wb_clk_i),
    .D(_0031_),
    .Q(\wb_io_override[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1007_ (.CLK(clknet_3_0__leaf_wb_clk_i),
    .D(_0032_),
    .Q(\wb_io_override[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1008_ (.CLK(clknet_3_0__leaf_wb_clk_i),
    .D(_0033_),
    .Q(\wb_io_override[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1009_ (.CLK(clknet_3_0__leaf_wb_clk_i),
    .D(_0034_),
    .Q(\wb_io_override[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1010_ (.CLK(clknet_3_0__leaf_wb_clk_i),
    .D(_0035_),
    .Q(\wb_io_override[4] ));
 sky130_fd_sc_hd__dfxtp_1 _1011_ (.CLK(clknet_3_0__leaf_wb_clk_i),
    .D(_0036_),
    .Q(\wb_io_override[5] ));
 sky130_fd_sc_hd__dfxtp_1 _1012_ (.CLK(clknet_3_0__leaf_wb_clk_i),
    .D(_0037_),
    .Q(\wb_io_override[6] ));
 sky130_fd_sc_hd__dfxtp_1 _1013_ (.CLK(clknet_3_1__leaf_wb_clk_i),
    .D(_0038_),
    .Q(\wb_io_override[7] ));
 sky130_fd_sc_hd__dfxtp_1 _1014_ (.CLK(clknet_3_0__leaf_wb_clk_i),
    .D(_0039_),
    .Q(\wb_io_override[8] ));
 sky130_fd_sc_hd__dfxtp_1 _1015_ (.CLK(clknet_3_0__leaf_wb_clk_i),
    .D(_0040_),
    .Q(\wb_io_override[9] ));
 sky130_fd_sc_hd__dfxtp_1 _1016_ (.CLK(clknet_3_0__leaf_wb_clk_i),
    .D(_0041_),
    .Q(\wb_io_override[10] ));
 sky130_fd_sc_hd__dfxtp_1 _1017_ (.CLK(clknet_3_2__leaf_wb_clk_i),
    .D(_0042_),
    .Q(\wb_io_override[11] ));
 sky130_fd_sc_hd__dfxtp_1 _1018_ (.CLK(clknet_3_3__leaf_wb_clk_i),
    .D(_0043_),
    .Q(\wb_io_override[12] ));
 sky130_fd_sc_hd__dfxtp_2 _1019_ (.CLK(clknet_3_4__leaf_wb_clk_i),
    .D(_0044_),
    .Q(\wb_io_override[13] ));
 sky130_fd_sc_hd__dfxtp_1 _1020_ (.CLK(clknet_3_2__leaf_wb_clk_i),
    .D(_0045_),
    .Q(\wb_io_override[14] ));
 sky130_fd_sc_hd__dfxtp_1 _1021_ (.CLK(clknet_3_3__leaf_wb_clk_i),
    .D(_0046_),
    .Q(\wb_io_override[15] ));
 sky130_fd_sc_hd__dfxtp_1 _1022_ (.CLK(clknet_3_0__leaf_wb_clk_i),
    .D(_0047_),
    .Q(\wb_io_override[16] ));
 sky130_fd_sc_hd__dfxtp_1 _1023_ (.CLK(clknet_3_1__leaf_wb_clk_i),
    .D(_0048_),
    .Q(\wb_io_override[17] ));
 sky130_fd_sc_hd__dfxtp_1 _1024_ (.CLK(clknet_3_3__leaf_wb_clk_i),
    .D(_0049_),
    .Q(\wb_io_override[18] ));
 sky130_fd_sc_hd__dfxtp_1 _1025_ (.CLK(clknet_3_1__leaf_wb_clk_i),
    .D(_0050_),
    .Q(\wb_io_override[19] ));
 sky130_fd_sc_hd__dfxtp_1 _1026_ (.CLK(clknet_3_0__leaf_wb_clk_i),
    .D(_0051_),
    .Q(\wb_io_override[20] ));
 sky130_fd_sc_hd__dfxtp_2 _1027_ (.CLK(clknet_3_6__leaf_wb_clk_i),
    .D(_0052_),
    .Q(\wb_io_override[21] ));
 sky130_fd_sc_hd__dfxtp_1 _1028_ (.CLK(clknet_3_1__leaf_wb_clk_i),
    .D(_0053_),
    .Q(\wb_io_override[22] ));
 sky130_fd_sc_hd__dfxtp_1 _1029_ (.CLK(clknet_3_2__leaf_wb_clk_i),
    .D(_0054_),
    .Q(\wb_io_override[23] ));
 sky130_fd_sc_hd__dfxtp_1 _1030_ (.CLK(clknet_3_2__leaf_wb_clk_i),
    .D(_0055_),
    .Q(\wb_io_override[24] ));
 sky130_fd_sc_hd__dfxtp_1 _1031_ (.CLK(clknet_3_2__leaf_wb_clk_i),
    .D(_0056_),
    .Q(\wb_io_override[25] ));
 sky130_fd_sc_hd__dfxtp_1 _1032_ (.CLK(clknet_3_2__leaf_wb_clk_i),
    .D(_0057_),
    .Q(\wb_io_override[26] ));
 sky130_fd_sc_hd__dfxtp_1 _1033_ (.CLK(clknet_3_2__leaf_wb_clk_i),
    .D(_0058_),
    .Q(\wb_io_override[27] ));
 sky130_fd_sc_hd__dfxtp_1 _1034_ (.CLK(clknet_3_0__leaf_wb_clk_i),
    .D(_0059_),
    .Q(\design_addr[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1035_ (.CLK(clknet_3_0__leaf_wb_clk_i),
    .D(_0060_),
    .Q(\design_addr[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1036_ (.CLK(clknet_3_0__leaf_wb_clk_i),
    .D(_0061_),
    .Q(\design_addr[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1037_ (.CLK(clknet_3_0__leaf_wb_clk_i),
    .D(_0062_),
    .Q(\design_addr[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1038_ (.CLK(clknet_3_5__leaf_wb_clk_i),
    .D(_0063_),
    .Q(net372));
 sky130_fd_sc_hd__dfxtp_1 _1039_ (.CLK(clknet_3_5__leaf_wb_clk_i),
    .D(_0064_),
    .Q(net383));
 sky130_fd_sc_hd__dfxtp_1 _1040_ (.CLK(clknet_3_5__leaf_wb_clk_i),
    .D(_0065_),
    .Q(net392));
 sky130_fd_sc_hd__dfxtp_1 _1041_ (.CLK(clknet_3_4__leaf_wb_clk_i),
    .D(_0066_),
    .Q(net393));
 sky130_fd_sc_hd__dfxtp_1 _1042_ (.CLK(clknet_3_5__leaf_wb_clk_i),
    .D(_0067_),
    .Q(net394));
 sky130_fd_sc_hd__dfxtp_1 _1043_ (.CLK(clknet_3_5__leaf_wb_clk_i),
    .D(_0068_),
    .Q(net395));
 sky130_fd_sc_hd__dfxtp_1 _1044_ (.CLK(clknet_3_4__leaf_wb_clk_i),
    .D(_0069_),
    .Q(net396));
 sky130_fd_sc_hd__dfxtp_1 _1045_ (.CLK(clknet_3_5__leaf_wb_clk_i),
    .D(_0070_),
    .Q(net397));
 sky130_fd_sc_hd__dfxtp_1 _1046_ (.CLK(clknet_3_6__leaf_wb_clk_i),
    .D(_0071_),
    .Q(net398));
 sky130_fd_sc_hd__dfxtp_1 _1047_ (.CLK(clknet_3_6__leaf_wb_clk_i),
    .D(_0072_),
    .Q(net399));
 sky130_fd_sc_hd__dfxtp_1 _1048_ (.CLK(clknet_3_4__leaf_wb_clk_i),
    .D(_0073_),
    .Q(net373));
 sky130_fd_sc_hd__dfxtp_1 _1049_ (.CLK(clknet_3_6__leaf_wb_clk_i),
    .D(_0074_),
    .Q(net374));
 sky130_fd_sc_hd__dfxtp_1 _1050_ (.CLK(clknet_3_6__leaf_wb_clk_i),
    .D(_0075_),
    .Q(net375));
 sky130_fd_sc_hd__dfxtp_2 _1051_ (.CLK(clknet_3_6__leaf_wb_clk_i),
    .D(_0076_),
    .Q(net376));
 sky130_fd_sc_hd__dfxtp_1 _1052_ (.CLK(clknet_3_6__leaf_wb_clk_i),
    .D(_0077_),
    .Q(net377));
 sky130_fd_sc_hd__dfxtp_1 _1053_ (.CLK(clknet_3_7__leaf_wb_clk_i),
    .D(_0078_),
    .Q(net378));
 sky130_fd_sc_hd__dfxtp_1 _1054_ (.CLK(clknet_3_7__leaf_wb_clk_i),
    .D(_0079_),
    .Q(net379));
 sky130_fd_sc_hd__dfxtp_1 _1055_ (.CLK(clknet_3_7__leaf_wb_clk_i),
    .D(_0080_),
    .Q(net380));
 sky130_fd_sc_hd__dfxtp_1 _1056_ (.CLK(clknet_3_7__leaf_wb_clk_i),
    .D(_0081_),
    .Q(net381));
 sky130_fd_sc_hd__dfxtp_1 _1057_ (.CLK(clknet_3_7__leaf_wb_clk_i),
    .D(_0082_),
    .Q(net382));
 sky130_fd_sc_hd__dfxtp_1 _1058_ (.CLK(clknet_3_7__leaf_wb_clk_i),
    .D(_0083_),
    .Q(net384));
 sky130_fd_sc_hd__dfxtp_2 _1059_ (.CLK(clknet_3_6__leaf_wb_clk_i),
    .D(_0084_),
    .Q(net385));
 sky130_fd_sc_hd__dfxtp_2 _1060_ (.CLK(clknet_3_4__leaf_wb_clk_i),
    .D(_0085_),
    .Q(net386));
 sky130_fd_sc_hd__dfxtp_2 _1061_ (.CLK(clknet_3_7__leaf_wb_clk_i),
    .D(_0086_),
    .Q(net387));
 sky130_fd_sc_hd__dfxtp_2 _1062_ (.CLK(clknet_3_7__leaf_wb_clk_i),
    .D(_0087_),
    .Q(net388));
 sky130_fd_sc_hd__dfxtp_2 _1063_ (.CLK(clknet_3_4__leaf_wb_clk_i),
    .D(_0088_),
    .Q(net389));
 sky130_fd_sc_hd__dfxtp_2 _1064_ (.CLK(clknet_3_5__leaf_wb_clk_i),
    .D(_0089_),
    .Q(net390));
 sky130_fd_sc_hd__dfxtp_2 _1065_ (.CLK(clknet_3_7__leaf_wb_clk_i),
    .D(_0090_),
    .Q(net391));
 sky130_fd_sc_hd__dfxtp_4 _1066_ (.CLK(net270),
    .D(net510),
    .Q(\wb_counter[0] ));
 sky130_fd_sc_hd__dfxtp_4 _1067_ (.CLK(net270),
    .D(net512),
    .Q(net337));
 sky130_fd_sc_hd__dfxtp_4 _1068_ (.CLK(net270),
    .D(net555),
    .Q(net348));
 sky130_fd_sc_hd__dfxtp_4 _1069_ (.CLK(net270),
    .D(net558),
    .Q(net357));
 sky130_fd_sc_hd__dfxtp_4 _1070_ (.CLK(net270),
    .D(net529),
    .Q(net358));
 sky130_fd_sc_hd__dfxtp_2 _1071_ (.CLK(net270),
    .D(net546),
    .Q(\wb_counter[5] ));
 sky130_fd_sc_hd__dfxtp_2 _1072_ (.CLK(net270),
    .D(net498),
    .Q(\wb_counter[6] ));
 sky130_fd_sc_hd__dfxtp_1 _1073_ (.CLK(net270),
    .D(net535),
    .Q(\wb_counter[7] ));
 sky130_fd_sc_hd__dfxtp_1 _1074_ (.CLK(net270),
    .D(net515),
    .Q(\wb_counter[8] ));
 sky130_fd_sc_hd__dfxtp_1 _1075_ (.CLK(net270),
    .D(net527),
    .Q(\wb_counter[9] ));
 sky130_fd_sc_hd__dfxtp_1 _1076_ (.CLK(net270),
    .D(net524),
    .Q(\wb_counter[10] ));
 sky130_fd_sc_hd__dfxtp_2 _1077_ (.CLK(net270),
    .D(net532),
    .Q(\wb_counter[11] ));
 sky130_fd_sc_hd__dfxtp_2 _1078_ (.CLK(net270),
    .D(net504),
    .Q(\wb_counter[12] ));
 sky130_fd_sc_hd__dfxtp_2 _1079_ (.CLK(net270),
    .D(net540),
    .Q(\wb_counter[13] ));
 sky130_fd_sc_hd__dfxtp_1 _1080_ (.CLK(net270),
    .D(net521),
    .Q(\wb_counter[14] ));
 sky130_fd_sc_hd__dfxtp_2 _1081_ (.CLK(net270),
    .D(net537),
    .Q(\wb_counter[15] ));
 sky130_fd_sc_hd__dfxtp_1 _1082_ (.CLK(net270),
    .D(net543),
    .Q(\wb_counter[16] ));
 sky130_fd_sc_hd__dfxtp_4 _1083_ (.CLK(net270),
    .D(net506),
    .Q(\wb_counter[17] ));
 sky130_fd_sc_hd__dfxtp_2 _1084_ (.CLK(net270),
    .D(net502),
    .Q(\wb_counter[18] ));
 sky130_fd_sc_hd__dfxtp_2 _1085_ (.CLK(net270),
    .D(net549),
    .Q(\wb_counter[19] ));
 sky130_fd_sc_hd__dfxtp_2 _1086_ (.CLK(net270),
    .D(net500),
    .Q(\wb_counter[20] ));
 sky130_fd_sc_hd__dfxtp_4 _1087_ (.CLK(net270),
    .D(net508),
    .Q(\wb_counter[21] ));
 sky130_fd_sc_hd__dfxtp_1 _1088_ (.CLK(net270),
    .D(net552),
    .Q(\wb_counter[22] ));
 sky130_fd_sc_hd__dfxtp_1 _1089_ (.CLK(net270),
    .D(net518),
    .Q(\wb_counter[23] ));
 sky130_fd_sc_hd__dfxtp_2 _1090_ (.CLK(clknet_3_1__leaf_wb_clk_i),
    .D(_0115_),
    .Q(wb_rst_override));
 sky130_fd_sc_hd__dfxtp_1 _1091_ (.CLK(clknet_3_0__leaf_wb_clk_i),
    .D(_0116_),
    .Q(wb_clk_override));
 sky130_fd_sc_hd__dfxtp_2 _1092_ (.CLK(clknet_3_1__leaf_wb_clk_i),
    .D(_0117_),
    .Q(wb_override));
 sky130_fd_sc_hd__conb_1 multiplexer_492 (.HI(net492));
 sky130_fd_sc_hd__conb_1 multiplexer_493 (.HI(net493));
 sky130_fd_sc_hd__conb_1 multiplexer_494 (.HI(net494));
 sky130_fd_sc_hd__conb_1 multiplexer_495 (.HI(net495));
 sky130_fd_sc_hd__conb_1 multiplexer_496 (.HI(net496));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_wb_clk_i (.A(wb_clk_i),
    .X(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__conb_1 multiplexer_478 (.LO(net478));
 sky130_fd_sc_hd__conb_1 multiplexer_479 (.LO(net479));
 sky130_fd_sc_hd__conb_1 multiplexer_480 (.LO(net480));
 sky130_fd_sc_hd__conb_1 multiplexer_481 (.LO(net481));
 sky130_fd_sc_hd__conb_1 multiplexer_482 (.LO(net482));
 sky130_fd_sc_hd__conb_1 multiplexer_483 (.LO(net483));
 sky130_fd_sc_hd__conb_1 multiplexer_484 (.LO(net484));
 sky130_fd_sc_hd__conb_1 multiplexer_485 (.LO(net485));
 sky130_fd_sc_hd__conb_1 multiplexer_486 (.LO(net486));
 sky130_fd_sc_hd__conb_1 multiplexer_487 (.LO(net487));
 sky130_fd_sc_hd__conb_1 multiplexer_488 (.LO(net488));
 sky130_fd_sc_hd__conb_1 multiplexer_489 (.LO(net489));
 sky130_fd_sc_hd__conb_1 multiplexer_490 (.LO(net490));
 sky130_fd_sc_hd__conb_1 multiplexer_491 (.HI(net491));
 sky130_fd_sc_hd__clkbuf_2 _1113_ (.A(net302),
    .X(net301));
 sky130_fd_sc_hd__clkbuf_2 _1114_ (.A(net307),
    .X(net306));
 sky130_fd_sc_hd__clkbuf_2 _1115_ (.A(net309),
    .X(net308));
 sky130_fd_sc_hd__clkbuf_2 _1116_ (.A(net311),
    .X(net310));
 sky130_fd_sc_hd__clkbuf_2 _1117_ (.A(net315),
    .X(net314));
 sky130_fd_sc_hd__clkbuf_2 _1118_ (.A(net415),
    .X(net316));
 sky130_fd_sc_hd__clkbuf_2 _1119_ (.A(net416),
    .X(net317));
 sky130_fd_sc_hd__clkbuf_2 _1120_ (.A(net416),
    .X(net318));
 sky130_fd_sc_hd__clkbuf_2 _1121_ (.A(net416),
    .X(net319));
 sky130_fd_sc_hd__clkbuf_2 _1122_ (.A(net416),
    .X(net320));
 sky130_fd_sc_hd__clkbuf_2 _1123_ (.A(net326),
    .X(net321));
 sky130_fd_sc_hd__clkbuf_2 _1124_ (.A(net416),
    .X(net322));
 sky130_fd_sc_hd__clkbuf_2 _1125_ (.A(net326),
    .X(net323));
 sky130_fd_sc_hd__clkbuf_2 _1126_ (.A(net416),
    .X(net324));
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__decap_3 PHY_166 ();
 sky130_fd_sc_hd__decap_3 PHY_167 ();
 sky130_fd_sc_hd__decap_3 PHY_168 ();
 sky130_fd_sc_hd__decap_3 PHY_169 ();
 sky130_fd_sc_hd__decap_3 PHY_170 ();
 sky130_fd_sc_hd__decap_3 PHY_171 ();
 sky130_fd_sc_hd__decap_3 PHY_172 ();
 sky130_fd_sc_hd__decap_3 PHY_173 ();
 sky130_fd_sc_hd__decap_3 PHY_174 ();
 sky130_fd_sc_hd__decap_3 PHY_175 ();
 sky130_fd_sc_hd__decap_3 PHY_176 ();
 sky130_fd_sc_hd__decap_3 PHY_177 ();
 sky130_fd_sc_hd__decap_3 PHY_178 ();
 sky130_fd_sc_hd__decap_3 PHY_179 ();
 sky130_fd_sc_hd__decap_3 PHY_180 ();
 sky130_fd_sc_hd__decap_3 PHY_181 ();
 sky130_fd_sc_hd__decap_3 PHY_182 ();
 sky130_fd_sc_hd__decap_3 PHY_183 ();
 sky130_fd_sc_hd__decap_3 PHY_184 ();
 sky130_fd_sc_hd__decap_3 PHY_185 ();
 sky130_fd_sc_hd__decap_3 PHY_186 ();
 sky130_fd_sc_hd__decap_3 PHY_187 ();
 sky130_fd_sc_hd__decap_3 PHY_188 ();
 sky130_fd_sc_hd__decap_3 PHY_189 ();
 sky130_fd_sc_hd__decap_3 PHY_190 ();
 sky130_fd_sc_hd__decap_3 PHY_191 ();
 sky130_fd_sc_hd__decap_3 PHY_192 ();
 sky130_fd_sc_hd__decap_3 PHY_193 ();
 sky130_fd_sc_hd__decap_3 PHY_194 ();
 sky130_fd_sc_hd__decap_3 PHY_195 ();
 sky130_fd_sc_hd__decap_3 PHY_196 ();
 sky130_fd_sc_hd__decap_3 PHY_197 ();
 sky130_fd_sc_hd__decap_3 PHY_198 ();
 sky130_fd_sc_hd__decap_3 PHY_199 ();
 sky130_fd_sc_hd__decap_3 PHY_200 ();
 sky130_fd_sc_hd__decap_3 PHY_201 ();
 sky130_fd_sc_hd__decap_3 PHY_202 ();
 sky130_fd_sc_hd__decap_3 PHY_203 ();
 sky130_fd_sc_hd__decap_3 PHY_204 ();
 sky130_fd_sc_hd__decap_3 PHY_205 ();
 sky130_fd_sc_hd__decap_3 PHY_206 ();
 sky130_fd_sc_hd__decap_3 PHY_207 ();
 sky130_fd_sc_hd__decap_3 PHY_208 ();
 sky130_fd_sc_hd__decap_3 PHY_209 ();
 sky130_fd_sc_hd__decap_3 PHY_210 ();
 sky130_fd_sc_hd__decap_3 PHY_211 ();
 sky130_fd_sc_hd__decap_3 PHY_212 ();
 sky130_fd_sc_hd__decap_3 PHY_213 ();
 sky130_fd_sc_hd__decap_3 PHY_214 ();
 sky130_fd_sc_hd__decap_3 PHY_215 ();
 sky130_fd_sc_hd__decap_3 PHY_216 ();
 sky130_fd_sc_hd__decap_3 PHY_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1438 ();
 sky130_fd_sc_hd__clkbuf_2 input1 (.A(dso_6502[0]),
    .X(net1));
 sky130_fd_sc_hd__buf_4 input2 (.A(dso_6502[10]),
    .X(net2));
 sky130_fd_sc_hd__buf_4 input3 (.A(dso_6502[11]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_2 input4 (.A(dso_6502[12]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_2 input5 (.A(dso_6502[13]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_4 input6 (.A(dso_6502[14]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_4 input7 (.A(dso_6502[15]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_4 input8 (.A(dso_6502[16]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_2 input9 (.A(dso_6502[17]),
    .X(net9));
 sky130_fd_sc_hd__buf_2 input10 (.A(dso_6502[18]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_2 input11 (.A(dso_6502[19]),
    .X(net11));
 sky130_fd_sc_hd__buf_2 input12 (.A(dso_6502[1]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_2 input13 (.A(dso_6502[20]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_2 input14 (.A(dso_6502[21]),
    .X(net14));
 sky130_fd_sc_hd__buf_2 input15 (.A(dso_6502[22]),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_2 input16 (.A(dso_6502[23]),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_2 input17 (.A(dso_6502[24]),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_2 input18 (.A(dso_6502[25]),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_2 input19 (.A(dso_6502[26]),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_2 input20 (.A(dso_6502[2]),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_4 input21 (.A(dso_6502[3]),
    .X(net21));
 sky130_fd_sc_hd__buf_2 input22 (.A(dso_6502[4]),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_4 input23 (.A(dso_6502[5]),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_4 input24 (.A(dso_6502[6]),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_2 input25 (.A(dso_6502[7]),
    .X(net25));
 sky130_fd_sc_hd__buf_4 input26 (.A(dso_6502[8]),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_4 input27 (.A(dso_6502[9]),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_2 input28 (.A(dso_LCD[0]),
    .X(net28));
 sky130_fd_sc_hd__clkbuf_2 input29 (.A(dso_LCD[1]),
    .X(net29));
 sky130_fd_sc_hd__clkbuf_2 input30 (.A(dso_LCD[2]),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_2 input31 (.A(dso_LCD[3]),
    .X(net31));
 sky130_fd_sc_hd__buf_2 input32 (.A(dso_LCD[4]),
    .X(net32));
 sky130_fd_sc_hd__clkbuf_4 input33 (.A(dso_LCD[5]),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_4 input34 (.A(dso_LCD[6]),
    .X(net34));
 sky130_fd_sc_hd__buf_4 input35 (.A(dso_LCD[7]),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_2 input36 (.A(dso_as1802[0]),
    .X(net36));
 sky130_fd_sc_hd__clkbuf_4 input37 (.A(dso_as1802[10]),
    .X(net37));
 sky130_fd_sc_hd__clkbuf_4 input38 (.A(dso_as1802[11]),
    .X(net38));
 sky130_fd_sc_hd__clkbuf_2 input39 (.A(dso_as1802[12]),
    .X(net39));
 sky130_fd_sc_hd__clkbuf_2 input40 (.A(dso_as1802[13]),
    .X(net40));
 sky130_fd_sc_hd__buf_2 input41 (.A(dso_as1802[14]),
    .X(net41));
 sky130_fd_sc_hd__clkbuf_4 input42 (.A(dso_as1802[15]),
    .X(net42));
 sky130_fd_sc_hd__buf_2 input43 (.A(dso_as1802[16]),
    .X(net43));
 sky130_fd_sc_hd__clkbuf_2 input44 (.A(dso_as1802[17]),
    .X(net44));
 sky130_fd_sc_hd__buf_2 input45 (.A(dso_as1802[18]),
    .X(net45));
 sky130_fd_sc_hd__clkbuf_2 input46 (.A(dso_as1802[19]),
    .X(net46));
 sky130_fd_sc_hd__buf_2 input47 (.A(dso_as1802[1]),
    .X(net47));
 sky130_fd_sc_hd__buf_2 input48 (.A(dso_as1802[20]),
    .X(net48));
 sky130_fd_sc_hd__clkbuf_2 input49 (.A(dso_as1802[21]),
    .X(net49));
 sky130_fd_sc_hd__buf_2 input50 (.A(dso_as1802[22]),
    .X(net50));
 sky130_fd_sc_hd__clkbuf_2 input51 (.A(dso_as1802[23]),
    .X(net51));
 sky130_fd_sc_hd__clkbuf_2 input52 (.A(dso_as1802[24]),
    .X(net52));
 sky130_fd_sc_hd__clkbuf_2 input53 (.A(dso_as1802[25]),
    .X(net53));
 sky130_fd_sc_hd__clkbuf_2 input54 (.A(dso_as1802[26]),
    .X(net54));
 sky130_fd_sc_hd__clkbuf_2 input55 (.A(dso_as1802[2]),
    .X(net55));
 sky130_fd_sc_hd__clkbuf_2 input56 (.A(dso_as1802[3]),
    .X(net56));
 sky130_fd_sc_hd__buf_2 input57 (.A(dso_as1802[4]),
    .X(net57));
 sky130_fd_sc_hd__clkbuf_4 input58 (.A(dso_as1802[5]),
    .X(net58));
 sky130_fd_sc_hd__buf_4 input59 (.A(dso_as1802[6]),
    .X(net59));
 sky130_fd_sc_hd__buf_2 input60 (.A(dso_as1802[7]),
    .X(net60));
 sky130_fd_sc_hd__clkbuf_4 input61 (.A(dso_as1802[8]),
    .X(net61));
 sky130_fd_sc_hd__clkbuf_4 input62 (.A(dso_as1802[9]),
    .X(net62));
 sky130_fd_sc_hd__buf_4 input63 (.A(dso_as2650[0]),
    .X(net63));
 sky130_fd_sc_hd__clkbuf_2 input64 (.A(dso_as2650[10]),
    .X(net64));
 sky130_fd_sc_hd__clkbuf_2 input65 (.A(dso_as2650[11]),
    .X(net65));
 sky130_fd_sc_hd__clkbuf_2 input66 (.A(dso_as2650[12]),
    .X(net66));
 sky130_fd_sc_hd__clkbuf_2 input67 (.A(dso_as2650[13]),
    .X(net67));
 sky130_fd_sc_hd__clkbuf_2 input68 (.A(dso_as2650[14]),
    .X(net68));
 sky130_fd_sc_hd__clkbuf_2 input69 (.A(dso_as2650[15]),
    .X(net69));
 sky130_fd_sc_hd__clkbuf_2 input70 (.A(dso_as2650[16]),
    .X(net70));
 sky130_fd_sc_hd__clkbuf_4 input71 (.A(dso_as2650[17]),
    .X(net71));
 sky130_fd_sc_hd__buf_2 input72 (.A(dso_as2650[18]),
    .X(net72));
 sky130_fd_sc_hd__clkbuf_4 input73 (.A(dso_as2650[19]),
    .X(net73));
 sky130_fd_sc_hd__clkbuf_4 input74 (.A(dso_as2650[1]),
    .X(net74));
 sky130_fd_sc_hd__buf_2 input75 (.A(dso_as2650[20]),
    .X(net75));
 sky130_fd_sc_hd__clkbuf_4 input76 (.A(dso_as2650[21]),
    .X(net76));
 sky130_fd_sc_hd__buf_2 input77 (.A(dso_as2650[22]),
    .X(net77));
 sky130_fd_sc_hd__buf_2 input78 (.A(dso_as2650[23]),
    .X(net78));
 sky130_fd_sc_hd__clkbuf_2 input79 (.A(dso_as2650[24]),
    .X(net79));
 sky130_fd_sc_hd__clkbuf_2 input80 (.A(dso_as2650[25]),
    .X(net80));
 sky130_fd_sc_hd__buf_2 input81 (.A(dso_as2650[26]),
    .X(net81));
 sky130_fd_sc_hd__clkbuf_2 input82 (.A(dso_as2650[2]),
    .X(net82));
 sky130_fd_sc_hd__clkbuf_2 input83 (.A(dso_as2650[3]),
    .X(net83));
 sky130_fd_sc_hd__clkbuf_2 input84 (.A(dso_as2650[4]),
    .X(net84));
 sky130_fd_sc_hd__clkbuf_2 input85 (.A(dso_as2650[5]),
    .X(net85));
 sky130_fd_sc_hd__clkbuf_2 input86 (.A(dso_as2650[6]),
    .X(net86));
 sky130_fd_sc_hd__clkbuf_2 input87 (.A(dso_as2650[7]),
    .X(net87));
 sky130_fd_sc_hd__clkbuf_2 input88 (.A(dso_as2650[8]),
    .X(net88));
 sky130_fd_sc_hd__clkbuf_2 input89 (.A(dso_as2650[9]),
    .X(net89));
 sky130_fd_sc_hd__clkbuf_4 input90 (.A(dso_as512512512[0]),
    .X(net90));
 sky130_fd_sc_hd__clkbuf_2 input91 (.A(dso_as512512512[10]),
    .X(net91));
 sky130_fd_sc_hd__clkbuf_2 input92 (.A(dso_as512512512[11]),
    .X(net92));
 sky130_fd_sc_hd__clkbuf_2 input93 (.A(dso_as512512512[12]),
    .X(net93));
 sky130_fd_sc_hd__clkbuf_2 input94 (.A(dso_as512512512[13]),
    .X(net94));
 sky130_fd_sc_hd__clkbuf_2 input95 (.A(dso_as512512512[14]),
    .X(net95));
 sky130_fd_sc_hd__buf_2 input96 (.A(dso_as512512512[15]),
    .X(net96));
 sky130_fd_sc_hd__buf_2 input97 (.A(dso_as512512512[16]),
    .X(net97));
 sky130_fd_sc_hd__clkbuf_4 input98 (.A(dso_as512512512[17]),
    .X(net98));
 sky130_fd_sc_hd__buf_2 input99 (.A(dso_as512512512[18]),
    .X(net99));
 sky130_fd_sc_hd__clkbuf_4 input100 (.A(dso_as512512512[19]),
    .X(net100));
 sky130_fd_sc_hd__buf_2 input101 (.A(dso_as512512512[1]),
    .X(net101));
 sky130_fd_sc_hd__clkbuf_2 input102 (.A(dso_as512512512[20]),
    .X(net102));
 sky130_fd_sc_hd__clkbuf_4 input103 (.A(dso_as512512512[21]),
    .X(net103));
 sky130_fd_sc_hd__buf_2 input104 (.A(dso_as512512512[22]),
    .X(net104));
 sky130_fd_sc_hd__clkbuf_4 input105 (.A(dso_as512512512[23]),
    .X(net105));
 sky130_fd_sc_hd__buf_2 input106 (.A(dso_as512512512[24]),
    .X(net106));
 sky130_fd_sc_hd__buf_2 input107 (.A(dso_as512512512[25]),
    .X(net107));
 sky130_fd_sc_hd__clkbuf_4 input108 (.A(dso_as512512512[26]),
    .X(net108));
 sky130_fd_sc_hd__clkbuf_4 input109 (.A(dso_as512512512[27]),
    .X(net109));
 sky130_fd_sc_hd__clkbuf_2 input110 (.A(dso_as512512512[2]),
    .X(net110));
 sky130_fd_sc_hd__clkbuf_2 input111 (.A(dso_as512512512[3]),
    .X(net111));
 sky130_fd_sc_hd__buf_2 input112 (.A(dso_as512512512[4]),
    .X(net112));
 sky130_fd_sc_hd__clkbuf_2 input113 (.A(dso_as512512512[5]),
    .X(net113));
 sky130_fd_sc_hd__clkbuf_2 input114 (.A(dso_as512512512[6]),
    .X(net114));
 sky130_fd_sc_hd__clkbuf_2 input115 (.A(dso_as512512512[7]),
    .X(net115));
 sky130_fd_sc_hd__clkbuf_2 input116 (.A(dso_as512512512[8]),
    .X(net116));
 sky130_fd_sc_hd__clkbuf_2 input117 (.A(dso_as512512512[9]),
    .X(net117));
 sky130_fd_sc_hd__buf_2 input118 (.A(dso_as5401[0]),
    .X(net118));
 sky130_fd_sc_hd__clkbuf_2 input119 (.A(dso_as5401[10]),
    .X(net119));
 sky130_fd_sc_hd__buf_2 input120 (.A(dso_as5401[11]),
    .X(net120));
 sky130_fd_sc_hd__clkbuf_4 input121 (.A(dso_as5401[12]),
    .X(net121));
 sky130_fd_sc_hd__clkbuf_2 input122 (.A(dso_as5401[13]),
    .X(net122));
 sky130_fd_sc_hd__clkbuf_2 input123 (.A(dso_as5401[14]),
    .X(net123));
 sky130_fd_sc_hd__clkbuf_2 input124 (.A(dso_as5401[15]),
    .X(net124));
 sky130_fd_sc_hd__clkbuf_2 input125 (.A(dso_as5401[16]),
    .X(net125));
 sky130_fd_sc_hd__clkbuf_2 input126 (.A(dso_as5401[17]),
    .X(net126));
 sky130_fd_sc_hd__clkbuf_2 input127 (.A(dso_as5401[18]),
    .X(net127));
 sky130_fd_sc_hd__clkbuf_2 input128 (.A(dso_as5401[19]),
    .X(net128));
 sky130_fd_sc_hd__clkbuf_2 input129 (.A(dso_as5401[1]),
    .X(net129));
 sky130_fd_sc_hd__clkbuf_2 input130 (.A(dso_as5401[20]),
    .X(net130));
 sky130_fd_sc_hd__clkbuf_2 input131 (.A(dso_as5401[21]),
    .X(net131));
 sky130_fd_sc_hd__buf_2 input132 (.A(dso_as5401[22]),
    .X(net132));
 sky130_fd_sc_hd__clkbuf_2 input133 (.A(dso_as5401[23]),
    .X(net133));
 sky130_fd_sc_hd__clkbuf_4 input134 (.A(dso_as5401[24]),
    .X(net134));
 sky130_fd_sc_hd__clkbuf_4 input135 (.A(dso_as5401[25]),
    .X(net135));
 sky130_fd_sc_hd__clkbuf_2 input136 (.A(dso_as5401[26]),
    .X(net136));
 sky130_fd_sc_hd__clkbuf_4 input137 (.A(dso_as5401[2]),
    .X(net137));
 sky130_fd_sc_hd__clkbuf_4 input138 (.A(dso_as5401[3]),
    .X(net138));
 sky130_fd_sc_hd__clkbuf_2 input139 (.A(dso_as5401[4]),
    .X(net139));
 sky130_fd_sc_hd__clkbuf_2 input140 (.A(dso_as5401[5]),
    .X(net140));
 sky130_fd_sc_hd__clkbuf_2 input141 (.A(dso_as5401[6]),
    .X(net141));
 sky130_fd_sc_hd__clkbuf_2 input142 (.A(dso_as5401[7]),
    .X(net142));
 sky130_fd_sc_hd__clkbuf_2 input143 (.A(dso_as5401[8]),
    .X(net143));
 sky130_fd_sc_hd__buf_2 input144 (.A(dso_as5401[9]),
    .X(net144));
 sky130_fd_sc_hd__clkbuf_2 input145 (.A(dso_counter[0]),
    .X(net145));
 sky130_fd_sc_hd__buf_4 input146 (.A(dso_counter[10]),
    .X(net146));
 sky130_fd_sc_hd__clkbuf_4 input147 (.A(dso_counter[11]),
    .X(net147));
 sky130_fd_sc_hd__clkbuf_2 input148 (.A(dso_counter[1]),
    .X(net148));
 sky130_fd_sc_hd__clkbuf_2 input149 (.A(dso_counter[2]),
    .X(net149));
 sky130_fd_sc_hd__clkbuf_2 input150 (.A(dso_counter[3]),
    .X(net150));
 sky130_fd_sc_hd__buf_2 input151 (.A(dso_counter[4]),
    .X(net151));
 sky130_fd_sc_hd__clkbuf_2 input152 (.A(dso_counter[5]),
    .X(net152));
 sky130_fd_sc_hd__clkbuf_4 input153 (.A(dso_counter[6]),
    .X(net153));
 sky130_fd_sc_hd__clkbuf_2 input154 (.A(dso_counter[7]),
    .X(net154));
 sky130_fd_sc_hd__buf_4 input155 (.A(dso_counter[8]),
    .X(net155));
 sky130_fd_sc_hd__clkbuf_4 input156 (.A(dso_counter[9]),
    .X(net156));
 sky130_fd_sc_hd__clkbuf_4 input157 (.A(dso_diceroll[0]),
    .X(net157));
 sky130_fd_sc_hd__buf_4 input158 (.A(dso_diceroll[1]),
    .X(net158));
 sky130_fd_sc_hd__clkbuf_2 input159 (.A(dso_diceroll[2]),
    .X(net159));
 sky130_fd_sc_hd__clkbuf_2 input160 (.A(dso_diceroll[3]),
    .X(net160));
 sky130_fd_sc_hd__clkbuf_2 input161 (.A(dso_diceroll[4]),
    .X(net161));
 sky130_fd_sc_hd__clkbuf_2 input162 (.A(dso_diceroll[5]),
    .X(net162));
 sky130_fd_sc_hd__clkbuf_2 input163 (.A(dso_diceroll[6]),
    .X(net163));
 sky130_fd_sc_hd__clkbuf_2 input164 (.A(dso_diceroll[7]),
    .X(net164));
 sky130_fd_sc_hd__clkbuf_2 input165 (.A(dso_mc14500[0]),
    .X(net165));
 sky130_fd_sc_hd__clkbuf_2 input166 (.A(dso_mc14500[1]),
    .X(net166));
 sky130_fd_sc_hd__clkbuf_2 input167 (.A(dso_mc14500[2]),
    .X(net167));
 sky130_fd_sc_hd__clkbuf_2 input168 (.A(dso_mc14500[3]),
    .X(net168));
 sky130_fd_sc_hd__clkbuf_2 input169 (.A(dso_mc14500[4]),
    .X(net169));
 sky130_fd_sc_hd__clkbuf_2 input170 (.A(dso_mc14500[5]),
    .X(net170));
 sky130_fd_sc_hd__clkbuf_2 input171 (.A(dso_mc14500[6]),
    .X(net171));
 sky130_fd_sc_hd__clkbuf_2 input172 (.A(dso_mc14500[7]),
    .X(net172));
 sky130_fd_sc_hd__clkbuf_2 input173 (.A(dso_mc14500[8]),
    .X(net173));
 sky130_fd_sc_hd__clkbuf_2 input174 (.A(dso_multiplier[0]),
    .X(net174));
 sky130_fd_sc_hd__clkbuf_2 input175 (.A(dso_multiplier[1]),
    .X(net175));
 sky130_fd_sc_hd__clkbuf_2 input176 (.A(dso_multiplier[2]),
    .X(net176));
 sky130_fd_sc_hd__clkbuf_2 input177 (.A(dso_multiplier[3]),
    .X(net177));
 sky130_fd_sc_hd__clkbuf_2 input178 (.A(dso_multiplier[4]),
    .X(net178));
 sky130_fd_sc_hd__clkbuf_2 input179 (.A(dso_multiplier[5]),
    .X(net179));
 sky130_fd_sc_hd__clkbuf_2 input180 (.A(dso_multiplier[6]),
    .X(net180));
 sky130_fd_sc_hd__clkbuf_2 input181 (.A(dso_multiplier[7]),
    .X(net181));
 sky130_fd_sc_hd__clkbuf_2 input182 (.A(dso_posit[0]),
    .X(net182));
 sky130_fd_sc_hd__clkbuf_2 input183 (.A(dso_posit[1]),
    .X(net183));
 sky130_fd_sc_hd__clkbuf_2 input184 (.A(dso_posit[2]),
    .X(net184));
 sky130_fd_sc_hd__clkbuf_2 input185 (.A(dso_posit[3]),
    .X(net185));
 sky130_fd_sc_hd__clkbuf_2 input186 (.A(dso_tbb1143[0]),
    .X(net186));
 sky130_fd_sc_hd__clkbuf_2 input187 (.A(dso_tbb1143[1]),
    .X(net187));
 sky130_fd_sc_hd__clkbuf_2 input188 (.A(dso_tbb1143[2]),
    .X(net188));
 sky130_fd_sc_hd__clkbuf_2 input189 (.A(dso_tbb1143[3]),
    .X(net189));
 sky130_fd_sc_hd__clkbuf_2 input190 (.A(dso_tbb1143[4]),
    .X(net190));
 sky130_fd_sc_hd__clkbuf_2 input191 (.A(dso_tbb1143[5]),
    .X(net191));
 sky130_fd_sc_hd__clkbuf_2 input192 (.A(dso_tbb1143[6]),
    .X(net192));
 sky130_fd_sc_hd__clkbuf_2 input193 (.A(dso_tbb1143[7]),
    .X(net193));
 sky130_fd_sc_hd__clkbuf_8 input194 (.A(dso_tune),
    .X(net194));
 sky130_fd_sc_hd__clkbuf_2 input195 (.A(io_in[0]),
    .X(net195));
 sky130_fd_sc_hd__clkbuf_2 input196 (.A(io_in[10]),
    .X(net196));
 sky130_fd_sc_hd__clkbuf_2 input197 (.A(io_in[11]),
    .X(net197));
 sky130_fd_sc_hd__clkbuf_2 input198 (.A(io_in[12]),
    .X(net198));
 sky130_fd_sc_hd__clkbuf_2 input199 (.A(io_in[13]),
    .X(net199));
 sky130_fd_sc_hd__clkbuf_2 input200 (.A(io_in[14]),
    .X(net200));
 sky130_fd_sc_hd__clkbuf_2 input201 (.A(io_in[15]),
    .X(net201));
 sky130_fd_sc_hd__clkbuf_2 input202 (.A(io_in[16]),
    .X(net202));
 sky130_fd_sc_hd__clkbuf_2 input203 (.A(io_in[17]),
    .X(net203));
 sky130_fd_sc_hd__clkbuf_2 input204 (.A(io_in[18]),
    .X(net204));
 sky130_fd_sc_hd__clkbuf_2 input205 (.A(io_in[19]),
    .X(net205));
 sky130_fd_sc_hd__clkbuf_2 input206 (.A(io_in[20]),
    .X(net206));
 sky130_fd_sc_hd__clkbuf_2 input207 (.A(io_in[21]),
    .X(net207));
 sky130_fd_sc_hd__clkbuf_2 input208 (.A(io_in[22]),
    .X(net208));
 sky130_fd_sc_hd__clkbuf_2 input209 (.A(io_in[23]),
    .X(net209));
 sky130_fd_sc_hd__clkbuf_2 input210 (.A(io_in[24]),
    .X(net210));
 sky130_fd_sc_hd__clkbuf_2 input211 (.A(io_in[25]),
    .X(net211));
 sky130_fd_sc_hd__clkbuf_2 input212 (.A(io_in[26]),
    .X(net212));
 sky130_fd_sc_hd__clkbuf_2 input213 (.A(io_in[27]),
    .X(net213));
 sky130_fd_sc_hd__clkbuf_2 input214 (.A(io_in[28]),
    .X(net214));
 sky130_fd_sc_hd__clkbuf_2 input215 (.A(io_in[29]),
    .X(net215));
 sky130_fd_sc_hd__clkbuf_2 input216 (.A(io_in[30]),
    .X(net216));
 sky130_fd_sc_hd__clkbuf_2 input217 (.A(io_in[31]),
    .X(net217));
 sky130_fd_sc_hd__clkbuf_2 input218 (.A(io_in[32]),
    .X(net218));
 sky130_fd_sc_hd__clkbuf_2 input219 (.A(io_in[33]),
    .X(net219));
 sky130_fd_sc_hd__clkbuf_2 input220 (.A(io_in[34]),
    .X(net220));
 sky130_fd_sc_hd__clkbuf_2 input221 (.A(io_in[35]),
    .X(net221));
 sky130_fd_sc_hd__clkbuf_2 input222 (.A(io_in[36]),
    .X(net222));
 sky130_fd_sc_hd__clkbuf_2 input223 (.A(io_in[37]),
    .X(net223));
 sky130_fd_sc_hd__clkbuf_2 input224 (.A(io_in[5]),
    .X(net224));
 sky130_fd_sc_hd__clkbuf_2 input225 (.A(io_in[6]),
    .X(net225));
 sky130_fd_sc_hd__clkbuf_2 input226 (.A(io_in[7]),
    .X(net226));
 sky130_fd_sc_hd__clkbuf_2 input227 (.A(io_in[8]),
    .X(net227));
 sky130_fd_sc_hd__clkbuf_2 input228 (.A(io_in[9]),
    .X(net228));
 sky130_fd_sc_hd__clkbuf_2 input229 (.A(oeb_6502),
    .X(net229));
 sky130_fd_sc_hd__clkbuf_2 input230 (.A(oeb_as1802),
    .X(net230));
 sky130_fd_sc_hd__clkbuf_4 input231 (.A(oeb_as2650),
    .X(net231));
 sky130_fd_sc_hd__buf_4 input232 (.A(oeb_as512512512),
    .X(net232));
 sky130_fd_sc_hd__buf_4 input233 (.A(oeb_as5401),
    .X(net233));
 sky130_fd_sc_hd__buf_2 input234 (.A(oeb_mc14500),
    .X(net234));
 sky130_fd_sc_hd__clkbuf_2 input235 (.A(wb_rst_i),
    .X(net235));
 sky130_fd_sc_hd__clkbuf_4 input236 (.A(wbs_adr_i[21]),
    .X(net236));
 sky130_fd_sc_hd__clkbuf_2 input237 (.A(wbs_adr_i[22]),
    .X(net237));
 sky130_fd_sc_hd__buf_4 input238 (.A(wbs_adr_i[23]),
    .X(net238));
 sky130_fd_sc_hd__clkbuf_2 input239 (.A(wbs_cyc_i),
    .X(net239));
 sky130_fd_sc_hd__buf_2 input240 (.A(wbs_dat_i[0]),
    .X(net240));
 sky130_fd_sc_hd__clkbuf_4 input241 (.A(wbs_dat_i[10]),
    .X(net241));
 sky130_fd_sc_hd__buf_2 input242 (.A(wbs_dat_i[11]),
    .X(net242));
 sky130_fd_sc_hd__buf_2 input243 (.A(wbs_dat_i[12]),
    .X(net243));
 sky130_fd_sc_hd__buf_2 input244 (.A(wbs_dat_i[13]),
    .X(net244));
 sky130_fd_sc_hd__clkbuf_4 input245 (.A(wbs_dat_i[14]),
    .X(net245));
 sky130_fd_sc_hd__clkbuf_4 input246 (.A(wbs_dat_i[15]),
    .X(net246));
 sky130_fd_sc_hd__clkbuf_4 input247 (.A(wbs_dat_i[16]),
    .X(net247));
 sky130_fd_sc_hd__clkbuf_4 input248 (.A(wbs_dat_i[17]),
    .X(net248));
 sky130_fd_sc_hd__clkbuf_4 input249 (.A(wbs_dat_i[18]),
    .X(net249));
 sky130_fd_sc_hd__clkbuf_4 input250 (.A(wbs_dat_i[19]),
    .X(net250));
 sky130_fd_sc_hd__clkbuf_4 input251 (.A(wbs_dat_i[1]),
    .X(net251));
 sky130_fd_sc_hd__buf_4 input252 (.A(wbs_dat_i[20]),
    .X(net252));
 sky130_fd_sc_hd__clkbuf_4 input253 (.A(wbs_dat_i[21]),
    .X(net253));
 sky130_fd_sc_hd__clkbuf_4 input254 (.A(wbs_dat_i[22]),
    .X(net254));
 sky130_fd_sc_hd__buf_4 input255 (.A(wbs_dat_i[23]),
    .X(net255));
 sky130_fd_sc_hd__clkbuf_4 input256 (.A(wbs_dat_i[24]),
    .X(net256));
 sky130_fd_sc_hd__clkbuf_4 input257 (.A(wbs_dat_i[25]),
    .X(net257));
 sky130_fd_sc_hd__clkbuf_4 input258 (.A(wbs_dat_i[26]),
    .X(net258));
 sky130_fd_sc_hd__clkbuf_4 input259 (.A(wbs_dat_i[27]),
    .X(net259));
 sky130_fd_sc_hd__clkbuf_4 input260 (.A(wbs_dat_i[2]),
    .X(net260));
 sky130_fd_sc_hd__clkbuf_4 input261 (.A(wbs_dat_i[3]),
    .X(net261));
 sky130_fd_sc_hd__clkbuf_4 input262 (.A(wbs_dat_i[4]),
    .X(net262));
 sky130_fd_sc_hd__clkbuf_4 input263 (.A(wbs_dat_i[5]),
    .X(net263));
 sky130_fd_sc_hd__clkbuf_4 input264 (.A(wbs_dat_i[6]),
    .X(net264));
 sky130_fd_sc_hd__clkbuf_4 input265 (.A(wbs_dat_i[7]),
    .X(net265));
 sky130_fd_sc_hd__clkbuf_4 input266 (.A(wbs_dat_i[8]),
    .X(net266));
 sky130_fd_sc_hd__clkbuf_4 input267 (.A(wbs_dat_i[9]),
    .X(net267));
 sky130_fd_sc_hd__clkbuf_2 input268 (.A(wbs_stb_i),
    .X(net268));
 sky130_fd_sc_hd__buf_2 input269 (.A(wbs_we_i),
    .X(net269));
 sky130_fd_sc_hd__clkbuf_2 output270 (.A(net270),
    .X(design_clk_o));
 sky130_fd_sc_hd__buf_4 output271 (.A(net271),
    .X(dsi_all[0]));
 sky130_fd_sc_hd__buf_4 output272 (.A(net272),
    .X(dsi_all[10]));
 sky130_fd_sc_hd__buf_4 output273 (.A(net273),
    .X(dsi_all[11]));
 sky130_fd_sc_hd__buf_4 output274 (.A(net274),
    .X(dsi_all[12]));
 sky130_fd_sc_hd__buf_4 output275 (.A(net275),
    .X(dsi_all[13]));
 sky130_fd_sc_hd__buf_4 output276 (.A(net276),
    .X(dsi_all[14]));
 sky130_fd_sc_hd__buf_4 output277 (.A(net277),
    .X(dsi_all[15]));
 sky130_fd_sc_hd__buf_4 output278 (.A(net278),
    .X(dsi_all[16]));
 sky130_fd_sc_hd__buf_4 output279 (.A(net279),
    .X(dsi_all[17]));
 sky130_fd_sc_hd__buf_4 output280 (.A(net280),
    .X(dsi_all[18]));
 sky130_fd_sc_hd__buf_4 output281 (.A(net281),
    .X(dsi_all[19]));
 sky130_fd_sc_hd__buf_4 output282 (.A(net282),
    .X(dsi_all[1]));
 sky130_fd_sc_hd__buf_4 output283 (.A(net283),
    .X(dsi_all[20]));
 sky130_fd_sc_hd__buf_4 output284 (.A(net284),
    .X(dsi_all[21]));
 sky130_fd_sc_hd__buf_4 output285 (.A(net285),
    .X(dsi_all[22]));
 sky130_fd_sc_hd__buf_4 output286 (.A(net286),
    .X(dsi_all[23]));
 sky130_fd_sc_hd__buf_4 output287 (.A(net287),
    .X(dsi_all[24]));
 sky130_fd_sc_hd__buf_4 output288 (.A(net288),
    .X(dsi_all[25]));
 sky130_fd_sc_hd__buf_4 output289 (.A(net289),
    .X(dsi_all[26]));
 sky130_fd_sc_hd__buf_4 output290 (.A(net290),
    .X(dsi_all[27]));
 sky130_fd_sc_hd__buf_4 output291 (.A(net291),
    .X(dsi_all[2]));
 sky130_fd_sc_hd__buf_4 output292 (.A(net292),
    .X(dsi_all[3]));
 sky130_fd_sc_hd__buf_4 output293 (.A(net293),
    .X(dsi_all[4]));
 sky130_fd_sc_hd__buf_4 output294 (.A(net294),
    .X(dsi_all[5]));
 sky130_fd_sc_hd__buf_4 output295 (.A(net295),
    .X(dsi_all[6]));
 sky130_fd_sc_hd__buf_4 output296 (.A(net296),
    .X(dsi_all[7]));
 sky130_fd_sc_hd__buf_4 output297 (.A(net297),
    .X(dsi_all[8]));
 sky130_fd_sc_hd__buf_4 output298 (.A(net298),
    .X(dsi_all[9]));
 sky130_fd_sc_hd__buf_4 output299 (.A(net299),
    .X(io_oeb[0]));
 sky130_fd_sc_hd__buf_4 output300 (.A(net300),
    .X(io_oeb[11]));
 sky130_fd_sc_hd__buf_4 output301 (.A(net301),
    .X(io_oeb[12]));
 sky130_fd_sc_hd__buf_4 output302 (.A(net302),
    .X(io_oeb[13]));
 sky130_fd_sc_hd__buf_4 output303 (.A(net303),
    .X(io_oeb[14]));
 sky130_fd_sc_hd__buf_4 output304 (.A(net304),
    .X(io_oeb[15]));
 sky130_fd_sc_hd__buf_4 output305 (.A(net305),
    .X(io_oeb[16]));
 sky130_fd_sc_hd__buf_4 output306 (.A(net306),
    .X(io_oeb[17]));
 sky130_fd_sc_hd__buf_4 output307 (.A(net307),
    .X(io_oeb[18]));
 sky130_fd_sc_hd__buf_4 output308 (.A(net308),
    .X(io_oeb[19]));
 sky130_fd_sc_hd__buf_4 output309 (.A(net309),
    .X(io_oeb[20]));
 sky130_fd_sc_hd__buf_4 output310 (.A(net310),
    .X(io_oeb[21]));
 sky130_fd_sc_hd__buf_4 output311 (.A(net311),
    .X(io_oeb[22]));
 sky130_fd_sc_hd__buf_4 output312 (.A(net312),
    .X(io_oeb[23]));
 sky130_fd_sc_hd__buf_4 output313 (.A(net313),
    .X(io_oeb[24]));
 sky130_fd_sc_hd__buf_4 output314 (.A(net314),
    .X(io_oeb[25]));
 sky130_fd_sc_hd__buf_4 output315 (.A(net315),
    .X(io_oeb[26]));
 sky130_fd_sc_hd__buf_4 output316 (.A(net316),
    .X(io_oeb[27]));
 sky130_fd_sc_hd__buf_4 output317 (.A(net317),
    .X(io_oeb[28]));
 sky130_fd_sc_hd__buf_4 output318 (.A(net318),
    .X(io_oeb[29]));
 sky130_fd_sc_hd__buf_4 output319 (.A(net319),
    .X(io_oeb[30]));
 sky130_fd_sc_hd__buf_4 output320 (.A(net320),
    .X(io_oeb[31]));
 sky130_fd_sc_hd__buf_4 output321 (.A(net321),
    .X(io_oeb[32]));
 sky130_fd_sc_hd__buf_4 output322 (.A(net322),
    .X(io_oeb[33]));
 sky130_fd_sc_hd__buf_4 output323 (.A(net323),
    .X(io_oeb[34]));
 sky130_fd_sc_hd__buf_4 output324 (.A(net324),
    .X(io_oeb[35]));
 sky130_fd_sc_hd__buf_4 output325 (.A(net416),
    .X(io_oeb[36]));
 sky130_fd_sc_hd__buf_4 output326 (.A(net326),
    .X(io_oeb[37]));
 sky130_fd_sc_hd__buf_4 output327 (.A(net327),
    .X(io_out[0]));
 sky130_fd_sc_hd__buf_4 output328 (.A(net328),
    .X(io_out[11]));
 sky130_fd_sc_hd__buf_4 output329 (.A(net329),
    .X(io_out[12]));
 sky130_fd_sc_hd__buf_4 output330 (.A(net330),
    .X(io_out[13]));
 sky130_fd_sc_hd__buf_4 output331 (.A(net331),
    .X(io_out[14]));
 sky130_fd_sc_hd__buf_4 output332 (.A(net332),
    .X(io_out[15]));
 sky130_fd_sc_hd__buf_4 output333 (.A(net333),
    .X(io_out[16]));
 sky130_fd_sc_hd__buf_4 output334 (.A(net334),
    .X(io_out[17]));
 sky130_fd_sc_hd__buf_4 output335 (.A(net335),
    .X(io_out[18]));
 sky130_fd_sc_hd__buf_4 output336 (.A(net336),
    .X(io_out[19]));
 sky130_fd_sc_hd__buf_4 output337 (.A(net337),
    .X(io_out[1]));
 sky130_fd_sc_hd__buf_4 output338 (.A(net338),
    .X(io_out[20]));
 sky130_fd_sc_hd__buf_4 output339 (.A(net339),
    .X(io_out[21]));
 sky130_fd_sc_hd__buf_4 output340 (.A(net340),
    .X(io_out[22]));
 sky130_fd_sc_hd__buf_4 output341 (.A(net341),
    .X(io_out[23]));
 sky130_fd_sc_hd__buf_4 output342 (.A(net342),
    .X(io_out[24]));
 sky130_fd_sc_hd__buf_4 output343 (.A(net343),
    .X(io_out[25]));
 sky130_fd_sc_hd__buf_4 output344 (.A(net344),
    .X(io_out[26]));
 sky130_fd_sc_hd__buf_4 output345 (.A(net345),
    .X(io_out[27]));
 sky130_fd_sc_hd__buf_4 output346 (.A(net346),
    .X(io_out[28]));
 sky130_fd_sc_hd__buf_4 output347 (.A(net347),
    .X(io_out[29]));
 sky130_fd_sc_hd__buf_4 output348 (.A(net348),
    .X(io_out[2]));
 sky130_fd_sc_hd__buf_4 output349 (.A(net349),
    .X(io_out[30]));
 sky130_fd_sc_hd__buf_4 output350 (.A(net350),
    .X(io_out[31]));
 sky130_fd_sc_hd__buf_4 output351 (.A(net351),
    .X(io_out[32]));
 sky130_fd_sc_hd__buf_4 output352 (.A(net352),
    .X(io_out[33]));
 sky130_fd_sc_hd__buf_4 output353 (.A(net353),
    .X(io_out[34]));
 sky130_fd_sc_hd__buf_4 output354 (.A(net354),
    .X(io_out[35]));
 sky130_fd_sc_hd__buf_4 output355 (.A(net355),
    .X(io_out[36]));
 sky130_fd_sc_hd__buf_4 output356 (.A(net356),
    .X(io_out[37]));
 sky130_fd_sc_hd__buf_4 output357 (.A(net357),
    .X(io_out[3]));
 sky130_fd_sc_hd__buf_4 output358 (.A(net358),
    .X(io_out[4]));
 sky130_fd_sc_hd__buf_4 output359 (.A(net359),
    .X(rst_6502));
 sky130_fd_sc_hd__buf_4 output360 (.A(net360),
    .X(rst_LCD));
 sky130_fd_sc_hd__buf_4 output361 (.A(net361),
    .X(rst_as1802));
 sky130_fd_sc_hd__buf_4 output362 (.A(net362),
    .X(rst_as2650));
 sky130_fd_sc_hd__buf_4 output363 (.A(net363),
    .X(rst_as512512512));
 sky130_fd_sc_hd__buf_4 output364 (.A(net364),
    .X(rst_as5401));
 sky130_fd_sc_hd__buf_4 output365 (.A(net365),
    .X(rst_counter));
 sky130_fd_sc_hd__buf_4 output366 (.A(net366),
    .X(rst_diceroll));
 sky130_fd_sc_hd__buf_4 output367 (.A(net367),
    .X(rst_mc14500));
 sky130_fd_sc_hd__buf_4 output368 (.A(net368),
    .X(rst_posit));
 sky130_fd_sc_hd__buf_4 output369 (.A(net369),
    .X(rst_tbb1143));
 sky130_fd_sc_hd__buf_4 output370 (.A(net370),
    .X(rst_tune));
 sky130_fd_sc_hd__buf_4 output371 (.A(net371),
    .X(wbs_ack_o));
 sky130_fd_sc_hd__buf_4 output372 (.A(net372),
    .X(wbs_dat_o[0]));
 sky130_fd_sc_hd__buf_4 output373 (.A(net373),
    .X(wbs_dat_o[10]));
 sky130_fd_sc_hd__buf_4 output374 (.A(net374),
    .X(wbs_dat_o[11]));
 sky130_fd_sc_hd__buf_4 output375 (.A(net375),
    .X(wbs_dat_o[12]));
 sky130_fd_sc_hd__buf_4 output376 (.A(net376),
    .X(wbs_dat_o[13]));
 sky130_fd_sc_hd__buf_4 output377 (.A(net377),
    .X(wbs_dat_o[14]));
 sky130_fd_sc_hd__buf_4 output378 (.A(net378),
    .X(wbs_dat_o[15]));
 sky130_fd_sc_hd__buf_4 output379 (.A(net379),
    .X(wbs_dat_o[16]));
 sky130_fd_sc_hd__buf_4 output380 (.A(net380),
    .X(wbs_dat_o[17]));
 sky130_fd_sc_hd__buf_4 output381 (.A(net381),
    .X(wbs_dat_o[18]));
 sky130_fd_sc_hd__buf_4 output382 (.A(net382),
    .X(wbs_dat_o[19]));
 sky130_fd_sc_hd__buf_4 output383 (.A(net383),
    .X(wbs_dat_o[1]));
 sky130_fd_sc_hd__buf_4 output384 (.A(net384),
    .X(wbs_dat_o[20]));
 sky130_fd_sc_hd__buf_4 output385 (.A(net385),
    .X(wbs_dat_o[21]));
 sky130_fd_sc_hd__buf_4 output386 (.A(net386),
    .X(wbs_dat_o[22]));
 sky130_fd_sc_hd__buf_4 output387 (.A(net387),
    .X(wbs_dat_o[23]));
 sky130_fd_sc_hd__buf_4 output388 (.A(net388),
    .X(wbs_dat_o[24]));
 sky130_fd_sc_hd__buf_4 output389 (.A(net389),
    .X(wbs_dat_o[25]));
 sky130_fd_sc_hd__buf_4 output390 (.A(net390),
    .X(wbs_dat_o[26]));
 sky130_fd_sc_hd__buf_4 output391 (.A(net391),
    .X(wbs_dat_o[27]));
 sky130_fd_sc_hd__buf_4 output392 (.A(net392),
    .X(wbs_dat_o[2]));
 sky130_fd_sc_hd__buf_4 output393 (.A(net393),
    .X(wbs_dat_o[3]));
 sky130_fd_sc_hd__buf_4 output394 (.A(net394),
    .X(wbs_dat_o[4]));
 sky130_fd_sc_hd__buf_4 output395 (.A(net395),
    .X(wbs_dat_o[5]));
 sky130_fd_sc_hd__buf_4 output396 (.A(net396),
    .X(wbs_dat_o[6]));
 sky130_fd_sc_hd__buf_4 output397 (.A(net397),
    .X(wbs_dat_o[7]));
 sky130_fd_sc_hd__buf_4 output398 (.A(net398),
    .X(wbs_dat_o[8]));
 sky130_fd_sc_hd__buf_4 output399 (.A(net399),
    .X(wbs_dat_o[9]));
 sky130_fd_sc_hd__buf_4 fanout400 (.A(_0421_),
    .X(net400));
 sky130_fd_sc_hd__clkbuf_4 fanout401 (.A(net402),
    .X(net401));
 sky130_fd_sc_hd__buf_4 fanout402 (.A(_0360_),
    .X(net402));
 sky130_fd_sc_hd__buf_4 fanout403 (.A(net404),
    .X(net403));
 sky130_fd_sc_hd__buf_4 fanout404 (.A(_0392_),
    .X(net404));
 sky130_fd_sc_hd__buf_4 fanout405 (.A(net406),
    .X(net405));
 sky130_fd_sc_hd__buf_4 fanout406 (.A(_0392_),
    .X(net406));
 sky130_fd_sc_hd__buf_6 fanout407 (.A(net408),
    .X(net407));
 sky130_fd_sc_hd__clkbuf_4 fanout408 (.A(net409),
    .X(net408));
 sky130_fd_sc_hd__buf_4 fanout409 (.A(net410),
    .X(net409));
 sky130_fd_sc_hd__buf_6 fanout410 (.A(_0386_),
    .X(net410));
 sky130_fd_sc_hd__buf_4 fanout411 (.A(net412),
    .X(net411));
 sky130_fd_sc_hd__buf_4 fanout412 (.A(_0361_),
    .X(net412));
 sky130_fd_sc_hd__buf_4 fanout413 (.A(_0361_),
    .X(net413));
 sky130_fd_sc_hd__buf_8 fanout414 (.A(_0212_),
    .X(net414));
 sky130_fd_sc_hd__buf_4 fanout415 (.A(net325),
    .X(net415));
 sky130_fd_sc_hd__buf_2 fanout416 (.A(net325),
    .X(net416));
 sky130_fd_sc_hd__buf_6 max_cap417 (.A(_0211_),
    .X(net417));
 sky130_fd_sc_hd__buf_8 fanout418 (.A(net419),
    .X(net418));
 sky130_fd_sc_hd__clkbuf_16 fanout419 (.A(net420),
    .X(net419));
 sky130_fd_sc_hd__buf_12 fanout420 (.A(_0202_),
    .X(net420));
 sky130_fd_sc_hd__clkbuf_8 fanout421 (.A(net422),
    .X(net421));
 sky130_fd_sc_hd__buf_6 fanout422 (.A(_0199_),
    .X(net422));
 sky130_fd_sc_hd__buf_6 fanout423 (.A(_0199_),
    .X(net423));
 sky130_fd_sc_hd__buf_2 fanout424 (.A(_0199_),
    .X(net424));
 sky130_fd_sc_hd__buf_6 fanout425 (.A(net426),
    .X(net425));
 sky130_fd_sc_hd__buf_6 fanout426 (.A(_0198_),
    .X(net426));
 sky130_fd_sc_hd__buf_6 fanout427 (.A(_0198_),
    .X(net427));
 sky130_fd_sc_hd__clkbuf_4 fanout428 (.A(_0198_),
    .X(net428));
 sky130_fd_sc_hd__buf_6 fanout429 (.A(_0196_),
    .X(net429));
 sky130_fd_sc_hd__buf_4 fanout430 (.A(_0196_),
    .X(net430));
 sky130_fd_sc_hd__buf_6 fanout431 (.A(_0196_),
    .X(net431));
 sky130_fd_sc_hd__buf_8 fanout432 (.A(_0195_),
    .X(net432));
 sky130_fd_sc_hd__buf_12 fanout433 (.A(_0194_),
    .X(net433));
 sky130_fd_sc_hd__buf_8 fanout434 (.A(_0193_),
    .X(net434));
 sky130_fd_sc_hd__buf_12 fanout435 (.A(_0187_),
    .X(net435));
 sky130_fd_sc_hd__clkbuf_4 fanout436 (.A(_0186_),
    .X(net436));
 sky130_fd_sc_hd__buf_8 fanout437 (.A(net440),
    .X(net437));
 sky130_fd_sc_hd__buf_6 fanout438 (.A(net440),
    .X(net438));
 sky130_fd_sc_hd__buf_4 fanout439 (.A(net440),
    .X(net439));
 sky130_fd_sc_hd__buf_6 fanout440 (.A(_0185_),
    .X(net440));
 sky130_fd_sc_hd__clkbuf_4 fanout441 (.A(net442),
    .X(net441));
 sky130_fd_sc_hd__buf_2 fanout442 (.A(net443),
    .X(net442));
 sky130_fd_sc_hd__buf_2 fanout443 (.A(net444),
    .X(net443));
 sky130_fd_sc_hd__clkbuf_4 fanout444 (.A(net445),
    .X(net444));
 sky130_fd_sc_hd__buf_4 fanout445 (.A(net446),
    .X(net445));
 sky130_fd_sc_hd__buf_4 fanout446 (.A(wb_override),
    .X(net446));
 sky130_fd_sc_hd__clkbuf_4 fanout447 (.A(net448),
    .X(net447));
 sky130_fd_sc_hd__buf_2 fanout448 (.A(wb_override),
    .X(net448));
 sky130_fd_sc_hd__buf_6 fanout449 (.A(net450),
    .X(net449));
 sky130_fd_sc_hd__clkbuf_4 fanout450 (.A(net451),
    .X(net450));
 sky130_fd_sc_hd__buf_4 fanout451 (.A(\design_addr[3] ),
    .X(net451));
 sky130_fd_sc_hd__buf_6 fanout452 (.A(net453),
    .X(net452));
 sky130_fd_sc_hd__clkbuf_4 fanout453 (.A(net454),
    .X(net453));
 sky130_fd_sc_hd__buf_4 fanout454 (.A(\design_addr[2] ),
    .X(net454));
 sky130_fd_sc_hd__clkbuf_8 fanout455 (.A(net457),
    .X(net455));
 sky130_fd_sc_hd__clkbuf_4 fanout456 (.A(net457),
    .X(net456));
 sky130_fd_sc_hd__clkbuf_8 fanout457 (.A(\design_addr[1] ),
    .X(net457));
 sky130_fd_sc_hd__buf_6 fanout458 (.A(net460),
    .X(net458));
 sky130_fd_sc_hd__buf_2 fanout459 (.A(net460),
    .X(net459));
 sky130_fd_sc_hd__buf_4 fanout460 (.A(\design_addr[0] ),
    .X(net460));
 sky130_fd_sc_hd__buf_4 fanout461 (.A(net462),
    .X(net461));
 sky130_fd_sc_hd__buf_6 fanout462 (.A(net467),
    .X(net462));
 sky130_fd_sc_hd__buf_4 fanout463 (.A(net464),
    .X(net463));
 sky130_fd_sc_hd__buf_2 fanout464 (.A(net467),
    .X(net464));
 sky130_fd_sc_hd__buf_4 fanout465 (.A(net466),
    .X(net465));
 sky130_fd_sc_hd__buf_4 fanout466 (.A(net467),
    .X(net466));
 sky130_fd_sc_hd__buf_4 fanout467 (.A(_0182_),
    .X(net467));
 sky130_fd_sc_hd__buf_8 fanout468 (.A(_0181_),
    .X(net468));
 sky130_fd_sc_hd__buf_6 fanout469 (.A(_0181_),
    .X(net469));
 sky130_fd_sc_hd__buf_4 fanout470 (.A(net238),
    .X(net470));
 sky130_fd_sc_hd__clkbuf_8 fanout471 (.A(net472),
    .X(net471));
 sky130_fd_sc_hd__buf_6 fanout472 (.A(net473),
    .X(net472));
 sky130_fd_sc_hd__buf_6 fanout473 (.A(net237),
    .X(net473));
 sky130_fd_sc_hd__buf_6 fanout474 (.A(net476),
    .X(net474));
 sky130_fd_sc_hd__clkbuf_4 fanout475 (.A(net476),
    .X(net475));
 sky130_fd_sc_hd__clkbuf_8 fanout476 (.A(net235),
    .X(net476));
 sky130_fd_sc_hd__conb_1 multiplexer_477 (.LO(net477));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_0__f_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_3_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_1__f_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_3_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_2__f_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_3_2__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_3__f_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_3_3__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_4__f_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_3_4__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_5__f_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_3_5__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_6__f_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_3_6__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_7__f_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_3_7__leaf_wb_clk_i));
 sky130_fd_sc_hd__bufbuf_16 hold1 (.A(net559),
    .X(net497));
 sky130_fd_sc_hd__bufbuf_16 hold2 (.A(_0097_),
    .X(net498));
 sky130_fd_sc_hd__bufbuf_16 hold3 (.A(net560),
    .X(net499));
 sky130_fd_sc_hd__bufbuf_16 hold4 (.A(_0111_),
    .X(net500));
 sky130_fd_sc_hd__bufbuf_16 hold5 (.A(net561),
    .X(net501));
 sky130_fd_sc_hd__bufbuf_16 hold6 (.A(net562),
    .X(net502));
 sky130_fd_sc_hd__bufbuf_16 hold7 (.A(net563),
    .X(net503));
 sky130_fd_sc_hd__bufbuf_16 hold8 (.A(_0103_),
    .X(net504));
 sky130_fd_sc_hd__bufbuf_16 hold9 (.A(net564),
    .X(net505));
 sky130_fd_sc_hd__bufbuf_16 hold10 (.A(_0108_),
    .X(net506));
 sky130_fd_sc_hd__bufbuf_16 hold11 (.A(net565),
    .X(net507));
 sky130_fd_sc_hd__bufbuf_16 hold12 (.A(_0112_),
    .X(net508));
 sky130_fd_sc_hd__bufbuf_16 hold13 (.A(net566),
    .X(net509));
 sky130_fd_sc_hd__bufbuf_16 hold14 (.A(_0091_),
    .X(net510));
 sky130_fd_sc_hd__bufbuf_16 hold15 (.A(net567),
    .X(net511));
 sky130_fd_sc_hd__bufbuf_16 hold16 (.A(_0092_),
    .X(net512));
 sky130_fd_sc_hd__bufbuf_16 hold17 (.A(\wb_counter[8] ),
    .X(net513));
 sky130_fd_sc_hd__bufbuf_16 hold18 (.A(_0175_),
    .X(net514));
 sky130_fd_sc_hd__bufbuf_16 hold19 (.A(_0099_),
    .X(net515));
 sky130_fd_sc_hd__bufbuf_16 hold20 (.A(\wb_counter[23] ),
    .X(net516));
 sky130_fd_sc_hd__bufbuf_16 hold21 (.A(_0172_),
    .X(net517));
 sky130_fd_sc_hd__bufbuf_16 hold22 (.A(_0114_),
    .X(net518));
 sky130_fd_sc_hd__bufbuf_16 hold23 (.A(\wb_counter[14] ),
    .X(net519));
 sky130_fd_sc_hd__bufbuf_16 hold24 (.A(_0173_),
    .X(net520));
 sky130_fd_sc_hd__bufbuf_16 hold25 (.A(_0105_),
    .X(net521));
 sky130_fd_sc_hd__bufbuf_16 hold26 (.A(\wb_counter[10] ),
    .X(net522));
 sky130_fd_sc_hd__bufbuf_16 hold27 (.A(_0155_),
    .X(net523));
 sky130_fd_sc_hd__bufbuf_16 hold28 (.A(_0101_),
    .X(net524));
 sky130_fd_sc_hd__bufbuf_16 hold29 (.A(\wb_counter[9] ),
    .X(net525));
 sky130_fd_sc_hd__bufbuf_16 hold30 (.A(_0153_),
    .X(net526));
 sky130_fd_sc_hd__bufbuf_16 hold31 (.A(_0100_),
    .X(net527));
 sky130_fd_sc_hd__bufbuf_16 hold32 (.A(net569),
    .X(net528));
 sky130_fd_sc_hd__bufbuf_16 hold33 (.A(_0095_),
    .X(net529));
 sky130_fd_sc_hd__bufbuf_16 hold34 (.A(\wb_counter[11] ),
    .X(net530));
 sky130_fd_sc_hd__bufbuf_16 hold35 (.A(_0157_),
    .X(net531));
 sky130_fd_sc_hd__bufbuf_16 hold36 (.A(_0102_),
    .X(net532));
 sky130_fd_sc_hd__bufbuf_16 hold37 (.A(\wb_counter[7] ),
    .X(net533));
 sky130_fd_sc_hd__bufbuf_16 hold38 (.A(_0150_),
    .X(net534));
 sky130_fd_sc_hd__bufbuf_16 hold39 (.A(_0098_),
    .X(net535));
 sky130_fd_sc_hd__bufbuf_16 hold40 (.A(net568),
    .X(net536));
 sky130_fd_sc_hd__bufbuf_16 hold41 (.A(_0106_),
    .X(net537));
 sky130_fd_sc_hd__bufbuf_16 hold42 (.A(\wb_counter[13] ),
    .X(net538));
 sky130_fd_sc_hd__bufbuf_16 hold43 (.A(_0159_),
    .X(net539));
 sky130_fd_sc_hd__bufbuf_16 hold44 (.A(_0104_),
    .X(net540));
 sky130_fd_sc_hd__bufbuf_16 hold45 (.A(\wb_counter[16] ),
    .X(net541));
 sky130_fd_sc_hd__bufbuf_16 hold46 (.A(_0163_),
    .X(net542));
 sky130_fd_sc_hd__bufbuf_16 hold47 (.A(_0107_),
    .X(net543));
 sky130_fd_sc_hd__bufbuf_16 hold48 (.A(\wb_counter[5] ),
    .X(net544));
 sky130_fd_sc_hd__bufbuf_16 hold49 (.A(_0147_),
    .X(net545));
 sky130_fd_sc_hd__bufbuf_16 hold50 (.A(_0096_),
    .X(net546));
 sky130_fd_sc_hd__bufbuf_16 hold51 (.A(\wb_counter[19] ),
    .X(net547));
 sky130_fd_sc_hd__bufbuf_16 hold52 (.A(_0166_),
    .X(net548));
 sky130_fd_sc_hd__bufbuf_16 hold53 (.A(_0110_),
    .X(net549));
 sky130_fd_sc_hd__bufbuf_16 hold54 (.A(\wb_counter[22] ),
    .X(net550));
 sky130_fd_sc_hd__bufbuf_16 hold55 (.A(_0169_),
    .X(net551));
 sky130_fd_sc_hd__bufbuf_16 hold56 (.A(_0113_),
    .X(net552));
 sky130_fd_sc_hd__bufbuf_16 hold57 (.A(net348),
    .X(net553));
 sky130_fd_sc_hd__bufbuf_16 hold58 (.A(_0143_),
    .X(net554));
 sky130_fd_sc_hd__bufbuf_16 hold59 (.A(_0093_),
    .X(net555));
 sky130_fd_sc_hd__bufbuf_16 hold60 (.A(net357),
    .X(net556));
 sky130_fd_sc_hd__bufbuf_16 hold61 (.A(_0144_),
    .X(net557));
 sky130_fd_sc_hd__bufbuf_16 hold62 (.A(_0094_),
    .X(net558));
 sky130_fd_sc_hd__bufbuf_16 hold63 (.A(\wb_counter[6] ),
    .X(net559));
 sky130_fd_sc_hd__bufbuf_16 hold64 (.A(\wb_counter[20] ),
    .X(net560));
 sky130_fd_sc_hd__bufbuf_16 hold65 (.A(\wb_counter[18] ),
    .X(net561));
 sky130_fd_sc_hd__bufbuf_16 hold66 (.A(_0109_),
    .X(net562));
 sky130_fd_sc_hd__bufbuf_16 hold67 (.A(\wb_counter[12] ),
    .X(net563));
 sky130_fd_sc_hd__bufbuf_16 hold68 (.A(\wb_counter[17] ),
    .X(net564));
 sky130_fd_sc_hd__bufbuf_16 hold69 (.A(\wb_counter[21] ),
    .X(net565));
 sky130_fd_sc_hd__bufbuf_16 hold70 (.A(\wb_counter[0] ),
    .X(net566));
 sky130_fd_sc_hd__bufbuf_16 hold71 (.A(net337),
    .X(net567));
 sky130_fd_sc_hd__bufbuf_16 hold72 (.A(\wb_counter[15] ),
    .X(net568));
 sky130_fd_sc_hd__bufbuf_16 hold73 (.A(net358),
    .X(net569));
 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(_0201_));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(_0429_));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(\wb_design_addr_override[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA_6 (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA_7 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA_8 (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA_9 (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA_10 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA_11 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA_12 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA_13 (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA_14 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA_15 (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA_16 (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA_17 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA_18 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA_19 (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA_20 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA_21 (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA_22 (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA_23 (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA_24 (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA_25 (.DIODE(net476));
 sky130_fd_sc_hd__diode_2 ANTENNA_26 (.DIODE(_0134_));
 sky130_fd_sc_hd__diode_2 ANTENNA_27 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA_28 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA_29 (.DIODE(net261));
 sky130_fd_sc_hd__fill_2 FILLER_0_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_487 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_239 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_322 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_375 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_431 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_583 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_115 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_383 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_571 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_602 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_264 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_425 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_593 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_160 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_228 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_264 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_350 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_379 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_406 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_124 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_238 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_287 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_312 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_348 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_367 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_476 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_159 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_273 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_322 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_142 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_267 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_322 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_328 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_210 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_340 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_394 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_407 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_422 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_290 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_300 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_428 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_602 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_341 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_430 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_403 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_215 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_292 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_339 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_383 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_398 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_156 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_270 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_208 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_327 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_299 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_344 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_158 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_188 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_351 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_208 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_602 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_157 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_319 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_269 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_352 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_450 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_300 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_358 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_329 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_409 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_592 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_604 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_292 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_551 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_602 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_404 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_386 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_400 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_360 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_443 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_452 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_542 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_570 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_580 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_602 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_156 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_199 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_216 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_244 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_226 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_271 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_576 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_347 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_351 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_590 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_600 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_210 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_246 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_13 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_198 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_203 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_170 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_216 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_364 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_382 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_216 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_455 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_198 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_235 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_173 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_256 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_351 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_623 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_36 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_234 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_235 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_565 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_388 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_623 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_10 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_11 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_437 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_493 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_567 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_11 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_66 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_292 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_325 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_572 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_580 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_623 ();
 assign io_oeb[10] = net496;
 assign io_oeb[1] = net477;
 assign io_oeb[2] = net478;
 assign io_oeb[3] = net479;
 assign io_oeb[4] = net480;
 assign io_oeb[5] = net491;
 assign io_oeb[6] = net492;
 assign io_oeb[7] = net493;
 assign io_oeb[8] = net494;
 assign io_oeb[9] = net495;
 assign io_out[10] = net486;
 assign io_out[5] = net481;
 assign io_out[6] = net482;
 assign io_out[7] = net483;
 assign io_out[8] = net484;
 assign io_out[9] = net485;
 assign wbs_dat_o[28] = net487;
 assign wbs_dat_o[29] = net488;
 assign wbs_dat_o[30] = net489;
 assign wbs_dat_o[31] = net490;
endmodule

