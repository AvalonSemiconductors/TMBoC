// This is the unpowered netlist.
module wrapped_as1802 (clk,
    io_oeb,
    rst,
    io_in,
    io_out);
 input clk;
 output io_oeb;
 input rst;
 input [12:0] io_in;
 output [26:0] io_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire _2477_;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire _2494_;
 wire _2495_;
 wire _2496_;
 wire _2497_;
 wire _2498_;
 wire _2499_;
 wire _2500_;
 wire _2501_;
 wire _2502_;
 wire _2503_;
 wire _2504_;
 wire _2505_;
 wire _2506_;
 wire _2507_;
 wire _2508_;
 wire _2509_;
 wire _2510_;
 wire _2511_;
 wire _2512_;
 wire _2513_;
 wire _2514_;
 wire _2515_;
 wire _2516_;
 wire _2517_;
 wire _2518_;
 wire _2519_;
 wire _2520_;
 wire _2521_;
 wire _2522_;
 wire _2523_;
 wire _2524_;
 wire _2525_;
 wire _2526_;
 wire _2527_;
 wire _2528_;
 wire _2529_;
 wire _2530_;
 wire _2531_;
 wire _2532_;
 wire _2533_;
 wire _2534_;
 wire _2535_;
 wire _2536_;
 wire _2537_;
 wire _2538_;
 wire _2539_;
 wire _2540_;
 wire _2541_;
 wire _2542_;
 wire _2543_;
 wire _2544_;
 wire _2545_;
 wire _2546_;
 wire _2547_;
 wire _2548_;
 wire _2549_;
 wire _2550_;
 wire _2551_;
 wire _2552_;
 wire _2553_;
 wire _2554_;
 wire _2555_;
 wire _2556_;
 wire _2557_;
 wire _2558_;
 wire _2559_;
 wire _2560_;
 wire _2561_;
 wire _2562_;
 wire _2563_;
 wire _2564_;
 wire _2565_;
 wire _2566_;
 wire _2567_;
 wire _2568_;
 wire _2569_;
 wire _2570_;
 wire _2571_;
 wire _2572_;
 wire _2573_;
 wire _2574_;
 wire _2575_;
 wire _2576_;
 wire _2577_;
 wire _2578_;
 wire _2579_;
 wire _2580_;
 wire _2581_;
 wire _2582_;
 wire _2583_;
 wire _2584_;
 wire _2585_;
 wire _2586_;
 wire _2587_;
 wire _2588_;
 wire _2589_;
 wire _2590_;
 wire _2591_;
 wire _2592_;
 wire _2593_;
 wire _2594_;
 wire _2595_;
 wire _2596_;
 wire _2597_;
 wire _2598_;
 wire _2599_;
 wire _2600_;
 wire _2601_;
 wire _2602_;
 wire _2603_;
 wire _2604_;
 wire _2605_;
 wire _2606_;
 wire _2607_;
 wire _2608_;
 wire _2609_;
 wire _2610_;
 wire _2611_;
 wire _2612_;
 wire _2613_;
 wire _2614_;
 wire _2615_;
 wire _2616_;
 wire _2617_;
 wire _2618_;
 wire _2619_;
 wire _2620_;
 wire _2621_;
 wire _2622_;
 wire _2623_;
 wire _2624_;
 wire _2625_;
 wire _2626_;
 wire _2627_;
 wire _2628_;
 wire _2629_;
 wire _2630_;
 wire _2631_;
 wire _2632_;
 wire _2633_;
 wire _2634_;
 wire _2635_;
 wire _2636_;
 wire _2637_;
 wire _2638_;
 wire _2639_;
 wire _2640_;
 wire _2641_;
 wire _2642_;
 wire _2643_;
 wire _2644_;
 wire _2645_;
 wire _2646_;
 wire _2647_;
 wire _2648_;
 wire _2649_;
 wire _2650_;
 wire _2651_;
 wire _2652_;
 wire _2653_;
 wire _2654_;
 wire _2655_;
 wire _2656_;
 wire _2657_;
 wire _2658_;
 wire _2659_;
 wire _2660_;
 wire _2661_;
 wire _2662_;
 wire _2663_;
 wire _2664_;
 wire _2665_;
 wire _2666_;
 wire _2667_;
 wire _2668_;
 wire _2669_;
 wire _2670_;
 wire _2671_;
 wire _2672_;
 wire _2673_;
 wire _2674_;
 wire _2675_;
 wire _2676_;
 wire _2677_;
 wire _2678_;
 wire _2679_;
 wire _2680_;
 wire _2681_;
 wire _2682_;
 wire _2683_;
 wire _2684_;
 wire _2685_;
 wire _2686_;
 wire _2687_;
 wire _2688_;
 wire _2689_;
 wire _2690_;
 wire _2691_;
 wire _2692_;
 wire _2693_;
 wire _2694_;
 wire _2695_;
 wire _2696_;
 wire _2697_;
 wire _2698_;
 wire _2699_;
 wire _2700_;
 wire _2701_;
 wire _2702_;
 wire _2703_;
 wire _2704_;
 wire _2705_;
 wire _2706_;
 wire _2707_;
 wire _2708_;
 wire _2709_;
 wire _2710_;
 wire _2711_;
 wire _2712_;
 wire _2713_;
 wire _2714_;
 wire _2715_;
 wire _2716_;
 wire _2717_;
 wire _2718_;
 wire _2719_;
 wire _2720_;
 wire _2721_;
 wire _2722_;
 wire \as1802.DF ;
 wire \as1802.D[0] ;
 wire \as1802.D[1] ;
 wire \as1802.D[2] ;
 wire \as1802.D[3] ;
 wire \as1802.D[4] ;
 wire \as1802.D[5] ;
 wire \as1802.D[6] ;
 wire \as1802.D[7] ;
 wire \as1802.EF_l[0] ;
 wire \as1802.EF_l[1] ;
 wire \as1802.EF_l[2] ;
 wire \as1802.EF_l[3] ;
 wire \as1802.IE ;
 wire \as1802.P[0] ;
 wire \as1802.P[1] ;
 wire \as1802.P[2] ;
 wire \as1802.P[3] ;
 wire \as1802.T[0] ;
 wire \as1802.T[1] ;
 wire \as1802.T[2] ;
 wire \as1802.T[3] ;
 wire \as1802.T[4] ;
 wire \as1802.T[5] ;
 wire \as1802.T[6] ;
 wire \as1802.T[7] ;
 wire \as1802.X[0] ;
 wire \as1802.X[1] ;
 wire \as1802.X[2] ;
 wire \as1802.X[3] ;
 wire \as1802.addr_buff[0] ;
 wire \as1802.addr_buff[10] ;
 wire \as1802.addr_buff[11] ;
 wire \as1802.addr_buff[12] ;
 wire \as1802.addr_buff[13] ;
 wire \as1802.addr_buff[14] ;
 wire \as1802.addr_buff[15] ;
 wire \as1802.addr_buff[1] ;
 wire \as1802.addr_buff[2] ;
 wire \as1802.addr_buff[3] ;
 wire \as1802.addr_buff[4] ;
 wire \as1802.addr_buff[5] ;
 wire \as1802.addr_buff[6] ;
 wire \as1802.addr_buff[7] ;
 wire \as1802.addr_buff[8] ;
 wire \as1802.addr_buff[9] ;
 wire \as1802.cond_inv ;
 wire \as1802.idle ;
 wire \as1802.instr_cycle[0] ;
 wire \as1802.instr_cycle[1] ;
 wire \as1802.instr_cycle[2] ;
 wire \as1802.instr_cycle[3] ;
 wire \as1802.instr_latch[0] ;
 wire \as1802.instr_latch[1] ;
 wire \as1802.instr_latch[2] ;
 wire \as1802.instr_latch[4] ;
 wire \as1802.instr_latch[5] ;
 wire \as1802.instr_latch[6] ;
 wire \as1802.instr_latch[7] ;
 wire \as1802.last_hi_addr[0] ;
 wire \as1802.last_hi_addr[1] ;
 wire \as1802.last_hi_addr[2] ;
 wire \as1802.last_hi_addr[3] ;
 wire \as1802.last_hi_addr[4] ;
 wire \as1802.last_hi_addr[5] ;
 wire \as1802.last_hi_addr[6] ;
 wire \as1802.last_hi_addr[7] ;
 wire \as1802.lda ;
 wire \as1802.mem_cycle[0] ;
 wire \as1802.mem_cycle[1] ;
 wire \as1802.mem_cycle[2] ;
 wire \as1802.mem_write ;
 wire \as1802.regs[0][0] ;
 wire \as1802.regs[0][10] ;
 wire \as1802.regs[0][11] ;
 wire \as1802.regs[0][12] ;
 wire \as1802.regs[0][13] ;
 wire \as1802.regs[0][14] ;
 wire \as1802.regs[0][15] ;
 wire \as1802.regs[0][1] ;
 wire \as1802.regs[0][2] ;
 wire \as1802.regs[0][3] ;
 wire \as1802.regs[0][4] ;
 wire \as1802.regs[0][5] ;
 wire \as1802.regs[0][6] ;
 wire \as1802.regs[0][7] ;
 wire \as1802.regs[0][8] ;
 wire \as1802.regs[0][9] ;
 wire \as1802.regs[10][0] ;
 wire \as1802.regs[10][10] ;
 wire \as1802.regs[10][11] ;
 wire \as1802.regs[10][12] ;
 wire \as1802.regs[10][13] ;
 wire \as1802.regs[10][14] ;
 wire \as1802.regs[10][15] ;
 wire \as1802.regs[10][1] ;
 wire \as1802.regs[10][2] ;
 wire \as1802.regs[10][3] ;
 wire \as1802.regs[10][4] ;
 wire \as1802.regs[10][5] ;
 wire \as1802.regs[10][6] ;
 wire \as1802.regs[10][7] ;
 wire \as1802.regs[10][8] ;
 wire \as1802.regs[10][9] ;
 wire \as1802.regs[11][0] ;
 wire \as1802.regs[11][10] ;
 wire \as1802.regs[11][11] ;
 wire \as1802.regs[11][12] ;
 wire \as1802.regs[11][13] ;
 wire \as1802.regs[11][14] ;
 wire \as1802.regs[11][15] ;
 wire \as1802.regs[11][1] ;
 wire \as1802.regs[11][2] ;
 wire \as1802.regs[11][3] ;
 wire \as1802.regs[11][4] ;
 wire \as1802.regs[11][5] ;
 wire \as1802.regs[11][6] ;
 wire \as1802.regs[11][7] ;
 wire \as1802.regs[11][8] ;
 wire \as1802.regs[11][9] ;
 wire \as1802.regs[12][0] ;
 wire \as1802.regs[12][10] ;
 wire \as1802.regs[12][11] ;
 wire \as1802.regs[12][12] ;
 wire \as1802.regs[12][13] ;
 wire \as1802.regs[12][14] ;
 wire \as1802.regs[12][15] ;
 wire \as1802.regs[12][1] ;
 wire \as1802.regs[12][2] ;
 wire \as1802.regs[12][3] ;
 wire \as1802.regs[12][4] ;
 wire \as1802.regs[12][5] ;
 wire \as1802.regs[12][6] ;
 wire \as1802.regs[12][7] ;
 wire \as1802.regs[12][8] ;
 wire \as1802.regs[12][9] ;
 wire \as1802.regs[13][0] ;
 wire \as1802.regs[13][10] ;
 wire \as1802.regs[13][11] ;
 wire \as1802.regs[13][12] ;
 wire \as1802.regs[13][13] ;
 wire \as1802.regs[13][14] ;
 wire \as1802.regs[13][15] ;
 wire \as1802.regs[13][1] ;
 wire \as1802.regs[13][2] ;
 wire \as1802.regs[13][3] ;
 wire \as1802.regs[13][4] ;
 wire \as1802.regs[13][5] ;
 wire \as1802.regs[13][6] ;
 wire \as1802.regs[13][7] ;
 wire \as1802.regs[13][8] ;
 wire \as1802.regs[13][9] ;
 wire \as1802.regs[14][0] ;
 wire \as1802.regs[14][10] ;
 wire \as1802.regs[14][11] ;
 wire \as1802.regs[14][12] ;
 wire \as1802.regs[14][13] ;
 wire \as1802.regs[14][14] ;
 wire \as1802.regs[14][15] ;
 wire \as1802.regs[14][1] ;
 wire \as1802.regs[14][2] ;
 wire \as1802.regs[14][3] ;
 wire \as1802.regs[14][4] ;
 wire \as1802.regs[14][5] ;
 wire \as1802.regs[14][6] ;
 wire \as1802.regs[14][7] ;
 wire \as1802.regs[14][8] ;
 wire \as1802.regs[14][9] ;
 wire \as1802.regs[15][0] ;
 wire \as1802.regs[15][10] ;
 wire \as1802.regs[15][11] ;
 wire \as1802.regs[15][12] ;
 wire \as1802.regs[15][13] ;
 wire \as1802.regs[15][14] ;
 wire \as1802.regs[15][15] ;
 wire \as1802.regs[15][1] ;
 wire \as1802.regs[15][2] ;
 wire \as1802.regs[15][3] ;
 wire \as1802.regs[15][4] ;
 wire \as1802.regs[15][5] ;
 wire \as1802.regs[15][6] ;
 wire \as1802.regs[15][7] ;
 wire \as1802.regs[15][8] ;
 wire \as1802.regs[15][9] ;
 wire \as1802.regs[1][0] ;
 wire \as1802.regs[1][10] ;
 wire \as1802.regs[1][11] ;
 wire \as1802.regs[1][12] ;
 wire \as1802.regs[1][13] ;
 wire \as1802.regs[1][14] ;
 wire \as1802.regs[1][15] ;
 wire \as1802.regs[1][1] ;
 wire \as1802.regs[1][2] ;
 wire \as1802.regs[1][3] ;
 wire \as1802.regs[1][4] ;
 wire \as1802.regs[1][5] ;
 wire \as1802.regs[1][6] ;
 wire \as1802.regs[1][7] ;
 wire \as1802.regs[1][8] ;
 wire \as1802.regs[1][9] ;
 wire \as1802.regs[2][0] ;
 wire \as1802.regs[2][10] ;
 wire \as1802.regs[2][11] ;
 wire \as1802.regs[2][12] ;
 wire \as1802.regs[2][13] ;
 wire \as1802.regs[2][14] ;
 wire \as1802.regs[2][15] ;
 wire \as1802.regs[2][1] ;
 wire \as1802.regs[2][2] ;
 wire \as1802.regs[2][3] ;
 wire \as1802.regs[2][4] ;
 wire \as1802.regs[2][5] ;
 wire \as1802.regs[2][6] ;
 wire \as1802.regs[2][7] ;
 wire \as1802.regs[2][8] ;
 wire \as1802.regs[2][9] ;
 wire \as1802.regs[3][0] ;
 wire \as1802.regs[3][10] ;
 wire \as1802.regs[3][11] ;
 wire \as1802.regs[3][12] ;
 wire \as1802.regs[3][13] ;
 wire \as1802.regs[3][14] ;
 wire \as1802.regs[3][15] ;
 wire \as1802.regs[3][1] ;
 wire \as1802.regs[3][2] ;
 wire \as1802.regs[3][3] ;
 wire \as1802.regs[3][4] ;
 wire \as1802.regs[3][5] ;
 wire \as1802.regs[3][6] ;
 wire \as1802.regs[3][7] ;
 wire \as1802.regs[3][8] ;
 wire \as1802.regs[3][9] ;
 wire \as1802.regs[4][0] ;
 wire \as1802.regs[4][10] ;
 wire \as1802.regs[4][11] ;
 wire \as1802.regs[4][12] ;
 wire \as1802.regs[4][13] ;
 wire \as1802.regs[4][14] ;
 wire \as1802.regs[4][15] ;
 wire \as1802.regs[4][1] ;
 wire \as1802.regs[4][2] ;
 wire \as1802.regs[4][3] ;
 wire \as1802.regs[4][4] ;
 wire \as1802.regs[4][5] ;
 wire \as1802.regs[4][6] ;
 wire \as1802.regs[4][7] ;
 wire \as1802.regs[4][8] ;
 wire \as1802.regs[4][9] ;
 wire \as1802.regs[5][0] ;
 wire \as1802.regs[5][10] ;
 wire \as1802.regs[5][11] ;
 wire \as1802.regs[5][12] ;
 wire \as1802.regs[5][13] ;
 wire \as1802.regs[5][14] ;
 wire \as1802.regs[5][15] ;
 wire \as1802.regs[5][1] ;
 wire \as1802.regs[5][2] ;
 wire \as1802.regs[5][3] ;
 wire \as1802.regs[5][4] ;
 wire \as1802.regs[5][5] ;
 wire \as1802.regs[5][6] ;
 wire \as1802.regs[5][7] ;
 wire \as1802.regs[5][8] ;
 wire \as1802.regs[5][9] ;
 wire \as1802.regs[6][0] ;
 wire \as1802.regs[6][10] ;
 wire \as1802.regs[6][11] ;
 wire \as1802.regs[6][12] ;
 wire \as1802.regs[6][13] ;
 wire \as1802.regs[6][14] ;
 wire \as1802.regs[6][15] ;
 wire \as1802.regs[6][1] ;
 wire \as1802.regs[6][2] ;
 wire \as1802.regs[6][3] ;
 wire \as1802.regs[6][4] ;
 wire \as1802.regs[6][5] ;
 wire \as1802.regs[6][6] ;
 wire \as1802.regs[6][7] ;
 wire \as1802.regs[6][8] ;
 wire \as1802.regs[6][9] ;
 wire \as1802.regs[7][0] ;
 wire \as1802.regs[7][10] ;
 wire \as1802.regs[7][11] ;
 wire \as1802.regs[7][12] ;
 wire \as1802.regs[7][13] ;
 wire \as1802.regs[7][14] ;
 wire \as1802.regs[7][15] ;
 wire \as1802.regs[7][1] ;
 wire \as1802.regs[7][2] ;
 wire \as1802.regs[7][3] ;
 wire \as1802.regs[7][4] ;
 wire \as1802.regs[7][5] ;
 wire \as1802.regs[7][6] ;
 wire \as1802.regs[7][7] ;
 wire \as1802.regs[7][8] ;
 wire \as1802.regs[7][9] ;
 wire \as1802.regs[8][0] ;
 wire \as1802.regs[8][10] ;
 wire \as1802.regs[8][11] ;
 wire \as1802.regs[8][12] ;
 wire \as1802.regs[8][13] ;
 wire \as1802.regs[8][14] ;
 wire \as1802.regs[8][15] ;
 wire \as1802.regs[8][1] ;
 wire \as1802.regs[8][2] ;
 wire \as1802.regs[8][3] ;
 wire \as1802.regs[8][4] ;
 wire \as1802.regs[8][5] ;
 wire \as1802.regs[8][6] ;
 wire \as1802.regs[8][7] ;
 wire \as1802.regs[8][8] ;
 wire \as1802.regs[8][9] ;
 wire \as1802.regs[9][0] ;
 wire \as1802.regs[9][10] ;
 wire \as1802.regs[9][11] ;
 wire \as1802.regs[9][12] ;
 wire \as1802.regs[9][13] ;
 wire \as1802.regs[9][14] ;
 wire \as1802.regs[9][15] ;
 wire \as1802.regs[9][1] ;
 wire \as1802.regs[9][2] ;
 wire \as1802.regs[9][3] ;
 wire \as1802.regs[9][4] ;
 wire \as1802.regs[9][5] ;
 wire \as1802.regs[9][6] ;
 wire \as1802.regs[9][7] ;
 wire \as1802.regs[9][8] ;
 wire \as1802.regs[9][9] ;
 wire \as1802.will_interrupt ;
 wire net18;
 wire net19;
 wire clknet_leaf_0_clk;
 wire net16;
 wire net17;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_45_clk;
 wire clknet_leaf_46_clk;
 wire clknet_leaf_47_clk;
 wire clknet_leaf_48_clk;
 wire clknet_leaf_49_clk;
 wire clknet_leaf_50_clk;
 wire clknet_0_clk;
 wire clknet_2_0__leaf_clk;
 wire clknet_2_1__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_3__leaf_clk;
 wire clknet_opt_1_0_clk;
 wire clknet_opt_2_0_clk;

 sky130_fd_sc_hd__buf_4 _2723_ (.A(net14),
    .X(_2456_));
 sky130_fd_sc_hd__clkinv_2 _2724_ (.A(_2456_),
    .Y(_2457_));
 sky130_fd_sc_hd__clkbuf_4 _2725_ (.A(_2457_),
    .X(_2458_));
 sky130_fd_sc_hd__or3_1 _2726_ (.A(\as1802.mem_cycle[2] ),
    .B(\as1802.mem_cycle[1] ),
    .C(\as1802.mem_cycle[0] ),
    .X(_2459_));
 sky130_fd_sc_hd__buf_2 _2727_ (.A(_2459_),
    .X(_2460_));
 sky130_fd_sc_hd__buf_4 _2728_ (.A(_2460_),
    .X(_2461_));
 sky130_fd_sc_hd__clkbuf_4 _2729_ (.A(_2461_),
    .X(_2462_));
 sky130_fd_sc_hd__xnor2_2 _2730_ (.A(\as1802.instr_latch[5] ),
    .B(\as1802.instr_latch[4] ),
    .Y(_2463_));
 sky130_fd_sc_hd__or3_2 _2731_ (.A(\as1802.instr_latch[7] ),
    .B(\as1802.instr_latch[6] ),
    .C(_2463_),
    .X(_2464_));
 sky130_fd_sc_hd__or4_1 _2732_ (.A(\as1802.instr_latch[5] ),
    .B(\as1802.instr_latch[4] ),
    .C(\as1802.instr_latch[7] ),
    .D(\as1802.instr_latch[6] ),
    .X(_2465_));
 sky130_fd_sc_hd__buf_2 _2733_ (.A(_2465_),
    .X(_2466_));
 sky130_fd_sc_hd__nor2_1 _2734_ (.A(net14),
    .B(_2460_),
    .Y(_2467_));
 sky130_fd_sc_hd__and3_1 _2735_ (.A(_2464_),
    .B(_2466_),
    .C(_2467_),
    .X(_2468_));
 sky130_fd_sc_hd__clkbuf_8 _2736_ (.A(\as1802.instr_latch[0] ),
    .X(_2469_));
 sky130_fd_sc_hd__nor2_4 _2737_ (.A(\as1802.instr_latch[1] ),
    .B(_2469_),
    .Y(_2470_));
 sky130_fd_sc_hd__a21o_1 _2738_ (.A1(\as1802.cond_inv ),
    .A2(_2470_),
    .B1(\as1802.instr_latch[2] ),
    .X(_2471_));
 sky130_fd_sc_hd__clkinv_2 _2739_ (.A(_2471_),
    .Y(_2472_));
 sky130_fd_sc_hd__clkbuf_4 _2740_ (.A(\as1802.instr_latch[5] ),
    .X(_2473_));
 sky130_fd_sc_hd__clkbuf_4 _2741_ (.A(\as1802.instr_latch[4] ),
    .X(_2474_));
 sky130_fd_sc_hd__or2_1 _2742_ (.A(_2473_),
    .B(_2474_),
    .X(_2475_));
 sky130_fd_sc_hd__clkbuf_4 _2743_ (.A(\as1802.instr_latch[7] ),
    .X(_2476_));
 sky130_fd_sc_hd__clkbuf_4 _2744_ (.A(\as1802.instr_latch[6] ),
    .X(_2477_));
 sky130_fd_sc_hd__nand2_2 _2745_ (.A(_2476_),
    .B(_2477_),
    .Y(_2478_));
 sky130_fd_sc_hd__nor2_1 _2746_ (.A(_2475_),
    .B(_2478_),
    .Y(_2479_));
 sky130_fd_sc_hd__clkbuf_4 _2747_ (.A(_2479_),
    .X(_2480_));
 sky130_fd_sc_hd__and3_1 _2748_ (.A(_2468_),
    .B(_2472_),
    .C(_2480_),
    .X(_2481_));
 sky130_fd_sc_hd__a32o_1 _2749_ (.A1(_2458_),
    .A2(\as1802.instr_cycle[3] ),
    .A3(_2462_),
    .B1(_2481_),
    .B2(\as1802.instr_cycle[1] ),
    .X(_0007_));
 sky130_fd_sc_hd__buf_2 _2750_ (.A(\as1802.instr_cycle[2] ),
    .X(_2482_));
 sky130_fd_sc_hd__or4_1 _2751_ (.A(\as1802.mem_cycle[2] ),
    .B(\as1802.mem_cycle[1] ),
    .C(\as1802.mem_cycle[0] ),
    .D(net14),
    .X(_2483_));
 sky130_fd_sc_hd__buf_2 _2752_ (.A(_2483_),
    .X(_2484_));
 sky130_fd_sc_hd__buf_4 _2753_ (.A(_2484_),
    .X(_2485_));
 sky130_fd_sc_hd__inv_2 _2754_ (.A(\as1802.instr_cycle[0] ),
    .Y(_2486_));
 sky130_fd_sc_hd__inv_2 _2755_ (.A(\as1802.idle ),
    .Y(_2487_));
 sky130_fd_sc_hd__nand2_1 _2756_ (.A(\as1802.IE ),
    .B(net12),
    .Y(_2488_));
 sky130_fd_sc_hd__nand2_1 _2757_ (.A(_2487_),
    .B(_2488_),
    .Y(_2489_));
 sky130_fd_sc_hd__or3_1 _2758_ (.A(\as1802.will_interrupt ),
    .B(_2486_),
    .C(_2489_),
    .X(_2490_));
 sky130_fd_sc_hd__nor2_1 _2759_ (.A(_2485_),
    .B(_2490_),
    .Y(_2491_));
 sky130_fd_sc_hd__a31o_1 _2760_ (.A1(_2482_),
    .A2(_2458_),
    .A3(_2462_),
    .B1(_2491_),
    .X(_0006_));
 sky130_fd_sc_hd__inv_2 _2761_ (.A(\as1802.cond_inv ),
    .Y(_2492_));
 sky130_fd_sc_hd__buf_4 _2762_ (.A(_2492_),
    .X(_2493_));
 sky130_fd_sc_hd__buf_4 _2763_ (.A(_2493_),
    .X(_2494_));
 sky130_fd_sc_hd__buf_2 _2764_ (.A(\as1802.instr_latch[2] ),
    .X(_2495_));
 sky130_fd_sc_hd__buf_4 _2765_ (.A(_2495_),
    .X(_2496_));
 sky130_fd_sc_hd__or2b_1 _2766_ (.A(_2469_),
    .B_N(\as1802.instr_latch[1] ),
    .X(_2497_));
 sky130_fd_sc_hd__or4_1 _2767_ (.A(\as1802.D[5] ),
    .B(\as1802.D[4] ),
    .C(\as1802.D[7] ),
    .D(\as1802.D[6] ),
    .X(_2498_));
 sky130_fd_sc_hd__or4_1 _2768_ (.A(\as1802.D[1] ),
    .B(\as1802.D[0] ),
    .C(\as1802.D[3] ),
    .D(\as1802.D[2] ),
    .X(_2499_));
 sky130_fd_sc_hd__nand2b_4 _2769_ (.A_N(\as1802.instr_latch[1] ),
    .B(_2469_),
    .Y(_2500_));
 sky130_fd_sc_hd__inv_2 _2770_ (.A(io_out[21]),
    .Y(_2501_));
 sky130_fd_sc_hd__o32a_1 _2771_ (.A1(_2497_),
    .A2(_2498_),
    .A3(_2499_),
    .B1(_2500_),
    .B2(_2501_),
    .X(_2502_));
 sky130_fd_sc_hd__inv_4 _2772_ (.A(\as1802.instr_latch[2] ),
    .Y(_2503_));
 sky130_fd_sc_hd__clkbuf_4 _2773_ (.A(\as1802.instr_latch[1] ),
    .X(_2504_));
 sky130_fd_sc_hd__nand2_2 _2774_ (.A(_2504_),
    .B(_2469_),
    .Y(_2505_));
 sky130_fd_sc_hd__nor2_4 _2775_ (.A(_2503_),
    .B(_2505_),
    .Y(_2506_));
 sky130_fd_sc_hd__nor2b_2 _2776_ (.A(_2469_),
    .B_N(_2504_),
    .Y(_2507_));
 sky130_fd_sc_hd__nor2_4 _2777_ (.A(_2503_),
    .B(_2500_),
    .Y(_2508_));
 sky130_fd_sc_hd__a32o_1 _2778_ (.A1(_2495_),
    .A2(\as1802.EF_l[2] ),
    .A3(_2507_),
    .B1(_2508_),
    .B2(\as1802.EF_l[1] ),
    .X(_2509_));
 sky130_fd_sc_hd__or2_1 _2779_ (.A(_2495_),
    .B(_2505_),
    .X(_2510_));
 sky130_fd_sc_hd__buf_4 _2780_ (.A(_2510_),
    .X(_2511_));
 sky130_fd_sc_hd__inv_2 _2781_ (.A(_2511_),
    .Y(_2512_));
 sky130_fd_sc_hd__inv_2 _2782_ (.A(\as1802.instr_latch[0] ),
    .Y(_2513_));
 sky130_fd_sc_hd__nand2_1 _2783_ (.A(_2513_),
    .B(_2495_),
    .Y(_2514_));
 sky130_fd_sc_hd__nor2_1 _2784_ (.A(_2504_),
    .B(_2514_),
    .Y(_2515_));
 sky130_fd_sc_hd__nor3_4 _2785_ (.A(\as1802.instr_latch[1] ),
    .B(_2469_),
    .C(\as1802.instr_latch[2] ),
    .Y(_2516_));
 sky130_fd_sc_hd__a221o_1 _2786_ (.A1(\as1802.DF ),
    .A2(_2512_),
    .B1(_2515_),
    .B2(\as1802.EF_l[0] ),
    .C1(_2516_),
    .X(_2517_));
 sky130_fd_sc_hd__a211o_1 _2787_ (.A1(\as1802.EF_l[3] ),
    .A2(_2506_),
    .B1(_2509_),
    .C1(_2517_),
    .X(_2518_));
 sky130_fd_sc_hd__o21ba_1 _2788_ (.A1(_2496_),
    .A2(_2502_),
    .B1_N(_2518_),
    .X(_2519_));
 sky130_fd_sc_hd__xnor2_2 _2789_ (.A(_2494_),
    .B(_2519_),
    .Y(_2520_));
 sky130_fd_sc_hd__nand2_2 _2790_ (.A(_2473_),
    .B(_2474_),
    .Y(_2521_));
 sky130_fd_sc_hd__or3_2 _2791_ (.A(_2476_),
    .B(_2477_),
    .C(_2521_),
    .X(_2522_));
 sky130_fd_sc_hd__nor3_1 _2792_ (.A(\as1802.instr_latch[5] ),
    .B(\as1802.instr_latch[7] ),
    .C(\as1802.instr_latch[6] ),
    .Y(_2523_));
 sky130_fd_sc_hd__or2_1 _2793_ (.A(_2460_),
    .B(_2523_),
    .X(_2524_));
 sky130_fd_sc_hd__nand2b_4 _2794_ (.A_N(\as1802.instr_latch[7] ),
    .B(_2477_),
    .Y(_2525_));
 sky130_fd_sc_hd__nor2_2 _2795_ (.A(_2521_),
    .B(_2525_),
    .Y(_2526_));
 sky130_fd_sc_hd__clkinv_2 _2796_ (.A(\as1802.instr_latch[1] ),
    .Y(_2527_));
 sky130_fd_sc_hd__a22o_1 _2797_ (.A1(_2527_),
    .A2(_2492_),
    .B1(_2497_),
    .B2(_2495_),
    .X(_2528_));
 sky130_fd_sc_hd__nand2_1 _2798_ (.A(_2526_),
    .B(_2528_),
    .Y(_2529_));
 sky130_fd_sc_hd__o32a_1 _2799_ (.A1(_2461_),
    .A2(_2520_),
    .A3(_2522_),
    .B1(_2524_),
    .B2(_2529_),
    .X(_2530_));
 sky130_fd_sc_hd__o21ai_1 _2800_ (.A1(_2498_),
    .A2(_2499_),
    .B1(_2507_),
    .Y(_2531_));
 sky130_fd_sc_hd__o22a_1 _2801_ (.A1(io_out[21]),
    .A2(_2500_),
    .B1(_2505_),
    .B2(\as1802.DF ),
    .X(_2532_));
 sky130_fd_sc_hd__clkbuf_4 _2802_ (.A(\as1802.cond_inv ),
    .X(_2533_));
 sky130_fd_sc_hd__xnor2_1 _2803_ (.A(\as1802.instr_latch[2] ),
    .B(_2533_),
    .Y(_2534_));
 sky130_fd_sc_hd__a21oi_1 _2804_ (.A1(_2531_),
    .A2(_2532_),
    .B1(_2534_),
    .Y(_2535_));
 sky130_fd_sc_hd__and2b_1 _2805_ (.A_N(_2502_),
    .B(_2534_),
    .X(_2536_));
 sky130_fd_sc_hd__nor2_1 _2806_ (.A(_2527_),
    .B(_2513_),
    .Y(_2537_));
 sky130_fd_sc_hd__a31o_1 _2807_ (.A1(\as1802.IE ),
    .A2(_2533_),
    .A3(_2470_),
    .B1(_2516_),
    .X(_2538_));
 sky130_fd_sc_hd__a31o_1 _2808_ (.A1(\as1802.DF ),
    .A2(_2537_),
    .A3(_2534_),
    .B1(_2538_),
    .X(_2539_));
 sky130_fd_sc_hd__or3_1 _2809_ (.A(_2535_),
    .B(_2536_),
    .C(_2539_),
    .X(_2540_));
 sky130_fd_sc_hd__a2bb2o_1 _2810_ (.A1_N(_2456_),
    .A2_N(_2530_),
    .B1(_2540_),
    .B2(_2481_),
    .X(_2541_));
 sky130_fd_sc_hd__nand2_2 _2811_ (.A(_2503_),
    .B(_2470_),
    .Y(_2542_));
 sky130_fd_sc_hd__nand2_2 _2812_ (.A(_2495_),
    .B(_2507_),
    .Y(_2543_));
 sky130_fd_sc_hd__nor2_1 _2813_ (.A(_2521_),
    .B(_2478_),
    .Y(_2544_));
 sky130_fd_sc_hd__and4_2 _2814_ (.A(\as1802.instr_cycle[2] ),
    .B(_2542_),
    .C(_2543_),
    .D(_2544_),
    .X(_2545_));
 sky130_fd_sc_hd__a32o_1 _2815_ (.A1(_2457_),
    .A2(\as1802.instr_cycle[1] ),
    .A3(_2462_),
    .B1(_2468_),
    .B2(_2545_),
    .X(_2546_));
 sky130_fd_sc_hd__a21o_1 _2816_ (.A1(_2482_),
    .A2(_2541_),
    .B1(_2546_),
    .X(_0005_));
 sky130_fd_sc_hd__nor3_4 _2817_ (.A(\as1802.mem_cycle[2] ),
    .B(\as1802.mem_cycle[1] ),
    .C(\as1802.mem_cycle[0] ),
    .Y(_2547_));
 sky130_fd_sc_hd__clkbuf_4 _2818_ (.A(_2547_),
    .X(_2548_));
 sky130_fd_sc_hd__nor2_2 _2819_ (.A(_2476_),
    .B(_2477_),
    .Y(_2549_));
 sky130_fd_sc_hd__and3_1 _2820_ (.A(_2473_),
    .B(_2474_),
    .C(_2549_),
    .X(_2550_));
 sky130_fd_sc_hd__buf_2 _2821_ (.A(_2550_),
    .X(_2551_));
 sky130_fd_sc_hd__or2_1 _2822_ (.A(_2521_),
    .B(_2525_),
    .X(_2552_));
 sky130_fd_sc_hd__buf_4 _2823_ (.A(_2552_),
    .X(_2553_));
 sky130_fd_sc_hd__clkbuf_4 _2824_ (.A(_2553_),
    .X(_2554_));
 sky130_fd_sc_hd__clkbuf_4 _2825_ (.A(_2533_),
    .X(_2555_));
 sky130_fd_sc_hd__buf_4 _2826_ (.A(_2555_),
    .X(_2556_));
 sky130_fd_sc_hd__nand2_2 _2827_ (.A(_2496_),
    .B(_2470_),
    .Y(_2557_));
 sky130_fd_sc_hd__nor2_1 _2828_ (.A(_2556_),
    .B(_2557_),
    .Y(_2558_));
 sky130_fd_sc_hd__a211o_1 _2829_ (.A1(_2471_),
    .A2(_2554_),
    .B1(_2558_),
    .C1(\as1802.instr_cycle[3] ),
    .X(_2559_));
 sky130_fd_sc_hd__and2b_1 _2830_ (.A_N(_2463_),
    .B(_2476_),
    .X(_2560_));
 sky130_fd_sc_hd__nand2b_4 _2831_ (.A_N(\as1802.instr_latch[6] ),
    .B(\as1802.instr_latch[7] ),
    .Y(_2561_));
 sky130_fd_sc_hd__nor2_2 _2832_ (.A(_2475_),
    .B(_2561_),
    .Y(_2562_));
 sky130_fd_sc_hd__nor2_4 _2833_ (.A(_2473_),
    .B(_2525_),
    .Y(_2563_));
 sky130_fd_sc_hd__a2111o_1 _2834_ (.A1(_2549_),
    .A2(_2521_),
    .B1(_2560_),
    .C1(_2562_),
    .D1(_2563_),
    .X(_2564_));
 sky130_fd_sc_hd__nand2_1 _2835_ (.A(_2482_),
    .B(_2543_),
    .Y(_2565_));
 sky130_fd_sc_hd__o21a_1 _2836_ (.A1(_2516_),
    .A2(_2565_),
    .B1(_2544_),
    .X(_2566_));
 sky130_fd_sc_hd__clkinv_2 _2837_ (.A(_2474_),
    .Y(_2567_));
 sky130_fd_sc_hd__nand2_1 _2838_ (.A(_2473_),
    .B(_2567_),
    .Y(_2568_));
 sky130_fd_sc_hd__nor2_2 _2839_ (.A(_2568_),
    .B(_2525_),
    .Y(_2569_));
 sky130_fd_sc_hd__nand2_4 _2840_ (.A(\as1802.instr_cycle[2] ),
    .B(_2528_),
    .Y(_2570_));
 sky130_fd_sc_hd__clkinv_2 _2841_ (.A(_2570_),
    .Y(_2571_));
 sky130_fd_sc_hd__nor2_2 _2842_ (.A(_2553_),
    .B(_2571_),
    .Y(_2572_));
 sky130_fd_sc_hd__or2_1 _2843_ (.A(_2569_),
    .B(_2572_),
    .X(_2573_));
 sky130_fd_sc_hd__a2111o_1 _2844_ (.A1(_2480_),
    .A2(_2559_),
    .B1(_2564_),
    .C1(_2566_),
    .D1(_2573_),
    .X(_2574_));
 sky130_fd_sc_hd__or3_1 _2845_ (.A(_2482_),
    .B(\as1802.instr_cycle[1] ),
    .C(\as1802.instr_cycle[3] ),
    .X(_2575_));
 sky130_fd_sc_hd__nand2_1 _2846_ (.A(_2482_),
    .B(_2481_),
    .Y(_2576_));
 sky130_fd_sc_hd__nor2_1 _2847_ (.A(\as1802.instr_cycle[1] ),
    .B(\as1802.instr_cycle[3] ),
    .Y(_2577_));
 sky130_fd_sc_hd__or2_1 _2848_ (.A(\as1802.will_interrupt ),
    .B(_2461_),
    .X(_2578_));
 sky130_fd_sc_hd__buf_2 _2849_ (.A(\as1802.instr_cycle[0] ),
    .X(_2579_));
 sky130_fd_sc_hd__clkbuf_4 _2850_ (.A(_2579_),
    .X(_2580_));
 sky130_fd_sc_hd__clkbuf_4 _2851_ (.A(_2580_),
    .X(_2581_));
 sky130_fd_sc_hd__o21ai_1 _2852_ (.A1(_2489_),
    .A2(_2578_),
    .B1(_2581_),
    .Y(_2582_));
 sky130_fd_sc_hd__or2_1 _2853_ (.A(_2475_),
    .B(_2525_),
    .X(_2583_));
 sky130_fd_sc_hd__or3b_1 _2854_ (.A(_2460_),
    .B(_2549_),
    .C_N(_2583_),
    .X(_2584_));
 sky130_fd_sc_hd__or2_1 _2855_ (.A(_2521_),
    .B(_2561_),
    .X(_2585_));
 sky130_fd_sc_hd__or3b_1 _2856_ (.A(_2584_),
    .B(_2585_),
    .C_N(_2575_),
    .X(_2586_));
 sky130_fd_sc_hd__o311a_1 _2857_ (.A1(_2461_),
    .A2(_2522_),
    .A3(_2577_),
    .B1(_2582_),
    .C1(_2586_),
    .X(_2587_));
 sky130_fd_sc_hd__o211ai_1 _2858_ (.A1(_2540_),
    .A2(_2576_),
    .B1(_2587_),
    .C1(_2457_),
    .Y(_2588_));
 sky130_fd_sc_hd__a31o_1 _2859_ (.A1(_2548_),
    .A2(_2574_),
    .A3(_2575_),
    .B1(_2588_),
    .X(_2589_));
 sky130_fd_sc_hd__a41o_1 _2860_ (.A1(_2482_),
    .A2(_2548_),
    .A3(_2520_),
    .A4(_2551_),
    .B1(_2589_),
    .X(_0004_));
 sky130_fd_sc_hd__inv_2 _2861_ (.A(net13),
    .Y(_0008_));
 sky130_fd_sc_hd__inv_2 _2862_ (.A(net2),
    .Y(_0009_));
 sky130_fd_sc_hd__clkinv_2 _2863_ (.A(net3),
    .Y(_0010_));
 sky130_fd_sc_hd__inv_2 _2864_ (.A(net4),
    .Y(_0011_));
 sky130_fd_sc_hd__inv_2 _2865_ (.A(\as1802.regs[2][0] ),
    .Y(_2590_));
 sky130_fd_sc_hd__nor2_4 _2866_ (.A(_2579_),
    .B(_2484_),
    .Y(_2591_));
 sky130_fd_sc_hd__nand2_4 _2867_ (.A(_2526_),
    .B(_2591_),
    .Y(_2592_));
 sky130_fd_sc_hd__or3_2 _2868_ (.A(_2504_),
    .B(_2495_),
    .C(_2493_),
    .X(_2593_));
 sky130_fd_sc_hd__or2_2 _2869_ (.A(_2513_),
    .B(_2593_),
    .X(_2594_));
 sky130_fd_sc_hd__nor2_1 _2870_ (.A(_2592_),
    .B(_2594_),
    .Y(_2595_));
 sky130_fd_sc_hd__clkbuf_4 _2871_ (.A(_2595_),
    .X(_2596_));
 sky130_fd_sc_hd__clkbuf_4 _2872_ (.A(_2596_),
    .X(_2597_));
 sky130_fd_sc_hd__or2_2 _2873_ (.A(\as1802.instr_cycle[0] ),
    .B(_2484_),
    .X(_2598_));
 sky130_fd_sc_hd__or2_1 _2874_ (.A(_2533_),
    .B(_2500_),
    .X(_2599_));
 sky130_fd_sc_hd__nand2_4 _2875_ (.A(_2503_),
    .B(_2507_),
    .Y(_2600_));
 sky130_fd_sc_hd__o32a_1 _2876_ (.A1(_2495_),
    .A2(_2571_),
    .A3(_2599_),
    .B1(_2600_),
    .B2(_2555_),
    .X(_2601_));
 sky130_fd_sc_hd__nor4_4 _2877_ (.A(\as1802.instr_latch[1] ),
    .B(\as1802.instr_latch[0] ),
    .C(\as1802.instr_latch[2] ),
    .D(\as1802.cond_inv ),
    .Y(_2602_));
 sky130_fd_sc_hd__and2_1 _2878_ (.A(_2573_),
    .B(_2602_),
    .X(_2603_));
 sky130_fd_sc_hd__o21ba_1 _2879_ (.A1(_2553_),
    .A2(_2601_),
    .B1_N(_2603_),
    .X(_2604_));
 sky130_fd_sc_hd__or3_1 _2880_ (.A(_2533_),
    .B(_2511_),
    .C(_2592_),
    .X(_2605_));
 sky130_fd_sc_hd__clkbuf_4 _2881_ (.A(_2605_),
    .X(_2606_));
 sky130_fd_sc_hd__o21a_2 _2882_ (.A1(_2598_),
    .A2(_2604_),
    .B1(_2606_),
    .X(_2607_));
 sky130_fd_sc_hd__or2_1 _2883_ (.A(_2464_),
    .B(_2598_),
    .X(_2608_));
 sky130_fd_sc_hd__buf_2 _2884_ (.A(_2608_),
    .X(_2609_));
 sky130_fd_sc_hd__nand2_2 _2885_ (.A(_2486_),
    .B(_2547_),
    .Y(_2610_));
 sky130_fd_sc_hd__or3_1 _2886_ (.A(\as1802.instr_latch[5] ),
    .B(_2567_),
    .C(_2561_),
    .X(_2611_));
 sky130_fd_sc_hd__or4b_1 _2887_ (.A(\as1802.instr_latch[5] ),
    .B(\as1802.instr_latch[4] ),
    .C(\as1802.instr_latch[6] ),
    .D_N(\as1802.instr_latch[7] ),
    .X(_2612_));
 sky130_fd_sc_hd__or4_1 _2888_ (.A(\as1802.instr_cycle[0] ),
    .B(_2459_),
    .C(_2523_),
    .D(_2612_),
    .X(_2613_));
 sky130_fd_sc_hd__or4b_1 _2889_ (.A(\as1802.instr_cycle[0] ),
    .B(\as1802.instr_latch[5] ),
    .C(\as1802.instr_latch[7] ),
    .D_N(\as1802.instr_latch[6] ),
    .X(_2614_));
 sky130_fd_sc_hd__o31a_1 _2890_ (.A1(\as1802.instr_cycle[0] ),
    .A2(_2466_),
    .A3(_2602_),
    .B1(_2614_),
    .X(_2615_));
 sky130_fd_sc_hd__o211a_4 _2891_ (.A1(_2610_),
    .A2(_2611_),
    .B1(_2613_),
    .C1(_2615_),
    .X(_2616_));
 sky130_fd_sc_hd__nand3_4 _2892_ (.A(\as1802.X[0] ),
    .B(_2609_),
    .C(_2616_),
    .Y(_2617_));
 sky130_fd_sc_hd__a21o_2 _2893_ (.A1(_2609_),
    .A2(_2616_),
    .B1(_2513_),
    .X(_2618_));
 sky130_fd_sc_hd__nand2_4 _2894_ (.A(_2617_),
    .B(_2618_),
    .Y(_2619_));
 sky130_fd_sc_hd__buf_2 _2895_ (.A(_2619_),
    .X(_2620_));
 sky130_fd_sc_hd__buf_2 _2896_ (.A(_2617_),
    .X(_2621_));
 sky130_fd_sc_hd__buf_2 _2897_ (.A(_2618_),
    .X(_2622_));
 sky130_fd_sc_hd__and3_1 _2898_ (.A(\as1802.regs[4][0] ),
    .B(_2621_),
    .C(_2622_),
    .X(_2623_));
 sky130_fd_sc_hd__and3_1 _2899_ (.A(\as1802.X[1] ),
    .B(_2609_),
    .C(_2616_),
    .X(_2624_));
 sky130_fd_sc_hd__a21oi_1 _2900_ (.A1(_2609_),
    .A2(_2616_),
    .B1(_2527_),
    .Y(_2625_));
 sky130_fd_sc_hd__or2_1 _2901_ (.A(_2624_),
    .B(_2625_),
    .X(_2626_));
 sky130_fd_sc_hd__buf_2 _2902_ (.A(_2626_),
    .X(_2627_));
 sky130_fd_sc_hd__a211o_1 _2903_ (.A1(\as1802.regs[5][0] ),
    .A2(_2620_),
    .B1(_2623_),
    .C1(_2627_),
    .X(_2628_));
 sky130_fd_sc_hd__buf_2 _2904_ (.A(_2619_),
    .X(_2629_));
 sky130_fd_sc_hd__and3_1 _2905_ (.A(\as1802.regs[6][0] ),
    .B(_2621_),
    .C(_2622_),
    .X(_2630_));
 sky130_fd_sc_hd__nor2_1 _2906_ (.A(_2624_),
    .B(_2625_),
    .Y(_2631_));
 sky130_fd_sc_hd__clkbuf_4 _2907_ (.A(_2631_),
    .X(_2632_));
 sky130_fd_sc_hd__a211o_1 _2908_ (.A1(\as1802.regs[7][0] ),
    .A2(_2629_),
    .B1(_2630_),
    .C1(_2632_),
    .X(_2633_));
 sky130_fd_sc_hd__inv_2 _2909_ (.A(\as1802.X[2] ),
    .Y(_2634_));
 sky130_fd_sc_hd__nand2_2 _2910_ (.A(_2609_),
    .B(_2616_),
    .Y(_2635_));
 sky130_fd_sc_hd__mux2_1 _2911_ (.A0(_2634_),
    .A1(_2503_),
    .S(_2635_),
    .X(_2636_));
 sky130_fd_sc_hd__clkbuf_4 _2912_ (.A(_2636_),
    .X(_2637_));
 sky130_fd_sc_hd__a21oi_1 _2913_ (.A1(_2628_),
    .A2(_2633_),
    .B1(_2637_),
    .Y(_2638_));
 sky130_fd_sc_hd__mux2_1 _2914_ (.A0(\as1802.X[3] ),
    .A1(\as1802.cond_inv ),
    .S(_2635_),
    .X(_2639_));
 sky130_fd_sc_hd__buf_6 _2915_ (.A(_2639_),
    .X(_2640_));
 sky130_fd_sc_hd__and3_1 _2916_ (.A(\as1802.regs[0][0] ),
    .B(_2621_),
    .C(_2622_),
    .X(_2641_));
 sky130_fd_sc_hd__clkbuf_4 _2917_ (.A(_2627_),
    .X(_2642_));
 sky130_fd_sc_hd__a211o_1 _2918_ (.A1(\as1802.regs[1][0] ),
    .A2(_2620_),
    .B1(_2641_),
    .C1(_2642_),
    .X(_2643_));
 sky130_fd_sc_hd__and3_1 _2919_ (.A(\as1802.regs[2][0] ),
    .B(_2621_),
    .C(_2622_),
    .X(_2644_));
 sky130_fd_sc_hd__clkbuf_4 _2920_ (.A(_2631_),
    .X(_2645_));
 sky130_fd_sc_hd__a211o_1 _2921_ (.A1(\as1802.regs[3][0] ),
    .A2(_2620_),
    .B1(_2644_),
    .C1(_2645_),
    .X(_2646_));
 sky130_fd_sc_hd__mux2_2 _2922_ (.A0(\as1802.X[2] ),
    .A1(\as1802.instr_latch[2] ),
    .S(_2635_),
    .X(_2647_));
 sky130_fd_sc_hd__clkbuf_4 _2923_ (.A(_2647_),
    .X(_2648_));
 sky130_fd_sc_hd__a21oi_1 _2924_ (.A1(_2643_),
    .A2(_2646_),
    .B1(_2648_),
    .Y(_2649_));
 sky130_fd_sc_hd__and3_1 _2925_ (.A(\as1802.regs[12][0] ),
    .B(_2621_),
    .C(_2622_),
    .X(_2650_));
 sky130_fd_sc_hd__a211o_1 _2926_ (.A1(\as1802.regs[13][0] ),
    .A2(_2620_),
    .B1(_2650_),
    .C1(_2642_),
    .X(_2651_));
 sky130_fd_sc_hd__and3_1 _2927_ (.A(\as1802.regs[14][0] ),
    .B(_2621_),
    .C(_2622_),
    .X(_2652_));
 sky130_fd_sc_hd__a211o_1 _2928_ (.A1(\as1802.regs[15][0] ),
    .A2(_2620_),
    .B1(_2652_),
    .C1(_2645_),
    .X(_2653_));
 sky130_fd_sc_hd__a21oi_1 _2929_ (.A1(_2651_),
    .A2(_2653_),
    .B1(_2637_),
    .Y(_2654_));
 sky130_fd_sc_hd__clkbuf_2 _2930_ (.A(_2617_),
    .X(_2655_));
 sky130_fd_sc_hd__buf_2 _2931_ (.A(_2655_),
    .X(_2656_));
 sky130_fd_sc_hd__buf_2 _2932_ (.A(_2618_),
    .X(_2657_));
 sky130_fd_sc_hd__buf_2 _2933_ (.A(_2657_),
    .X(_2658_));
 sky130_fd_sc_hd__a21o_1 _2934_ (.A1(_2656_),
    .A2(_2658_),
    .B1(\as1802.regs[9][0] ),
    .X(_2659_));
 sky130_fd_sc_hd__o211a_1 _2935_ (.A1(\as1802.regs[8][0] ),
    .A2(_2620_),
    .B1(_2659_),
    .C1(_2645_),
    .X(_2660_));
 sky130_fd_sc_hd__a21o_1 _2936_ (.A1(_2656_),
    .A2(_2658_),
    .B1(\as1802.regs[11][0] ),
    .X(_2661_));
 sky130_fd_sc_hd__o211a_1 _2937_ (.A1(\as1802.regs[10][0] ),
    .A2(_2620_),
    .B1(_2661_),
    .C1(_2642_),
    .X(_2662_));
 sky130_fd_sc_hd__o31ai_1 _2938_ (.A1(_2648_),
    .A2(_2660_),
    .A3(_2662_),
    .B1(_2640_),
    .Y(_2663_));
 sky130_fd_sc_hd__o32a_1 _2939_ (.A1(_2638_),
    .A2(_2640_),
    .A3(_2649_),
    .B1(_2654_),
    .B2(_2663_),
    .X(_2664_));
 sky130_fd_sc_hd__clkbuf_4 _2940_ (.A(_2664_),
    .X(_2665_));
 sky130_fd_sc_hd__inv_2 _2941_ (.A(_0003_),
    .Y(_2666_));
 sky130_fd_sc_hd__buf_4 _2942_ (.A(_2666_),
    .X(_2667_));
 sky130_fd_sc_hd__buf_4 _2943_ (.A(_0000_),
    .X(_2668_));
 sky130_fd_sc_hd__buf_4 _2944_ (.A(_2668_),
    .X(_2669_));
 sky130_fd_sc_hd__buf_4 _2945_ (.A(_2669_),
    .X(_2670_));
 sky130_fd_sc_hd__clkbuf_4 _2946_ (.A(_0001_),
    .X(_2671_));
 sky130_fd_sc_hd__clkbuf_4 _2947_ (.A(_2671_),
    .X(_2672_));
 sky130_fd_sc_hd__clkbuf_4 _2948_ (.A(_2672_),
    .X(_2673_));
 sky130_fd_sc_hd__clkbuf_4 _2949_ (.A(_2673_),
    .X(_2674_));
 sky130_fd_sc_hd__mux4_1 _2950_ (.A0(\as1802.regs[0][0] ),
    .A1(\as1802.regs[1][0] ),
    .A2(\as1802.regs[2][0] ),
    .A3(\as1802.regs[3][0] ),
    .S0(_2670_),
    .S1(_2674_),
    .X(_2675_));
 sky130_fd_sc_hd__mux4_1 _2951_ (.A0(\as1802.regs[4][0] ),
    .A1(\as1802.regs[5][0] ),
    .A2(\as1802.regs[6][0] ),
    .A3(\as1802.regs[7][0] ),
    .S0(_2670_),
    .S1(_2673_),
    .X(_2676_));
 sky130_fd_sc_hd__buf_4 _2952_ (.A(_0002_),
    .X(_2677_));
 sky130_fd_sc_hd__buf_4 _2953_ (.A(_2677_),
    .X(_2678_));
 sky130_fd_sc_hd__mux2_1 _2954_ (.A0(_2675_),
    .A1(_2676_),
    .S(_2678_),
    .X(_2679_));
 sky130_fd_sc_hd__mux4_1 _2955_ (.A0(\as1802.regs[8][0] ),
    .A1(\as1802.regs[9][0] ),
    .A2(\as1802.regs[10][0] ),
    .A3(\as1802.regs[11][0] ),
    .S0(_2670_),
    .S1(_2674_),
    .X(_2680_));
 sky130_fd_sc_hd__buf_4 _2956_ (.A(_2670_),
    .X(_2681_));
 sky130_fd_sc_hd__inv_2 _2957_ (.A(\as1802.regs[13][0] ),
    .Y(_2682_));
 sky130_fd_sc_hd__clkbuf_4 _2958_ (.A(_2670_),
    .X(_2683_));
 sky130_fd_sc_hd__nor2_1 _2959_ (.A(_2683_),
    .B(\as1802.regs[12][0] ),
    .Y(_2684_));
 sky130_fd_sc_hd__clkbuf_4 _2960_ (.A(_2673_),
    .X(_2685_));
 sky130_fd_sc_hd__a211oi_1 _2961_ (.A1(_2681_),
    .A2(_2682_),
    .B1(_2684_),
    .C1(_2685_),
    .Y(_2686_));
 sky130_fd_sc_hd__mux2_1 _2962_ (.A0(\as1802.regs[14][0] ),
    .A1(\as1802.regs[15][0] ),
    .S(_2670_),
    .X(_2687_));
 sky130_fd_sc_hd__inv_2 _2963_ (.A(_0002_),
    .Y(_2688_));
 sky130_fd_sc_hd__buf_4 _2964_ (.A(_2688_),
    .X(_2689_));
 sky130_fd_sc_hd__a21o_1 _2965_ (.A1(_2685_),
    .A2(_2687_),
    .B1(_2689_),
    .X(_2690_));
 sky130_fd_sc_hd__buf_8 _2966_ (.A(_0003_),
    .X(_2691_));
 sky130_fd_sc_hd__o221ai_1 _2967_ (.A1(_2678_),
    .A2(_2680_),
    .B1(_2686_),
    .B2(_2690_),
    .C1(_2691_),
    .Y(_2692_));
 sky130_fd_sc_hd__a21bo_1 _2968_ (.A1(_2667_),
    .A2(_2679_),
    .B1_N(_2692_),
    .X(_2693_));
 sky130_fd_sc_hd__buf_4 _2969_ (.A(_2693_),
    .X(_2694_));
 sky130_fd_sc_hd__nand2_4 _2970_ (.A(_2533_),
    .B(_2694_),
    .Y(_2695_));
 sky130_fd_sc_hd__clkbuf_4 _2971_ (.A(_2694_),
    .X(_2696_));
 sky130_fd_sc_hd__or2_1 _2972_ (.A(_2533_),
    .B(_2696_),
    .X(_2697_));
 sky130_fd_sc_hd__and2_1 _2973_ (.A(_2695_),
    .B(_2697_),
    .X(_2698_));
 sky130_fd_sc_hd__or4b_2 _2974_ (.A(_2579_),
    .B(_2479_),
    .C(_2542_),
    .D_N(_2544_),
    .X(_2699_));
 sky130_fd_sc_hd__or2_2 _2975_ (.A(_2485_),
    .B(_2699_),
    .X(_2700_));
 sky130_fd_sc_hd__clkbuf_4 _2976_ (.A(_2700_),
    .X(_2701_));
 sky130_fd_sc_hd__buf_4 _2977_ (.A(io_out[0]),
    .X(_2702_));
 sky130_fd_sc_hd__or4bb_1 _2978_ (.A(_2473_),
    .B(_2474_),
    .C_N(\as1802.instr_latch[7] ),
    .D_N(_2477_),
    .X(_2703_));
 sky130_fd_sc_hd__clkbuf_4 _2979_ (.A(_2703_),
    .X(_2704_));
 sky130_fd_sc_hd__or2_1 _2980_ (.A(_2579_),
    .B(_2704_),
    .X(_2705_));
 sky130_fd_sc_hd__or4_2 _2981_ (.A(\as1802.instr_cycle[2] ),
    .B(_2484_),
    .C(_2471_),
    .D(_2705_),
    .X(_2706_));
 sky130_fd_sc_hd__nor2_1 _2982_ (.A(\as1802.instr_cycle[1] ),
    .B(_2706_),
    .Y(_2707_));
 sky130_fd_sc_hd__nor4_1 _2983_ (.A(_2579_),
    .B(\as1802.instr_cycle[2] ),
    .C(_2471_),
    .D(_2704_),
    .Y(_2708_));
 sky130_fd_sc_hd__or2b_1 _2984_ (.A(\as1802.instr_cycle[1] ),
    .B_N(_2708_),
    .X(_2709_));
 sky130_fd_sc_hd__nor2_2 _2985_ (.A(_2485_),
    .B(_2709_),
    .Y(_2710_));
 sky130_fd_sc_hd__nor2_1 _2986_ (.A(_2579_),
    .B(_2704_),
    .Y(_2711_));
 sky130_fd_sc_hd__mux2_2 _2987_ (.A0(_2495_),
    .A1(_2533_),
    .S(_2470_),
    .X(_2712_));
 sky130_fd_sc_hd__and2_1 _2988_ (.A(_2711_),
    .B(_2712_),
    .X(_2713_));
 sky130_fd_sc_hd__o31ai_2 _2989_ (.A1(_2535_),
    .A2(_2536_),
    .A3(_2539_),
    .B1(_2713_),
    .Y(_2714_));
 sky130_fd_sc_hd__nand2_1 _2990_ (.A(_2486_),
    .B(\as1802.instr_cycle[2] ),
    .Y(_2715_));
 sky130_fd_sc_hd__or3_1 _2991_ (.A(_2471_),
    .B(_2704_),
    .C(_2715_),
    .X(_2716_));
 sky130_fd_sc_hd__or4_2 _2992_ (.A(_2535_),
    .B(_2536_),
    .C(_2539_),
    .D(_2716_),
    .X(_2717_));
 sky130_fd_sc_hd__a21oi_4 _2993_ (.A1(_2714_),
    .A2(_2717_),
    .B1(_2484_),
    .Y(_2718_));
 sky130_fd_sc_hd__clkbuf_4 _2994_ (.A(_2718_),
    .X(_2719_));
 sky130_fd_sc_hd__inv_2 _2995_ (.A(_2694_),
    .Y(_2720_));
 sky130_fd_sc_hd__or3_1 _2996_ (.A(_2579_),
    .B(\as1802.instr_cycle[2] ),
    .C(_2522_),
    .X(_2721_));
 sky130_fd_sc_hd__or2_2 _2997_ (.A(_2484_),
    .B(_2721_),
    .X(_2722_));
 sky130_fd_sc_hd__mux2_1 _2998_ (.A0(_2702_),
    .A1(_2720_),
    .S(_2722_),
    .X(_0359_));
 sky130_fd_sc_hd__or2_1 _2999_ (.A(_2570_),
    .B(_2592_),
    .X(_0360_));
 sky130_fd_sc_hd__buf_2 _3000_ (.A(_0360_),
    .X(_0361_));
 sky130_fd_sc_hd__mux2_1 _3001_ (.A0(_2698_),
    .A1(_0359_),
    .S(_0361_),
    .X(_0362_));
 sky130_fd_sc_hd__xnor2_1 _3002_ (.A(_2719_),
    .B(_0362_),
    .Y(_0363_));
 sky130_fd_sc_hd__nor2_1 _3003_ (.A(_2710_),
    .B(_0363_),
    .Y(_0364_));
 sky130_fd_sc_hd__nor2_2 _3004_ (.A(_2485_),
    .B(_2699_),
    .Y(_0365_));
 sky130_fd_sc_hd__clkbuf_4 _3005_ (.A(_0365_),
    .X(_0366_));
 sky130_fd_sc_hd__a211o_1 _3006_ (.A1(_2702_),
    .A2(_2707_),
    .B1(_0364_),
    .C1(_0366_),
    .X(_0367_));
 sky130_fd_sc_hd__and3_1 _3007_ (.A(_2533_),
    .B(_2545_),
    .C(_2591_),
    .X(_0368_));
 sky130_fd_sc_hd__buf_2 _3008_ (.A(_0368_),
    .X(_0369_));
 sky130_fd_sc_hd__o211a_1 _3009_ (.A1(_2522_),
    .A2(_2715_),
    .B1(_2699_),
    .C1(_2490_),
    .X(_0370_));
 sky130_fd_sc_hd__o21ai_1 _3010_ (.A1(_2485_),
    .A2(_0370_),
    .B1(_0361_),
    .Y(_0371_));
 sky130_fd_sc_hd__nand2_1 _3011_ (.A(\as1802.instr_cycle[2] ),
    .B(_2711_),
    .Y(_0372_));
 sky130_fd_sc_hd__nor4b_4 _3012_ (.A(_2485_),
    .B(_2712_),
    .C(_0372_),
    .D_N(_2540_),
    .Y(_0373_));
 sky130_fd_sc_hd__or4_1 _3013_ (.A(_2718_),
    .B(_0369_),
    .C(_0371_),
    .D(_0373_),
    .X(_0374_));
 sky130_fd_sc_hd__nor2_2 _3014_ (.A(_2484_),
    .B(_2721_),
    .Y(_0375_));
 sky130_fd_sc_hd__or3_1 _3015_ (.A(_0374_),
    .B(_0375_),
    .C(_2710_),
    .X(_0376_));
 sky130_fd_sc_hd__inv_2 _3016_ (.A(_2706_),
    .Y(_0377_));
 sky130_fd_sc_hd__and2_1 _3017_ (.A(\as1802.instr_cycle[1] ),
    .B(_0377_),
    .X(_0378_));
 sky130_fd_sc_hd__or2_2 _3018_ (.A(_0376_),
    .B(_0378_),
    .X(_0379_));
 sky130_fd_sc_hd__buf_4 _3019_ (.A(_0379_),
    .X(_0380_));
 sky130_fd_sc_hd__o211a_1 _3020_ (.A1(_2698_),
    .A2(_2701_),
    .B1(_0367_),
    .C1(_0380_),
    .X(_0381_));
 sky130_fd_sc_hd__buf_4 _3021_ (.A(\as1802.D[0] ),
    .X(_0382_));
 sky130_fd_sc_hd__or2_2 _3022_ (.A(_2568_),
    .B(_2561_),
    .X(_0383_));
 sky130_fd_sc_hd__nor2_4 _3023_ (.A(_2598_),
    .B(_0383_),
    .Y(_0384_));
 sky130_fd_sc_hd__or3_2 _3024_ (.A(_2579_),
    .B(_2584_),
    .C(_2585_),
    .X(_0385_));
 sky130_fd_sc_hd__nor2_2 _3025_ (.A(net14),
    .B(_0385_),
    .Y(_0386_));
 sky130_fd_sc_hd__a21oi_1 _3026_ (.A1(_2464_),
    .A2(_2583_),
    .B1(_2598_),
    .Y(_0387_));
 sky130_fd_sc_hd__or2_2 _3027_ (.A(_0386_),
    .B(_0387_),
    .X(_0388_));
 sky130_fd_sc_hd__nor2_2 _3028_ (.A(_2592_),
    .B(_2601_),
    .Y(_0389_));
 sky130_fd_sc_hd__a21oi_4 _3029_ (.A1(_2591_),
    .A2(_2603_),
    .B1(_0389_),
    .Y(_0390_));
 sky130_fd_sc_hd__nand2_2 _3030_ (.A(_2606_),
    .B(_0390_),
    .Y(_0391_));
 sky130_fd_sc_hd__a221o_1 _3031_ (.A1(_0382_),
    .A2(_0384_),
    .B1(_0388_),
    .B2(_2665_),
    .C1(_0391_),
    .X(_0392_));
 sky130_fd_sc_hd__o22a_1 _3032_ (.A1(_2607_),
    .A2(_2665_),
    .B1(_0381_),
    .B2(_0392_),
    .X(_0393_));
 sky130_fd_sc_hd__a21o_1 _3033_ (.A1(_2590_),
    .A2(_2597_),
    .B1(_0393_),
    .X(_0394_));
 sky130_fd_sc_hd__buf_2 _3034_ (.A(_0394_),
    .X(_0395_));
 sky130_fd_sc_hd__or2_1 _3035_ (.A(_0384_),
    .B(_0388_),
    .X(_0396_));
 sky130_fd_sc_hd__buf_2 _3036_ (.A(_0396_),
    .X(_0397_));
 sky130_fd_sc_hd__a221o_1 _3037_ (.A1(_2504_),
    .A2(_0397_),
    .B1(_0391_),
    .B2(\as1802.X[1] ),
    .C1(_2595_),
    .X(_0398_));
 sky130_fd_sc_hd__a21oi_2 _3038_ (.A1(\as1802.P[1] ),
    .A2(_0380_),
    .B1(_0398_),
    .Y(_0399_));
 sky130_fd_sc_hd__a22o_1 _3039_ (.A1(\as1802.P[0] ),
    .A2(_0379_),
    .B1(_0397_),
    .B2(_2469_),
    .X(_0400_));
 sky130_fd_sc_hd__mux2_2 _3040_ (.A0(\as1802.X[0] ),
    .A1(_0400_),
    .S(_2607_),
    .X(_0401_));
 sky130_fd_sc_hd__and2b_1 _3041_ (.A_N(_0399_),
    .B(_0401_),
    .X(_0402_));
 sky130_fd_sc_hd__inv_2 _3042_ (.A(_2607_),
    .Y(_0403_));
 sky130_fd_sc_hd__a221o_1 _3043_ (.A1(\as1802.P[3] ),
    .A2(_0379_),
    .B1(_0397_),
    .B2(_2556_),
    .C1(_0403_),
    .X(_0404_));
 sky130_fd_sc_hd__o21ai_1 _3044_ (.A1(\as1802.X[3] ),
    .A2(_2607_),
    .B1(_0404_),
    .Y(_0405_));
 sky130_fd_sc_hd__a22o_1 _3045_ (.A1(\as1802.P[2] ),
    .A2(_0379_),
    .B1(_0397_),
    .B2(_2496_),
    .X(_0406_));
 sky130_fd_sc_hd__or2_1 _3046_ (.A(_0403_),
    .B(_0406_),
    .X(_0407_));
 sky130_fd_sc_hd__o21ai_1 _3047_ (.A1(\as1802.X[2] ),
    .A2(_2607_),
    .B1(_0407_),
    .Y(_0408_));
 sky130_fd_sc_hd__nor2_2 _3048_ (.A(_0405_),
    .B(_0408_),
    .Y(_0409_));
 sky130_fd_sc_hd__or4_1 _3049_ (.A(_2456_),
    .B(_0376_),
    .C(_0384_),
    .D(_0387_),
    .X(_0410_));
 sky130_fd_sc_hd__or3_2 _3050_ (.A(_2596_),
    .B(_0391_),
    .C(_0410_),
    .X(_0411_));
 sky130_fd_sc_hd__and3_1 _3051_ (.A(_0402_),
    .B(_0409_),
    .C(_0411_),
    .X(_0412_));
 sky130_fd_sc_hd__buf_4 _3052_ (.A(_0412_),
    .X(_0413_));
 sky130_fd_sc_hd__mux2_1 _3053_ (.A0(\as1802.regs[15][0] ),
    .A1(_0395_),
    .S(_0413_),
    .X(_0414_));
 sky130_fd_sc_hd__clkbuf_1 _3054_ (.A(_0414_),
    .X(_0012_));
 sky130_fd_sc_hd__or2_2 _3055_ (.A(_2592_),
    .B(_2594_),
    .X(_0415_));
 sky130_fd_sc_hd__clkbuf_4 _3056_ (.A(_0415_),
    .X(_0416_));
 sky130_fd_sc_hd__and2_1 _3057_ (.A(\as1802.regs[2][0] ),
    .B(\as1802.regs[2][1] ),
    .X(_0417_));
 sky130_fd_sc_hd__nor2_1 _3058_ (.A(\as1802.regs[2][0] ),
    .B(\as1802.regs[2][1] ),
    .Y(_0418_));
 sky130_fd_sc_hd__mux2_1 _3059_ (.A0(\as1802.regs[6][1] ),
    .A1(\as1802.regs[7][1] ),
    .S(_2619_),
    .X(_0419_));
 sky130_fd_sc_hd__clkbuf_4 _3060_ (.A(_2619_),
    .X(_0420_));
 sky130_fd_sc_hd__and3_1 _3061_ (.A(\as1802.regs[4][1] ),
    .B(_2617_),
    .C(_2618_),
    .X(_0421_));
 sky130_fd_sc_hd__a211o_1 _3062_ (.A1(\as1802.regs[5][1] ),
    .A2(_0420_),
    .B1(_0421_),
    .C1(_2627_),
    .X(_0422_));
 sky130_fd_sc_hd__o211a_1 _3063_ (.A1(_2645_),
    .A2(_0419_),
    .B1(_0422_),
    .C1(_2647_),
    .X(_0423_));
 sky130_fd_sc_hd__mux2_1 _3064_ (.A0(\as1802.regs[0][1] ),
    .A1(\as1802.regs[1][1] ),
    .S(_2619_),
    .X(_0424_));
 sky130_fd_sc_hd__and3_1 _3065_ (.A(\as1802.regs[2][1] ),
    .B(_2617_),
    .C(_2618_),
    .X(_0425_));
 sky130_fd_sc_hd__a211o_1 _3066_ (.A1(\as1802.regs[3][1] ),
    .A2(_0420_),
    .B1(_0425_),
    .C1(_2632_),
    .X(_0426_));
 sky130_fd_sc_hd__o211a_1 _3067_ (.A1(_2642_),
    .A2(_0424_),
    .B1(_0426_),
    .C1(_2636_),
    .X(_0427_));
 sky130_fd_sc_hd__mux2_1 _3068_ (.A0(\as1802.regs[8][1] ),
    .A1(\as1802.regs[9][1] ),
    .S(_2619_),
    .X(_0428_));
 sky130_fd_sc_hd__and3_1 _3069_ (.A(\as1802.regs[10][1] ),
    .B(_2655_),
    .C(_2657_),
    .X(_0429_));
 sky130_fd_sc_hd__a211o_1 _3070_ (.A1(\as1802.regs[11][1] ),
    .A2(_2629_),
    .B1(_0429_),
    .C1(_2632_),
    .X(_0430_));
 sky130_fd_sc_hd__o211a_1 _3071_ (.A1(_2642_),
    .A2(_0428_),
    .B1(_0430_),
    .C1(_2637_),
    .X(_0431_));
 sky130_fd_sc_hd__and3_1 _3072_ (.A(\as1802.regs[12][1] ),
    .B(_2655_),
    .C(_2657_),
    .X(_0432_));
 sky130_fd_sc_hd__a211o_1 _3073_ (.A1(\as1802.regs[13][1] ),
    .A2(_0420_),
    .B1(_0432_),
    .C1(_2627_),
    .X(_0433_));
 sky130_fd_sc_hd__and3_1 _3074_ (.A(\as1802.regs[14][1] ),
    .B(_2655_),
    .C(_2657_),
    .X(_0434_));
 sky130_fd_sc_hd__a211o_1 _3075_ (.A1(\as1802.regs[15][1] ),
    .A2(_0420_),
    .B1(_0434_),
    .C1(_2632_),
    .X(_0435_));
 sky130_fd_sc_hd__inv_2 _3076_ (.A(\as1802.X[3] ),
    .Y(_0436_));
 sky130_fd_sc_hd__mux2_8 _3077_ (.A0(_0436_),
    .A1(_2492_),
    .S(_2635_),
    .X(_0437_));
 sky130_fd_sc_hd__a31o_1 _3078_ (.A1(_2647_),
    .A2(_0433_),
    .A3(_0435_),
    .B1(_0437_),
    .X(_0438_));
 sky130_fd_sc_hd__o32ai_4 _3079_ (.A1(_2640_),
    .A2(_0423_),
    .A3(_0427_),
    .B1(_0431_),
    .B2(_0438_),
    .Y(_0439_));
 sky130_fd_sc_hd__nor2_1 _3080_ (.A(_2665_),
    .B(_0439_),
    .Y(_0440_));
 sky130_fd_sc_hd__nand2_1 _3081_ (.A(_2665_),
    .B(_0439_),
    .Y(_0441_));
 sky130_fd_sc_hd__and2b_1 _3082_ (.A_N(_0440_),
    .B(_0441_),
    .X(_0442_));
 sky130_fd_sc_hd__or3_1 _3083_ (.A(_2579_),
    .B(_2476_),
    .C(_2568_),
    .X(_0443_));
 sky130_fd_sc_hd__or2_2 _3084_ (.A(_2477_),
    .B(_0443_),
    .X(_0444_));
 sky130_fd_sc_hd__or2_1 _3085_ (.A(_2485_),
    .B(_0444_),
    .X(_0445_));
 sky130_fd_sc_hd__buf_2 _3086_ (.A(_0445_),
    .X(_0446_));
 sky130_fd_sc_hd__clkbuf_4 _3087_ (.A(_0446_),
    .X(_0447_));
 sky130_fd_sc_hd__nand2_1 _3088_ (.A(_2493_),
    .B(_2516_),
    .Y(_0448_));
 sky130_fd_sc_hd__nor2_1 _3089_ (.A(_2580_),
    .B(_0448_),
    .Y(_0449_));
 sky130_fd_sc_hd__a31o_2 _3090_ (.A1(_2467_),
    .A2(_2573_),
    .A3(_0449_),
    .B1(_0389_),
    .X(_0450_));
 sky130_fd_sc_hd__a21o_1 _3091_ (.A1(_0388_),
    .A2(_0447_),
    .B1(_0450_),
    .X(_0451_));
 sky130_fd_sc_hd__buf_4 _3092_ (.A(\as1802.D[1] ),
    .X(_0452_));
 sky130_fd_sc_hd__buf_4 _3093_ (.A(_2555_),
    .X(_0453_));
 sky130_fd_sc_hd__nor3_4 _3094_ (.A(_0453_),
    .B(_2511_),
    .C(_2592_),
    .Y(_0454_));
 sky130_fd_sc_hd__nor2_4 _3095_ (.A(_2485_),
    .B(_0444_),
    .Y(_0455_));
 sky130_fd_sc_hd__nor2_1 _3096_ (.A(_0454_),
    .B(_0455_),
    .Y(_0456_));
 sky130_fd_sc_hd__nor2_1 _3097_ (.A(_0442_),
    .B(_0456_),
    .Y(_0457_));
 sky130_fd_sc_hd__clkbuf_4 _3098_ (.A(_0000_),
    .X(_0458_));
 sky130_fd_sc_hd__and2b_1 _3099_ (.A_N(_0458_),
    .B(\as1802.regs[10][1] ),
    .X(_0459_));
 sky130_fd_sc_hd__a21bo_1 _3100_ (.A1(_0458_),
    .A2(\as1802.regs[11][1] ),
    .B1_N(_2671_),
    .X(_0460_));
 sky130_fd_sc_hd__mux2_1 _3101_ (.A0(\as1802.regs[8][1] ),
    .A1(\as1802.regs[9][1] ),
    .S(_0458_),
    .X(_0461_));
 sky130_fd_sc_hd__o221a_1 _3102_ (.A1(_0459_),
    .A2(_0460_),
    .B1(_0461_),
    .B2(_2672_),
    .C1(_2689_),
    .X(_0462_));
 sky130_fd_sc_hd__mux4_1 _3103_ (.A0(\as1802.regs[12][1] ),
    .A1(\as1802.regs[13][1] ),
    .A2(\as1802.regs[14][1] ),
    .A3(\as1802.regs[15][1] ),
    .S0(_2668_),
    .S1(_2671_),
    .X(_0463_));
 sky130_fd_sc_hd__a21o_1 _3104_ (.A1(_2677_),
    .A2(_0463_),
    .B1(_2666_),
    .X(_0464_));
 sky130_fd_sc_hd__mux4_1 _3105_ (.A0(\as1802.regs[0][1] ),
    .A1(\as1802.regs[1][1] ),
    .A2(\as1802.regs[2][1] ),
    .A3(\as1802.regs[3][1] ),
    .S0(_2668_),
    .S1(_2671_),
    .X(_0465_));
 sky130_fd_sc_hd__mux4_1 _3106_ (.A0(\as1802.regs[4][1] ),
    .A1(\as1802.regs[5][1] ),
    .A2(\as1802.regs[6][1] ),
    .A3(\as1802.regs[7][1] ),
    .S0(_2668_),
    .S1(_0001_),
    .X(_0466_));
 sky130_fd_sc_hd__mux2_1 _3107_ (.A0(_0465_),
    .A1(_0466_),
    .S(_2677_),
    .X(_0467_));
 sky130_fd_sc_hd__o22a_1 _3108_ (.A1(_0462_),
    .A2(_0464_),
    .B1(_0467_),
    .B2(_0003_),
    .X(_0468_));
 sky130_fd_sc_hd__buf_2 _3109_ (.A(_0468_),
    .X(_0469_));
 sky130_fd_sc_hd__nand2_1 _3110_ (.A(_2695_),
    .B(_0469_),
    .Y(_0470_));
 sky130_fd_sc_hd__or2_1 _3111_ (.A(_2695_),
    .B(_0469_),
    .X(_0471_));
 sky130_fd_sc_hd__nand2_1 _3112_ (.A(_0470_),
    .B(_0471_),
    .Y(_0472_));
 sky130_fd_sc_hd__a21o_2 _3113_ (.A1(_2714_),
    .A2(_2717_),
    .B1(_2485_),
    .X(_0473_));
 sky130_fd_sc_hd__buf_4 _3114_ (.A(io_out[1]),
    .X(_0474_));
 sky130_fd_sc_hd__xor2_1 _3115_ (.A(_2694_),
    .B(_0469_),
    .X(_0475_));
 sky130_fd_sc_hd__mux2_1 _3116_ (.A0(_0474_),
    .A1(_0475_),
    .S(_2722_),
    .X(_0476_));
 sky130_fd_sc_hd__mux2_1 _3117_ (.A0(_0472_),
    .A1(_0476_),
    .S(_0361_),
    .X(_0477_));
 sky130_fd_sc_hd__nor2_1 _3118_ (.A(_0473_),
    .B(_0469_),
    .Y(_0478_));
 sky130_fd_sc_hd__a211o_1 _3119_ (.A1(_0473_),
    .A2(_0477_),
    .B1(_0478_),
    .C1(_2707_),
    .X(_0479_));
 sky130_fd_sc_hd__or2_2 _3120_ (.A(\as1802.instr_cycle[1] ),
    .B(_2706_),
    .X(_0480_));
 sky130_fd_sc_hd__or2_1 _3121_ (.A(_0474_),
    .B(_0480_),
    .X(_0481_));
 sky130_fd_sc_hd__a21o_1 _3122_ (.A1(_0479_),
    .A2(_0481_),
    .B1(_0365_),
    .X(_0482_));
 sky130_fd_sc_hd__o211a_1 _3123_ (.A1(_2701_),
    .A2(_0472_),
    .B1(_0482_),
    .C1(_0379_),
    .X(_0483_));
 sky130_fd_sc_hd__a2111o_1 _3124_ (.A1(_0452_),
    .A2(_0384_),
    .B1(_2596_),
    .C1(_0457_),
    .D1(_0483_),
    .X(_0484_));
 sky130_fd_sc_hd__a21o_1 _3125_ (.A1(_0442_),
    .A2(_0451_),
    .B1(_0484_),
    .X(_0485_));
 sky130_fd_sc_hd__o31a_2 _3126_ (.A1(_0416_),
    .A2(_0417_),
    .A3(_0418_),
    .B1(_0485_),
    .X(_0486_));
 sky130_fd_sc_hd__buf_2 _3127_ (.A(_0486_),
    .X(_0487_));
 sky130_fd_sc_hd__mux2_1 _3128_ (.A0(\as1802.regs[15][1] ),
    .A1(_0487_),
    .S(_0413_),
    .X(_0488_));
 sky130_fd_sc_hd__clkbuf_1 _3129_ (.A(_0488_),
    .X(_0013_));
 sky130_fd_sc_hd__inv_2 _3130_ (.A(_0450_),
    .Y(_0489_));
 sky130_fd_sc_hd__mux2_1 _3131_ (.A0(\as1802.regs[12][2] ),
    .A1(\as1802.regs[13][2] ),
    .S(_2619_),
    .X(_0490_));
 sky130_fd_sc_hd__and3_1 _3132_ (.A(\as1802.regs[14][2] ),
    .B(_2617_),
    .C(_2618_),
    .X(_0491_));
 sky130_fd_sc_hd__a211o_1 _3133_ (.A1(\as1802.regs[15][2] ),
    .A2(_0420_),
    .B1(_0491_),
    .C1(_2631_),
    .X(_0492_));
 sky130_fd_sc_hd__o211a_1 _3134_ (.A1(_2642_),
    .A2(_0490_),
    .B1(_0492_),
    .C1(_2647_),
    .X(_0493_));
 sky130_fd_sc_hd__mux2_1 _3135_ (.A0(\as1802.regs[8][2] ),
    .A1(\as1802.regs[9][2] ),
    .S(_2619_),
    .X(_0494_));
 sky130_fd_sc_hd__and3_1 _3136_ (.A(\as1802.regs[10][2] ),
    .B(_2617_),
    .C(_2618_),
    .X(_0495_));
 sky130_fd_sc_hd__a211o_1 _3137_ (.A1(\as1802.regs[11][2] ),
    .A2(_0420_),
    .B1(_0495_),
    .C1(_2632_),
    .X(_0496_));
 sky130_fd_sc_hd__o211a_1 _3138_ (.A1(_2642_),
    .A2(_0494_),
    .B1(_0496_),
    .C1(_2636_),
    .X(_0497_));
 sky130_fd_sc_hd__mux2_1 _3139_ (.A0(\as1802.regs[0][2] ),
    .A1(\as1802.regs[1][2] ),
    .S(_2619_),
    .X(_0498_));
 sky130_fd_sc_hd__and3_1 _3140_ (.A(\as1802.regs[2][2] ),
    .B(_2655_),
    .C(_2657_),
    .X(_0499_));
 sky130_fd_sc_hd__a211o_1 _3141_ (.A1(\as1802.regs[3][2] ),
    .A2(_0420_),
    .B1(_0499_),
    .C1(_2632_),
    .X(_0500_));
 sky130_fd_sc_hd__o211a_1 _3142_ (.A1(_2642_),
    .A2(_0498_),
    .B1(_0500_),
    .C1(_2636_),
    .X(_0501_));
 sky130_fd_sc_hd__and3_1 _3143_ (.A(\as1802.regs[4][2] ),
    .B(_2655_),
    .C(_2657_),
    .X(_0502_));
 sky130_fd_sc_hd__a211o_1 _3144_ (.A1(\as1802.regs[5][2] ),
    .A2(_0420_),
    .B1(_0502_),
    .C1(_2627_),
    .X(_0503_));
 sky130_fd_sc_hd__and3_1 _3145_ (.A(\as1802.regs[6][2] ),
    .B(_2655_),
    .C(_2657_),
    .X(_0504_));
 sky130_fd_sc_hd__a211o_1 _3146_ (.A1(\as1802.regs[7][2] ),
    .A2(_0420_),
    .B1(_0504_),
    .C1(_2632_),
    .X(_0505_));
 sky130_fd_sc_hd__a31o_1 _3147_ (.A1(_2647_),
    .A2(_0503_),
    .A3(_0505_),
    .B1(_2640_),
    .X(_0506_));
 sky130_fd_sc_hd__o32ai_4 _3148_ (.A1(_0437_),
    .A2(_0493_),
    .A3(_0497_),
    .B1(_0501_),
    .B2(_0506_),
    .Y(_0507_));
 sky130_fd_sc_hd__xor2_1 _3149_ (.A(_0440_),
    .B(_0507_),
    .X(_0508_));
 sky130_fd_sc_hd__mux4_1 _3150_ (.A0(\as1802.regs[12][2] ),
    .A1(\as1802.regs[13][2] ),
    .A2(\as1802.regs[14][2] ),
    .A3(\as1802.regs[15][2] ),
    .S0(_2668_),
    .S1(_2671_),
    .X(_0509_));
 sky130_fd_sc_hd__nand2_1 _3151_ (.A(_2677_),
    .B(_0509_),
    .Y(_0510_));
 sky130_fd_sc_hd__and2b_1 _3152_ (.A_N(_0458_),
    .B(\as1802.regs[10][2] ),
    .X(_0511_));
 sky130_fd_sc_hd__a21bo_1 _3153_ (.A1(_2669_),
    .A2(\as1802.regs[11][2] ),
    .B1_N(_2671_),
    .X(_0512_));
 sky130_fd_sc_hd__mux2_1 _3154_ (.A0(\as1802.regs[8][2] ),
    .A1(\as1802.regs[9][2] ),
    .S(_0458_),
    .X(_0513_));
 sky130_fd_sc_hd__o221ai_4 _3155_ (.A1(_0511_),
    .A2(_0512_),
    .B1(_0513_),
    .B2(_2672_),
    .C1(_2689_),
    .Y(_0514_));
 sky130_fd_sc_hd__mux4_1 _3156_ (.A0(\as1802.regs[0][2] ),
    .A1(\as1802.regs[1][2] ),
    .A2(\as1802.regs[2][2] ),
    .A3(\as1802.regs[3][2] ),
    .S0(_0458_),
    .S1(_2671_),
    .X(_0515_));
 sky130_fd_sc_hd__nand2_1 _3157_ (.A(_2689_),
    .B(_0515_),
    .Y(_0516_));
 sky130_fd_sc_hd__mux4_1 _3158_ (.A0(\as1802.regs[4][2] ),
    .A1(\as1802.regs[5][2] ),
    .A2(\as1802.regs[6][2] ),
    .A3(\as1802.regs[7][2] ),
    .S0(_2668_),
    .S1(_2671_),
    .X(_0517_));
 sky130_fd_sc_hd__a21oi_2 _3159_ (.A1(_2677_),
    .A2(_0517_),
    .B1(_0003_),
    .Y(_0518_));
 sky130_fd_sc_hd__a32oi_4 _3160_ (.A1(_0003_),
    .A2(_0510_),
    .A3(_0514_),
    .B1(_0516_),
    .B2(_0518_),
    .Y(_0519_));
 sky130_fd_sc_hd__and2_1 _3161_ (.A(_0468_),
    .B(_0519_),
    .X(_0520_));
 sky130_fd_sc_hd__a21oi_1 _3162_ (.A1(_2694_),
    .A2(_0469_),
    .B1(_0519_),
    .Y(_0521_));
 sky130_fd_sc_hd__a21o_1 _3163_ (.A1(_2694_),
    .A2(_0520_),
    .B1(_0521_),
    .X(_0522_));
 sky130_fd_sc_hd__a32o_1 _3164_ (.A1(_2691_),
    .A2(_0510_),
    .A3(_0514_),
    .B1(_0516_),
    .B2(_0518_),
    .X(_0523_));
 sky130_fd_sc_hd__nor2_1 _3165_ (.A(_0469_),
    .B(_0519_),
    .Y(_0524_));
 sky130_fd_sc_hd__or2_1 _3166_ (.A(_0520_),
    .B(_0524_),
    .X(_0525_));
 sky130_fd_sc_hd__mux2_1 _3167_ (.A0(_0523_),
    .A1(_0525_),
    .S(_0470_),
    .X(_0526_));
 sky130_fd_sc_hd__clkinv_2 _3168_ (.A(io_out[2]),
    .Y(_0527_));
 sky130_fd_sc_hd__mux2_1 _3169_ (.A0(_0527_),
    .A1(_0522_),
    .S(_2722_),
    .X(_0528_));
 sky130_fd_sc_hd__nor2_4 _3170_ (.A(_2570_),
    .B(_2592_),
    .Y(_0529_));
 sky130_fd_sc_hd__mux2_1 _3171_ (.A0(_0528_),
    .A1(_0526_),
    .S(_0529_),
    .X(_0530_));
 sky130_fd_sc_hd__or2_1 _3172_ (.A(_0473_),
    .B(_0525_),
    .X(_0531_));
 sky130_fd_sc_hd__o211a_1 _3173_ (.A1(_2719_),
    .A2(_0530_),
    .B1(_0531_),
    .C1(_0480_),
    .X(_0532_));
 sky130_fd_sc_hd__a211o_1 _3174_ (.A1(_0527_),
    .A2(_2707_),
    .B1(_0365_),
    .C1(_0532_),
    .X(_0533_));
 sky130_fd_sc_hd__nand3_2 _3175_ (.A(_0453_),
    .B(_2545_),
    .C(_2591_),
    .Y(_0534_));
 sky130_fd_sc_hd__o211a_1 _3176_ (.A1(_2701_),
    .A2(_0526_),
    .B1(_0533_),
    .C1(_0534_),
    .X(_0535_));
 sky130_fd_sc_hd__buf_2 _3177_ (.A(_0378_),
    .X(_0536_));
 sky130_fd_sc_hd__nor2_2 _3178_ (.A(_0376_),
    .B(_0536_),
    .Y(_0537_));
 sky130_fd_sc_hd__a211o_1 _3179_ (.A1(_0369_),
    .A2(_0522_),
    .B1(_0535_),
    .C1(_0537_),
    .X(_0538_));
 sky130_fd_sc_hd__buf_4 _3180_ (.A(\as1802.D[2] ),
    .X(_0539_));
 sky130_fd_sc_hd__a21oi_1 _3181_ (.A1(_0539_),
    .A2(_0384_),
    .B1(_2596_),
    .Y(_0540_));
 sky130_fd_sc_hd__o211a_1 _3182_ (.A1(_0489_),
    .A2(_0508_),
    .B1(_0538_),
    .C1(_0540_),
    .X(_0541_));
 sky130_fd_sc_hd__inv_2 _3183_ (.A(_0388_),
    .Y(_0542_));
 sky130_fd_sc_hd__xnor2_1 _3184_ (.A(_0441_),
    .B(_0507_),
    .Y(_0543_));
 sky130_fd_sc_hd__o32a_1 _3185_ (.A1(_0542_),
    .A2(_0455_),
    .A3(_0508_),
    .B1(_0543_),
    .B2(_0456_),
    .X(_0544_));
 sky130_fd_sc_hd__o21ai_1 _3186_ (.A1(\as1802.regs[2][0] ),
    .A2(\as1802.regs[2][1] ),
    .B1(\as1802.regs[2][2] ),
    .Y(_0545_));
 sky130_fd_sc_hd__or3_1 _3187_ (.A(\as1802.regs[2][0] ),
    .B(\as1802.regs[2][1] ),
    .C(\as1802.regs[2][2] ),
    .X(_0546_));
 sky130_fd_sc_hd__and3_1 _3188_ (.A(_2597_),
    .B(_0545_),
    .C(_0546_),
    .X(_0547_));
 sky130_fd_sc_hd__a21oi_4 _3189_ (.A1(_0541_),
    .A2(_0544_),
    .B1(_0547_),
    .Y(_0548_));
 sky130_fd_sc_hd__buf_2 _3190_ (.A(_0548_),
    .X(_0549_));
 sky130_fd_sc_hd__mux2_1 _3191_ (.A0(\as1802.regs[15][2] ),
    .A1(_0549_),
    .S(_0413_),
    .X(_0550_));
 sky130_fd_sc_hd__clkbuf_1 _3192_ (.A(_0550_),
    .X(_0014_));
 sky130_fd_sc_hd__mux2_1 _3193_ (.A0(\as1802.regs[6][3] ),
    .A1(\as1802.regs[7][3] ),
    .S(_0420_),
    .X(_0551_));
 sky130_fd_sc_hd__and3_1 _3194_ (.A(\as1802.regs[4][3] ),
    .B(_2655_),
    .C(_2657_),
    .X(_0552_));
 sky130_fd_sc_hd__a211o_1 _3195_ (.A1(\as1802.regs[5][3] ),
    .A2(_2629_),
    .B1(_0552_),
    .C1(_2627_),
    .X(_0553_));
 sky130_fd_sc_hd__o211a_1 _3196_ (.A1(_2645_),
    .A2(_0551_),
    .B1(_0553_),
    .C1(_2648_),
    .X(_0554_));
 sky130_fd_sc_hd__and3_1 _3197_ (.A(\as1802.regs[0][3] ),
    .B(_2655_),
    .C(_2657_),
    .X(_0555_));
 sky130_fd_sc_hd__a211o_1 _3198_ (.A1(\as1802.regs[1][3] ),
    .A2(_2629_),
    .B1(_0555_),
    .C1(_2627_),
    .X(_0556_));
 sky130_fd_sc_hd__and3_1 _3199_ (.A(\as1802.regs[2][3] ),
    .B(_2655_),
    .C(_2657_),
    .X(_0557_));
 sky130_fd_sc_hd__a211o_1 _3200_ (.A1(\as1802.regs[3][3] ),
    .A2(_2629_),
    .B1(_0557_),
    .C1(_2632_),
    .X(_0558_));
 sky130_fd_sc_hd__a31o_1 _3201_ (.A1(_2637_),
    .A2(_0556_),
    .A3(_0558_),
    .B1(_2640_),
    .X(_0559_));
 sky130_fd_sc_hd__clkbuf_4 _3202_ (.A(_2627_),
    .X(_0560_));
 sky130_fd_sc_hd__mux2_1 _3203_ (.A0(\as1802.regs[12][3] ),
    .A1(\as1802.regs[13][3] ),
    .S(_2629_),
    .X(_0561_));
 sky130_fd_sc_hd__and3_1 _3204_ (.A(\as1802.regs[14][3] ),
    .B(_2621_),
    .C(_2622_),
    .X(_0562_));
 sky130_fd_sc_hd__a211o_1 _3205_ (.A1(\as1802.regs[15][3] ),
    .A2(_2629_),
    .B1(_0562_),
    .C1(_2632_),
    .X(_0563_));
 sky130_fd_sc_hd__o211a_1 _3206_ (.A1(_0560_),
    .A2(_0561_),
    .B1(_0563_),
    .C1(_2648_),
    .X(_0564_));
 sky130_fd_sc_hd__and3_1 _3207_ (.A(\as1802.regs[10][3] ),
    .B(_2621_),
    .C(_2622_),
    .X(_0565_));
 sky130_fd_sc_hd__a211o_1 _3208_ (.A1(\as1802.regs[11][3] ),
    .A2(_2629_),
    .B1(_0565_),
    .C1(_2632_),
    .X(_0566_));
 sky130_fd_sc_hd__and3_1 _3209_ (.A(\as1802.regs[8][3] ),
    .B(_2621_),
    .C(_2622_),
    .X(_0567_));
 sky130_fd_sc_hd__a211o_1 _3210_ (.A1(\as1802.regs[9][3] ),
    .A2(_2629_),
    .B1(_0567_),
    .C1(_2627_),
    .X(_0568_));
 sky130_fd_sc_hd__a31o_1 _3211_ (.A1(_2637_),
    .A2(_0566_),
    .A3(_0568_),
    .B1(_0437_),
    .X(_0569_));
 sky130_fd_sc_hd__o22ai_4 _3212_ (.A1(_0554_),
    .A2(_0559_),
    .B1(_0564_),
    .B2(_0569_),
    .Y(_0570_));
 sky130_fd_sc_hd__and4_2 _3213_ (.A(_2664_),
    .B(_0439_),
    .C(_0507_),
    .D(_0570_),
    .X(_0571_));
 sky130_fd_sc_hd__a31o_1 _3214_ (.A1(_2665_),
    .A2(_0439_),
    .A3(_0507_),
    .B1(_0570_),
    .X(_0572_));
 sky130_fd_sc_hd__and2b_1 _3215_ (.A_N(_0571_),
    .B(_0572_),
    .X(_0573_));
 sky130_fd_sc_hd__nor2_1 _3216_ (.A(_2606_),
    .B(_0573_),
    .Y(_0574_));
 sky130_fd_sc_hd__a31o_4 _3217_ (.A1(_2573_),
    .A2(_2591_),
    .A3(_2602_),
    .B1(_0389_),
    .X(_0575_));
 sky130_fd_sc_hd__or4_1 _3218_ (.A(_2664_),
    .B(_0439_),
    .C(_0507_),
    .D(_0570_),
    .X(_0576_));
 sky130_fd_sc_hd__o31ai_1 _3219_ (.A1(_2665_),
    .A2(_0439_),
    .A3(_0507_),
    .B1(_0570_),
    .Y(_0577_));
 sky130_fd_sc_hd__and2_1 _3220_ (.A(_0576_),
    .B(_0577_),
    .X(_0578_));
 sky130_fd_sc_hd__buf_4 _3221_ (.A(\as1802.D[3] ),
    .X(_0579_));
 sky130_fd_sc_hd__or2_2 _3222_ (.A(_2598_),
    .B(_0383_),
    .X(_0580_));
 sky130_fd_sc_hd__nor2_1 _3223_ (.A(_0446_),
    .B(_0573_),
    .Y(_0581_));
 sky130_fd_sc_hd__a211o_1 _3224_ (.A1(_0446_),
    .A2(_0578_),
    .B1(_0581_),
    .C1(_0384_),
    .X(_0582_));
 sky130_fd_sc_hd__o211a_1 _3225_ (.A1(_0579_),
    .A2(_0580_),
    .B1(_0397_),
    .C1(_0582_),
    .X(_0583_));
 sky130_fd_sc_hd__and2b_1 _3226_ (.A_N(_0458_),
    .B(\as1802.regs[10][3] ),
    .X(_0584_));
 sky130_fd_sc_hd__a21bo_1 _3227_ (.A1(_0458_),
    .A2(\as1802.regs[11][3] ),
    .B1_N(_0001_),
    .X(_0585_));
 sky130_fd_sc_hd__mux2_1 _3228_ (.A0(\as1802.regs[8][3] ),
    .A1(\as1802.regs[9][3] ),
    .S(_2668_),
    .X(_0586_));
 sky130_fd_sc_hd__o221a_1 _3229_ (.A1(_0584_),
    .A2(_0585_),
    .B1(_0586_),
    .B2(_2672_),
    .C1(_2688_),
    .X(_0587_));
 sky130_fd_sc_hd__mux4_1 _3230_ (.A0(\as1802.regs[12][3] ),
    .A1(\as1802.regs[13][3] ),
    .A2(\as1802.regs[14][3] ),
    .A3(\as1802.regs[15][3] ),
    .S0(_2668_),
    .S1(_2671_),
    .X(_0588_));
 sky130_fd_sc_hd__a21o_1 _3231_ (.A1(_2677_),
    .A2(_0588_),
    .B1(_2666_),
    .X(_0589_));
 sky130_fd_sc_hd__mux4_1 _3232_ (.A0(\as1802.regs[0][3] ),
    .A1(\as1802.regs[1][3] ),
    .A2(\as1802.regs[2][3] ),
    .A3(\as1802.regs[3][3] ),
    .S0(_0000_),
    .S1(_0001_),
    .X(_0590_));
 sky130_fd_sc_hd__mux4_1 _3233_ (.A0(\as1802.regs[4][3] ),
    .A1(\as1802.regs[5][3] ),
    .A2(\as1802.regs[6][3] ),
    .A3(\as1802.regs[7][3] ),
    .S0(_0000_),
    .S1(_0001_),
    .X(_0591_));
 sky130_fd_sc_hd__mux2_1 _3234_ (.A0(_0590_),
    .A1(_0591_),
    .S(_2677_),
    .X(_0592_));
 sky130_fd_sc_hd__o22a_4 _3235_ (.A1(_0587_),
    .A2(_0589_),
    .B1(_0592_),
    .B2(_0003_),
    .X(_0593_));
 sky130_fd_sc_hd__and3_1 _3236_ (.A(_0469_),
    .B(_0519_),
    .C(_0593_),
    .X(_0594_));
 sky130_fd_sc_hd__nor2_1 _3237_ (.A(_0520_),
    .B(_0593_),
    .Y(_0595_));
 sky130_fd_sc_hd__nor2_1 _3238_ (.A(_0594_),
    .B(_0595_),
    .Y(_0596_));
 sky130_fd_sc_hd__mux2_1 _3239_ (.A0(_0596_),
    .A1(_0593_),
    .S(_2695_),
    .X(_0597_));
 sky130_fd_sc_hd__a21o_1 _3240_ (.A1(_2694_),
    .A2(_0520_),
    .B1(_0593_),
    .X(_0598_));
 sky130_fd_sc_hd__a21bo_1 _3241_ (.A1(_2696_),
    .A2(_0594_),
    .B1_N(_0598_),
    .X(_0599_));
 sky130_fd_sc_hd__nor2_1 _3242_ (.A(_0375_),
    .B(_0599_),
    .Y(_0600_));
 sky130_fd_sc_hd__a21o_1 _3243_ (.A1(io_out[3]),
    .A2(_0375_),
    .B1(_0529_),
    .X(_0601_));
 sky130_fd_sc_hd__o221a_1 _3244_ (.A1(_0361_),
    .A2(_0597_),
    .B1(_0600_),
    .B2(_0601_),
    .C1(_0473_),
    .X(_0602_));
 sky130_fd_sc_hd__a211o_1 _3245_ (.A1(_2719_),
    .A2(_0596_),
    .B1(_0602_),
    .C1(_2707_),
    .X(_0603_));
 sky130_fd_sc_hd__o211a_1 _3246_ (.A1(io_out[3]),
    .A2(_0480_),
    .B1(_2700_),
    .C1(_0603_),
    .X(_0604_));
 sky130_fd_sc_hd__a211o_1 _3247_ (.A1(_0366_),
    .A2(_0597_),
    .B1(_0604_),
    .C1(_0369_),
    .X(_0605_));
 sky130_fd_sc_hd__nand2_1 _3248_ (.A(_0369_),
    .B(_0599_),
    .Y(_0606_));
 sky130_fd_sc_hd__a31o_1 _3249_ (.A1(_0380_),
    .A2(_0605_),
    .A3(_0606_),
    .B1(_2596_),
    .X(_0607_));
 sky130_fd_sc_hd__a211o_1 _3250_ (.A1(_0575_),
    .A2(_0578_),
    .B1(_0583_),
    .C1(_0607_),
    .X(_0608_));
 sky130_fd_sc_hd__and2_1 _3251_ (.A(\as1802.regs[2][3] ),
    .B(_0546_),
    .X(_0609_));
 sky130_fd_sc_hd__or2_1 _3252_ (.A(\as1802.regs[2][3] ),
    .B(_0546_),
    .X(_0610_));
 sky130_fd_sc_hd__or3b_1 _3253_ (.A(_0609_),
    .B(_0416_),
    .C_N(_0610_),
    .X(_0611_));
 sky130_fd_sc_hd__o21a_2 _3254_ (.A1(_0574_),
    .A2(_0608_),
    .B1(_0611_),
    .X(_0612_));
 sky130_fd_sc_hd__buf_2 _3255_ (.A(_0612_),
    .X(_0613_));
 sky130_fd_sc_hd__mux2_1 _3256_ (.A0(\as1802.regs[15][3] ),
    .A1(_0613_),
    .S(_0413_),
    .X(_0614_));
 sky130_fd_sc_hd__clkbuf_1 _3257_ (.A(_0614_),
    .X(_0015_));
 sky130_fd_sc_hd__nand2_1 _3258_ (.A(\as1802.regs[2][4] ),
    .B(_0610_),
    .Y(_0615_));
 sky130_fd_sc_hd__or2_1 _3259_ (.A(\as1802.regs[2][4] ),
    .B(_0610_),
    .X(_0616_));
 sky130_fd_sc_hd__clkbuf_4 _3260_ (.A(_0560_),
    .X(_0617_));
 sky130_fd_sc_hd__clkbuf_4 _3261_ (.A(_2629_),
    .X(_0618_));
 sky130_fd_sc_hd__mux2_1 _3262_ (.A0(\as1802.regs[4][4] ),
    .A1(\as1802.regs[5][4] ),
    .S(_0618_),
    .X(_0619_));
 sky130_fd_sc_hd__clkbuf_4 _3263_ (.A(_2620_),
    .X(_0620_));
 sky130_fd_sc_hd__and3_1 _3264_ (.A(\as1802.regs[6][4] ),
    .B(_2656_),
    .C(_2658_),
    .X(_0621_));
 sky130_fd_sc_hd__a211o_1 _3265_ (.A1(\as1802.regs[7][4] ),
    .A2(_0620_),
    .B1(_0621_),
    .C1(_2645_),
    .X(_0622_));
 sky130_fd_sc_hd__o211a_1 _3266_ (.A1(_0617_),
    .A2(_0619_),
    .B1(_0622_),
    .C1(_2648_),
    .X(_0623_));
 sky130_fd_sc_hd__mux2_1 _3267_ (.A0(\as1802.regs[0][4] ),
    .A1(\as1802.regs[1][4] ),
    .S(_0618_),
    .X(_0624_));
 sky130_fd_sc_hd__clkbuf_2 _3268_ (.A(_2621_),
    .X(_0625_));
 sky130_fd_sc_hd__buf_2 _3269_ (.A(_2622_),
    .X(_0626_));
 sky130_fd_sc_hd__and3_1 _3270_ (.A(\as1802.regs[2][4] ),
    .B(_0625_),
    .C(_0626_),
    .X(_0627_));
 sky130_fd_sc_hd__clkbuf_4 _3271_ (.A(_2645_),
    .X(_0628_));
 sky130_fd_sc_hd__a211o_1 _3272_ (.A1(\as1802.regs[3][4] ),
    .A2(_0620_),
    .B1(_0627_),
    .C1(_0628_),
    .X(_0629_));
 sky130_fd_sc_hd__o211a_1 _3273_ (.A1(_0617_),
    .A2(_0624_),
    .B1(_0629_),
    .C1(_2637_),
    .X(_0630_));
 sky130_fd_sc_hd__mux2_1 _3274_ (.A0(\as1802.regs[8][4] ),
    .A1(\as1802.regs[9][4] ),
    .S(_0620_),
    .X(_0631_));
 sky130_fd_sc_hd__clkbuf_4 _3275_ (.A(_0618_),
    .X(_0632_));
 sky130_fd_sc_hd__and3_1 _3276_ (.A(\as1802.regs[10][4] ),
    .B(_0625_),
    .C(_0626_),
    .X(_0633_));
 sky130_fd_sc_hd__a211o_1 _3277_ (.A1(\as1802.regs[11][4] ),
    .A2(_0632_),
    .B1(_0633_),
    .C1(_0628_),
    .X(_0634_));
 sky130_fd_sc_hd__o211a_1 _3278_ (.A1(_0617_),
    .A2(_0631_),
    .B1(_0634_),
    .C1(_2637_),
    .X(_0635_));
 sky130_fd_sc_hd__buf_4 _3279_ (.A(_2648_),
    .X(_0636_));
 sky130_fd_sc_hd__mux2_1 _3280_ (.A0(\as1802.regs[12][4] ),
    .A1(\as1802.regs[13][4] ),
    .S(_2620_),
    .X(_0637_));
 sky130_fd_sc_hd__or2_1 _3281_ (.A(_0560_),
    .B(_0637_),
    .X(_0638_));
 sky130_fd_sc_hd__mux2_1 _3282_ (.A0(\as1802.regs[14][4] ),
    .A1(\as1802.regs[15][4] ),
    .S(_2620_),
    .X(_0639_));
 sky130_fd_sc_hd__or2_1 _3283_ (.A(_0628_),
    .B(_0639_),
    .X(_0640_));
 sky130_fd_sc_hd__a31o_1 _3284_ (.A1(_0636_),
    .A2(_0638_),
    .A3(_0640_),
    .B1(_0437_),
    .X(_0641_));
 sky130_fd_sc_hd__o32ai_4 _3285_ (.A1(_2640_),
    .A2(_0623_),
    .A3(_0630_),
    .B1(_0635_),
    .B2(_0641_),
    .Y(_0642_));
 sky130_fd_sc_hd__nor2_1 _3286_ (.A(_0576_),
    .B(_0642_),
    .Y(_0643_));
 sky130_fd_sc_hd__and2_1 _3287_ (.A(_0576_),
    .B(_0642_),
    .X(_0644_));
 sky130_fd_sc_hd__nor2_1 _3288_ (.A(_0643_),
    .B(_0644_),
    .Y(_0645_));
 sky130_fd_sc_hd__buf_4 _3289_ (.A(\as1802.D[4] ),
    .X(_0646_));
 sky130_fd_sc_hd__clkbuf_4 _3290_ (.A(_0397_),
    .X(_0647_));
 sky130_fd_sc_hd__buf_6 _3291_ (.A(_2640_),
    .X(_0648_));
 sky130_fd_sc_hd__o32a_2 _3292_ (.A1(_0648_),
    .A2(_0623_),
    .A3(_0630_),
    .B1(_0635_),
    .B2(_0641_),
    .X(_0649_));
 sky130_fd_sc_hd__xnor2_1 _3293_ (.A(_0571_),
    .B(_0649_),
    .Y(_0650_));
 sky130_fd_sc_hd__nor2_1 _3294_ (.A(_0446_),
    .B(_0650_),
    .Y(_0651_));
 sky130_fd_sc_hd__a211o_1 _3295_ (.A1(_0447_),
    .A2(_0645_),
    .B1(_0651_),
    .C1(_0384_),
    .X(_0652_));
 sky130_fd_sc_hd__o211a_1 _3296_ (.A1(_0646_),
    .A2(_0580_),
    .B1(_0647_),
    .C1(_0652_),
    .X(_0653_));
 sky130_fd_sc_hd__and2b_1 _3297_ (.A_N(_0458_),
    .B(\as1802.regs[10][4] ),
    .X(_0654_));
 sky130_fd_sc_hd__a21bo_1 _3298_ (.A1(_0458_),
    .A2(\as1802.regs[11][4] ),
    .B1_N(_0001_),
    .X(_0655_));
 sky130_fd_sc_hd__mux2_1 _3299_ (.A0(\as1802.regs[8][4] ),
    .A1(\as1802.regs[9][4] ),
    .S(_2668_),
    .X(_0656_));
 sky130_fd_sc_hd__o221a_1 _3300_ (.A1(_0654_),
    .A2(_0655_),
    .B1(_0656_),
    .B2(_2672_),
    .C1(_2688_),
    .X(_0657_));
 sky130_fd_sc_hd__mux4_1 _3301_ (.A0(\as1802.regs[12][4] ),
    .A1(\as1802.regs[13][4] ),
    .A2(\as1802.regs[14][4] ),
    .A3(\as1802.regs[15][4] ),
    .S0(_2668_),
    .S1(_2671_),
    .X(_0658_));
 sky130_fd_sc_hd__a21o_1 _3302_ (.A1(_2677_),
    .A2(_0658_),
    .B1(_2666_),
    .X(_0659_));
 sky130_fd_sc_hd__mux4_1 _3303_ (.A0(\as1802.regs[0][4] ),
    .A1(\as1802.regs[1][4] ),
    .A2(\as1802.regs[2][4] ),
    .A3(\as1802.regs[3][4] ),
    .S0(_0000_),
    .S1(_0001_),
    .X(_0660_));
 sky130_fd_sc_hd__mux4_1 _3304_ (.A0(\as1802.regs[4][4] ),
    .A1(\as1802.regs[5][4] ),
    .A2(\as1802.regs[6][4] ),
    .A3(\as1802.regs[7][4] ),
    .S0(_0000_),
    .S1(_0001_),
    .X(_0661_));
 sky130_fd_sc_hd__mux2_1 _3305_ (.A0(_0660_),
    .A1(_0661_),
    .S(_2677_),
    .X(_0662_));
 sky130_fd_sc_hd__o22a_2 _3306_ (.A1(_0657_),
    .A2(_0659_),
    .B1(_0662_),
    .B2(_0003_),
    .X(_0663_));
 sky130_fd_sc_hd__and4_1 _3307_ (.A(_0468_),
    .B(_0519_),
    .C(_0593_),
    .D(_0663_),
    .X(_0664_));
 sky130_fd_sc_hd__clkbuf_2 _3308_ (.A(_0664_),
    .X(_0665_));
 sky130_fd_sc_hd__nor2_1 _3309_ (.A(_0594_),
    .B(_0663_),
    .Y(_0666_));
 sky130_fd_sc_hd__nor2_1 _3310_ (.A(_0665_),
    .B(_0666_),
    .Y(_0667_));
 sky130_fd_sc_hd__mux2_1 _3311_ (.A0(_0667_),
    .A1(_0663_),
    .S(_2695_),
    .X(_0668_));
 sky130_fd_sc_hd__a21oi_1 _3312_ (.A1(_2694_),
    .A2(_0594_),
    .B1(_0663_),
    .Y(_0669_));
 sky130_fd_sc_hd__a21oi_1 _3313_ (.A1(_2696_),
    .A2(_0665_),
    .B1(_0669_),
    .Y(_0670_));
 sky130_fd_sc_hd__or2_1 _3314_ (.A(io_out[4]),
    .B(_2722_),
    .X(_0671_));
 sky130_fd_sc_hd__o211a_1 _3315_ (.A1(_0375_),
    .A2(_0670_),
    .B1(_0671_),
    .C1(_0361_),
    .X(_0672_));
 sky130_fd_sc_hd__a211o_1 _3316_ (.A1(_0529_),
    .A2(_0668_),
    .B1(_0672_),
    .C1(_2719_),
    .X(_0673_));
 sky130_fd_sc_hd__or4b_2 _3317_ (.A(_2485_),
    .B(_2712_),
    .C(_0372_),
    .D_N(_2540_),
    .X(_0674_));
 sky130_fd_sc_hd__o211a_1 _3318_ (.A1(_0473_),
    .A2(_0667_),
    .B1(_0673_),
    .C1(_0674_),
    .X(_0675_));
 sky130_fd_sc_hd__a211o_1 _3319_ (.A1(_0373_),
    .A2(_0670_),
    .B1(_0675_),
    .C1(_2710_),
    .X(_0676_));
 sky130_fd_sc_hd__o211a_1 _3320_ (.A1(io_out[4]),
    .A2(_0480_),
    .B1(_2701_),
    .C1(_0676_),
    .X(_0677_));
 sky130_fd_sc_hd__a21oi_1 _3321_ (.A1(_0366_),
    .A2(_0668_),
    .B1(_0677_),
    .Y(_0678_));
 sky130_fd_sc_hd__or2_1 _3322_ (.A(_2606_),
    .B(_0650_),
    .X(_0679_));
 sky130_fd_sc_hd__o211ai_1 _3323_ (.A1(_0537_),
    .A2(_0678_),
    .B1(_0679_),
    .C1(_0416_),
    .Y(_0680_));
 sky130_fd_sc_hd__a211oi_2 _3324_ (.A1(_0575_),
    .A2(_0645_),
    .B1(_0653_),
    .C1(_0680_),
    .Y(_0681_));
 sky130_fd_sc_hd__a31oi_4 _3325_ (.A1(_2597_),
    .A2(_0615_),
    .A3(_0616_),
    .B1(_0681_),
    .Y(_0682_));
 sky130_fd_sc_hd__buf_2 _3326_ (.A(_0682_),
    .X(_0683_));
 sky130_fd_sc_hd__mux2_1 _3327_ (.A0(\as1802.regs[15][4] ),
    .A1(_0683_),
    .S(_0413_),
    .X(_0684_));
 sky130_fd_sc_hd__clkbuf_1 _3328_ (.A(_0684_),
    .X(_0016_));
 sky130_fd_sc_hd__clkbuf_4 _3329_ (.A(_2645_),
    .X(_0685_));
 sky130_fd_sc_hd__mux2_1 _3330_ (.A0(\as1802.regs[6][5] ),
    .A1(\as1802.regs[7][5] ),
    .S(_0618_),
    .X(_0686_));
 sky130_fd_sc_hd__and3_1 _3331_ (.A(\as1802.regs[4][5] ),
    .B(_2656_),
    .C(_2658_),
    .X(_0687_));
 sky130_fd_sc_hd__a211o_1 _3332_ (.A1(\as1802.regs[5][5] ),
    .A2(_0618_),
    .B1(_0687_),
    .C1(_0560_),
    .X(_0688_));
 sky130_fd_sc_hd__o211ai_1 _3333_ (.A1(_0685_),
    .A2(_0686_),
    .B1(_0688_),
    .C1(_2648_),
    .Y(_0689_));
 sky130_fd_sc_hd__and3_1 _3334_ (.A(\as1802.regs[0][5] ),
    .B(_2656_),
    .C(_2658_),
    .X(_0690_));
 sky130_fd_sc_hd__a211oi_1 _3335_ (.A1(\as1802.regs[1][5] ),
    .A2(_0620_),
    .B1(_0690_),
    .C1(_0560_),
    .Y(_0691_));
 sky130_fd_sc_hd__and3_1 _3336_ (.A(\as1802.X[0] ),
    .B(_2609_),
    .C(_2616_),
    .X(_0692_));
 sky130_fd_sc_hd__a21oi_2 _3337_ (.A1(_2609_),
    .A2(_2616_),
    .B1(_2513_),
    .Y(_0693_));
 sky130_fd_sc_hd__o21ai_1 _3338_ (.A1(_0692_),
    .A2(_0693_),
    .B1(\as1802.regs[3][5] ),
    .Y(_0694_));
 sky130_fd_sc_hd__or3b_1 _3339_ (.A(_0692_),
    .B(_0693_),
    .C_N(\as1802.regs[2][5] ),
    .X(_0695_));
 sky130_fd_sc_hd__a31o_1 _3340_ (.A1(_0560_),
    .A2(_0694_),
    .A3(_0695_),
    .B1(_2648_),
    .X(_0696_));
 sky130_fd_sc_hd__o21a_1 _3341_ (.A1(_0691_),
    .A2(_0696_),
    .B1(_0437_),
    .X(_0697_));
 sky130_fd_sc_hd__and3_1 _3342_ (.A(\as1802.regs[12][5] ),
    .B(_2656_),
    .C(_2658_),
    .X(_0698_));
 sky130_fd_sc_hd__a211o_1 _3343_ (.A1(\as1802.regs[13][5] ),
    .A2(_0618_),
    .B1(_0698_),
    .C1(_2642_),
    .X(_0699_));
 sky130_fd_sc_hd__and3_1 _3344_ (.A(\as1802.regs[14][5] ),
    .B(_2656_),
    .C(_2658_),
    .X(_0700_));
 sky130_fd_sc_hd__a211o_1 _3345_ (.A1(\as1802.regs[15][5] ),
    .A2(_0618_),
    .B1(_0700_),
    .C1(_2645_),
    .X(_0701_));
 sky130_fd_sc_hd__and3_1 _3346_ (.A(\as1802.regs[10][5] ),
    .B(_2656_),
    .C(_2658_),
    .X(_0702_));
 sky130_fd_sc_hd__a211o_1 _3347_ (.A1(\as1802.regs[11][5] ),
    .A2(_0618_),
    .B1(_0702_),
    .C1(_2645_),
    .X(_0703_));
 sky130_fd_sc_hd__and3_1 _3348_ (.A(\as1802.regs[8][5] ),
    .B(_2656_),
    .C(_2658_),
    .X(_0704_));
 sky130_fd_sc_hd__o21a_1 _3349_ (.A1(_0692_),
    .A2(_0693_),
    .B1(\as1802.regs[9][5] ),
    .X(_0705_));
 sky130_fd_sc_hd__o31a_1 _3350_ (.A1(_2642_),
    .A2(_0704_),
    .A3(_0705_),
    .B1(_2637_),
    .X(_0706_));
 sky130_fd_sc_hd__a32o_1 _3351_ (.A1(_2648_),
    .A2(_0699_),
    .A3(_0701_),
    .B1(_0703_),
    .B2(_0706_),
    .X(_0707_));
 sky130_fd_sc_hd__buf_6 _3352_ (.A(_0437_),
    .X(_0708_));
 sky130_fd_sc_hd__o2bb2a_2 _3353_ (.A1_N(_0689_),
    .A2_N(_0697_),
    .B1(_0707_),
    .B2(_0708_),
    .X(_0709_));
 sky130_fd_sc_hd__clkinv_2 _3354_ (.A(_0709_),
    .Y(_0710_));
 sky130_fd_sc_hd__and3_1 _3355_ (.A(_0571_),
    .B(_0642_),
    .C(_0710_),
    .X(_0711_));
 sky130_fd_sc_hd__a21oi_1 _3356_ (.A1(_0571_),
    .A2(_0642_),
    .B1(_0710_),
    .Y(_0712_));
 sky130_fd_sc_hd__or2_1 _3357_ (.A(_0711_),
    .B(_0712_),
    .X(_0713_));
 sky130_fd_sc_hd__xnor2_1 _3358_ (.A(_0643_),
    .B(_0710_),
    .Y(_0714_));
 sky130_fd_sc_hd__mux2_1 _3359_ (.A0(_0713_),
    .A1(_0714_),
    .S(_0447_),
    .X(_0715_));
 sky130_fd_sc_hd__clkbuf_4 _3360_ (.A(\as1802.D[5] ),
    .X(_0716_));
 sky130_fd_sc_hd__o21a_1 _3361_ (.A1(_0716_),
    .A2(_0580_),
    .B1(_0647_),
    .X(_0717_));
 sky130_fd_sc_hd__o21ai_1 _3362_ (.A1(_0384_),
    .A2(_0715_),
    .B1(_0717_),
    .Y(_0718_));
 sky130_fd_sc_hd__clkbuf_4 _3363_ (.A(_2669_),
    .X(_0719_));
 sky130_fd_sc_hd__and2b_1 _3364_ (.A_N(_0719_),
    .B(\as1802.regs[10][5] ),
    .X(_0720_));
 sky130_fd_sc_hd__a21bo_1 _3365_ (.A1(_0719_),
    .A2(\as1802.regs[11][5] ),
    .B1_N(_2673_),
    .X(_0721_));
 sky130_fd_sc_hd__mux2_1 _3366_ (.A0(\as1802.regs[8][5] ),
    .A1(\as1802.regs[9][5] ),
    .S(_0719_),
    .X(_0722_));
 sky130_fd_sc_hd__o221a_1 _3367_ (.A1(_0720_),
    .A2(_0721_),
    .B1(_0722_),
    .B2(_2674_),
    .C1(_2689_),
    .X(_0723_));
 sky130_fd_sc_hd__mux4_1 _3368_ (.A0(\as1802.regs[12][5] ),
    .A1(\as1802.regs[13][5] ),
    .A2(\as1802.regs[14][5] ),
    .A3(\as1802.regs[15][5] ),
    .S0(_0719_),
    .S1(_2673_),
    .X(_0724_));
 sky130_fd_sc_hd__a21o_1 _3369_ (.A1(_2678_),
    .A2(_0724_),
    .B1(_2666_),
    .X(_0725_));
 sky130_fd_sc_hd__mux4_1 _3370_ (.A0(\as1802.regs[0][5] ),
    .A1(\as1802.regs[1][5] ),
    .A2(\as1802.regs[2][5] ),
    .A3(\as1802.regs[3][5] ),
    .S0(_2669_),
    .S1(_2672_),
    .X(_0726_));
 sky130_fd_sc_hd__mux4_1 _3371_ (.A0(\as1802.regs[4][5] ),
    .A1(\as1802.regs[5][5] ),
    .A2(\as1802.regs[6][5] ),
    .A3(\as1802.regs[7][5] ),
    .S0(_2669_),
    .S1(_2672_),
    .X(_0727_));
 sky130_fd_sc_hd__mux2_1 _3372_ (.A0(_0726_),
    .A1(_0727_),
    .S(_2678_),
    .X(_0728_));
 sky130_fd_sc_hd__o22a_4 _3373_ (.A1(_0723_),
    .A2(_0725_),
    .B1(_0728_),
    .B2(_0003_),
    .X(_0729_));
 sky130_fd_sc_hd__nand2_1 _3374_ (.A(_0665_),
    .B(_0729_),
    .Y(_0730_));
 sky130_fd_sc_hd__or2_1 _3375_ (.A(_0665_),
    .B(_0729_),
    .X(_0731_));
 sky130_fd_sc_hd__and2_1 _3376_ (.A(_0730_),
    .B(_0731_),
    .X(_0732_));
 sky130_fd_sc_hd__mux2_1 _3377_ (.A0(_0732_),
    .A1(_0729_),
    .S(_2695_),
    .X(_0733_));
 sky130_fd_sc_hd__nor2_1 _3378_ (.A(_2720_),
    .B(_0730_),
    .Y(_0734_));
 sky130_fd_sc_hd__a21oi_1 _3379_ (.A1(_2696_),
    .A2(_0665_),
    .B1(_0729_),
    .Y(_0735_));
 sky130_fd_sc_hd__nor2_1 _3380_ (.A(_0734_),
    .B(_0735_),
    .Y(_0736_));
 sky130_fd_sc_hd__or2_1 _3381_ (.A(io_out[5]),
    .B(_2722_),
    .X(_0737_));
 sky130_fd_sc_hd__o211a_1 _3382_ (.A1(_0375_),
    .A2(_0736_),
    .B1(_0737_),
    .C1(_0361_),
    .X(_0738_));
 sky130_fd_sc_hd__a211o_1 _3383_ (.A1(_0529_),
    .A2(_0733_),
    .B1(_0738_),
    .C1(_2719_),
    .X(_0739_));
 sky130_fd_sc_hd__o211a_1 _3384_ (.A1(_0473_),
    .A2(_0732_),
    .B1(_0739_),
    .C1(_0674_),
    .X(_0740_));
 sky130_fd_sc_hd__a211o_1 _3385_ (.A1(_0373_),
    .A2(_0736_),
    .B1(_0740_),
    .C1(_2710_),
    .X(_0741_));
 sky130_fd_sc_hd__o211a_1 _3386_ (.A1(io_out[5]),
    .A2(_0480_),
    .B1(_2701_),
    .C1(_0741_),
    .X(_0742_));
 sky130_fd_sc_hd__a21o_1 _3387_ (.A1(_0366_),
    .A2(_0733_),
    .B1(_0742_),
    .X(_0743_));
 sky130_fd_sc_hd__a221o_1 _3388_ (.A1(_0454_),
    .A2(_0713_),
    .B1(_0714_),
    .B2(_0575_),
    .C1(_2596_),
    .X(_0744_));
 sky130_fd_sc_hd__a21oi_2 _3389_ (.A1(_0380_),
    .A2(_0743_),
    .B1(_0744_),
    .Y(_0745_));
 sky130_fd_sc_hd__nand2_1 _3390_ (.A(\as1802.regs[2][5] ),
    .B(_0616_),
    .Y(_0746_));
 sky130_fd_sc_hd__or2_1 _3391_ (.A(\as1802.regs[2][5] ),
    .B(_0616_),
    .X(_0747_));
 sky130_fd_sc_hd__and3_1 _3392_ (.A(_2597_),
    .B(_0746_),
    .C(_0747_),
    .X(_0748_));
 sky130_fd_sc_hd__a21oi_4 _3393_ (.A1(_0718_),
    .A2(_0745_),
    .B1(_0748_),
    .Y(_0749_));
 sky130_fd_sc_hd__buf_2 _3394_ (.A(_0749_),
    .X(_0750_));
 sky130_fd_sc_hd__mux2_1 _3395_ (.A0(\as1802.regs[15][5] ),
    .A1(_0750_),
    .S(_0413_),
    .X(_0751_));
 sky130_fd_sc_hd__clkbuf_1 _3396_ (.A(_0751_),
    .X(_0017_));
 sky130_fd_sc_hd__and2b_1 _3397_ (.A_N(_0719_),
    .B(\as1802.regs[10][6] ),
    .X(_0752_));
 sky130_fd_sc_hd__a21bo_1 _3398_ (.A1(_0719_),
    .A2(\as1802.regs[11][6] ),
    .B1_N(_2673_),
    .X(_0753_));
 sky130_fd_sc_hd__mux2_1 _3399_ (.A0(\as1802.regs[8][6] ),
    .A1(\as1802.regs[9][6] ),
    .S(_0719_),
    .X(_0754_));
 sky130_fd_sc_hd__o221a_1 _3400_ (.A1(_0752_),
    .A2(_0753_),
    .B1(_0754_),
    .B2(_2674_),
    .C1(_2689_),
    .X(_0755_));
 sky130_fd_sc_hd__mux4_1 _3401_ (.A0(\as1802.regs[12][6] ),
    .A1(\as1802.regs[13][6] ),
    .A2(\as1802.regs[14][6] ),
    .A3(\as1802.regs[15][6] ),
    .S0(_2669_),
    .S1(_2673_),
    .X(_0756_));
 sky130_fd_sc_hd__a21o_1 _3402_ (.A1(_2678_),
    .A2(_0756_),
    .B1(_2666_),
    .X(_0757_));
 sky130_fd_sc_hd__mux4_1 _3403_ (.A0(\as1802.regs[0][6] ),
    .A1(\as1802.regs[1][6] ),
    .A2(\as1802.regs[2][6] ),
    .A3(\as1802.regs[3][6] ),
    .S0(_2669_),
    .S1(_2672_),
    .X(_0758_));
 sky130_fd_sc_hd__mux4_1 _3404_ (.A0(\as1802.regs[4][6] ),
    .A1(\as1802.regs[5][6] ),
    .A2(\as1802.regs[6][6] ),
    .A3(\as1802.regs[7][6] ),
    .S0(_2669_),
    .S1(_2672_),
    .X(_0759_));
 sky130_fd_sc_hd__mux2_1 _3405_ (.A0(_0758_),
    .A1(_0759_),
    .S(_2677_),
    .X(_0760_));
 sky130_fd_sc_hd__o22a_4 _3406_ (.A1(_0755_),
    .A2(_0757_),
    .B1(_0760_),
    .B2(_0003_),
    .X(_0761_));
 sky130_fd_sc_hd__xor2_1 _3407_ (.A(_0730_),
    .B(_0761_),
    .X(_0762_));
 sky130_fd_sc_hd__inv_2 _3408_ (.A(_0762_),
    .Y(_0763_));
 sky130_fd_sc_hd__mux2_1 _3409_ (.A0(_0763_),
    .A1(_0761_),
    .S(_2695_),
    .X(_0764_));
 sky130_fd_sc_hd__xor2_1 _3410_ (.A(_0734_),
    .B(_0761_),
    .X(_0765_));
 sky130_fd_sc_hd__or2_1 _3411_ (.A(io_out[6]),
    .B(_2722_),
    .X(_0766_));
 sky130_fd_sc_hd__o211a_1 _3412_ (.A1(_0375_),
    .A2(_0765_),
    .B1(_0766_),
    .C1(_0361_),
    .X(_0767_));
 sky130_fd_sc_hd__a211o_1 _3413_ (.A1(_0529_),
    .A2(_0764_),
    .B1(_0767_),
    .C1(_2719_),
    .X(_0768_));
 sky130_fd_sc_hd__o211a_1 _3414_ (.A1(_0473_),
    .A2(_0763_),
    .B1(_0768_),
    .C1(_0674_),
    .X(_0769_));
 sky130_fd_sc_hd__a211o_1 _3415_ (.A1(_0373_),
    .A2(_0765_),
    .B1(_0769_),
    .C1(_2710_),
    .X(_0770_));
 sky130_fd_sc_hd__o211a_1 _3416_ (.A1(io_out[6]),
    .A2(_0480_),
    .B1(_2701_),
    .C1(_0770_),
    .X(_0771_));
 sky130_fd_sc_hd__a21o_1 _3417_ (.A1(_0366_),
    .A2(_0764_),
    .B1(_0771_),
    .X(_0772_));
 sky130_fd_sc_hd__mux2_1 _3418_ (.A0(\as1802.regs[0][6] ),
    .A1(\as1802.regs[1][6] ),
    .S(_0618_),
    .X(_0773_));
 sky130_fd_sc_hd__and3_1 _3419_ (.A(\as1802.regs[2][6] ),
    .B(_0625_),
    .C(_0626_),
    .X(_0774_));
 sky130_fd_sc_hd__a211o_1 _3420_ (.A1(\as1802.regs[3][6] ),
    .A2(_0620_),
    .B1(_0774_),
    .C1(_0628_),
    .X(_0775_));
 sky130_fd_sc_hd__o211a_1 _3421_ (.A1(_0617_),
    .A2(_0773_),
    .B1(_0775_),
    .C1(_2637_),
    .X(_0776_));
 sky130_fd_sc_hd__and3_1 _3422_ (.A(\as1802.regs[4][6] ),
    .B(_0625_),
    .C(_0626_),
    .X(_0777_));
 sky130_fd_sc_hd__a211o_1 _3423_ (.A1(\as1802.regs[5][6] ),
    .A2(_0620_),
    .B1(_0777_),
    .C1(_0560_),
    .X(_0778_));
 sky130_fd_sc_hd__and3_1 _3424_ (.A(\as1802.regs[6][6] ),
    .B(_0625_),
    .C(_0626_),
    .X(_0779_));
 sky130_fd_sc_hd__a211o_1 _3425_ (.A1(\as1802.regs[7][6] ),
    .A2(_0620_),
    .B1(_0779_),
    .C1(_0628_),
    .X(_0780_));
 sky130_fd_sc_hd__a31o_1 _3426_ (.A1(_2648_),
    .A2(_0778_),
    .A3(_0780_),
    .B1(_2640_),
    .X(_0781_));
 sky130_fd_sc_hd__mux2_1 _3427_ (.A0(\as1802.regs[8][6] ),
    .A1(\as1802.regs[9][6] ),
    .S(_0620_),
    .X(_0782_));
 sky130_fd_sc_hd__and3_1 _3428_ (.A(\as1802.regs[10][6] ),
    .B(_0625_),
    .C(_0626_),
    .X(_0783_));
 sky130_fd_sc_hd__a211o_1 _3429_ (.A1(\as1802.regs[11][6] ),
    .A2(_0632_),
    .B1(_0783_),
    .C1(_0628_),
    .X(_0784_));
 sky130_fd_sc_hd__clkbuf_4 _3430_ (.A(_2637_),
    .X(_0785_));
 sky130_fd_sc_hd__o211a_1 _3431_ (.A1(_0617_),
    .A2(_0782_),
    .B1(_0784_),
    .C1(_0785_),
    .X(_0786_));
 sky130_fd_sc_hd__and3_1 _3432_ (.A(\as1802.regs[14][6] ),
    .B(_0625_),
    .C(_0626_),
    .X(_0787_));
 sky130_fd_sc_hd__a211o_1 _3433_ (.A1(\as1802.regs[15][6] ),
    .A2(_0632_),
    .B1(_0787_),
    .C1(_0628_),
    .X(_0788_));
 sky130_fd_sc_hd__and3_1 _3434_ (.A(\as1802.regs[12][6] ),
    .B(_0625_),
    .C(_0626_),
    .X(_0789_));
 sky130_fd_sc_hd__a211o_1 _3435_ (.A1(\as1802.regs[13][6] ),
    .A2(_0632_),
    .B1(_0789_),
    .C1(_0560_),
    .X(_0790_));
 sky130_fd_sc_hd__a31o_1 _3436_ (.A1(_0636_),
    .A2(_0788_),
    .A3(_0790_),
    .B1(_0437_),
    .X(_0791_));
 sky130_fd_sc_hd__o22a_4 _3437_ (.A1(_0776_),
    .A2(_0781_),
    .B1(_0786_),
    .B2(_0791_),
    .X(_0792_));
 sky130_fd_sc_hd__xnor2_1 _3438_ (.A(_0711_),
    .B(_0792_),
    .Y(_0793_));
 sky130_fd_sc_hd__or3_1 _3439_ (.A(_0576_),
    .B(_0642_),
    .C(_0710_),
    .X(_0794_));
 sky130_fd_sc_hd__xor2_1 _3440_ (.A(_0794_),
    .B(_0792_),
    .X(_0795_));
 sky130_fd_sc_hd__mux2_1 _3441_ (.A0(_0793_),
    .A1(_0795_),
    .S(_0446_),
    .X(_0796_));
 sky130_fd_sc_hd__buf_4 _3442_ (.A(\as1802.D[6] ),
    .X(_0797_));
 sky130_fd_sc_hd__o21ai_1 _3443_ (.A1(_0797_),
    .A2(_0580_),
    .B1(_0397_),
    .Y(_0798_));
 sky130_fd_sc_hd__a21oi_1 _3444_ (.A1(_0580_),
    .A2(_0796_),
    .B1(_0798_),
    .Y(_0799_));
 sky130_fd_sc_hd__a211o_1 _3445_ (.A1(_0380_),
    .A2(_0772_),
    .B1(_0799_),
    .C1(_0403_),
    .X(_0800_));
 sky130_fd_sc_hd__a221oi_1 _3446_ (.A1(_0454_),
    .A2(_0793_),
    .B1(_0795_),
    .B2(_0450_),
    .C1(_2597_),
    .Y(_0801_));
 sky130_fd_sc_hd__or2_1 _3447_ (.A(\as1802.regs[2][6] ),
    .B(_0747_),
    .X(_0802_));
 sky130_fd_sc_hd__nand2_1 _3448_ (.A(\as1802.regs[2][6] ),
    .B(_0747_),
    .Y(_0803_));
 sky130_fd_sc_hd__nand2_1 _3449_ (.A(_0802_),
    .B(_0803_),
    .Y(_0804_));
 sky130_fd_sc_hd__a22o_2 _3450_ (.A1(_0800_),
    .A2(_0801_),
    .B1(_0804_),
    .B2(_2597_),
    .X(_0805_));
 sky130_fd_sc_hd__buf_2 _3451_ (.A(_0805_),
    .X(_0806_));
 sky130_fd_sc_hd__mux2_1 _3452_ (.A0(\as1802.regs[15][6] ),
    .A1(_0806_),
    .S(_0413_),
    .X(_0807_));
 sky130_fd_sc_hd__clkbuf_1 _3453_ (.A(_0807_),
    .X(_0018_));
 sky130_fd_sc_hd__or2_1 _3454_ (.A(\as1802.regs[2][7] ),
    .B(_0802_),
    .X(_0808_));
 sky130_fd_sc_hd__a21oi_1 _3455_ (.A1(\as1802.regs[2][7] ),
    .A2(_0802_),
    .B1(_0416_),
    .Y(_0809_));
 sky130_fd_sc_hd__or4b_1 _3456_ (.A(_0649_),
    .B(_0709_),
    .C(_0792_),
    .D_N(_0571_),
    .X(_0810_));
 sky130_fd_sc_hd__mux2_1 _3457_ (.A0(\as1802.regs[6][7] ),
    .A1(\as1802.regs[7][7] ),
    .S(_0620_),
    .X(_0811_));
 sky130_fd_sc_hd__and3_1 _3458_ (.A(\as1802.regs[4][7] ),
    .B(_0625_),
    .C(_0626_),
    .X(_0812_));
 sky130_fd_sc_hd__a211o_1 _3459_ (.A1(\as1802.regs[5][7] ),
    .A2(_0632_),
    .B1(_0812_),
    .C1(_0560_),
    .X(_0813_));
 sky130_fd_sc_hd__o211a_1 _3460_ (.A1(_0685_),
    .A2(_0811_),
    .B1(_0813_),
    .C1(_0636_),
    .X(_0814_));
 sky130_fd_sc_hd__mux2_1 _3461_ (.A0(\as1802.regs[0][7] ),
    .A1(\as1802.regs[1][7] ),
    .S(_0620_),
    .X(_0815_));
 sky130_fd_sc_hd__and3_1 _3462_ (.A(\as1802.regs[2][7] ),
    .B(_0625_),
    .C(_0626_),
    .X(_0816_));
 sky130_fd_sc_hd__a211o_1 _3463_ (.A1(\as1802.regs[3][7] ),
    .A2(_0632_),
    .B1(_0816_),
    .C1(_0628_),
    .X(_0817_));
 sky130_fd_sc_hd__o211a_1 _3464_ (.A1(_0617_),
    .A2(_0815_),
    .B1(_0817_),
    .C1(_0785_),
    .X(_0818_));
 sky130_fd_sc_hd__mux2_1 _3465_ (.A0(\as1802.regs[8][7] ),
    .A1(\as1802.regs[9][7] ),
    .S(_0632_),
    .X(_0819_));
 sky130_fd_sc_hd__buf_4 _3466_ (.A(_0618_),
    .X(_0820_));
 sky130_fd_sc_hd__buf_2 _3467_ (.A(_2656_),
    .X(_0821_));
 sky130_fd_sc_hd__buf_2 _3468_ (.A(_2658_),
    .X(_0822_));
 sky130_fd_sc_hd__and3_1 _3469_ (.A(\as1802.regs[10][7] ),
    .B(_0821_),
    .C(_0822_),
    .X(_0823_));
 sky130_fd_sc_hd__a211o_1 _3470_ (.A1(\as1802.regs[11][7] ),
    .A2(_0820_),
    .B1(_0823_),
    .C1(_0628_),
    .X(_0824_));
 sky130_fd_sc_hd__o211a_1 _3471_ (.A1(_0617_),
    .A2(_0819_),
    .B1(_0824_),
    .C1(_0785_),
    .X(_0825_));
 sky130_fd_sc_hd__and3_1 _3472_ (.A(\as1802.regs[12][7] ),
    .B(_0821_),
    .C(_0822_),
    .X(_0826_));
 sky130_fd_sc_hd__a211o_1 _3473_ (.A1(\as1802.regs[13][7] ),
    .A2(_0820_),
    .B1(_0826_),
    .C1(_0560_),
    .X(_0827_));
 sky130_fd_sc_hd__and3_1 _3474_ (.A(\as1802.regs[14][7] ),
    .B(_0821_),
    .C(_0822_),
    .X(_0828_));
 sky130_fd_sc_hd__a211o_1 _3475_ (.A1(\as1802.regs[15][7] ),
    .A2(_0632_),
    .B1(_0828_),
    .C1(_0628_),
    .X(_0829_));
 sky130_fd_sc_hd__a31o_1 _3476_ (.A1(_0636_),
    .A2(_0827_),
    .A3(_0829_),
    .B1(_0708_),
    .X(_0830_));
 sky130_fd_sc_hd__o32ai_4 _3477_ (.A1(_2640_),
    .A2(_0814_),
    .A3(_0818_),
    .B1(_0825_),
    .B2(_0830_),
    .Y(_0831_));
 sky130_fd_sc_hd__clkinv_2 _3478_ (.A(_0831_),
    .Y(_0832_));
 sky130_fd_sc_hd__nor3b_1 _3479_ (.A(_0709_),
    .B(_0792_),
    .C_N(_0831_),
    .Y(_0833_));
 sky130_fd_sc_hd__and3_1 _3480_ (.A(_0571_),
    .B(_0642_),
    .C(_0833_),
    .X(_0834_));
 sky130_fd_sc_hd__a21o_1 _3481_ (.A1(_0810_),
    .A2(_0832_),
    .B1(_0834_),
    .X(_0835_));
 sky130_fd_sc_hd__or4b_1 _3482_ (.A(_0576_),
    .B(_0642_),
    .C(_0710_),
    .D_N(_0792_),
    .X(_0836_));
 sky130_fd_sc_hd__buf_2 _3483_ (.A(_0836_),
    .X(_0837_));
 sky130_fd_sc_hd__xnor2_1 _3484_ (.A(_0837_),
    .B(_0832_),
    .Y(_0838_));
 sky130_fd_sc_hd__mux2_1 _3485_ (.A0(_0835_),
    .A1(_0838_),
    .S(_0446_),
    .X(_0839_));
 sky130_fd_sc_hd__inv_2 _3486_ (.A(\as1802.D[7] ),
    .Y(_0840_));
 sky130_fd_sc_hd__nand2_1 _3487_ (.A(_0840_),
    .B(_0384_),
    .Y(_0841_));
 sky130_fd_sc_hd__o211a_1 _3488_ (.A1(_0384_),
    .A2(_0839_),
    .B1(_0841_),
    .C1(_0397_),
    .X(_0842_));
 sky130_fd_sc_hd__and2_1 _3489_ (.A(_0454_),
    .B(_0835_),
    .X(_0843_));
 sky130_fd_sc_hd__and2b_1 _3490_ (.A_N(_0719_),
    .B(\as1802.regs[10][7] ),
    .X(_0844_));
 sky130_fd_sc_hd__a21bo_1 _3491_ (.A1(_2670_),
    .A2(\as1802.regs[11][7] ),
    .B1_N(_2673_),
    .X(_0845_));
 sky130_fd_sc_hd__mux2_1 _3492_ (.A0(\as1802.regs[8][7] ),
    .A1(\as1802.regs[9][7] ),
    .S(_0719_),
    .X(_0846_));
 sky130_fd_sc_hd__o221a_1 _3493_ (.A1(_0844_),
    .A2(_0845_),
    .B1(_0846_),
    .B2(_2674_),
    .C1(_2689_),
    .X(_0847_));
 sky130_fd_sc_hd__mux4_1 _3494_ (.A0(\as1802.regs[12][7] ),
    .A1(\as1802.regs[13][7] ),
    .A2(\as1802.regs[14][7] ),
    .A3(\as1802.regs[15][7] ),
    .S0(_0719_),
    .S1(_2673_),
    .X(_0848_));
 sky130_fd_sc_hd__a21o_1 _3495_ (.A1(_2678_),
    .A2(_0848_),
    .B1(_2667_),
    .X(_0849_));
 sky130_fd_sc_hd__mux4_1 _3496_ (.A0(\as1802.regs[4][7] ),
    .A1(\as1802.regs[5][7] ),
    .A2(\as1802.regs[6][7] ),
    .A3(\as1802.regs[7][7] ),
    .S0(_2669_),
    .S1(_2673_),
    .X(_0850_));
 sky130_fd_sc_hd__mux4_1 _3497_ (.A0(\as1802.regs[0][7] ),
    .A1(\as1802.regs[1][7] ),
    .A2(\as1802.regs[2][7] ),
    .A3(\as1802.regs[3][7] ),
    .S0(_2669_),
    .S1(_2672_),
    .X(_0851_));
 sky130_fd_sc_hd__mux2_1 _3498_ (.A0(_0850_),
    .A1(_0851_),
    .S(_2689_),
    .X(_0852_));
 sky130_fd_sc_hd__o22a_4 _3499_ (.A1(_0847_),
    .A2(_0849_),
    .B1(_0852_),
    .B2(_0003_),
    .X(_0853_));
 sky130_fd_sc_hd__and4_1 _3500_ (.A(_0665_),
    .B(_0729_),
    .C(_0761_),
    .D(_0853_),
    .X(_0854_));
 sky130_fd_sc_hd__clkbuf_2 _3501_ (.A(_0854_),
    .X(_0855_));
 sky130_fd_sc_hd__a31o_1 _3502_ (.A1(_0665_),
    .A2(_0729_),
    .A3(_0761_),
    .B1(_0853_),
    .X(_0856_));
 sky130_fd_sc_hd__and2b_1 _3503_ (.A_N(_0855_),
    .B(_0856_),
    .X(_0857_));
 sky130_fd_sc_hd__mux2_1 _3504_ (.A0(_0857_),
    .A1(_0853_),
    .S(_2695_),
    .X(_0858_));
 sky130_fd_sc_hd__a41o_1 _3505_ (.A1(_2693_),
    .A2(_0665_),
    .A3(_0729_),
    .A4(_0761_),
    .B1(_0853_),
    .X(_0859_));
 sky130_fd_sc_hd__a21boi_1 _3506_ (.A1(_2694_),
    .A2(_0855_),
    .B1_N(_0859_),
    .Y(_0860_));
 sky130_fd_sc_hd__or2_1 _3507_ (.A(io_out[7]),
    .B(_2722_),
    .X(_0861_));
 sky130_fd_sc_hd__o21a_1 _3508_ (.A1(_0375_),
    .A2(_0860_),
    .B1(_0361_),
    .X(_0862_));
 sky130_fd_sc_hd__a221o_1 _3509_ (.A1(_0861_),
    .A2(_0862_),
    .B1(_0858_),
    .B2(_0529_),
    .C1(_2719_),
    .X(_0863_));
 sky130_fd_sc_hd__o211a_1 _3510_ (.A1(_0473_),
    .A2(_0857_),
    .B1(_0863_),
    .C1(_0674_),
    .X(_0864_));
 sky130_fd_sc_hd__a211o_1 _3511_ (.A1(_0373_),
    .A2(_0860_),
    .B1(_0864_),
    .C1(_2710_),
    .X(_0865_));
 sky130_fd_sc_hd__o211a_1 _3512_ (.A1(io_out[7]),
    .A2(_0480_),
    .B1(_2700_),
    .C1(_0865_),
    .X(_0866_));
 sky130_fd_sc_hd__a21o_1 _3513_ (.A1(_0366_),
    .A2(_0858_),
    .B1(_0866_),
    .X(_0867_));
 sky130_fd_sc_hd__a221o_1 _3514_ (.A1(_0450_),
    .A2(_0838_),
    .B1(_0867_),
    .B2(_0380_),
    .C1(_2596_),
    .X(_0868_));
 sky130_fd_sc_hd__or3_1 _3515_ (.A(_0842_),
    .B(_0843_),
    .C(_0868_),
    .X(_0869_));
 sky130_fd_sc_hd__a21boi_4 _3516_ (.A1(_0808_),
    .A2(_0809_),
    .B1_N(_0869_),
    .Y(_0870_));
 sky130_fd_sc_hd__buf_2 _3517_ (.A(_0870_),
    .X(_0871_));
 sky130_fd_sc_hd__mux2_1 _3518_ (.A0(\as1802.regs[15][7] ),
    .A1(_0871_),
    .S(_0413_),
    .X(_0872_));
 sky130_fd_sc_hd__clkbuf_1 _3519_ (.A(_0872_),
    .X(_0019_));
 sky130_fd_sc_hd__a21oi_1 _3520_ (.A1(\as1802.regs[2][8] ),
    .A2(_0808_),
    .B1(_0416_),
    .Y(_0873_));
 sky130_fd_sc_hd__or2_1 _3521_ (.A(\as1802.regs[2][8] ),
    .B(_0808_),
    .X(_0874_));
 sky130_fd_sc_hd__nor2_1 _3522_ (.A(_0837_),
    .B(_0831_),
    .Y(_0875_));
 sky130_fd_sc_hd__clkbuf_4 _3523_ (.A(_0617_),
    .X(_0876_));
 sky130_fd_sc_hd__buf_4 _3524_ (.A(_0632_),
    .X(_0877_));
 sky130_fd_sc_hd__mux2_1 _3525_ (.A0(\as1802.regs[12][8] ),
    .A1(\as1802.regs[13][8] ),
    .S(_0877_),
    .X(_0878_));
 sky130_fd_sc_hd__clkbuf_4 _3526_ (.A(_0820_),
    .X(_0879_));
 sky130_fd_sc_hd__clkbuf_2 _3527_ (.A(_0821_),
    .X(_0880_));
 sky130_fd_sc_hd__clkbuf_2 _3528_ (.A(_0822_),
    .X(_0881_));
 sky130_fd_sc_hd__and3_1 _3529_ (.A(\as1802.regs[14][8] ),
    .B(_0880_),
    .C(_0881_),
    .X(_0882_));
 sky130_fd_sc_hd__clkbuf_4 _3530_ (.A(_0685_),
    .X(_0883_));
 sky130_fd_sc_hd__a211o_1 _3531_ (.A1(\as1802.regs[15][8] ),
    .A2(_0879_),
    .B1(_0882_),
    .C1(_0883_),
    .X(_0884_));
 sky130_fd_sc_hd__o211a_1 _3532_ (.A1(_0876_),
    .A2(_0878_),
    .B1(_0884_),
    .C1(_0636_),
    .X(_0885_));
 sky130_fd_sc_hd__mux2_1 _3533_ (.A0(\as1802.regs[8][8] ),
    .A1(\as1802.regs[9][8] ),
    .S(_0877_),
    .X(_0886_));
 sky130_fd_sc_hd__and3_1 _3534_ (.A(\as1802.regs[10][8] ),
    .B(_0880_),
    .C(_0881_),
    .X(_0887_));
 sky130_fd_sc_hd__a211o_1 _3535_ (.A1(\as1802.regs[11][8] ),
    .A2(_0879_),
    .B1(_0887_),
    .C1(_0883_),
    .X(_0888_));
 sky130_fd_sc_hd__o211a_1 _3536_ (.A1(_0876_),
    .A2(_0886_),
    .B1(_0888_),
    .C1(_0785_),
    .X(_0889_));
 sky130_fd_sc_hd__buf_4 _3537_ (.A(_0632_),
    .X(_0890_));
 sky130_fd_sc_hd__mux2_1 _3538_ (.A0(\as1802.regs[0][8] ),
    .A1(\as1802.regs[1][8] ),
    .S(_0890_),
    .X(_0891_));
 sky130_fd_sc_hd__buf_4 _3539_ (.A(_0820_),
    .X(_0892_));
 sky130_fd_sc_hd__and3_1 _3540_ (.A(\as1802.regs[2][8] ),
    .B(_0880_),
    .C(_0881_),
    .X(_0893_));
 sky130_fd_sc_hd__a211o_1 _3541_ (.A1(\as1802.regs[3][8] ),
    .A2(_0892_),
    .B1(_0893_),
    .C1(_0883_),
    .X(_0894_));
 sky130_fd_sc_hd__o211a_1 _3542_ (.A1(_0876_),
    .A2(_0891_),
    .B1(_0894_),
    .C1(_0785_),
    .X(_0895_));
 sky130_fd_sc_hd__clkbuf_4 _3543_ (.A(_0636_),
    .X(_0896_));
 sky130_fd_sc_hd__and3_1 _3544_ (.A(\as1802.regs[4][8] ),
    .B(_0880_),
    .C(_0881_),
    .X(_0897_));
 sky130_fd_sc_hd__buf_4 _3545_ (.A(_0617_),
    .X(_0898_));
 sky130_fd_sc_hd__a211o_1 _3546_ (.A1(\as1802.regs[5][8] ),
    .A2(_0879_),
    .B1(_0897_),
    .C1(_0898_),
    .X(_0899_));
 sky130_fd_sc_hd__and3_1 _3547_ (.A(\as1802.regs[6][8] ),
    .B(_0880_),
    .C(_0881_),
    .X(_0900_));
 sky130_fd_sc_hd__a211o_1 _3548_ (.A1(\as1802.regs[7][8] ),
    .A2(_0879_),
    .B1(_0900_),
    .C1(_0883_),
    .X(_0901_));
 sky130_fd_sc_hd__a31o_1 _3549_ (.A1(_0896_),
    .A2(_0899_),
    .A3(_0901_),
    .B1(_0648_),
    .X(_0902_));
 sky130_fd_sc_hd__o32ai_4 _3550_ (.A1(_0708_),
    .A2(_0885_),
    .A3(_0889_),
    .B1(_0895_),
    .B2(_0902_),
    .Y(_0903_));
 sky130_fd_sc_hd__buf_4 _3551_ (.A(_0903_),
    .X(_0904_));
 sky130_fd_sc_hd__xnor2_1 _3552_ (.A(_0875_),
    .B(_0904_),
    .Y(_0905_));
 sky130_fd_sc_hd__xor2_1 _3553_ (.A(_0834_),
    .B(_0904_),
    .X(_0906_));
 sky130_fd_sc_hd__nand2_1 _3554_ (.A(_2696_),
    .B(_0855_),
    .Y(_0907_));
 sky130_fd_sc_hd__and2b_1 _3555_ (.A_N(_2683_),
    .B(\as1802.regs[10][8] ),
    .X(_0908_));
 sky130_fd_sc_hd__a21bo_1 _3556_ (.A1(_2681_),
    .A2(\as1802.regs[11][8] ),
    .B1_N(_2685_),
    .X(_0909_));
 sky130_fd_sc_hd__mux2_1 _3557_ (.A0(\as1802.regs[8][8] ),
    .A1(\as1802.regs[9][8] ),
    .S(_2683_),
    .X(_0910_));
 sky130_fd_sc_hd__buf_4 _3558_ (.A(_2685_),
    .X(_0911_));
 sky130_fd_sc_hd__buf_4 _3559_ (.A(_2689_),
    .X(_0912_));
 sky130_fd_sc_hd__o221a_1 _3560_ (.A1(_0908_),
    .A2(_0909_),
    .B1(_0910_),
    .B2(_0911_),
    .C1(_0912_),
    .X(_0913_));
 sky130_fd_sc_hd__mux4_1 _3561_ (.A0(\as1802.regs[12][8] ),
    .A1(\as1802.regs[13][8] ),
    .A2(\as1802.regs[14][8] ),
    .A3(\as1802.regs[15][8] ),
    .S0(_2683_),
    .S1(_2685_),
    .X(_0914_));
 sky130_fd_sc_hd__a21o_1 _3562_ (.A1(_2678_),
    .A2(_0914_),
    .B1(_2667_),
    .X(_0915_));
 sky130_fd_sc_hd__mux4_1 _3563_ (.A0(\as1802.regs[0][8] ),
    .A1(\as1802.regs[1][8] ),
    .A2(\as1802.regs[2][8] ),
    .A3(\as1802.regs[3][8] ),
    .S0(_2683_),
    .S1(_2674_),
    .X(_0916_));
 sky130_fd_sc_hd__mux4_1 _3564_ (.A0(\as1802.regs[4][8] ),
    .A1(\as1802.regs[5][8] ),
    .A2(\as1802.regs[6][8] ),
    .A3(\as1802.regs[7][8] ),
    .S0(_2670_),
    .S1(_2674_),
    .X(_0917_));
 sky130_fd_sc_hd__mux2_1 _3565_ (.A0(_0916_),
    .A1(_0917_),
    .S(_2678_),
    .X(_0918_));
 sky130_fd_sc_hd__o22ai_4 _3566_ (.A1(_0913_),
    .A2(_0915_),
    .B1(_0918_),
    .B2(_2691_),
    .Y(_0919_));
 sky130_fd_sc_hd__inv_2 _3567_ (.A(_0919_),
    .Y(_0920_));
 sky130_fd_sc_hd__xnor2_1 _3568_ (.A(_0907_),
    .B(_0920_),
    .Y(_0921_));
 sky130_fd_sc_hd__a21oi_4 _3569_ (.A1(_2493_),
    .A2(_0529_),
    .B1(_2718_),
    .Y(_0922_));
 sky130_fd_sc_hd__and3_1 _3570_ (.A(_2718_),
    .B(_0855_),
    .C(_0920_),
    .X(_0923_));
 sky130_fd_sc_hd__o2bb2a_1 _3571_ (.A1_N(_2718_),
    .A2_N(_0855_),
    .B1(_0919_),
    .B2(_0922_),
    .X(_0924_));
 sky130_fd_sc_hd__o2bb2a_1 _3572_ (.A1_N(_0921_),
    .A2_N(_0922_),
    .B1(_0923_),
    .B2(_0924_),
    .X(_0925_));
 sky130_fd_sc_hd__nor2_1 _3573_ (.A(_0378_),
    .B(_0925_),
    .Y(_0926_));
 sky130_fd_sc_hd__a211o_1 _3574_ (.A1(_2702_),
    .A2(_0536_),
    .B1(_0365_),
    .C1(_0926_),
    .X(_0927_));
 sky130_fd_sc_hd__nor2_1 _3575_ (.A(_2555_),
    .B(_0919_),
    .Y(_0928_));
 sky130_fd_sc_hd__a211o_1 _3576_ (.A1(_2555_),
    .A2(_0921_),
    .B1(_0928_),
    .C1(_2700_),
    .X(_0929_));
 sky130_fd_sc_hd__a21o_1 _3577_ (.A1(_0927_),
    .A2(_0929_),
    .B1(_0369_),
    .X(_0930_));
 sky130_fd_sc_hd__o211ai_1 _3578_ (.A1(_0534_),
    .A2(_0921_),
    .B1(_0930_),
    .C1(_0380_),
    .Y(_0931_));
 sky130_fd_sc_hd__o211a_1 _3579_ (.A1(_2606_),
    .A2(_0906_),
    .B1(_0931_),
    .C1(_0415_),
    .X(_0932_));
 sky130_fd_sc_hd__a21bo_1 _3580_ (.A1(_0575_),
    .A2(_0905_),
    .B1_N(_0932_),
    .X(_0933_));
 sky130_fd_sc_hd__or2_1 _3581_ (.A(net14),
    .B(_0385_),
    .X(_0934_));
 sky130_fd_sc_hd__clkbuf_4 _3582_ (.A(_0934_),
    .X(_0935_));
 sky130_fd_sc_hd__nor2_1 _3583_ (.A(_0446_),
    .B(_0906_),
    .Y(_0936_));
 sky130_fd_sc_hd__a211o_1 _3584_ (.A1(_0447_),
    .A2(_0905_),
    .B1(_0936_),
    .C1(_0386_),
    .X(_0937_));
 sky130_fd_sc_hd__o211a_1 _3585_ (.A1(_0382_),
    .A2(_0935_),
    .B1(_0647_),
    .C1(_0937_),
    .X(_0938_));
 sky130_fd_sc_hd__o2bb2a_2 _3586_ (.A1_N(_0873_),
    .A2_N(_0874_),
    .B1(_0933_),
    .B2(_0938_),
    .X(_0939_));
 sky130_fd_sc_hd__buf_2 _3587_ (.A(_0939_),
    .X(_0940_));
 sky130_fd_sc_hd__nor2_2 _3588_ (.A(_0399_),
    .B(_0401_),
    .Y(_0941_));
 sky130_fd_sc_hd__o21a_1 _3589_ (.A1(\as1802.X[2] ),
    .A2(_2607_),
    .B1(_0407_),
    .X(_0942_));
 sky130_fd_sc_hd__nor2_2 _3590_ (.A(_0405_),
    .B(_0942_),
    .Y(_0943_));
 sky130_fd_sc_hd__or4_1 _3591_ (.A(_2456_),
    .B(_0374_),
    .C(_0536_),
    .D(_0388_),
    .X(_0944_));
 sky130_fd_sc_hd__or3_2 _3592_ (.A(_2595_),
    .B(_0391_),
    .C(_0944_),
    .X(_0945_));
 sky130_fd_sc_hd__and3_1 _3593_ (.A(_0941_),
    .B(_0943_),
    .C(_0945_),
    .X(_0946_));
 sky130_fd_sc_hd__buf_4 _3594_ (.A(_0946_),
    .X(_0947_));
 sky130_fd_sc_hd__mux2_1 _3595_ (.A0(\as1802.regs[10][8] ),
    .A1(_0940_),
    .S(_0947_),
    .X(_0948_));
 sky130_fd_sc_hd__clkbuf_1 _3596_ (.A(_0948_),
    .X(_0020_));
 sky130_fd_sc_hd__a21oi_1 _3597_ (.A1(\as1802.regs[2][9] ),
    .A2(_0874_),
    .B1(_0416_),
    .Y(_0949_));
 sky130_fd_sc_hd__or2_1 _3598_ (.A(\as1802.regs[2][9] ),
    .B(_0874_),
    .X(_0950_));
 sky130_fd_sc_hd__mux2_1 _3599_ (.A0(\as1802.regs[0][9] ),
    .A1(\as1802.regs[1][9] ),
    .S(_0820_),
    .X(_0951_));
 sky130_fd_sc_hd__and3_1 _3600_ (.A(\as1802.regs[2][9] ),
    .B(_0821_),
    .C(_0822_),
    .X(_0952_));
 sky130_fd_sc_hd__a211o_1 _3601_ (.A1(\as1802.regs[3][9] ),
    .A2(_0890_),
    .B1(_0952_),
    .C1(_0685_),
    .X(_0953_));
 sky130_fd_sc_hd__o211a_1 _3602_ (.A1(_0898_),
    .A2(_0951_),
    .B1(_0953_),
    .C1(_0785_),
    .X(_0954_));
 sky130_fd_sc_hd__and3_1 _3603_ (.A(\as1802.regs[4][9] ),
    .B(_0821_),
    .C(_0822_),
    .X(_0955_));
 sky130_fd_sc_hd__a211o_1 _3604_ (.A1(\as1802.regs[5][9] ),
    .A2(_0890_),
    .B1(_0955_),
    .C1(_0617_),
    .X(_0956_));
 sky130_fd_sc_hd__and3_1 _3605_ (.A(\as1802.regs[6][9] ),
    .B(_0821_),
    .C(_0822_),
    .X(_0957_));
 sky130_fd_sc_hd__a211o_1 _3606_ (.A1(\as1802.regs[7][9] ),
    .A2(_0890_),
    .B1(_0957_),
    .C1(_0685_),
    .X(_0958_));
 sky130_fd_sc_hd__a31o_1 _3607_ (.A1(_0636_),
    .A2(_0956_),
    .A3(_0958_),
    .B1(_0648_),
    .X(_0959_));
 sky130_fd_sc_hd__mux2_1 _3608_ (.A0(\as1802.regs[12][9] ),
    .A1(\as1802.regs[13][9] ),
    .S(_0877_),
    .X(_0960_));
 sky130_fd_sc_hd__and3_1 _3609_ (.A(\as1802.regs[14][9] ),
    .B(_0880_),
    .C(_0881_),
    .X(_0961_));
 sky130_fd_sc_hd__a211o_1 _3610_ (.A1(\as1802.regs[15][9] ),
    .A2(_0879_),
    .B1(_0961_),
    .C1(_0685_),
    .X(_0962_));
 sky130_fd_sc_hd__o211a_1 _3611_ (.A1(_0876_),
    .A2(_0960_),
    .B1(_0962_),
    .C1(_0636_),
    .X(_0963_));
 sky130_fd_sc_hd__and3_1 _3612_ (.A(\as1802.regs[10][9] ),
    .B(_0880_),
    .C(_0881_),
    .X(_0964_));
 sky130_fd_sc_hd__a211o_1 _3613_ (.A1(\as1802.regs[11][9] ),
    .A2(_0879_),
    .B1(_0964_),
    .C1(_0685_),
    .X(_0965_));
 sky130_fd_sc_hd__and3_1 _3614_ (.A(\as1802.regs[8][9] ),
    .B(_0880_),
    .C(_0881_),
    .X(_0966_));
 sky130_fd_sc_hd__a211o_1 _3615_ (.A1(\as1802.regs[9][9] ),
    .A2(_0879_),
    .B1(_0966_),
    .C1(_0898_),
    .X(_0967_));
 sky130_fd_sc_hd__a31o_1 _3616_ (.A1(_0785_),
    .A2(_0965_),
    .A3(_0967_),
    .B1(_0708_),
    .X(_0968_));
 sky130_fd_sc_hd__o22ai_4 _3617_ (.A1(_0954_),
    .A2(_0959_),
    .B1(_0963_),
    .B2(_0968_),
    .Y(_0969_));
 sky130_fd_sc_hd__o31a_1 _3618_ (.A1(_0837_),
    .A2(_0831_),
    .A3(_0904_),
    .B1(_0969_),
    .X(_0970_));
 sky130_fd_sc_hd__or4_1 _3619_ (.A(_0837_),
    .B(_0831_),
    .C(_0904_),
    .D(_0969_),
    .X(_0971_));
 sky130_fd_sc_hd__and2b_1 _3620_ (.A_N(_0970_),
    .B(_0971_),
    .X(_0972_));
 sky130_fd_sc_hd__and4_1 _3621_ (.A(_0571_),
    .B(_0642_),
    .C(_0833_),
    .D(_0903_),
    .X(_0973_));
 sky130_fd_sc_hd__buf_2 _3622_ (.A(_0973_),
    .X(_0974_));
 sky130_fd_sc_hd__xnor2_1 _3623_ (.A(_0974_),
    .B(_0969_),
    .Y(_0975_));
 sky130_fd_sc_hd__a21o_2 _3624_ (.A1(_2493_),
    .A2(_0529_),
    .B1(_2718_),
    .X(_0976_));
 sky130_fd_sc_hd__clkbuf_4 _3625_ (.A(_2683_),
    .X(_0977_));
 sky130_fd_sc_hd__and2b_1 _3626_ (.A_N(_0977_),
    .B(\as1802.regs[10][9] ),
    .X(_0978_));
 sky130_fd_sc_hd__a21bo_1 _3627_ (.A1(_0977_),
    .A2(\as1802.regs[11][9] ),
    .B1_N(_2685_),
    .X(_0979_));
 sky130_fd_sc_hd__mux2_1 _3628_ (.A0(\as1802.regs[8][9] ),
    .A1(\as1802.regs[9][9] ),
    .S(_0977_),
    .X(_0980_));
 sky130_fd_sc_hd__clkbuf_4 _3629_ (.A(_2685_),
    .X(_0981_));
 sky130_fd_sc_hd__o221a_1 _3630_ (.A1(_0978_),
    .A2(_0979_),
    .B1(_0980_),
    .B2(_0981_),
    .C1(_0912_),
    .X(_0982_));
 sky130_fd_sc_hd__buf_4 _3631_ (.A(_2678_),
    .X(_0983_));
 sky130_fd_sc_hd__mux4_1 _3632_ (.A0(\as1802.regs[12][9] ),
    .A1(\as1802.regs[13][9] ),
    .A2(\as1802.regs[14][9] ),
    .A3(\as1802.regs[15][9] ),
    .S0(_2681_),
    .S1(_0911_),
    .X(_0984_));
 sky130_fd_sc_hd__a21o_1 _3633_ (.A1(_0983_),
    .A2(_0984_),
    .B1(_2667_),
    .X(_0985_));
 sky130_fd_sc_hd__mux4_1 _3634_ (.A0(\as1802.regs[0][9] ),
    .A1(\as1802.regs[1][9] ),
    .A2(\as1802.regs[2][9] ),
    .A3(\as1802.regs[3][9] ),
    .S0(_2681_),
    .S1(_2685_),
    .X(_0986_));
 sky130_fd_sc_hd__mux4_1 _3635_ (.A0(\as1802.regs[4][9] ),
    .A1(\as1802.regs[5][9] ),
    .A2(\as1802.regs[6][9] ),
    .A3(\as1802.regs[7][9] ),
    .S0(_2681_),
    .S1(_2685_),
    .X(_0987_));
 sky130_fd_sc_hd__mux2_1 _3636_ (.A0(_0986_),
    .A1(_0987_),
    .S(_0983_),
    .X(_0988_));
 sky130_fd_sc_hd__o22a_2 _3637_ (.A1(_0982_),
    .A2(_0985_),
    .B1(_0988_),
    .B2(_2691_),
    .X(_0989_));
 sky130_fd_sc_hd__a31o_1 _3638_ (.A1(_2696_),
    .A2(_0855_),
    .A3(_0920_),
    .B1(_0989_),
    .X(_0990_));
 sky130_fd_sc_hd__nand4_1 _3639_ (.A(_2694_),
    .B(_0855_),
    .C(_0920_),
    .D(_0989_),
    .Y(_0991_));
 sky130_fd_sc_hd__and2_1 _3640_ (.A(_0990_),
    .B(_0991_),
    .X(_0992_));
 sky130_fd_sc_hd__nand2_2 _3641_ (.A(\as1802.instr_cycle[1] ),
    .B(_0377_),
    .Y(_0993_));
 sky130_fd_sc_hd__o31a_1 _3642_ (.A1(_0922_),
    .A2(_0923_),
    .A3(_0989_),
    .B1(_0993_),
    .X(_0994_));
 sky130_fd_sc_hd__nand2_1 _3643_ (.A(_0923_),
    .B(_0989_),
    .Y(_0995_));
 sky130_fd_sc_hd__o211a_1 _3644_ (.A1(_0976_),
    .A2(_0992_),
    .B1(_0994_),
    .C1(_0995_),
    .X(_0996_));
 sky130_fd_sc_hd__a211o_1 _3645_ (.A1(_0474_),
    .A2(_0536_),
    .B1(_0365_),
    .C1(_0996_),
    .X(_0997_));
 sky130_fd_sc_hd__inv_2 _3646_ (.A(_0989_),
    .Y(_0998_));
 sky130_fd_sc_hd__nor2_1 _3647_ (.A(_2555_),
    .B(_0998_),
    .Y(_0999_));
 sky130_fd_sc_hd__a211o_1 _3648_ (.A1(_0453_),
    .A2(_0992_),
    .B1(_0999_),
    .C1(_2700_),
    .X(_1000_));
 sky130_fd_sc_hd__and3_1 _3649_ (.A(_0379_),
    .B(_0997_),
    .C(_1000_),
    .X(_1001_));
 sky130_fd_sc_hd__or2_1 _3650_ (.A(_2596_),
    .B(_1001_),
    .X(_1002_));
 sky130_fd_sc_hd__a221o_1 _3651_ (.A1(_0450_),
    .A2(_0972_),
    .B1(_0975_),
    .B2(_0454_),
    .C1(_1002_),
    .X(_1003_));
 sky130_fd_sc_hd__mux2_1 _3652_ (.A0(_0972_),
    .A1(_0975_),
    .S(_0455_),
    .X(_1004_));
 sky130_fd_sc_hd__or2_1 _3653_ (.A(_0452_),
    .B(_0935_),
    .X(_1005_));
 sky130_fd_sc_hd__o211a_1 _3654_ (.A1(_0386_),
    .A2(_1004_),
    .B1(_1005_),
    .C1(_0647_),
    .X(_1006_));
 sky130_fd_sc_hd__o2bb2a_2 _3655_ (.A1_N(_0949_),
    .A2_N(_0950_),
    .B1(_1003_),
    .B2(_1006_),
    .X(_1007_));
 sky130_fd_sc_hd__buf_2 _3656_ (.A(_1007_),
    .X(_1008_));
 sky130_fd_sc_hd__mux2_1 _3657_ (.A0(\as1802.regs[10][9] ),
    .A1(_1008_),
    .S(_0947_),
    .X(_1009_));
 sky130_fd_sc_hd__clkbuf_1 _3658_ (.A(_1009_),
    .X(_0021_));
 sky130_fd_sc_hd__xnor2_1 _3659_ (.A(\as1802.regs[2][10] ),
    .B(_0950_),
    .Y(_1010_));
 sky130_fd_sc_hd__mux2_1 _3660_ (.A0(\as1802.regs[0][10] ),
    .A1(\as1802.regs[1][10] ),
    .S(_0879_),
    .X(_1011_));
 sky130_fd_sc_hd__buf_2 _3661_ (.A(_0821_),
    .X(_1012_));
 sky130_fd_sc_hd__buf_2 _3662_ (.A(_0822_),
    .X(_1013_));
 sky130_fd_sc_hd__and3_1 _3663_ (.A(\as1802.regs[2][10] ),
    .B(_1012_),
    .C(_1013_),
    .X(_1014_));
 sky130_fd_sc_hd__a211o_1 _3664_ (.A1(\as1802.regs[3][10] ),
    .A2(_0892_),
    .B1(_1014_),
    .C1(_0883_),
    .X(_1015_));
 sky130_fd_sc_hd__o211a_1 _3665_ (.A1(_0876_),
    .A2(_1011_),
    .B1(_1015_),
    .C1(_0785_),
    .X(_1016_));
 sky130_fd_sc_hd__and3_1 _3666_ (.A(\as1802.regs[6][10] ),
    .B(_0880_),
    .C(_0881_),
    .X(_1017_));
 sky130_fd_sc_hd__a211o_1 _3667_ (.A1(\as1802.regs[7][10] ),
    .A2(_0892_),
    .B1(_1017_),
    .C1(_0883_),
    .X(_1018_));
 sky130_fd_sc_hd__and3_1 _3668_ (.A(\as1802.regs[4][10] ),
    .B(_0880_),
    .C(_0881_),
    .X(_1019_));
 sky130_fd_sc_hd__a211o_1 _3669_ (.A1(\as1802.regs[5][10] ),
    .A2(_0892_),
    .B1(_1019_),
    .C1(_0898_),
    .X(_1020_));
 sky130_fd_sc_hd__a31o_1 _3670_ (.A1(_0896_),
    .A2(_1018_),
    .A3(_1020_),
    .B1(_0648_),
    .X(_1021_));
 sky130_fd_sc_hd__mux2_1 _3671_ (.A0(\as1802.regs[8][10] ),
    .A1(\as1802.regs[9][10] ),
    .S(_0879_),
    .X(_1022_));
 sky130_fd_sc_hd__and3_1 _3672_ (.A(\as1802.regs[10][10] ),
    .B(_1012_),
    .C(_1013_),
    .X(_1023_));
 sky130_fd_sc_hd__a211o_1 _3673_ (.A1(\as1802.regs[11][10] ),
    .A2(_0892_),
    .B1(_1023_),
    .C1(_0883_),
    .X(_1024_));
 sky130_fd_sc_hd__clkbuf_4 _3674_ (.A(_0785_),
    .X(_1025_));
 sky130_fd_sc_hd__o211a_1 _3675_ (.A1(_0876_),
    .A2(_1022_),
    .B1(_1024_),
    .C1(_1025_),
    .X(_1026_));
 sky130_fd_sc_hd__mux2_1 _3676_ (.A0(\as1802.regs[14][10] ),
    .A1(\as1802.regs[15][10] ),
    .S(_0820_),
    .X(_1027_));
 sky130_fd_sc_hd__mux2_1 _3677_ (.A0(\as1802.regs[12][10] ),
    .A1(\as1802.regs[13][10] ),
    .S(_0820_),
    .X(_1028_));
 sky130_fd_sc_hd__mux2_1 _3678_ (.A0(_1027_),
    .A1(_1028_),
    .S(_0883_),
    .X(_1029_));
 sky130_fd_sc_hd__a21o_1 _3679_ (.A1(_0896_),
    .A2(_1029_),
    .B1(_0708_),
    .X(_1030_));
 sky130_fd_sc_hd__o22a_1 _3680_ (.A1(_1016_),
    .A2(_1021_),
    .B1(_1026_),
    .B2(_1030_),
    .X(_1031_));
 sky130_fd_sc_hd__clkbuf_4 _3681_ (.A(_1031_),
    .X(_1032_));
 sky130_fd_sc_hd__xnor2_1 _3682_ (.A(_0971_),
    .B(_1032_),
    .Y(_1033_));
 sky130_fd_sc_hd__inv_2 _3683_ (.A(_0969_),
    .Y(_1034_));
 sky130_fd_sc_hd__nor2_1 _3684_ (.A(_1034_),
    .B(_1032_),
    .Y(_1035_));
 sky130_fd_sc_hd__nand2_1 _3685_ (.A(_0974_),
    .B(_1035_),
    .Y(_1036_));
 sky130_fd_sc_hd__a21bo_1 _3686_ (.A1(_0974_),
    .A2(_0969_),
    .B1_N(_1032_),
    .X(_1037_));
 sky130_fd_sc_hd__a21oi_1 _3687_ (.A1(_1036_),
    .A2(_1037_),
    .B1(_0447_),
    .Y(_1038_));
 sky130_fd_sc_hd__a211o_1 _3688_ (.A1(_0447_),
    .A2(_1033_),
    .B1(_1038_),
    .C1(_0386_),
    .X(_1039_));
 sky130_fd_sc_hd__or2_1 _3689_ (.A(_0539_),
    .B(_0935_),
    .X(_1040_));
 sky130_fd_sc_hd__and2b_1 _3690_ (.A_N(_2683_),
    .B(\as1802.regs[10][10] ),
    .X(_1041_));
 sky130_fd_sc_hd__a21bo_1 _3691_ (.A1(_2683_),
    .A2(\as1802.regs[11][10] ),
    .B1_N(_2674_),
    .X(_1042_));
 sky130_fd_sc_hd__mux2_1 _3692_ (.A0(\as1802.regs[8][10] ),
    .A1(\as1802.regs[9][10] ),
    .S(_2683_),
    .X(_1043_));
 sky130_fd_sc_hd__o221a_1 _3693_ (.A1(_1041_),
    .A2(_1042_),
    .B1(_1043_),
    .B2(_0911_),
    .C1(_0912_),
    .X(_1044_));
 sky130_fd_sc_hd__mux4_1 _3694_ (.A0(\as1802.regs[12][10] ),
    .A1(\as1802.regs[13][10] ),
    .A2(\as1802.regs[14][10] ),
    .A3(\as1802.regs[15][10] ),
    .S0(_2683_),
    .S1(_2685_),
    .X(_1045_));
 sky130_fd_sc_hd__a21o_1 _3695_ (.A1(_2678_),
    .A2(_1045_),
    .B1(_2667_),
    .X(_1046_));
 sky130_fd_sc_hd__mux4_1 _3696_ (.A0(\as1802.regs[4][10] ),
    .A1(\as1802.regs[5][10] ),
    .A2(\as1802.regs[6][10] ),
    .A3(\as1802.regs[7][10] ),
    .S0(_2670_),
    .S1(_2674_),
    .X(_1047_));
 sky130_fd_sc_hd__mux4_1 _3697_ (.A0(\as1802.regs[0][10] ),
    .A1(\as1802.regs[1][10] ),
    .A2(\as1802.regs[2][10] ),
    .A3(\as1802.regs[3][10] ),
    .S0(_2670_),
    .S1(_2674_),
    .X(_1048_));
 sky130_fd_sc_hd__mux2_1 _3698_ (.A0(_1047_),
    .A1(_1048_),
    .S(_2689_),
    .X(_1049_));
 sky130_fd_sc_hd__o22ai_4 _3699_ (.A1(_1044_),
    .A2(_1046_),
    .B1(_1049_),
    .B2(_2691_),
    .Y(_1050_));
 sky130_fd_sc_hd__nand2_1 _3700_ (.A(_0991_),
    .B(_1050_),
    .Y(_1051_));
 sky130_fd_sc_hd__inv_2 _3701_ (.A(_1050_),
    .Y(_1052_));
 sky130_fd_sc_hd__and4_1 _3702_ (.A(_0855_),
    .B(_0920_),
    .C(_0989_),
    .D(_1052_),
    .X(_1053_));
 sky130_fd_sc_hd__nand2_1 _3703_ (.A(_2696_),
    .B(_1053_),
    .Y(_1054_));
 sky130_fd_sc_hd__and2_1 _3704_ (.A(_1051_),
    .B(_1054_),
    .X(_1055_));
 sky130_fd_sc_hd__nand2_1 _3705_ (.A(_0922_),
    .B(_1055_),
    .Y(_1056_));
 sky130_fd_sc_hd__a221o_1 _3706_ (.A1(_0995_),
    .A2(_1050_),
    .B1(_1053_),
    .B2(_2719_),
    .C1(_0922_),
    .X(_1057_));
 sky130_fd_sc_hd__a21oi_1 _3707_ (.A1(_1056_),
    .A2(_1057_),
    .B1(_0536_),
    .Y(_1058_));
 sky130_fd_sc_hd__a211o_1 _3708_ (.A1(io_out[2]),
    .A2(_0536_),
    .B1(_0365_),
    .C1(_1058_),
    .X(_1059_));
 sky130_fd_sc_hd__nor2_1 _3709_ (.A(_0453_),
    .B(_1050_),
    .Y(_1060_));
 sky130_fd_sc_hd__a211o_1 _3710_ (.A1(_0453_),
    .A2(_1055_),
    .B1(_1060_),
    .C1(_2701_),
    .X(_1061_));
 sky130_fd_sc_hd__a21o_1 _3711_ (.A1(_1059_),
    .A2(_1061_),
    .B1(_0369_),
    .X(_1062_));
 sky130_fd_sc_hd__or4bb_1 _3712_ (.A(_1055_),
    .B(_2598_),
    .C_N(_2545_),
    .D_N(_2556_),
    .X(_1063_));
 sky130_fd_sc_hd__a31o_1 _3713_ (.A1(_0380_),
    .A2(_1062_),
    .A3(_1063_),
    .B1(_0391_),
    .X(_1064_));
 sky130_fd_sc_hd__a31o_1 _3714_ (.A1(_0647_),
    .A2(_1039_),
    .A3(_1040_),
    .B1(_1064_),
    .X(_1065_));
 sky130_fd_sc_hd__and3_1 _3715_ (.A(_0454_),
    .B(_1036_),
    .C(_1037_),
    .X(_1066_));
 sky130_fd_sc_hd__o21ba_1 _3716_ (.A1(_0390_),
    .A2(_1033_),
    .B1_N(_1066_),
    .X(_1067_));
 sky130_fd_sc_hd__a22o_2 _3717_ (.A1(_2597_),
    .A2(_1010_),
    .B1(_1065_),
    .B2(_1067_),
    .X(_1068_));
 sky130_fd_sc_hd__buf_2 _3718_ (.A(_1068_),
    .X(_1069_));
 sky130_fd_sc_hd__mux2_1 _3719_ (.A0(\as1802.regs[10][10] ),
    .A1(_1069_),
    .S(_0947_),
    .X(_1070_));
 sky130_fd_sc_hd__clkbuf_1 _3720_ (.A(_1070_),
    .X(_0022_));
 sky130_fd_sc_hd__nor2_1 _3721_ (.A(_0904_),
    .B(_0969_),
    .Y(_1071_));
 sky130_fd_sc_hd__and4b_1 _3722_ (.A_N(_0837_),
    .B(_0832_),
    .C(_1071_),
    .D(_1032_),
    .X(_1072_));
 sky130_fd_sc_hd__mux2_1 _3723_ (.A0(\as1802.regs[4][11] ),
    .A1(\as1802.regs[5][11] ),
    .S(_0892_),
    .X(_1073_));
 sky130_fd_sc_hd__buf_4 _3724_ (.A(_0877_),
    .X(_1074_));
 sky130_fd_sc_hd__and3_1 _3725_ (.A(\as1802.regs[6][11] ),
    .B(_1012_),
    .C(_1013_),
    .X(_1075_));
 sky130_fd_sc_hd__a211o_1 _3726_ (.A1(\as1802.regs[7][11] ),
    .A2(_1074_),
    .B1(_1075_),
    .C1(_0883_),
    .X(_1076_));
 sky130_fd_sc_hd__o211a_1 _3727_ (.A1(_0876_),
    .A2(_1073_),
    .B1(_1076_),
    .C1(_0896_),
    .X(_1077_));
 sky130_fd_sc_hd__mux2_1 _3728_ (.A0(\as1802.regs[0][11] ),
    .A1(\as1802.regs[1][11] ),
    .S(_0892_),
    .X(_1078_));
 sky130_fd_sc_hd__and3_1 _3729_ (.A(\as1802.regs[2][11] ),
    .B(_1012_),
    .C(_1013_),
    .X(_1079_));
 sky130_fd_sc_hd__a211o_1 _3730_ (.A1(\as1802.regs[3][11] ),
    .A2(_1074_),
    .B1(_1079_),
    .C1(_0883_),
    .X(_1080_));
 sky130_fd_sc_hd__o211a_1 _3731_ (.A1(_0876_),
    .A2(_1078_),
    .B1(_1080_),
    .C1(_1025_),
    .X(_1081_));
 sky130_fd_sc_hd__clkbuf_4 _3732_ (.A(_0898_),
    .X(_1082_));
 sky130_fd_sc_hd__mux2_1 _3733_ (.A0(\as1802.regs[8][11] ),
    .A1(\as1802.regs[9][11] ),
    .S(_0892_),
    .X(_1083_));
 sky130_fd_sc_hd__and3_1 _3734_ (.A(\as1802.regs[10][11] ),
    .B(_1012_),
    .C(_1013_),
    .X(_1084_));
 sky130_fd_sc_hd__clkbuf_4 _3735_ (.A(_0685_),
    .X(_1085_));
 sky130_fd_sc_hd__a211o_1 _3736_ (.A1(\as1802.regs[11][11] ),
    .A2(_1074_),
    .B1(_1084_),
    .C1(_1085_),
    .X(_1086_));
 sky130_fd_sc_hd__o211a_1 _3737_ (.A1(_1082_),
    .A2(_1083_),
    .B1(_1086_),
    .C1(_1025_),
    .X(_1087_));
 sky130_fd_sc_hd__mux2_1 _3738_ (.A0(\as1802.regs[12][11] ),
    .A1(\as1802.regs[13][11] ),
    .S(_0820_),
    .X(_1088_));
 sky130_fd_sc_hd__or2_1 _3739_ (.A(_0898_),
    .B(_1088_),
    .X(_1089_));
 sky130_fd_sc_hd__mux2_1 _3740_ (.A0(\as1802.regs[14][11] ),
    .A1(\as1802.regs[15][11] ),
    .S(_0820_),
    .X(_1090_));
 sky130_fd_sc_hd__or2_1 _3741_ (.A(_1085_),
    .B(_1090_),
    .X(_1091_));
 sky130_fd_sc_hd__a31o_1 _3742_ (.A1(_0896_),
    .A2(_1089_),
    .A3(_1091_),
    .B1(_0708_),
    .X(_1092_));
 sky130_fd_sc_hd__o32a_4 _3743_ (.A1(_0648_),
    .A2(_1077_),
    .A3(_1081_),
    .B1(_1087_),
    .B2(_1092_),
    .X(_1093_));
 sky130_fd_sc_hd__nand3_1 _3744_ (.A(_1034_),
    .B(_1031_),
    .C(_1093_),
    .Y(_1094_));
 sky130_fd_sc_hd__or4_2 _3745_ (.A(_0837_),
    .B(_0831_),
    .C(_0904_),
    .D(_1094_),
    .X(_1095_));
 sky130_fd_sc_hd__o21a_1 _3746_ (.A1(_1072_),
    .A2(_1093_),
    .B1(_1095_),
    .X(_1096_));
 sky130_fd_sc_hd__nor3_2 _3747_ (.A(_1034_),
    .B(_1032_),
    .C(_1093_),
    .Y(_1097_));
 sky130_fd_sc_hd__and2_1 _3748_ (.A(_0974_),
    .B(_1097_),
    .X(_1098_));
 sky130_fd_sc_hd__o32ai_4 _3749_ (.A1(_0648_),
    .A2(_1077_),
    .A3(_1081_),
    .B1(_1087_),
    .B2(_1092_),
    .Y(_1099_));
 sky130_fd_sc_hd__a21oi_1 _3750_ (.A1(_0974_),
    .A2(_1035_),
    .B1(_1099_),
    .Y(_1100_));
 sky130_fd_sc_hd__o31a_1 _3751_ (.A1(_0447_),
    .A2(_1098_),
    .A3(_1100_),
    .B1(_0935_),
    .X(_1101_));
 sky130_fd_sc_hd__o21ai_1 _3752_ (.A1(_0455_),
    .A2(_1096_),
    .B1(_1101_),
    .Y(_1102_));
 sky130_fd_sc_hd__nand2_1 _3753_ (.A(_0579_),
    .B(_0386_),
    .Y(_1103_));
 sky130_fd_sc_hd__and2b_1 _3754_ (.A_N(_0977_),
    .B(\as1802.regs[10][11] ),
    .X(_1104_));
 sky130_fd_sc_hd__clkbuf_4 _3755_ (.A(_2681_),
    .X(_1105_));
 sky130_fd_sc_hd__a21bo_1 _3756_ (.A1(_1105_),
    .A2(\as1802.regs[11][11] ),
    .B1_N(_0911_),
    .X(_1106_));
 sky130_fd_sc_hd__mux2_1 _3757_ (.A0(\as1802.regs[8][11] ),
    .A1(\as1802.regs[9][11] ),
    .S(_0977_),
    .X(_1107_));
 sky130_fd_sc_hd__o221a_1 _3758_ (.A1(_1104_),
    .A2(_1106_),
    .B1(_1107_),
    .B2(_0981_),
    .C1(_0912_),
    .X(_1108_));
 sky130_fd_sc_hd__mux4_1 _3759_ (.A0(\as1802.regs[12][11] ),
    .A1(\as1802.regs[13][11] ),
    .A2(\as1802.regs[14][11] ),
    .A3(\as1802.regs[15][11] ),
    .S0(_0977_),
    .S1(_0911_),
    .X(_1109_));
 sky130_fd_sc_hd__a21o_1 _3760_ (.A1(_0983_),
    .A2(_1109_),
    .B1(_2667_),
    .X(_1110_));
 sky130_fd_sc_hd__mux4_1 _3761_ (.A0(\as1802.regs[4][11] ),
    .A1(\as1802.regs[5][11] ),
    .A2(\as1802.regs[6][11] ),
    .A3(\as1802.regs[7][11] ),
    .S0(_2681_),
    .S1(_0911_),
    .X(_1111_));
 sky130_fd_sc_hd__mux4_1 _3762_ (.A0(\as1802.regs[0][11] ),
    .A1(\as1802.regs[1][11] ),
    .A2(\as1802.regs[2][11] ),
    .A3(\as1802.regs[3][11] ),
    .S0(_2681_),
    .S1(_0911_),
    .X(_1112_));
 sky130_fd_sc_hd__mux2_1 _3763_ (.A0(_1111_),
    .A1(_1112_),
    .S(_0912_),
    .X(_1113_));
 sky130_fd_sc_hd__o22a_2 _3764_ (.A1(_1108_),
    .A2(_1110_),
    .B1(_1113_),
    .B2(_2691_),
    .X(_1114_));
 sky130_fd_sc_hd__clkinv_2 _3765_ (.A(_1114_),
    .Y(_1115_));
 sky130_fd_sc_hd__xnor2_1 _3766_ (.A(_1054_),
    .B(_1115_),
    .Y(_1116_));
 sky130_fd_sc_hd__nor2_1 _3767_ (.A(_0922_),
    .B(_1114_),
    .Y(_1117_));
 sky130_fd_sc_hd__nand2_1 _3768_ (.A(_2718_),
    .B(_1053_),
    .Y(_1118_));
 sky130_fd_sc_hd__nor2_1 _3769_ (.A(_1118_),
    .B(_1115_),
    .Y(_1119_));
 sky130_fd_sc_hd__a221o_1 _3770_ (.A1(_0922_),
    .A2(_1116_),
    .B1(_1117_),
    .B2(_1118_),
    .C1(_1119_),
    .X(_1120_));
 sky130_fd_sc_hd__nand2_1 _3771_ (.A(_0993_),
    .B(_1120_),
    .Y(_1121_));
 sky130_fd_sc_hd__o211a_1 _3772_ (.A1(io_out[3]),
    .A2(_0993_),
    .B1(_2701_),
    .C1(_1121_),
    .X(_1122_));
 sky130_fd_sc_hd__nand2_1 _3773_ (.A(_2556_),
    .B(_1116_),
    .Y(_1123_));
 sky130_fd_sc_hd__or2_1 _3774_ (.A(_2555_),
    .B(_1114_),
    .X(_1124_));
 sky130_fd_sc_hd__a31o_1 _3775_ (.A1(_0366_),
    .A2(_1123_),
    .A3(_1124_),
    .B1(_0369_),
    .X(_1125_));
 sky130_fd_sc_hd__o2bb2a_1 _3776_ (.A1_N(_0369_),
    .A2_N(_1116_),
    .B1(_1122_),
    .B2(_1125_),
    .X(_1126_));
 sky130_fd_sc_hd__a21oi_1 _3777_ (.A1(_0380_),
    .A2(_1126_),
    .B1(_0647_),
    .Y(_1127_));
 sky130_fd_sc_hd__a31o_1 _3778_ (.A1(_0647_),
    .A2(_1102_),
    .A3(_1103_),
    .B1(_1127_),
    .X(_1128_));
 sky130_fd_sc_hd__o21a_1 _3779_ (.A1(_1098_),
    .A2(_1100_),
    .B1(_0454_),
    .X(_1129_));
 sky130_fd_sc_hd__a211oi_2 _3780_ (.A1(_0575_),
    .A2(_1096_),
    .B1(_1129_),
    .C1(_2597_),
    .Y(_1130_));
 sky130_fd_sc_hd__or3_1 _3781_ (.A(\as1802.regs[2][10] ),
    .B(\as1802.regs[2][11] ),
    .C(_0950_),
    .X(_1131_));
 sky130_fd_sc_hd__o21ai_1 _3782_ (.A1(\as1802.regs[2][10] ),
    .A2(_0950_),
    .B1(\as1802.regs[2][11] ),
    .Y(_1132_));
 sky130_fd_sc_hd__and3_1 _3783_ (.A(_2597_),
    .B(_1131_),
    .C(_1132_),
    .X(_1133_));
 sky130_fd_sc_hd__a21oi_4 _3784_ (.A1(_1128_),
    .A2(_1130_),
    .B1(_1133_),
    .Y(_1134_));
 sky130_fd_sc_hd__buf_2 _3785_ (.A(_1134_),
    .X(_1135_));
 sky130_fd_sc_hd__mux2_1 _3786_ (.A0(\as1802.regs[10][11] ),
    .A1(_1135_),
    .S(_0947_),
    .X(_1136_));
 sky130_fd_sc_hd__clkbuf_1 _3787_ (.A(_1136_),
    .X(_0023_));
 sky130_fd_sc_hd__mux2_1 _3788_ (.A0(\as1802.regs[0][12] ),
    .A1(\as1802.regs[1][12] ),
    .S(_1074_),
    .X(_1137_));
 sky130_fd_sc_hd__clkbuf_4 _3789_ (.A(_0879_),
    .X(_1138_));
 sky130_fd_sc_hd__and3_1 _3790_ (.A(\as1802.regs[2][12] ),
    .B(_1012_),
    .C(_1013_),
    .X(_1139_));
 sky130_fd_sc_hd__a211o_1 _3791_ (.A1(\as1802.regs[3][12] ),
    .A2(_1138_),
    .B1(_1139_),
    .C1(_1085_),
    .X(_1140_));
 sky130_fd_sc_hd__o211a_1 _3792_ (.A1(_1082_),
    .A2(_1137_),
    .B1(_1140_),
    .C1(_1025_),
    .X(_1141_));
 sky130_fd_sc_hd__mux2_1 _3793_ (.A0(\as1802.regs[4][12] ),
    .A1(\as1802.regs[5][12] ),
    .S(_0877_),
    .X(_1142_));
 sky130_fd_sc_hd__mux2_1 _3794_ (.A0(\as1802.regs[6][12] ),
    .A1(\as1802.regs[7][12] ),
    .S(_0877_),
    .X(_1143_));
 sky130_fd_sc_hd__mux2_1 _3795_ (.A0(_1142_),
    .A1(_1143_),
    .S(_0898_),
    .X(_1144_));
 sky130_fd_sc_hd__a21o_1 _3796_ (.A1(_0896_),
    .A2(_1144_),
    .B1(_0648_),
    .X(_1145_));
 sky130_fd_sc_hd__mux2_1 _3797_ (.A0(\as1802.regs[12][12] ),
    .A1(\as1802.regs[13][12] ),
    .S(_0820_),
    .X(_1146_));
 sky130_fd_sc_hd__and3_1 _3798_ (.A(\as1802.regs[14][12] ),
    .B(_0821_),
    .C(_0822_),
    .X(_1147_));
 sky130_fd_sc_hd__a211o_1 _3799_ (.A1(\as1802.regs[15][12] ),
    .A2(_0890_),
    .B1(_1147_),
    .C1(_0685_),
    .X(_1148_));
 sky130_fd_sc_hd__o211a_1 _3800_ (.A1(_0898_),
    .A2(_1146_),
    .B1(_1148_),
    .C1(_0636_),
    .X(_1149_));
 sky130_fd_sc_hd__mux2_1 _3801_ (.A0(\as1802.regs[8][12] ),
    .A1(\as1802.regs[9][12] ),
    .S(_0877_),
    .X(_1150_));
 sky130_fd_sc_hd__and3_1 _3802_ (.A(\as1802.regs[10][12] ),
    .B(_0821_),
    .C(_0822_),
    .X(_1151_));
 sky130_fd_sc_hd__a211o_1 _3803_ (.A1(\as1802.regs[11][12] ),
    .A2(_0890_),
    .B1(_1151_),
    .C1(_0685_),
    .X(_1152_));
 sky130_fd_sc_hd__o211a_1 _3804_ (.A1(_0876_),
    .A2(_1150_),
    .B1(_1152_),
    .C1(_0785_),
    .X(_1153_));
 sky130_fd_sc_hd__or3_1 _3805_ (.A(_0708_),
    .B(_1149_),
    .C(_1153_),
    .X(_1154_));
 sky130_fd_sc_hd__o21ai_4 _3806_ (.A1(_1141_),
    .A2(_1145_),
    .B1(_1154_),
    .Y(_1155_));
 sky130_fd_sc_hd__xnor2_1 _3807_ (.A(_1095_),
    .B(_1155_),
    .Y(_1156_));
 sky130_fd_sc_hd__xor2_1 _3808_ (.A(_1098_),
    .B(_1155_),
    .X(_1157_));
 sky130_fd_sc_hd__mux2_1 _3809_ (.A0(_1156_),
    .A1(_1157_),
    .S(_0455_),
    .X(_1158_));
 sky130_fd_sc_hd__o21ai_1 _3810_ (.A1(_0646_),
    .A2(_0935_),
    .B1(_0647_),
    .Y(_1159_));
 sky130_fd_sc_hd__a21o_1 _3811_ (.A1(_0935_),
    .A2(_1158_),
    .B1(_1159_),
    .X(_1160_));
 sky130_fd_sc_hd__and2b_1 _3812_ (.A_N(_0977_),
    .B(\as1802.regs[10][12] ),
    .X(_1161_));
 sky130_fd_sc_hd__a21bo_1 _3813_ (.A1(_1105_),
    .A2(\as1802.regs[11][12] ),
    .B1_N(_0911_),
    .X(_1162_));
 sky130_fd_sc_hd__mux2_1 _3814_ (.A0(\as1802.regs[8][12] ),
    .A1(\as1802.regs[9][12] ),
    .S(_0977_),
    .X(_1163_));
 sky130_fd_sc_hd__o221a_1 _3815_ (.A1(_1161_),
    .A2(_1162_),
    .B1(_1163_),
    .B2(_0981_),
    .C1(_0912_),
    .X(_1164_));
 sky130_fd_sc_hd__mux4_1 _3816_ (.A0(\as1802.regs[12][12] ),
    .A1(\as1802.regs[13][12] ),
    .A2(\as1802.regs[14][12] ),
    .A3(\as1802.regs[15][12] ),
    .S0(_0977_),
    .S1(_0981_),
    .X(_1165_));
 sky130_fd_sc_hd__a21o_1 _3817_ (.A1(_0983_),
    .A2(_1165_),
    .B1(_2667_),
    .X(_1166_));
 sky130_fd_sc_hd__mux4_1 _3818_ (.A0(\as1802.regs[0][12] ),
    .A1(\as1802.regs[1][12] ),
    .A2(\as1802.regs[2][12] ),
    .A3(\as1802.regs[3][12] ),
    .S0(_2681_),
    .S1(_0911_),
    .X(_1167_));
 sky130_fd_sc_hd__mux4_1 _3819_ (.A0(\as1802.regs[4][12] ),
    .A1(\as1802.regs[5][12] ),
    .A2(\as1802.regs[6][12] ),
    .A3(\as1802.regs[7][12] ),
    .S0(_2681_),
    .S1(_0911_),
    .X(_1168_));
 sky130_fd_sc_hd__mux2_1 _3820_ (.A0(_1167_),
    .A1(_1168_),
    .S(_0983_),
    .X(_1169_));
 sky130_fd_sc_hd__o22a_2 _3821_ (.A1(_1164_),
    .A2(_1166_),
    .B1(_1169_),
    .B2(_2691_),
    .X(_1170_));
 sky130_fd_sc_hd__inv_2 _3822_ (.A(_1170_),
    .Y(_1171_));
 sky130_fd_sc_hd__a31o_1 _3823_ (.A1(_2696_),
    .A2(_1053_),
    .A3(_1114_),
    .B1(_1170_),
    .X(_1172_));
 sky130_fd_sc_hd__nand2_1 _3824_ (.A(_1114_),
    .B(_1170_),
    .Y(_1173_));
 sky130_fd_sc_hd__or3_1 _3825_ (.A(_0991_),
    .B(_1050_),
    .C(_1173_),
    .X(_1174_));
 sky130_fd_sc_hd__nand2_1 _3826_ (.A(_1172_),
    .B(_1174_),
    .Y(_1175_));
 sky130_fd_sc_hd__mux2_1 _3827_ (.A0(_1171_),
    .A1(_1175_),
    .S(_0453_),
    .X(_1176_));
 sky130_fd_sc_hd__a31o_1 _3828_ (.A1(_2719_),
    .A2(_1053_),
    .A3(_1114_),
    .B1(_1170_),
    .X(_1177_));
 sky130_fd_sc_hd__nand2_1 _3829_ (.A(_0976_),
    .B(_1177_),
    .Y(_1178_));
 sky130_fd_sc_hd__nor2_1 _3830_ (.A(_1118_),
    .B(_1173_),
    .Y(_1179_));
 sky130_fd_sc_hd__o22a_1 _3831_ (.A1(_1178_),
    .A2(_1179_),
    .B1(_1175_),
    .B2(_0976_),
    .X(_1180_));
 sky130_fd_sc_hd__nor2_1 _3832_ (.A(_0536_),
    .B(_1180_),
    .Y(_1181_));
 sky130_fd_sc_hd__a211o_1 _3833_ (.A1(io_out[4]),
    .A2(_0536_),
    .B1(_0365_),
    .C1(_1181_),
    .X(_1182_));
 sky130_fd_sc_hd__a21bo_1 _3834_ (.A1(_0366_),
    .A2(_1176_),
    .B1_N(_1182_),
    .X(_1183_));
 sky130_fd_sc_hd__o21a_1 _3835_ (.A1(_0537_),
    .A2(_1183_),
    .B1(_0416_),
    .X(_1184_));
 sky130_fd_sc_hd__o221a_1 _3836_ (.A1(_0489_),
    .A2(_1156_),
    .B1(_1157_),
    .B2(_2606_),
    .C1(_1184_),
    .X(_1185_));
 sky130_fd_sc_hd__or2_1 _3837_ (.A(\as1802.regs[2][12] ),
    .B(_1131_),
    .X(_1186_));
 sky130_fd_sc_hd__a21oi_1 _3838_ (.A1(\as1802.regs[2][12] ),
    .A2(_1131_),
    .B1(_0416_),
    .Y(_1187_));
 sky130_fd_sc_hd__a22oi_4 _3839_ (.A1(_1160_),
    .A2(_1185_),
    .B1(_1186_),
    .B2(_1187_),
    .Y(_1188_));
 sky130_fd_sc_hd__buf_2 _3840_ (.A(_1188_),
    .X(_1189_));
 sky130_fd_sc_hd__mux2_1 _3841_ (.A0(\as1802.regs[10][12] ),
    .A1(_1189_),
    .S(_0947_),
    .X(_1190_));
 sky130_fd_sc_hd__clkbuf_1 _3842_ (.A(_1190_),
    .X(_0024_));
 sky130_fd_sc_hd__or2_1 _3843_ (.A(\as1802.regs[2][13] ),
    .B(_1186_),
    .X(_1191_));
 sky130_fd_sc_hd__a21oi_1 _3844_ (.A1(\as1802.regs[2][13] ),
    .A2(_1186_),
    .B1(_0416_),
    .Y(_1192_));
 sky130_fd_sc_hd__nand3_1 _3845_ (.A(_1071_),
    .B(_1031_),
    .C(_1093_),
    .Y(_1193_));
 sky130_fd_sc_hd__or4_1 _3846_ (.A(_0837_),
    .B(_0831_),
    .C(_1193_),
    .D(_1155_),
    .X(_1194_));
 sky130_fd_sc_hd__mux2_1 _3847_ (.A0(\as1802.regs[4][13] ),
    .A1(\as1802.regs[5][13] ),
    .S(_1074_),
    .X(_1195_));
 sky130_fd_sc_hd__and3_1 _3848_ (.A(\as1802.regs[6][13] ),
    .B(_1012_),
    .C(_1013_),
    .X(_1196_));
 sky130_fd_sc_hd__a211o_1 _3849_ (.A1(\as1802.regs[7][13] ),
    .A2(_1138_),
    .B1(_1196_),
    .C1(_1085_),
    .X(_1197_));
 sky130_fd_sc_hd__o211a_1 _3850_ (.A1(_1082_),
    .A2(_1195_),
    .B1(_1197_),
    .C1(_0896_),
    .X(_1198_));
 sky130_fd_sc_hd__mux2_1 _3851_ (.A0(\as1802.regs[0][13] ),
    .A1(\as1802.regs[1][13] ),
    .S(_0890_),
    .X(_1199_));
 sky130_fd_sc_hd__mux2_1 _3852_ (.A0(\as1802.regs[2][13] ),
    .A1(\as1802.regs[3][13] ),
    .S(_0877_),
    .X(_1200_));
 sky130_fd_sc_hd__mux2_1 _3853_ (.A0(_1199_),
    .A1(_1200_),
    .S(_0898_),
    .X(_1201_));
 sky130_fd_sc_hd__a21o_1 _3854_ (.A1(_1025_),
    .A2(_1201_),
    .B1(_0648_),
    .X(_1202_));
 sky130_fd_sc_hd__mux2_1 _3855_ (.A0(\as1802.regs[8][13] ),
    .A1(\as1802.regs[9][13] ),
    .S(_0877_),
    .X(_1203_));
 sky130_fd_sc_hd__mux2_1 _3856_ (.A0(\as1802.regs[10][13] ),
    .A1(\as1802.regs[11][13] ),
    .S(_0877_),
    .X(_1204_));
 sky130_fd_sc_hd__mux2_1 _3857_ (.A0(_1203_),
    .A1(_1204_),
    .S(_0898_),
    .X(_1205_));
 sky130_fd_sc_hd__mux2_1 _3858_ (.A0(\as1802.regs[14][13] ),
    .A1(\as1802.regs[15][13] ),
    .S(_0890_),
    .X(_1206_));
 sky130_fd_sc_hd__or2_1 _3859_ (.A(_1085_),
    .B(_1206_),
    .X(_1207_));
 sky130_fd_sc_hd__mux2_1 _3860_ (.A0(\as1802.regs[12][13] ),
    .A1(\as1802.regs[13][13] ),
    .S(_0890_),
    .X(_1208_));
 sky130_fd_sc_hd__o21a_1 _3861_ (.A1(_0876_),
    .A2(_1208_),
    .B1(_0636_),
    .X(_1209_));
 sky130_fd_sc_hd__a22o_1 _3862_ (.A1(_1025_),
    .A2(_1205_),
    .B1(_1207_),
    .B2(_1209_),
    .X(_1210_));
 sky130_fd_sc_hd__o22ai_4 _3863_ (.A1(_1198_),
    .A2(_1202_),
    .B1(_1210_),
    .B2(_0708_),
    .Y(_1211_));
 sky130_fd_sc_hd__or2_1 _3864_ (.A(_1155_),
    .B(_1211_),
    .X(_1212_));
 sky130_fd_sc_hd__nor4_2 _3865_ (.A(_0837_),
    .B(_0831_),
    .C(_1193_),
    .D(_1212_),
    .Y(_1213_));
 sky130_fd_sc_hd__a211o_1 _3866_ (.A1(_1194_),
    .A2(_1211_),
    .B1(_1213_),
    .C1(_0455_),
    .X(_1214_));
 sky130_fd_sc_hd__and2_1 _3867_ (.A(_1155_),
    .B(_1211_),
    .X(_1215_));
 sky130_fd_sc_hd__nand3_1 _3868_ (.A(_0974_),
    .B(_1097_),
    .C(_1215_),
    .Y(_1216_));
 sky130_fd_sc_hd__a31o_1 _3869_ (.A1(_0974_),
    .A2(_1097_),
    .A3(_1155_),
    .B1(_1211_),
    .X(_1217_));
 sky130_fd_sc_hd__a21o_1 _3870_ (.A1(_1216_),
    .A2(_1217_),
    .B1(_0446_),
    .X(_1218_));
 sky130_fd_sc_hd__o21ai_1 _3871_ (.A1(_0716_),
    .A2(_0934_),
    .B1(_0397_),
    .Y(_1219_));
 sky130_fd_sc_hd__a31o_1 _3872_ (.A1(_0935_),
    .A2(_1214_),
    .A3(_1218_),
    .B1(_1219_),
    .X(_1220_));
 sky130_fd_sc_hd__a21o_1 _3873_ (.A1(_1216_),
    .A2(_1217_),
    .B1(_2606_),
    .X(_1221_));
 sky130_fd_sc_hd__mux4_1 _3874_ (.A0(\as1802.regs[0][13] ),
    .A1(\as1802.regs[1][13] ),
    .A2(\as1802.regs[2][13] ),
    .A3(\as1802.regs[3][13] ),
    .S0(_1105_),
    .S1(_0981_),
    .X(_1222_));
 sky130_fd_sc_hd__mux4_1 _3875_ (.A0(\as1802.regs[4][13] ),
    .A1(\as1802.regs[5][13] ),
    .A2(\as1802.regs[6][13] ),
    .A3(\as1802.regs[7][13] ),
    .S0(_1105_),
    .S1(_0981_),
    .X(_1223_));
 sky130_fd_sc_hd__mux2_1 _3876_ (.A0(_1222_),
    .A1(_1223_),
    .S(_0983_),
    .X(_1224_));
 sky130_fd_sc_hd__buf_4 _3877_ (.A(_0977_),
    .X(_1225_));
 sky130_fd_sc_hd__clkbuf_4 _3878_ (.A(_0981_),
    .X(_1226_));
 sky130_fd_sc_hd__mux4_1 _3879_ (.A0(\as1802.regs[12][13] ),
    .A1(\as1802.regs[13][13] ),
    .A2(\as1802.regs[14][13] ),
    .A3(\as1802.regs[15][13] ),
    .S0(_1225_),
    .S1(_1226_),
    .X(_1227_));
 sky130_fd_sc_hd__and2b_1 _3880_ (.A_N(_1105_),
    .B(\as1802.regs[10][13] ),
    .X(_1228_));
 sky130_fd_sc_hd__a21bo_1 _3881_ (.A1(_1105_),
    .A2(\as1802.regs[11][13] ),
    .B1_N(_0981_),
    .X(_1229_));
 sky130_fd_sc_hd__mux2_1 _3882_ (.A0(\as1802.regs[8][13] ),
    .A1(\as1802.regs[9][13] ),
    .S(_1105_),
    .X(_1230_));
 sky130_fd_sc_hd__o221a_1 _3883_ (.A1(_1228_),
    .A2(_1229_),
    .B1(_1230_),
    .B2(_1226_),
    .C1(_0912_),
    .X(_1231_));
 sky130_fd_sc_hd__a211o_1 _3884_ (.A1(_0983_),
    .A2(_1227_),
    .B1(_1231_),
    .C1(_2667_),
    .X(_1232_));
 sky130_fd_sc_hd__o21ai_4 _3885_ (.A1(_2691_),
    .A2(_1224_),
    .B1(_1232_),
    .Y(_1233_));
 sky130_fd_sc_hd__xnor2_1 _3886_ (.A(_1174_),
    .B(_1233_),
    .Y(_1234_));
 sky130_fd_sc_hd__mux2_1 _3887_ (.A0(_1233_),
    .A1(_1234_),
    .S(_2555_),
    .X(_1235_));
 sky130_fd_sc_hd__o211a_1 _3888_ (.A1(_1118_),
    .A2(_1173_),
    .B1(_1233_),
    .C1(_0976_),
    .X(_1236_));
 sky130_fd_sc_hd__nor3_1 _3889_ (.A(_1118_),
    .B(_1173_),
    .C(_1233_),
    .Y(_1237_));
 sky130_fd_sc_hd__a211o_1 _3890_ (.A1(_0922_),
    .A2(_1234_),
    .B1(_1236_),
    .C1(_1237_),
    .X(_1238_));
 sky130_fd_sc_hd__o21ai_1 _3891_ (.A1(io_out[5]),
    .A2(_0993_),
    .B1(_2700_),
    .Y(_1239_));
 sky130_fd_sc_hd__a21o_1 _3892_ (.A1(_0993_),
    .A2(_1238_),
    .B1(_1239_),
    .X(_1240_));
 sky130_fd_sc_hd__o211a_1 _3893_ (.A1(_2700_),
    .A2(_1235_),
    .B1(_1240_),
    .C1(_0534_),
    .X(_1241_));
 sky130_fd_sc_hd__a211o_1 _3894_ (.A1(_0369_),
    .A2(_1234_),
    .B1(_1241_),
    .C1(_0537_),
    .X(_1242_));
 sky130_fd_sc_hd__and3_1 _3895_ (.A(_0415_),
    .B(_1221_),
    .C(_1242_),
    .X(_1243_));
 sky130_fd_sc_hd__a211o_1 _3896_ (.A1(_1194_),
    .A2(_1211_),
    .B1(_1213_),
    .C1(_0390_),
    .X(_1244_));
 sky130_fd_sc_hd__and3_1 _3897_ (.A(_1220_),
    .B(_1243_),
    .C(_1244_),
    .X(_1245_));
 sky130_fd_sc_hd__a21oi_4 _3898_ (.A1(_1191_),
    .A2(_1192_),
    .B1(_1245_),
    .Y(_1246_));
 sky130_fd_sc_hd__buf_2 _3899_ (.A(_1246_),
    .X(_1247_));
 sky130_fd_sc_hd__mux2_1 _3900_ (.A0(\as1802.regs[10][13] ),
    .A1(_1247_),
    .S(_0947_),
    .X(_1248_));
 sky130_fd_sc_hd__clkbuf_1 _3901_ (.A(_1248_),
    .X(_0025_));
 sky130_fd_sc_hd__mux2_1 _3902_ (.A0(\as1802.regs[4][14] ),
    .A1(\as1802.regs[5][14] ),
    .S(_1138_),
    .X(_1249_));
 sky130_fd_sc_hd__and3_1 _3903_ (.A(\as1802.regs[6][14] ),
    .B(_1012_),
    .C(_1013_),
    .X(_1250_));
 sky130_fd_sc_hd__a211o_1 _3904_ (.A1(\as1802.regs[7][14] ),
    .A2(_1138_),
    .B1(_1250_),
    .C1(_1085_),
    .X(_1251_));
 sky130_fd_sc_hd__o211a_1 _3905_ (.A1(_1082_),
    .A2(_1249_),
    .B1(_1251_),
    .C1(_0896_),
    .X(_1252_));
 sky130_fd_sc_hd__mux2_1 _3906_ (.A0(\as1802.regs[0][14] ),
    .A1(\as1802.regs[1][14] ),
    .S(_1138_),
    .X(_1253_));
 sky130_fd_sc_hd__and3_1 _3907_ (.A(\as1802.regs[2][14] ),
    .B(_1012_),
    .C(_1013_),
    .X(_1254_));
 sky130_fd_sc_hd__a211o_1 _3908_ (.A1(\as1802.regs[3][14] ),
    .A2(_1138_),
    .B1(_1254_),
    .C1(_1085_),
    .X(_1255_));
 sky130_fd_sc_hd__o211a_1 _3909_ (.A1(_1082_),
    .A2(_1253_),
    .B1(_1255_),
    .C1(_1025_),
    .X(_1256_));
 sky130_fd_sc_hd__mux2_1 _3910_ (.A0(\as1802.regs[14][14] ),
    .A1(\as1802.regs[15][14] ),
    .S(_1138_),
    .X(_1257_));
 sky130_fd_sc_hd__mux2_1 _3911_ (.A0(\as1802.regs[12][14] ),
    .A1(\as1802.regs[13][14] ),
    .S(_1138_),
    .X(_1258_));
 sky130_fd_sc_hd__mux2_1 _3912_ (.A0(_1257_),
    .A1(_1258_),
    .S(_1085_),
    .X(_1259_));
 sky130_fd_sc_hd__mux2_1 _3913_ (.A0(\as1802.regs[8][14] ),
    .A1(\as1802.regs[9][14] ),
    .S(_1138_),
    .X(_1260_));
 sky130_fd_sc_hd__and3_1 _3914_ (.A(\as1802.regs[10][14] ),
    .B(_1012_),
    .C(_1013_),
    .X(_1261_));
 sky130_fd_sc_hd__a211o_1 _3915_ (.A1(\as1802.regs[11][14] ),
    .A2(_1138_),
    .B1(_1261_),
    .C1(_1085_),
    .X(_1262_));
 sky130_fd_sc_hd__o211a_1 _3916_ (.A1(_1082_),
    .A2(_1260_),
    .B1(_1262_),
    .C1(_1025_),
    .X(_1263_));
 sky130_fd_sc_hd__a211o_1 _3917_ (.A1(_0896_),
    .A2(_1259_),
    .B1(_1263_),
    .C1(_0708_),
    .X(_1264_));
 sky130_fd_sc_hd__o31ai_4 _3918_ (.A1(_0648_),
    .A2(_1252_),
    .A3(_1256_),
    .B1(_1264_),
    .Y(_1265_));
 sky130_fd_sc_hd__xnor2_1 _3919_ (.A(_1213_),
    .B(_1265_),
    .Y(_1266_));
 sky130_fd_sc_hd__nand4_2 _3920_ (.A(_0974_),
    .B(_1097_),
    .C(_1215_),
    .D(_1265_),
    .Y(_1267_));
 sky130_fd_sc_hd__a31o_1 _3921_ (.A1(_0974_),
    .A2(_1097_),
    .A3(_1215_),
    .B1(_1265_),
    .X(_1268_));
 sky130_fd_sc_hd__a21oi_1 _3922_ (.A1(_1267_),
    .A2(_1268_),
    .B1(_2606_),
    .Y(_1269_));
 sky130_fd_sc_hd__a211o_1 _3923_ (.A1(_0575_),
    .A2(_1266_),
    .B1(_1269_),
    .C1(_2596_),
    .X(_1270_));
 sky130_fd_sc_hd__or2_1 _3924_ (.A(_1174_),
    .B(_1233_),
    .X(_1271_));
 sky130_fd_sc_hd__mux4_1 _3925_ (.A0(\as1802.regs[0][14] ),
    .A1(\as1802.regs[1][14] ),
    .A2(\as1802.regs[2][14] ),
    .A3(\as1802.regs[3][14] ),
    .S0(_1225_),
    .S1(_1226_),
    .X(_1272_));
 sky130_fd_sc_hd__mux4_1 _3926_ (.A0(\as1802.regs[4][14] ),
    .A1(\as1802.regs[5][14] ),
    .A2(\as1802.regs[6][14] ),
    .A3(\as1802.regs[7][14] ),
    .S0(_1105_),
    .S1(_0981_),
    .X(_1273_));
 sky130_fd_sc_hd__mux2_1 _3927_ (.A0(_1272_),
    .A1(_1273_),
    .S(_0983_),
    .X(_1274_));
 sky130_fd_sc_hd__mux4_1 _3928_ (.A0(\as1802.regs[12][14] ),
    .A1(\as1802.regs[13][14] ),
    .A2(\as1802.regs[14][14] ),
    .A3(\as1802.regs[15][14] ),
    .S0(_1225_),
    .S1(_1226_),
    .X(_1275_));
 sky130_fd_sc_hd__and2b_1 _3929_ (.A_N(_1105_),
    .B(\as1802.regs[10][14] ),
    .X(_1276_));
 sky130_fd_sc_hd__a21bo_1 _3930_ (.A1(_1225_),
    .A2(\as1802.regs[11][14] ),
    .B1_N(_0981_),
    .X(_1277_));
 sky130_fd_sc_hd__mux2_1 _3931_ (.A0(\as1802.regs[8][14] ),
    .A1(\as1802.regs[9][14] ),
    .S(_1105_),
    .X(_1278_));
 sky130_fd_sc_hd__o221a_1 _3932_ (.A1(_1276_),
    .A2(_1277_),
    .B1(_1278_),
    .B2(_1226_),
    .C1(_0912_),
    .X(_1279_));
 sky130_fd_sc_hd__a211o_1 _3933_ (.A1(_0983_),
    .A2(_1275_),
    .B1(_1279_),
    .C1(_2667_),
    .X(_1280_));
 sky130_fd_sc_hd__o21ai_4 _3934_ (.A1(_2691_),
    .A2(_1274_),
    .B1(_1280_),
    .Y(_1281_));
 sky130_fd_sc_hd__xor2_1 _3935_ (.A(_1271_),
    .B(_1281_),
    .X(_1282_));
 sky130_fd_sc_hd__nor2_1 _3936_ (.A(_1237_),
    .B(_1281_),
    .Y(_1283_));
 sky130_fd_sc_hd__nand2_1 _3937_ (.A(_1237_),
    .B(_1281_),
    .Y(_1284_));
 sky130_fd_sc_hd__or3b_1 _3938_ (.A(_0922_),
    .B(_1283_),
    .C_N(_1284_),
    .X(_1285_));
 sky130_fd_sc_hd__o211a_1 _3939_ (.A1(_0976_),
    .A2(_1282_),
    .B1(_1285_),
    .C1(_0993_),
    .X(_1286_));
 sky130_fd_sc_hd__a211o_1 _3940_ (.A1(io_out[6]),
    .A2(_0536_),
    .B1(_0366_),
    .C1(_1286_),
    .X(_1287_));
 sky130_fd_sc_hd__clkbuf_4 _3941_ (.A(_0453_),
    .X(_1288_));
 sky130_fd_sc_hd__nor2_1 _3942_ (.A(_1288_),
    .B(_1281_),
    .Y(_1289_));
 sky130_fd_sc_hd__a211o_1 _3943_ (.A1(_1288_),
    .A2(_1282_),
    .B1(_1289_),
    .C1(_2701_),
    .X(_1290_));
 sky130_fd_sc_hd__a21oi_1 _3944_ (.A1(_1267_),
    .A2(_1268_),
    .B1(_0447_),
    .Y(_1291_));
 sky130_fd_sc_hd__a211o_1 _3945_ (.A1(_0447_),
    .A2(_1266_),
    .B1(_1291_),
    .C1(_0386_),
    .X(_1292_));
 sky130_fd_sc_hd__o21a_1 _3946_ (.A1(_0797_),
    .A2(_0935_),
    .B1(_0647_),
    .X(_1293_));
 sky130_fd_sc_hd__a32o_1 _3947_ (.A1(_0380_),
    .A2(_1287_),
    .A3(_1290_),
    .B1(_1292_),
    .B2(_1293_),
    .X(_1294_));
 sky130_fd_sc_hd__or2_1 _3948_ (.A(\as1802.regs[2][14] ),
    .B(_1191_),
    .X(_1295_));
 sky130_fd_sc_hd__nand2_1 _3949_ (.A(\as1802.regs[2][14] ),
    .B(_1191_),
    .Y(_1296_));
 sky130_fd_sc_hd__and3_1 _3950_ (.A(_2596_),
    .B(_1295_),
    .C(_1296_),
    .X(_1297_));
 sky130_fd_sc_hd__o21ba_2 _3951_ (.A1(_1270_),
    .A2(_1294_),
    .B1_N(_1297_),
    .X(_1298_));
 sky130_fd_sc_hd__buf_2 _3952_ (.A(_1298_),
    .X(_1299_));
 sky130_fd_sc_hd__mux2_1 _3953_ (.A0(\as1802.regs[10][14] ),
    .A1(_1299_),
    .S(_0947_),
    .X(_1300_));
 sky130_fd_sc_hd__clkbuf_1 _3954_ (.A(_1300_),
    .X(_0026_));
 sky130_fd_sc_hd__mux2_1 _3955_ (.A0(\as1802.regs[4][15] ),
    .A1(\as1802.regs[5][15] ),
    .S(_1074_),
    .X(_1301_));
 sky130_fd_sc_hd__mux2_1 _3956_ (.A0(\as1802.regs[6][15] ),
    .A1(\as1802.regs[7][15] ),
    .S(_0892_),
    .X(_1302_));
 sky130_fd_sc_hd__mux2_1 _3957_ (.A0(_1301_),
    .A1(_1302_),
    .S(_1082_),
    .X(_1303_));
 sky130_fd_sc_hd__mux2_1 _3958_ (.A0(\as1802.regs[0][15] ),
    .A1(\as1802.regs[1][15] ),
    .S(_1074_),
    .X(_1304_));
 sky130_fd_sc_hd__mux2_1 _3959_ (.A0(\as1802.regs[2][15] ),
    .A1(\as1802.regs[3][15] ),
    .S(_0892_),
    .X(_1305_));
 sky130_fd_sc_hd__mux2_1 _3960_ (.A0(_1304_),
    .A1(_1305_),
    .S(_1082_),
    .X(_1306_));
 sky130_fd_sc_hd__mux2_1 _3961_ (.A0(_1303_),
    .A1(_1306_),
    .S(_1025_),
    .X(_1307_));
 sky130_fd_sc_hd__mux2_1 _3962_ (.A0(\as1802.regs[8][15] ),
    .A1(\as1802.regs[9][15] ),
    .S(_1074_),
    .X(_1308_));
 sky130_fd_sc_hd__mux2_1 _3963_ (.A0(\as1802.regs[10][15] ),
    .A1(\as1802.regs[11][15] ),
    .S(_1074_),
    .X(_1309_));
 sky130_fd_sc_hd__mux2_1 _3964_ (.A0(_1308_),
    .A1(_1309_),
    .S(_1082_),
    .X(_1310_));
 sky130_fd_sc_hd__mux2_1 _3965_ (.A0(\as1802.regs[12][15] ),
    .A1(\as1802.regs[13][15] ),
    .S(_1074_),
    .X(_1311_));
 sky130_fd_sc_hd__mux2_1 _3966_ (.A0(\as1802.regs[14][15] ),
    .A1(\as1802.regs[15][15] ),
    .S(_0890_),
    .X(_1312_));
 sky130_fd_sc_hd__or2_1 _3967_ (.A(_1085_),
    .B(_1312_),
    .X(_1313_));
 sky130_fd_sc_hd__o211a_1 _3968_ (.A1(_1082_),
    .A2(_1311_),
    .B1(_1313_),
    .C1(_0896_),
    .X(_1314_));
 sky130_fd_sc_hd__a211o_1 _3969_ (.A1(_1025_),
    .A2(_1310_),
    .B1(_1314_),
    .C1(_0708_),
    .X(_1315_));
 sky130_fd_sc_hd__o21ai_4 _3970_ (.A1(_0648_),
    .A2(_1307_),
    .B1(_1315_),
    .Y(_1316_));
 sky130_fd_sc_hd__inv_2 _3971_ (.A(_1316_),
    .Y(_1317_));
 sky130_fd_sc_hd__o31ai_1 _3972_ (.A1(_1095_),
    .A2(_1212_),
    .A3(_1265_),
    .B1(_1317_),
    .Y(_1318_));
 sky130_fd_sc_hd__or4_1 _3973_ (.A(_1095_),
    .B(_1212_),
    .C(_1265_),
    .D(_1317_),
    .X(_1319_));
 sky130_fd_sc_hd__a21oi_1 _3974_ (.A1(_1318_),
    .A2(_1319_),
    .B1(_0455_),
    .Y(_1320_));
 sky130_fd_sc_hd__xnor2_1 _3975_ (.A(_1267_),
    .B(_1316_),
    .Y(_1321_));
 sky130_fd_sc_hd__o21ai_1 _3976_ (.A1(_0447_),
    .A2(_1321_),
    .B1(_0935_),
    .Y(_1322_));
 sky130_fd_sc_hd__o221ai_4 _3977_ (.A1(\as1802.D[7] ),
    .A2(_0935_),
    .B1(_1320_),
    .B2(_1322_),
    .C1(_0647_),
    .Y(_1323_));
 sky130_fd_sc_hd__and2b_1 _3978_ (.A_N(_1225_),
    .B(\as1802.regs[10][15] ),
    .X(_1324_));
 sky130_fd_sc_hd__a21bo_1 _3979_ (.A1(_1225_),
    .A2(\as1802.regs[11][15] ),
    .B1_N(_1226_),
    .X(_1325_));
 sky130_fd_sc_hd__mux2_1 _3980_ (.A0(\as1802.regs[8][15] ),
    .A1(\as1802.regs[9][15] ),
    .S(_1225_),
    .X(_1326_));
 sky130_fd_sc_hd__o221a_1 _3981_ (.A1(_1324_),
    .A2(_1325_),
    .B1(_1326_),
    .B2(_1226_),
    .C1(_0912_),
    .X(_1327_));
 sky130_fd_sc_hd__mux4_1 _3982_ (.A0(\as1802.regs[12][15] ),
    .A1(\as1802.regs[13][15] ),
    .A2(\as1802.regs[14][15] ),
    .A3(\as1802.regs[15][15] ),
    .S0(_1225_),
    .S1(_1226_),
    .X(_1328_));
 sky130_fd_sc_hd__a21o_1 _3983_ (.A1(_0983_),
    .A2(_1328_),
    .B1(_2667_),
    .X(_1329_));
 sky130_fd_sc_hd__mux4_1 _3984_ (.A0(\as1802.regs[4][15] ),
    .A1(\as1802.regs[5][15] ),
    .A2(\as1802.regs[6][15] ),
    .A3(\as1802.regs[7][15] ),
    .S0(_1225_),
    .S1(_1226_),
    .X(_1330_));
 sky130_fd_sc_hd__mux4_1 _3985_ (.A0(\as1802.regs[0][15] ),
    .A1(\as1802.regs[1][15] ),
    .A2(\as1802.regs[2][15] ),
    .A3(\as1802.regs[3][15] ),
    .S0(_1225_),
    .S1(_1226_),
    .X(_1331_));
 sky130_fd_sc_hd__mux2_1 _3986_ (.A0(_1330_),
    .A1(_1331_),
    .S(_0912_),
    .X(_1332_));
 sky130_fd_sc_hd__o22a_2 _3987_ (.A1(_1327_),
    .A2(_1329_),
    .B1(_1332_),
    .B2(_2691_),
    .X(_1333_));
 sky130_fd_sc_hd__inv_2 _3988_ (.A(_1333_),
    .Y(_1334_));
 sky130_fd_sc_hd__nor2_1 _3989_ (.A(_1233_),
    .B(_1281_),
    .Y(_1335_));
 sky130_fd_sc_hd__and4_1 _3990_ (.A(_1053_),
    .B(_1114_),
    .C(_1170_),
    .D(_1335_),
    .X(_1336_));
 sky130_fd_sc_hd__xnor2_1 _3991_ (.A(_1334_),
    .B(_1336_),
    .Y(_1337_));
 sky130_fd_sc_hd__mux2_1 _3992_ (.A0(_1333_),
    .A1(_1337_),
    .S(_2696_),
    .X(_1338_));
 sky130_fd_sc_hd__mux2_1 _3993_ (.A0(_1333_),
    .A1(_1338_),
    .S(_2556_),
    .X(_1339_));
 sky130_fd_sc_hd__a21oi_1 _3994_ (.A1(io_out[7]),
    .A2(_0536_),
    .B1(_0366_),
    .Y(_1340_));
 sky130_fd_sc_hd__mux2_1 _3995_ (.A0(_1333_),
    .A1(_1337_),
    .S(_2719_),
    .X(_1341_));
 sky130_fd_sc_hd__mux2_1 _3996_ (.A0(_1338_),
    .A1(_1341_),
    .S(_0976_),
    .X(_1342_));
 sky130_fd_sc_hd__nand2_1 _3997_ (.A(_0993_),
    .B(_1342_),
    .Y(_1343_));
 sky130_fd_sc_hd__a2bb2o_1 _3998_ (.A1_N(_2701_),
    .A2_N(_1339_),
    .B1(_1340_),
    .B2(_1343_),
    .X(_1344_));
 sky130_fd_sc_hd__a21o_1 _3999_ (.A1(_1318_),
    .A2(_1319_),
    .B1(_0390_),
    .X(_1345_));
 sky130_fd_sc_hd__a21o_1 _4000_ (.A1(_0390_),
    .A2(_1321_),
    .B1(_2606_),
    .X(_1346_));
 sky130_fd_sc_hd__o2111a_1 _4001_ (.A1(_0537_),
    .A2(_1344_),
    .B1(_1345_),
    .C1(_1346_),
    .D1(_0416_),
    .X(_1347_));
 sky130_fd_sc_hd__nand2_1 _4002_ (.A(\as1802.regs[2][15] ),
    .B(_1295_),
    .Y(_1348_));
 sky130_fd_sc_hd__or2_1 _4003_ (.A(\as1802.regs[2][15] ),
    .B(_1295_),
    .X(_1349_));
 sky130_fd_sc_hd__and3_1 _4004_ (.A(_2597_),
    .B(_1348_),
    .C(_1349_),
    .X(_1350_));
 sky130_fd_sc_hd__a21oi_4 _4005_ (.A1(_1323_),
    .A2(_1347_),
    .B1(_1350_),
    .Y(_1351_));
 sky130_fd_sc_hd__buf_2 _4006_ (.A(_1351_),
    .X(_1352_));
 sky130_fd_sc_hd__mux2_1 _4007_ (.A0(\as1802.regs[10][15] ),
    .A1(_1352_),
    .S(_0947_),
    .X(_1353_));
 sky130_fd_sc_hd__clkbuf_1 _4008_ (.A(_1353_),
    .X(_0027_));
 sky130_fd_sc_hd__clkbuf_2 _4009_ (.A(_0945_),
    .X(_1354_));
 sky130_fd_sc_hd__and2b_1 _4010_ (.A_N(_0401_),
    .B(_0399_),
    .X(_1355_));
 sky130_fd_sc_hd__o21a_1 _4011_ (.A1(\as1802.X[3] ),
    .A2(_2607_),
    .B1(_0404_),
    .X(_1356_));
 sky130_fd_sc_hd__nor2_2 _4012_ (.A(_1356_),
    .B(_0942_),
    .Y(_1357_));
 sky130_fd_sc_hd__and3_1 _4013_ (.A(_1354_),
    .B(_1355_),
    .C(_1357_),
    .X(_1358_));
 sky130_fd_sc_hd__buf_4 _4014_ (.A(_1358_),
    .X(_1359_));
 sky130_fd_sc_hd__mux2_1 _4015_ (.A0(\as1802.regs[0][8] ),
    .A1(_0940_),
    .S(_1359_),
    .X(_1360_));
 sky130_fd_sc_hd__clkbuf_1 _4016_ (.A(_1360_),
    .X(_0028_));
 sky130_fd_sc_hd__mux2_1 _4017_ (.A0(\as1802.regs[0][9] ),
    .A1(_1008_),
    .S(_1359_),
    .X(_1361_));
 sky130_fd_sc_hd__clkbuf_1 _4018_ (.A(_1361_),
    .X(_0029_));
 sky130_fd_sc_hd__mux2_1 _4019_ (.A0(\as1802.regs[0][10] ),
    .A1(_1069_),
    .S(_1359_),
    .X(_1362_));
 sky130_fd_sc_hd__clkbuf_1 _4020_ (.A(_1362_),
    .X(_0030_));
 sky130_fd_sc_hd__mux2_1 _4021_ (.A0(\as1802.regs[0][11] ),
    .A1(_1135_),
    .S(_1359_),
    .X(_1363_));
 sky130_fd_sc_hd__clkbuf_1 _4022_ (.A(_1363_),
    .X(_0031_));
 sky130_fd_sc_hd__mux2_1 _4023_ (.A0(\as1802.regs[0][12] ),
    .A1(_1189_),
    .S(_1359_),
    .X(_1364_));
 sky130_fd_sc_hd__clkbuf_1 _4024_ (.A(_1364_),
    .X(_0032_));
 sky130_fd_sc_hd__mux2_1 _4025_ (.A0(\as1802.regs[0][13] ),
    .A1(_1247_),
    .S(_1359_),
    .X(_1365_));
 sky130_fd_sc_hd__clkbuf_1 _4026_ (.A(_1365_),
    .X(_0033_));
 sky130_fd_sc_hd__mux2_1 _4027_ (.A0(\as1802.regs[0][14] ),
    .A1(_1299_),
    .S(_1359_),
    .X(_1366_));
 sky130_fd_sc_hd__clkbuf_1 _4028_ (.A(_1366_),
    .X(_0034_));
 sky130_fd_sc_hd__mux2_1 _4029_ (.A0(\as1802.regs[0][15] ),
    .A1(_1352_),
    .S(_1359_),
    .X(_1367_));
 sky130_fd_sc_hd__clkbuf_1 _4030_ (.A(_1367_),
    .X(_0035_));
 sky130_fd_sc_hd__and3_1 _4031_ (.A(_0943_),
    .B(_1354_),
    .C(_1355_),
    .X(_1368_));
 sky130_fd_sc_hd__buf_4 _4032_ (.A(_1368_),
    .X(_1369_));
 sky130_fd_sc_hd__mux2_1 _4033_ (.A0(\as1802.regs[8][8] ),
    .A1(_0940_),
    .S(_1369_),
    .X(_1370_));
 sky130_fd_sc_hd__clkbuf_1 _4034_ (.A(_1370_),
    .X(_0036_));
 sky130_fd_sc_hd__mux2_1 _4035_ (.A0(\as1802.regs[8][9] ),
    .A1(_1008_),
    .S(_1369_),
    .X(_1371_));
 sky130_fd_sc_hd__clkbuf_1 _4036_ (.A(_1371_),
    .X(_0037_));
 sky130_fd_sc_hd__mux2_1 _4037_ (.A0(\as1802.regs[8][10] ),
    .A1(_1069_),
    .S(_1369_),
    .X(_1372_));
 sky130_fd_sc_hd__clkbuf_1 _4038_ (.A(_1372_),
    .X(_0038_));
 sky130_fd_sc_hd__mux2_1 _4039_ (.A0(\as1802.regs[8][11] ),
    .A1(_1135_),
    .S(_1369_),
    .X(_1373_));
 sky130_fd_sc_hd__clkbuf_1 _4040_ (.A(_1373_),
    .X(_0039_));
 sky130_fd_sc_hd__mux2_1 _4041_ (.A0(\as1802.regs[8][12] ),
    .A1(_1189_),
    .S(_1369_),
    .X(_1374_));
 sky130_fd_sc_hd__clkbuf_1 _4042_ (.A(_1374_),
    .X(_0040_));
 sky130_fd_sc_hd__mux2_1 _4043_ (.A0(\as1802.regs[8][13] ),
    .A1(_1247_),
    .S(_1369_),
    .X(_1375_));
 sky130_fd_sc_hd__clkbuf_1 _4044_ (.A(_1375_),
    .X(_0041_));
 sky130_fd_sc_hd__mux2_1 _4045_ (.A0(\as1802.regs[8][14] ),
    .A1(_1299_),
    .S(_1369_),
    .X(_1376_));
 sky130_fd_sc_hd__clkbuf_1 _4046_ (.A(_1376_),
    .X(_0042_));
 sky130_fd_sc_hd__mux2_1 _4047_ (.A0(\as1802.regs[8][15] ),
    .A1(_1352_),
    .S(_1369_),
    .X(_1377_));
 sky130_fd_sc_hd__clkbuf_1 _4048_ (.A(_1377_),
    .X(_0043_));
 sky130_fd_sc_hd__nor2_2 _4049_ (.A(_1356_),
    .B(_0408_),
    .Y(_1378_));
 sky130_fd_sc_hd__and3_1 _4050_ (.A(_1354_),
    .B(_1355_),
    .C(_1378_),
    .X(_1379_));
 sky130_fd_sc_hd__buf_4 _4051_ (.A(_1379_),
    .X(_1380_));
 sky130_fd_sc_hd__mux2_1 _4052_ (.A0(\as1802.regs[4][8] ),
    .A1(_0940_),
    .S(_1380_),
    .X(_1381_));
 sky130_fd_sc_hd__clkbuf_1 _4053_ (.A(_1381_),
    .X(_0044_));
 sky130_fd_sc_hd__mux2_1 _4054_ (.A0(\as1802.regs[4][9] ),
    .A1(_1008_),
    .S(_1380_),
    .X(_1382_));
 sky130_fd_sc_hd__clkbuf_1 _4055_ (.A(_1382_),
    .X(_0045_));
 sky130_fd_sc_hd__mux2_1 _4056_ (.A0(\as1802.regs[4][10] ),
    .A1(_1069_),
    .S(_1380_),
    .X(_1383_));
 sky130_fd_sc_hd__clkbuf_1 _4057_ (.A(_1383_),
    .X(_0046_));
 sky130_fd_sc_hd__mux2_1 _4058_ (.A0(\as1802.regs[4][11] ),
    .A1(_1135_),
    .S(_1380_),
    .X(_1384_));
 sky130_fd_sc_hd__clkbuf_1 _4059_ (.A(_1384_),
    .X(_0047_));
 sky130_fd_sc_hd__mux2_1 _4060_ (.A0(\as1802.regs[4][12] ),
    .A1(_1189_),
    .S(_1380_),
    .X(_1385_));
 sky130_fd_sc_hd__clkbuf_1 _4061_ (.A(_1385_),
    .X(_0048_));
 sky130_fd_sc_hd__mux2_1 _4062_ (.A0(\as1802.regs[4][13] ),
    .A1(_1247_),
    .S(_1380_),
    .X(_1386_));
 sky130_fd_sc_hd__clkbuf_1 _4063_ (.A(_1386_),
    .X(_0049_));
 sky130_fd_sc_hd__mux2_1 _4064_ (.A0(\as1802.regs[4][14] ),
    .A1(_1299_),
    .S(_1380_),
    .X(_1387_));
 sky130_fd_sc_hd__clkbuf_1 _4065_ (.A(_1387_),
    .X(_0050_));
 sky130_fd_sc_hd__mux2_1 _4066_ (.A0(\as1802.regs[4][15] ),
    .A1(_1352_),
    .S(_1380_),
    .X(_1388_));
 sky130_fd_sc_hd__clkbuf_1 _4067_ (.A(_1388_),
    .X(_0051_));
 sky130_fd_sc_hd__and2_1 _4068_ (.A(_0399_),
    .B(_0401_),
    .X(_1389_));
 sky130_fd_sc_hd__and3_1 _4069_ (.A(_1354_),
    .B(_1378_),
    .C(_1389_),
    .X(_1390_));
 sky130_fd_sc_hd__buf_4 _4070_ (.A(_1390_),
    .X(_1391_));
 sky130_fd_sc_hd__mux2_1 _4071_ (.A0(\as1802.regs[5][8] ),
    .A1(_0940_),
    .S(_1391_),
    .X(_1392_));
 sky130_fd_sc_hd__clkbuf_1 _4072_ (.A(_1392_),
    .X(_0052_));
 sky130_fd_sc_hd__mux2_1 _4073_ (.A0(\as1802.regs[5][9] ),
    .A1(_1008_),
    .S(_1391_),
    .X(_1393_));
 sky130_fd_sc_hd__clkbuf_1 _4074_ (.A(_1393_),
    .X(_0053_));
 sky130_fd_sc_hd__mux2_1 _4075_ (.A0(\as1802.regs[5][10] ),
    .A1(_1069_),
    .S(_1391_),
    .X(_1394_));
 sky130_fd_sc_hd__clkbuf_1 _4076_ (.A(_1394_),
    .X(_0054_));
 sky130_fd_sc_hd__mux2_1 _4077_ (.A0(\as1802.regs[5][11] ),
    .A1(_1135_),
    .S(_1391_),
    .X(_1395_));
 sky130_fd_sc_hd__clkbuf_1 _4078_ (.A(_1395_),
    .X(_0055_));
 sky130_fd_sc_hd__mux2_1 _4079_ (.A0(\as1802.regs[5][12] ),
    .A1(_1189_),
    .S(_1391_),
    .X(_1396_));
 sky130_fd_sc_hd__clkbuf_1 _4080_ (.A(_1396_),
    .X(_0056_));
 sky130_fd_sc_hd__mux2_1 _4081_ (.A0(\as1802.regs[5][13] ),
    .A1(_1247_),
    .S(_1391_),
    .X(_1397_));
 sky130_fd_sc_hd__clkbuf_1 _4082_ (.A(_1397_),
    .X(_0057_));
 sky130_fd_sc_hd__mux2_1 _4083_ (.A0(\as1802.regs[5][14] ),
    .A1(_1299_),
    .S(_1391_),
    .X(_1398_));
 sky130_fd_sc_hd__clkbuf_1 _4084_ (.A(_1398_),
    .X(_0058_));
 sky130_fd_sc_hd__mux2_1 _4085_ (.A0(\as1802.regs[5][15] ),
    .A1(_1352_),
    .S(_1391_),
    .X(_1399_));
 sky130_fd_sc_hd__clkbuf_1 _4086_ (.A(_1399_),
    .X(_0059_));
 sky130_fd_sc_hd__and3_1 _4087_ (.A(_0402_),
    .B(_1354_),
    .C(_1378_),
    .X(_1400_));
 sky130_fd_sc_hd__buf_4 _4088_ (.A(_1400_),
    .X(_1401_));
 sky130_fd_sc_hd__mux2_1 _4089_ (.A0(\as1802.regs[7][8] ),
    .A1(_0940_),
    .S(_1401_),
    .X(_1402_));
 sky130_fd_sc_hd__clkbuf_1 _4090_ (.A(_1402_),
    .X(_0060_));
 sky130_fd_sc_hd__mux2_1 _4091_ (.A0(\as1802.regs[7][9] ),
    .A1(_1008_),
    .S(_1401_),
    .X(_1403_));
 sky130_fd_sc_hd__clkbuf_1 _4092_ (.A(_1403_),
    .X(_0061_));
 sky130_fd_sc_hd__mux2_1 _4093_ (.A0(\as1802.regs[7][10] ),
    .A1(_1069_),
    .S(_1401_),
    .X(_1404_));
 sky130_fd_sc_hd__clkbuf_1 _4094_ (.A(_1404_),
    .X(_0062_));
 sky130_fd_sc_hd__mux2_1 _4095_ (.A0(\as1802.regs[7][11] ),
    .A1(_1135_),
    .S(_1401_),
    .X(_1405_));
 sky130_fd_sc_hd__clkbuf_1 _4096_ (.A(_1405_),
    .X(_0063_));
 sky130_fd_sc_hd__mux2_1 _4097_ (.A0(\as1802.regs[7][12] ),
    .A1(_1189_),
    .S(_1401_),
    .X(_1406_));
 sky130_fd_sc_hd__clkbuf_1 _4098_ (.A(_1406_),
    .X(_0064_));
 sky130_fd_sc_hd__mux2_1 _4099_ (.A0(\as1802.regs[7][13] ),
    .A1(_1247_),
    .S(_1401_),
    .X(_1407_));
 sky130_fd_sc_hd__clkbuf_1 _4100_ (.A(_1407_),
    .X(_0065_));
 sky130_fd_sc_hd__mux2_1 _4101_ (.A0(\as1802.regs[7][14] ),
    .A1(_1299_),
    .S(_1401_),
    .X(_1408_));
 sky130_fd_sc_hd__clkbuf_1 _4102_ (.A(_1408_),
    .X(_0066_));
 sky130_fd_sc_hd__mux2_1 _4103_ (.A0(\as1802.regs[7][15] ),
    .A1(_1352_),
    .S(_1401_),
    .X(_1409_));
 sky130_fd_sc_hd__clkbuf_1 _4104_ (.A(_1409_),
    .X(_0067_));
 sky130_fd_sc_hd__and3_1 _4105_ (.A(_0941_),
    .B(_1354_),
    .C(_1378_),
    .X(_1410_));
 sky130_fd_sc_hd__buf_4 _4106_ (.A(_1410_),
    .X(_1411_));
 sky130_fd_sc_hd__mux2_1 _4107_ (.A0(\as1802.regs[6][8] ),
    .A1(_0940_),
    .S(_1411_),
    .X(_1412_));
 sky130_fd_sc_hd__clkbuf_1 _4108_ (.A(_1412_),
    .X(_0068_));
 sky130_fd_sc_hd__mux2_1 _4109_ (.A0(\as1802.regs[6][9] ),
    .A1(_1008_),
    .S(_1411_),
    .X(_1413_));
 sky130_fd_sc_hd__clkbuf_1 _4110_ (.A(_1413_),
    .X(_0069_));
 sky130_fd_sc_hd__mux2_1 _4111_ (.A0(\as1802.regs[6][10] ),
    .A1(_1069_),
    .S(_1411_),
    .X(_1414_));
 sky130_fd_sc_hd__clkbuf_1 _4112_ (.A(_1414_),
    .X(_0070_));
 sky130_fd_sc_hd__mux2_1 _4113_ (.A0(\as1802.regs[6][11] ),
    .A1(_1135_),
    .S(_1411_),
    .X(_1415_));
 sky130_fd_sc_hd__clkbuf_1 _4114_ (.A(_1415_),
    .X(_0071_));
 sky130_fd_sc_hd__mux2_1 _4115_ (.A0(\as1802.regs[6][12] ),
    .A1(_1189_),
    .S(_1411_),
    .X(_1416_));
 sky130_fd_sc_hd__clkbuf_1 _4116_ (.A(_1416_),
    .X(_0072_));
 sky130_fd_sc_hd__mux2_1 _4117_ (.A0(\as1802.regs[6][13] ),
    .A1(_1247_),
    .S(_1411_),
    .X(_1417_));
 sky130_fd_sc_hd__clkbuf_1 _4118_ (.A(_1417_),
    .X(_0073_));
 sky130_fd_sc_hd__mux2_1 _4119_ (.A0(\as1802.regs[6][14] ),
    .A1(_1299_),
    .S(_1411_),
    .X(_1418_));
 sky130_fd_sc_hd__clkbuf_1 _4120_ (.A(_1418_),
    .X(_0074_));
 sky130_fd_sc_hd__mux2_1 _4121_ (.A0(\as1802.regs[6][15] ),
    .A1(_1352_),
    .S(_1411_),
    .X(_1419_));
 sky130_fd_sc_hd__clkbuf_1 _4122_ (.A(_1419_),
    .X(_0075_));
 sky130_fd_sc_hd__and3_1 _4123_ (.A(_0402_),
    .B(_1354_),
    .C(_1357_),
    .X(_1420_));
 sky130_fd_sc_hd__buf_4 _4124_ (.A(_1420_),
    .X(_1421_));
 sky130_fd_sc_hd__mux2_1 _4125_ (.A0(\as1802.regs[3][8] ),
    .A1(_0940_),
    .S(_1421_),
    .X(_1422_));
 sky130_fd_sc_hd__clkbuf_1 _4126_ (.A(_1422_),
    .X(_0076_));
 sky130_fd_sc_hd__mux2_1 _4127_ (.A0(\as1802.regs[3][9] ),
    .A1(_1008_),
    .S(_1421_),
    .X(_1423_));
 sky130_fd_sc_hd__clkbuf_1 _4128_ (.A(_1423_),
    .X(_0077_));
 sky130_fd_sc_hd__mux2_1 _4129_ (.A0(\as1802.regs[3][10] ),
    .A1(_1069_),
    .S(_1421_),
    .X(_1424_));
 sky130_fd_sc_hd__clkbuf_1 _4130_ (.A(_1424_),
    .X(_0078_));
 sky130_fd_sc_hd__mux2_1 _4131_ (.A0(\as1802.regs[3][11] ),
    .A1(_1135_),
    .S(_1421_),
    .X(_1425_));
 sky130_fd_sc_hd__clkbuf_1 _4132_ (.A(_1425_),
    .X(_0079_));
 sky130_fd_sc_hd__mux2_1 _4133_ (.A0(\as1802.regs[3][12] ),
    .A1(_1189_),
    .S(_1421_),
    .X(_1426_));
 sky130_fd_sc_hd__clkbuf_1 _4134_ (.A(_1426_),
    .X(_0080_));
 sky130_fd_sc_hd__mux2_1 _4135_ (.A0(\as1802.regs[3][13] ),
    .A1(_1247_),
    .S(_1421_),
    .X(_1427_));
 sky130_fd_sc_hd__clkbuf_1 _4136_ (.A(_1427_),
    .X(_0081_));
 sky130_fd_sc_hd__mux2_1 _4137_ (.A0(\as1802.regs[3][14] ),
    .A1(_1299_),
    .S(_1421_),
    .X(_1428_));
 sky130_fd_sc_hd__clkbuf_1 _4138_ (.A(_1428_),
    .X(_0082_));
 sky130_fd_sc_hd__mux2_1 _4139_ (.A0(\as1802.regs[3][15] ),
    .A1(_1352_),
    .S(_1421_),
    .X(_1429_));
 sky130_fd_sc_hd__clkbuf_1 _4140_ (.A(_1429_),
    .X(_0083_));
 sky130_fd_sc_hd__clkbuf_2 _4141_ (.A(_0411_),
    .X(_1430_));
 sky130_fd_sc_hd__and3_1 _4142_ (.A(_1430_),
    .B(_0943_),
    .C(_1389_),
    .X(_1431_));
 sky130_fd_sc_hd__buf_4 _4143_ (.A(_1431_),
    .X(_1432_));
 sky130_fd_sc_hd__mux2_1 _4144_ (.A0(\as1802.regs[9][0] ),
    .A1(_0395_),
    .S(_1432_),
    .X(_1433_));
 sky130_fd_sc_hd__clkbuf_1 _4145_ (.A(_1433_),
    .X(_0084_));
 sky130_fd_sc_hd__mux2_1 _4146_ (.A0(\as1802.regs[9][1] ),
    .A1(_0487_),
    .S(_1432_),
    .X(_1434_));
 sky130_fd_sc_hd__clkbuf_1 _4147_ (.A(_1434_),
    .X(_0085_));
 sky130_fd_sc_hd__mux2_1 _4148_ (.A0(\as1802.regs[9][2] ),
    .A1(_0549_),
    .S(_1432_),
    .X(_1435_));
 sky130_fd_sc_hd__clkbuf_1 _4149_ (.A(_1435_),
    .X(_0086_));
 sky130_fd_sc_hd__mux2_1 _4150_ (.A0(\as1802.regs[9][3] ),
    .A1(_0613_),
    .S(_1432_),
    .X(_1436_));
 sky130_fd_sc_hd__clkbuf_1 _4151_ (.A(_1436_),
    .X(_0087_));
 sky130_fd_sc_hd__mux2_1 _4152_ (.A0(\as1802.regs[9][4] ),
    .A1(_0683_),
    .S(_1432_),
    .X(_1437_));
 sky130_fd_sc_hd__clkbuf_1 _4153_ (.A(_1437_),
    .X(_0088_));
 sky130_fd_sc_hd__mux2_1 _4154_ (.A0(\as1802.regs[9][5] ),
    .A1(_0750_),
    .S(_1432_),
    .X(_1438_));
 sky130_fd_sc_hd__clkbuf_1 _4155_ (.A(_1438_),
    .X(_0089_));
 sky130_fd_sc_hd__mux2_1 _4156_ (.A0(\as1802.regs[9][6] ),
    .A1(_0806_),
    .S(_1432_),
    .X(_1439_));
 sky130_fd_sc_hd__clkbuf_1 _4157_ (.A(_1439_),
    .X(_0090_));
 sky130_fd_sc_hd__mux2_1 _4158_ (.A0(\as1802.regs[9][7] ),
    .A1(_0871_),
    .S(_1432_),
    .X(_1440_));
 sky130_fd_sc_hd__clkbuf_1 _4159_ (.A(_1440_),
    .X(_0091_));
 sky130_fd_sc_hd__and3_1 _4160_ (.A(_1430_),
    .B(_0943_),
    .C(_1355_),
    .X(_1441_));
 sky130_fd_sc_hd__buf_4 _4161_ (.A(_1441_),
    .X(_1442_));
 sky130_fd_sc_hd__mux2_1 _4162_ (.A0(\as1802.regs[8][0] ),
    .A1(_0395_),
    .S(_1442_),
    .X(_1443_));
 sky130_fd_sc_hd__clkbuf_1 _4163_ (.A(_1443_),
    .X(_0092_));
 sky130_fd_sc_hd__mux2_1 _4164_ (.A0(\as1802.regs[8][1] ),
    .A1(_0487_),
    .S(_1442_),
    .X(_1444_));
 sky130_fd_sc_hd__clkbuf_1 _4165_ (.A(_1444_),
    .X(_0093_));
 sky130_fd_sc_hd__mux2_1 _4166_ (.A0(\as1802.regs[8][2] ),
    .A1(_0549_),
    .S(_1442_),
    .X(_1445_));
 sky130_fd_sc_hd__clkbuf_1 _4167_ (.A(_1445_),
    .X(_0094_));
 sky130_fd_sc_hd__mux2_1 _4168_ (.A0(\as1802.regs[8][3] ),
    .A1(_0613_),
    .S(_1442_),
    .X(_1446_));
 sky130_fd_sc_hd__clkbuf_1 _4169_ (.A(_1446_),
    .X(_0095_));
 sky130_fd_sc_hd__mux2_1 _4170_ (.A0(\as1802.regs[8][4] ),
    .A1(_0683_),
    .S(_1442_),
    .X(_1447_));
 sky130_fd_sc_hd__clkbuf_1 _4171_ (.A(_1447_),
    .X(_0096_));
 sky130_fd_sc_hd__mux2_1 _4172_ (.A0(\as1802.regs[8][5] ),
    .A1(_0750_),
    .S(_1442_),
    .X(_1448_));
 sky130_fd_sc_hd__clkbuf_1 _4173_ (.A(_1448_),
    .X(_0097_));
 sky130_fd_sc_hd__mux2_1 _4174_ (.A0(\as1802.regs[8][6] ),
    .A1(_0806_),
    .S(_1442_),
    .X(_1449_));
 sky130_fd_sc_hd__clkbuf_1 _4175_ (.A(_1449_),
    .X(_0098_));
 sky130_fd_sc_hd__mux2_1 _4176_ (.A0(\as1802.regs[8][7] ),
    .A1(_0871_),
    .S(_1442_),
    .X(_1450_));
 sky130_fd_sc_hd__clkbuf_1 _4177_ (.A(_1450_),
    .X(_0099_));
 sky130_fd_sc_hd__and3_1 _4178_ (.A(_0402_),
    .B(_1430_),
    .C(_1378_),
    .X(_1451_));
 sky130_fd_sc_hd__buf_4 _4179_ (.A(_1451_),
    .X(_1452_));
 sky130_fd_sc_hd__mux2_1 _4180_ (.A0(\as1802.regs[7][0] ),
    .A1(_0395_),
    .S(_1452_),
    .X(_1453_));
 sky130_fd_sc_hd__clkbuf_1 _4181_ (.A(_1453_),
    .X(_0100_));
 sky130_fd_sc_hd__mux2_1 _4182_ (.A0(\as1802.regs[7][1] ),
    .A1(_0487_),
    .S(_1452_),
    .X(_1454_));
 sky130_fd_sc_hd__clkbuf_1 _4183_ (.A(_1454_),
    .X(_0101_));
 sky130_fd_sc_hd__mux2_1 _4184_ (.A0(\as1802.regs[7][2] ),
    .A1(_0549_),
    .S(_1452_),
    .X(_1455_));
 sky130_fd_sc_hd__clkbuf_1 _4185_ (.A(_1455_),
    .X(_0102_));
 sky130_fd_sc_hd__mux2_1 _4186_ (.A0(\as1802.regs[7][3] ),
    .A1(_0613_),
    .S(_1452_),
    .X(_1456_));
 sky130_fd_sc_hd__clkbuf_1 _4187_ (.A(_1456_),
    .X(_0103_));
 sky130_fd_sc_hd__mux2_1 _4188_ (.A0(\as1802.regs[7][4] ),
    .A1(_0683_),
    .S(_1452_),
    .X(_1457_));
 sky130_fd_sc_hd__clkbuf_1 _4189_ (.A(_1457_),
    .X(_0104_));
 sky130_fd_sc_hd__mux2_1 _4190_ (.A0(\as1802.regs[7][5] ),
    .A1(_0750_),
    .S(_1452_),
    .X(_1458_));
 sky130_fd_sc_hd__clkbuf_1 _4191_ (.A(_1458_),
    .X(_0105_));
 sky130_fd_sc_hd__mux2_1 _4192_ (.A0(\as1802.regs[7][6] ),
    .A1(_0806_),
    .S(_1452_),
    .X(_1459_));
 sky130_fd_sc_hd__clkbuf_1 _4193_ (.A(_1459_),
    .X(_0106_));
 sky130_fd_sc_hd__mux2_1 _4194_ (.A0(\as1802.regs[7][7] ),
    .A1(_0871_),
    .S(_1452_),
    .X(_1460_));
 sky130_fd_sc_hd__clkbuf_1 _4195_ (.A(_1460_),
    .X(_0107_));
 sky130_fd_sc_hd__and3_1 _4196_ (.A(_1430_),
    .B(_0941_),
    .C(_1378_),
    .X(_1461_));
 sky130_fd_sc_hd__buf_4 _4197_ (.A(_1461_),
    .X(_1462_));
 sky130_fd_sc_hd__mux2_1 _4198_ (.A0(\as1802.regs[6][0] ),
    .A1(_0395_),
    .S(_1462_),
    .X(_1463_));
 sky130_fd_sc_hd__clkbuf_1 _4199_ (.A(_1463_),
    .X(_0108_));
 sky130_fd_sc_hd__mux2_1 _4200_ (.A0(\as1802.regs[6][1] ),
    .A1(_0487_),
    .S(_1462_),
    .X(_1464_));
 sky130_fd_sc_hd__clkbuf_1 _4201_ (.A(_1464_),
    .X(_0109_));
 sky130_fd_sc_hd__mux2_1 _4202_ (.A0(\as1802.regs[6][2] ),
    .A1(_0549_),
    .S(_1462_),
    .X(_1465_));
 sky130_fd_sc_hd__clkbuf_1 _4203_ (.A(_1465_),
    .X(_0110_));
 sky130_fd_sc_hd__mux2_1 _4204_ (.A0(\as1802.regs[6][3] ),
    .A1(_0613_),
    .S(_1462_),
    .X(_1466_));
 sky130_fd_sc_hd__clkbuf_1 _4205_ (.A(_1466_),
    .X(_0111_));
 sky130_fd_sc_hd__mux2_1 _4206_ (.A0(\as1802.regs[6][4] ),
    .A1(_0683_),
    .S(_1462_),
    .X(_1467_));
 sky130_fd_sc_hd__clkbuf_1 _4207_ (.A(_1467_),
    .X(_0112_));
 sky130_fd_sc_hd__mux2_1 _4208_ (.A0(\as1802.regs[6][5] ),
    .A1(_0750_),
    .S(_1462_),
    .X(_1468_));
 sky130_fd_sc_hd__clkbuf_1 _4209_ (.A(_1468_),
    .X(_0113_));
 sky130_fd_sc_hd__mux2_1 _4210_ (.A0(\as1802.regs[6][6] ),
    .A1(_0806_),
    .S(_1462_),
    .X(_1469_));
 sky130_fd_sc_hd__clkbuf_1 _4211_ (.A(_1469_),
    .X(_0114_));
 sky130_fd_sc_hd__mux2_1 _4212_ (.A0(\as1802.regs[6][7] ),
    .A1(_0871_),
    .S(_1462_),
    .X(_1470_));
 sky130_fd_sc_hd__clkbuf_1 _4213_ (.A(_1470_),
    .X(_0115_));
 sky130_fd_sc_hd__o31a_1 _4214_ (.A1(_2580_),
    .A2(_2476_),
    .A3(_2463_),
    .B1(_2547_),
    .X(_1471_));
 sky130_fd_sc_hd__or2_1 _4215_ (.A(_2529_),
    .B(_2715_),
    .X(_1472_));
 sky130_fd_sc_hd__nand2_1 _4216_ (.A(_1471_),
    .B(_1472_),
    .Y(_1473_));
 sky130_fd_sc_hd__nor2_1 _4217_ (.A(_2476_),
    .B(_2475_),
    .Y(_1474_));
 sky130_fd_sc_hd__nand2_2 _4218_ (.A(_2486_),
    .B(_2522_),
    .Y(_1475_));
 sky130_fd_sc_hd__nand2_2 _4219_ (.A(\as1802.will_interrupt ),
    .B(_2580_),
    .Y(_1476_));
 sky130_fd_sc_hd__o21a_1 _4220_ (.A1(_1474_),
    .A2(_1475_),
    .B1(_1476_),
    .X(_1477_));
 sky130_fd_sc_hd__nor2_1 _4221_ (.A(_1473_),
    .B(_1477_),
    .Y(_1478_));
 sky130_fd_sc_hd__or2_1 _4222_ (.A(\as1802.IE ),
    .B(_1476_),
    .X(_1479_));
 sky130_fd_sc_hd__o2111a_1 _4223_ (.A1(_2581_),
    .A2(_2561_),
    .B1(_2705_),
    .C1(_1478_),
    .D1(_1479_),
    .X(_1480_));
 sky130_fd_sc_hd__nor2_1 _4224_ (.A(_2579_),
    .B(_2553_),
    .Y(_1481_));
 sky130_fd_sc_hd__nand2_2 _4225_ (.A(_2570_),
    .B(_1481_),
    .Y(_1482_));
 sky130_fd_sc_hd__a31o_1 _4226_ (.A1(_2527_),
    .A2(_2503_),
    .A3(_2494_),
    .B1(_1482_),
    .X(_1483_));
 sky130_fd_sc_hd__o211a_1 _4227_ (.A1(_2473_),
    .A2(_2478_),
    .B1(_2585_),
    .C1(_2486_),
    .X(_1484_));
 sky130_fd_sc_hd__a21o_1 _4228_ (.A1(_2473_),
    .A2(_2474_),
    .B1(_2477_),
    .X(_1485_));
 sky130_fd_sc_hd__nand3_1 _4229_ (.A(_2476_),
    .B(_1484_),
    .C(_1485_),
    .Y(_1486_));
 sky130_fd_sc_hd__and3_1 _4230_ (.A(_1480_),
    .B(_1483_),
    .C(_1486_),
    .X(_1487_));
 sky130_fd_sc_hd__buf_2 _4231_ (.A(_1487_),
    .X(_1488_));
 sky130_fd_sc_hd__clkbuf_4 _4232_ (.A(_2581_),
    .X(_1489_));
 sky130_fd_sc_hd__clkbuf_4 _4233_ (.A(_2526_),
    .X(_1490_));
 sky130_fd_sc_hd__buf_4 _4234_ (.A(_1490_),
    .X(_1491_));
 sky130_fd_sc_hd__mux2_1 _4235_ (.A0(_2469_),
    .A1(_2702_),
    .S(_1491_),
    .X(_1492_));
 sky130_fd_sc_hd__or3b_1 _4236_ (.A(_1489_),
    .B(_1492_),
    .C_N(_1488_),
    .X(_1493_));
 sky130_fd_sc_hd__clkbuf_4 _4237_ (.A(_2457_),
    .X(_1494_));
 sky130_fd_sc_hd__o211a_1 _4238_ (.A1(\as1802.P[0] ),
    .A2(_1488_),
    .B1(_1493_),
    .C1(_1494_),
    .X(_0116_));
 sky130_fd_sc_hd__buf_2 _4239_ (.A(_2554_),
    .X(_1495_));
 sky130_fd_sc_hd__buf_4 _4240_ (.A(_1495_),
    .X(_1496_));
 sky130_fd_sc_hd__nand2_1 _4241_ (.A(_2504_),
    .B(_1496_),
    .Y(_1497_));
 sky130_fd_sc_hd__o2bb2a_1 _4242_ (.A1_N(_0474_),
    .A2_N(_1481_),
    .B1(_1497_),
    .B2(_1489_),
    .X(_1498_));
 sky130_fd_sc_hd__clkbuf_4 _4243_ (.A(_2456_),
    .X(_1499_));
 sky130_fd_sc_hd__a21oi_1 _4244_ (.A1(_1488_),
    .A2(_1498_),
    .B1(_1499_),
    .Y(_1500_));
 sky130_fd_sc_hd__o21a_1 _4245_ (.A1(\as1802.P[1] ),
    .A2(_1488_),
    .B1(_1500_),
    .X(_0117_));
 sky130_fd_sc_hd__nor2_1 _4246_ (.A(io_out[2]),
    .B(_1496_),
    .Y(_1501_));
 sky130_fd_sc_hd__nor2_1 _4247_ (.A(_2496_),
    .B(_1491_),
    .Y(_1502_));
 sky130_fd_sc_hd__o31ai_1 _4248_ (.A1(_1489_),
    .A2(_1501_),
    .A3(_1502_),
    .B1(_1488_),
    .Y(_1503_));
 sky130_fd_sc_hd__o211a_1 _4249_ (.A1(\as1802.P[2] ),
    .A2(_1488_),
    .B1(_1503_),
    .C1(_1494_),
    .X(_0118_));
 sky130_fd_sc_hd__buf_2 _4250_ (.A(_2457_),
    .X(_1504_));
 sky130_fd_sc_hd__a21oi_1 _4251_ (.A1(_2494_),
    .A2(_2554_),
    .B1(_2581_),
    .Y(_1505_));
 sky130_fd_sc_hd__o21a_1 _4252_ (.A1(io_out[3]),
    .A2(_1495_),
    .B1(_1505_),
    .X(_1506_));
 sky130_fd_sc_hd__mux2_1 _4253_ (.A0(\as1802.P[3] ),
    .A1(_1506_),
    .S(_1488_),
    .X(_1507_));
 sky130_fd_sc_hd__and2_1 _4254_ (.A(_1504_),
    .B(_1507_),
    .X(_1508_));
 sky130_fd_sc_hd__clkbuf_1 _4255_ (.A(_1508_),
    .X(_0119_));
 sky130_fd_sc_hd__and3_1 _4256_ (.A(_1430_),
    .B(_1378_),
    .C(_1389_),
    .X(_1509_));
 sky130_fd_sc_hd__buf_4 _4257_ (.A(_1509_),
    .X(_1510_));
 sky130_fd_sc_hd__mux2_1 _4258_ (.A0(\as1802.regs[5][0] ),
    .A1(_0395_),
    .S(_1510_),
    .X(_1511_));
 sky130_fd_sc_hd__clkbuf_1 _4259_ (.A(_1511_),
    .X(_0120_));
 sky130_fd_sc_hd__mux2_1 _4260_ (.A0(\as1802.regs[5][1] ),
    .A1(_0487_),
    .S(_1510_),
    .X(_1512_));
 sky130_fd_sc_hd__clkbuf_1 _4261_ (.A(_1512_),
    .X(_0121_));
 sky130_fd_sc_hd__mux2_1 _4262_ (.A0(\as1802.regs[5][2] ),
    .A1(_0549_),
    .S(_1510_),
    .X(_1513_));
 sky130_fd_sc_hd__clkbuf_1 _4263_ (.A(_1513_),
    .X(_0122_));
 sky130_fd_sc_hd__mux2_1 _4264_ (.A0(\as1802.regs[5][3] ),
    .A1(_0613_),
    .S(_1510_),
    .X(_1514_));
 sky130_fd_sc_hd__clkbuf_1 _4265_ (.A(_1514_),
    .X(_0123_));
 sky130_fd_sc_hd__mux2_1 _4266_ (.A0(\as1802.regs[5][4] ),
    .A1(_0683_),
    .S(_1510_),
    .X(_1515_));
 sky130_fd_sc_hd__clkbuf_1 _4267_ (.A(_1515_),
    .X(_0124_));
 sky130_fd_sc_hd__mux2_1 _4268_ (.A0(\as1802.regs[5][5] ),
    .A1(_0750_),
    .S(_1510_),
    .X(_1516_));
 sky130_fd_sc_hd__clkbuf_1 _4269_ (.A(_1516_),
    .X(_0125_));
 sky130_fd_sc_hd__mux2_1 _4270_ (.A0(\as1802.regs[5][6] ),
    .A1(_0806_),
    .S(_1510_),
    .X(_1517_));
 sky130_fd_sc_hd__clkbuf_1 _4271_ (.A(_1517_),
    .X(_0126_));
 sky130_fd_sc_hd__mux2_1 _4272_ (.A0(\as1802.regs[5][7] ),
    .A1(_0871_),
    .S(_1510_),
    .X(_1518_));
 sky130_fd_sc_hd__clkbuf_1 _4273_ (.A(_1518_),
    .X(_0127_));
 sky130_fd_sc_hd__and3_1 _4274_ (.A(_1430_),
    .B(_1355_),
    .C(_1378_),
    .X(_1519_));
 sky130_fd_sc_hd__buf_4 _4275_ (.A(_1519_),
    .X(_1520_));
 sky130_fd_sc_hd__mux2_1 _4276_ (.A0(\as1802.regs[4][0] ),
    .A1(_0395_),
    .S(_1520_),
    .X(_1521_));
 sky130_fd_sc_hd__clkbuf_1 _4277_ (.A(_1521_),
    .X(_0128_));
 sky130_fd_sc_hd__mux2_1 _4278_ (.A0(\as1802.regs[4][1] ),
    .A1(_0487_),
    .S(_1520_),
    .X(_1522_));
 sky130_fd_sc_hd__clkbuf_1 _4279_ (.A(_1522_),
    .X(_0129_));
 sky130_fd_sc_hd__mux2_1 _4280_ (.A0(\as1802.regs[4][2] ),
    .A1(_0549_),
    .S(_1520_),
    .X(_1523_));
 sky130_fd_sc_hd__clkbuf_1 _4281_ (.A(_1523_),
    .X(_0130_));
 sky130_fd_sc_hd__mux2_1 _4282_ (.A0(\as1802.regs[4][3] ),
    .A1(_0613_),
    .S(_1520_),
    .X(_1524_));
 sky130_fd_sc_hd__clkbuf_1 _4283_ (.A(_1524_),
    .X(_0131_));
 sky130_fd_sc_hd__mux2_1 _4284_ (.A0(\as1802.regs[4][4] ),
    .A1(_0683_),
    .S(_1520_),
    .X(_1525_));
 sky130_fd_sc_hd__clkbuf_1 _4285_ (.A(_1525_),
    .X(_0132_));
 sky130_fd_sc_hd__mux2_1 _4286_ (.A0(\as1802.regs[4][5] ),
    .A1(_0750_),
    .S(_1520_),
    .X(_1526_));
 sky130_fd_sc_hd__clkbuf_1 _4287_ (.A(_1526_),
    .X(_0133_));
 sky130_fd_sc_hd__mux2_1 _4288_ (.A0(\as1802.regs[4][6] ),
    .A1(_0806_),
    .S(_1520_),
    .X(_1527_));
 sky130_fd_sc_hd__clkbuf_1 _4289_ (.A(_1527_),
    .X(_0134_));
 sky130_fd_sc_hd__mux2_1 _4290_ (.A0(\as1802.regs[4][7] ),
    .A1(_0871_),
    .S(_1520_),
    .X(_1528_));
 sky130_fd_sc_hd__clkbuf_1 _4291_ (.A(_1528_),
    .X(_0135_));
 sky130_fd_sc_hd__and3_1 _4292_ (.A(_0402_),
    .B(_0411_),
    .C(_1357_),
    .X(_1529_));
 sky130_fd_sc_hd__buf_4 _4293_ (.A(_1529_),
    .X(_1530_));
 sky130_fd_sc_hd__mux2_1 _4294_ (.A0(\as1802.regs[3][0] ),
    .A1(_0395_),
    .S(_1530_),
    .X(_1531_));
 sky130_fd_sc_hd__clkbuf_1 _4295_ (.A(_1531_),
    .X(_0136_));
 sky130_fd_sc_hd__mux2_1 _4296_ (.A0(\as1802.regs[3][1] ),
    .A1(_0487_),
    .S(_1530_),
    .X(_1532_));
 sky130_fd_sc_hd__clkbuf_1 _4297_ (.A(_1532_),
    .X(_0137_));
 sky130_fd_sc_hd__mux2_1 _4298_ (.A0(\as1802.regs[3][2] ),
    .A1(_0549_),
    .S(_1530_),
    .X(_1533_));
 sky130_fd_sc_hd__clkbuf_1 _4299_ (.A(_1533_),
    .X(_0138_));
 sky130_fd_sc_hd__mux2_1 _4300_ (.A0(\as1802.regs[3][3] ),
    .A1(_0613_),
    .S(_1530_),
    .X(_1534_));
 sky130_fd_sc_hd__clkbuf_1 _4301_ (.A(_1534_),
    .X(_0139_));
 sky130_fd_sc_hd__mux2_1 _4302_ (.A0(\as1802.regs[3][4] ),
    .A1(_0683_),
    .S(_1530_),
    .X(_1535_));
 sky130_fd_sc_hd__clkbuf_1 _4303_ (.A(_1535_),
    .X(_0140_));
 sky130_fd_sc_hd__mux2_1 _4304_ (.A0(\as1802.regs[3][5] ),
    .A1(_0750_),
    .S(_1530_),
    .X(_1536_));
 sky130_fd_sc_hd__clkbuf_1 _4305_ (.A(_1536_),
    .X(_0141_));
 sky130_fd_sc_hd__mux2_1 _4306_ (.A0(\as1802.regs[3][6] ),
    .A1(_0806_),
    .S(_1530_),
    .X(_1537_));
 sky130_fd_sc_hd__clkbuf_1 _4307_ (.A(_1537_),
    .X(_0142_));
 sky130_fd_sc_hd__mux2_1 _4308_ (.A0(\as1802.regs[3][7] ),
    .A1(_0871_),
    .S(_1530_),
    .X(_1538_));
 sky130_fd_sc_hd__clkbuf_1 _4309_ (.A(_1538_),
    .X(_0143_));
 sky130_fd_sc_hd__and3_1 _4310_ (.A(_1430_),
    .B(_0941_),
    .C(_1357_),
    .X(_1539_));
 sky130_fd_sc_hd__buf_4 _4311_ (.A(_1539_),
    .X(_1540_));
 sky130_fd_sc_hd__mux2_1 _4312_ (.A0(\as1802.regs[2][0] ),
    .A1(_0395_),
    .S(_1540_),
    .X(_1541_));
 sky130_fd_sc_hd__clkbuf_1 _4313_ (.A(_1541_),
    .X(_0144_));
 sky130_fd_sc_hd__mux2_1 _4314_ (.A0(\as1802.regs[2][1] ),
    .A1(_0487_),
    .S(_1540_),
    .X(_1542_));
 sky130_fd_sc_hd__clkbuf_1 _4315_ (.A(_1542_),
    .X(_0145_));
 sky130_fd_sc_hd__mux2_1 _4316_ (.A0(\as1802.regs[2][2] ),
    .A1(_0549_),
    .S(_1540_),
    .X(_1543_));
 sky130_fd_sc_hd__clkbuf_1 _4317_ (.A(_1543_),
    .X(_0146_));
 sky130_fd_sc_hd__mux2_1 _4318_ (.A0(\as1802.regs[2][3] ),
    .A1(_0613_),
    .S(_1540_),
    .X(_1544_));
 sky130_fd_sc_hd__clkbuf_1 _4319_ (.A(_1544_),
    .X(_0147_));
 sky130_fd_sc_hd__mux2_1 _4320_ (.A0(\as1802.regs[2][4] ),
    .A1(_0683_),
    .S(_1540_),
    .X(_1545_));
 sky130_fd_sc_hd__clkbuf_1 _4321_ (.A(_1545_),
    .X(_0148_));
 sky130_fd_sc_hd__mux2_1 _4322_ (.A0(\as1802.regs[2][5] ),
    .A1(_0750_),
    .S(_1540_),
    .X(_1546_));
 sky130_fd_sc_hd__clkbuf_1 _4323_ (.A(_1546_),
    .X(_0149_));
 sky130_fd_sc_hd__mux2_1 _4324_ (.A0(\as1802.regs[2][6] ),
    .A1(_0806_),
    .S(_1540_),
    .X(_1547_));
 sky130_fd_sc_hd__clkbuf_1 _4325_ (.A(_1547_),
    .X(_0150_));
 sky130_fd_sc_hd__mux2_1 _4326_ (.A0(\as1802.regs[2][7] ),
    .A1(_0871_),
    .S(_1540_),
    .X(_1548_));
 sky130_fd_sc_hd__clkbuf_1 _4327_ (.A(_1548_),
    .X(_0151_));
 sky130_fd_sc_hd__and3_1 _4328_ (.A(_1430_),
    .B(_1357_),
    .C(_1389_),
    .X(_1549_));
 sky130_fd_sc_hd__buf_4 _4329_ (.A(_1549_),
    .X(_1550_));
 sky130_fd_sc_hd__mux2_1 _4330_ (.A0(\as1802.regs[1][0] ),
    .A1(_0395_),
    .S(_1550_),
    .X(_1551_));
 sky130_fd_sc_hd__clkbuf_1 _4331_ (.A(_1551_),
    .X(_0152_));
 sky130_fd_sc_hd__mux2_1 _4332_ (.A0(\as1802.regs[1][1] ),
    .A1(_0487_),
    .S(_1550_),
    .X(_1552_));
 sky130_fd_sc_hd__clkbuf_1 _4333_ (.A(_1552_),
    .X(_0153_));
 sky130_fd_sc_hd__mux2_1 _4334_ (.A0(\as1802.regs[1][2] ),
    .A1(_0549_),
    .S(_1550_),
    .X(_1553_));
 sky130_fd_sc_hd__clkbuf_1 _4335_ (.A(_1553_),
    .X(_0154_));
 sky130_fd_sc_hd__mux2_1 _4336_ (.A0(\as1802.regs[1][3] ),
    .A1(_0613_),
    .S(_1550_),
    .X(_1554_));
 sky130_fd_sc_hd__clkbuf_1 _4337_ (.A(_1554_),
    .X(_0155_));
 sky130_fd_sc_hd__mux2_1 _4338_ (.A0(\as1802.regs[1][4] ),
    .A1(_0683_),
    .S(_1550_),
    .X(_1555_));
 sky130_fd_sc_hd__clkbuf_1 _4339_ (.A(_1555_),
    .X(_0156_));
 sky130_fd_sc_hd__mux2_1 _4340_ (.A0(\as1802.regs[1][5] ),
    .A1(_0750_),
    .S(_1550_),
    .X(_1556_));
 sky130_fd_sc_hd__clkbuf_1 _4341_ (.A(_1556_),
    .X(_0157_));
 sky130_fd_sc_hd__mux2_1 _4342_ (.A0(\as1802.regs[1][6] ),
    .A1(_0806_),
    .S(_1550_),
    .X(_1557_));
 sky130_fd_sc_hd__clkbuf_1 _4343_ (.A(_1557_),
    .X(_0158_));
 sky130_fd_sc_hd__mux2_1 _4344_ (.A0(\as1802.regs[1][7] ),
    .A1(_0871_),
    .S(_1550_),
    .X(_1558_));
 sky130_fd_sc_hd__clkbuf_1 _4345_ (.A(_1558_),
    .X(_0159_));
 sky130_fd_sc_hd__and3_1 _4346_ (.A(_0402_),
    .B(_0409_),
    .C(_0945_),
    .X(_1559_));
 sky130_fd_sc_hd__buf_4 _4347_ (.A(_1559_),
    .X(_1560_));
 sky130_fd_sc_hd__mux2_1 _4348_ (.A0(\as1802.regs[15][8] ),
    .A1(_0940_),
    .S(_1560_),
    .X(_1561_));
 sky130_fd_sc_hd__clkbuf_1 _4349_ (.A(_1561_),
    .X(_0160_));
 sky130_fd_sc_hd__mux2_1 _4350_ (.A0(\as1802.regs[15][9] ),
    .A1(_1008_),
    .S(_1560_),
    .X(_1562_));
 sky130_fd_sc_hd__clkbuf_1 _4351_ (.A(_1562_),
    .X(_0161_));
 sky130_fd_sc_hd__mux2_1 _4352_ (.A0(\as1802.regs[15][10] ),
    .A1(_1069_),
    .S(_1560_),
    .X(_1563_));
 sky130_fd_sc_hd__clkbuf_1 _4353_ (.A(_1563_),
    .X(_0162_));
 sky130_fd_sc_hd__mux2_1 _4354_ (.A0(\as1802.regs[15][11] ),
    .A1(_1135_),
    .S(_1560_),
    .X(_1564_));
 sky130_fd_sc_hd__clkbuf_1 _4355_ (.A(_1564_),
    .X(_0163_));
 sky130_fd_sc_hd__mux2_1 _4356_ (.A0(\as1802.regs[15][12] ),
    .A1(_1189_),
    .S(_1560_),
    .X(_1565_));
 sky130_fd_sc_hd__clkbuf_1 _4357_ (.A(_1565_),
    .X(_0164_));
 sky130_fd_sc_hd__mux2_1 _4358_ (.A0(\as1802.regs[15][13] ),
    .A1(_1247_),
    .S(_1560_),
    .X(_1566_));
 sky130_fd_sc_hd__clkbuf_1 _4359_ (.A(_1566_),
    .X(_0165_));
 sky130_fd_sc_hd__mux2_1 _4360_ (.A0(\as1802.regs[15][14] ),
    .A1(_1299_),
    .S(_1560_),
    .X(_1567_));
 sky130_fd_sc_hd__clkbuf_1 _4361_ (.A(_1567_),
    .X(_0166_));
 sky130_fd_sc_hd__mux2_1 _4362_ (.A0(\as1802.regs[15][15] ),
    .A1(_1352_),
    .S(_1560_),
    .X(_1568_));
 sky130_fd_sc_hd__clkbuf_1 _4363_ (.A(_1568_),
    .X(_0167_));
 sky130_fd_sc_hd__and3_1 _4364_ (.A(_0409_),
    .B(_0411_),
    .C(_0941_),
    .X(_1569_));
 sky130_fd_sc_hd__buf_4 _4365_ (.A(_1569_),
    .X(_1570_));
 sky130_fd_sc_hd__mux2_1 _4366_ (.A0(\as1802.regs[14][0] ),
    .A1(_0394_),
    .S(_1570_),
    .X(_1571_));
 sky130_fd_sc_hd__clkbuf_1 _4367_ (.A(_1571_),
    .X(_0168_));
 sky130_fd_sc_hd__mux2_1 _4368_ (.A0(\as1802.regs[14][1] ),
    .A1(_0486_),
    .S(_1570_),
    .X(_1572_));
 sky130_fd_sc_hd__clkbuf_1 _4369_ (.A(_1572_),
    .X(_0169_));
 sky130_fd_sc_hd__mux2_1 _4370_ (.A0(\as1802.regs[14][2] ),
    .A1(_0548_),
    .S(_1570_),
    .X(_1573_));
 sky130_fd_sc_hd__clkbuf_1 _4371_ (.A(_1573_),
    .X(_0170_));
 sky130_fd_sc_hd__mux2_1 _4372_ (.A0(\as1802.regs[14][3] ),
    .A1(_0612_),
    .S(_1570_),
    .X(_1574_));
 sky130_fd_sc_hd__clkbuf_1 _4373_ (.A(_1574_),
    .X(_0171_));
 sky130_fd_sc_hd__mux2_1 _4374_ (.A0(\as1802.regs[14][4] ),
    .A1(_0682_),
    .S(_1570_),
    .X(_1575_));
 sky130_fd_sc_hd__clkbuf_1 _4375_ (.A(_1575_),
    .X(_0172_));
 sky130_fd_sc_hd__mux2_1 _4376_ (.A0(\as1802.regs[14][5] ),
    .A1(_0749_),
    .S(_1570_),
    .X(_1576_));
 sky130_fd_sc_hd__clkbuf_1 _4377_ (.A(_1576_),
    .X(_0173_));
 sky130_fd_sc_hd__mux2_1 _4378_ (.A0(\as1802.regs[14][6] ),
    .A1(_0805_),
    .S(_1570_),
    .X(_1577_));
 sky130_fd_sc_hd__clkbuf_1 _4379_ (.A(_1577_),
    .X(_0174_));
 sky130_fd_sc_hd__mux2_1 _4380_ (.A0(\as1802.regs[14][7] ),
    .A1(_0870_),
    .S(_1570_),
    .X(_1578_));
 sky130_fd_sc_hd__clkbuf_1 _4381_ (.A(_1578_),
    .X(_0175_));
 sky130_fd_sc_hd__and3_1 _4382_ (.A(_0409_),
    .B(_0411_),
    .C(_1389_),
    .X(_1579_));
 sky130_fd_sc_hd__buf_4 _4383_ (.A(_1579_),
    .X(_1580_));
 sky130_fd_sc_hd__mux2_1 _4384_ (.A0(\as1802.regs[13][0] ),
    .A1(_0394_),
    .S(_1580_),
    .X(_1581_));
 sky130_fd_sc_hd__clkbuf_1 _4385_ (.A(_1581_),
    .X(_0176_));
 sky130_fd_sc_hd__mux2_1 _4386_ (.A0(\as1802.regs[13][1] ),
    .A1(_0486_),
    .S(_1580_),
    .X(_1582_));
 sky130_fd_sc_hd__clkbuf_1 _4387_ (.A(_1582_),
    .X(_0177_));
 sky130_fd_sc_hd__mux2_1 _4388_ (.A0(\as1802.regs[13][2] ),
    .A1(_0548_),
    .S(_1580_),
    .X(_1583_));
 sky130_fd_sc_hd__clkbuf_1 _4389_ (.A(_1583_),
    .X(_0178_));
 sky130_fd_sc_hd__mux2_1 _4390_ (.A0(\as1802.regs[13][3] ),
    .A1(_0612_),
    .S(_1580_),
    .X(_1584_));
 sky130_fd_sc_hd__clkbuf_1 _4391_ (.A(_1584_),
    .X(_0179_));
 sky130_fd_sc_hd__mux2_1 _4392_ (.A0(\as1802.regs[13][4] ),
    .A1(_0682_),
    .S(_1580_),
    .X(_1585_));
 sky130_fd_sc_hd__clkbuf_1 _4393_ (.A(_1585_),
    .X(_0180_));
 sky130_fd_sc_hd__mux2_1 _4394_ (.A0(\as1802.regs[13][5] ),
    .A1(_0749_),
    .S(_1580_),
    .X(_1586_));
 sky130_fd_sc_hd__clkbuf_1 _4395_ (.A(_1586_),
    .X(_0181_));
 sky130_fd_sc_hd__mux2_1 _4396_ (.A0(\as1802.regs[13][6] ),
    .A1(_0805_),
    .S(_1580_),
    .X(_1587_));
 sky130_fd_sc_hd__clkbuf_1 _4397_ (.A(_1587_),
    .X(_0182_));
 sky130_fd_sc_hd__mux2_1 _4398_ (.A0(\as1802.regs[13][7] ),
    .A1(_0870_),
    .S(_1580_),
    .X(_1588_));
 sky130_fd_sc_hd__clkbuf_1 _4399_ (.A(_1588_),
    .X(_0183_));
 sky130_fd_sc_hd__and3_1 _4400_ (.A(_0409_),
    .B(_1354_),
    .C(_1355_),
    .X(_1589_));
 sky130_fd_sc_hd__buf_4 _4401_ (.A(_1589_),
    .X(_1590_));
 sky130_fd_sc_hd__mux2_1 _4402_ (.A0(\as1802.regs[12][8] ),
    .A1(_0940_),
    .S(_1590_),
    .X(_1591_));
 sky130_fd_sc_hd__clkbuf_1 _4403_ (.A(_1591_),
    .X(_0184_));
 sky130_fd_sc_hd__mux2_1 _4404_ (.A0(\as1802.regs[12][9] ),
    .A1(_1008_),
    .S(_1590_),
    .X(_1592_));
 sky130_fd_sc_hd__clkbuf_1 _4405_ (.A(_1592_),
    .X(_0185_));
 sky130_fd_sc_hd__mux2_1 _4406_ (.A0(\as1802.regs[12][10] ),
    .A1(_1069_),
    .S(_1590_),
    .X(_1593_));
 sky130_fd_sc_hd__clkbuf_1 _4407_ (.A(_1593_),
    .X(_0186_));
 sky130_fd_sc_hd__mux2_1 _4408_ (.A0(\as1802.regs[12][11] ),
    .A1(_1135_),
    .S(_1590_),
    .X(_1594_));
 sky130_fd_sc_hd__clkbuf_1 _4409_ (.A(_1594_),
    .X(_0187_));
 sky130_fd_sc_hd__mux2_1 _4410_ (.A0(\as1802.regs[12][12] ),
    .A1(_1189_),
    .S(_1590_),
    .X(_1595_));
 sky130_fd_sc_hd__clkbuf_1 _4411_ (.A(_1595_),
    .X(_0188_));
 sky130_fd_sc_hd__mux2_1 _4412_ (.A0(\as1802.regs[12][13] ),
    .A1(_1247_),
    .S(_1590_),
    .X(_1596_));
 sky130_fd_sc_hd__clkbuf_1 _4413_ (.A(_1596_),
    .X(_0189_));
 sky130_fd_sc_hd__mux2_1 _4414_ (.A0(\as1802.regs[12][14] ),
    .A1(_1299_),
    .S(_1590_),
    .X(_1597_));
 sky130_fd_sc_hd__clkbuf_1 _4415_ (.A(_1597_),
    .X(_0190_));
 sky130_fd_sc_hd__mux2_1 _4416_ (.A0(\as1802.regs[12][15] ),
    .A1(_1352_),
    .S(_1590_),
    .X(_1598_));
 sky130_fd_sc_hd__clkbuf_1 _4417_ (.A(_1598_),
    .X(_0191_));
 sky130_fd_sc_hd__and3_1 _4418_ (.A(_0402_),
    .B(_0411_),
    .C(_0943_),
    .X(_1599_));
 sky130_fd_sc_hd__buf_4 _4419_ (.A(_1599_),
    .X(_1600_));
 sky130_fd_sc_hd__mux2_1 _4420_ (.A0(\as1802.regs[11][0] ),
    .A1(_0394_),
    .S(_1600_),
    .X(_1601_));
 sky130_fd_sc_hd__clkbuf_1 _4421_ (.A(_1601_),
    .X(_0192_));
 sky130_fd_sc_hd__mux2_1 _4422_ (.A0(\as1802.regs[11][1] ),
    .A1(_0486_),
    .S(_1600_),
    .X(_1602_));
 sky130_fd_sc_hd__clkbuf_1 _4423_ (.A(_1602_),
    .X(_0193_));
 sky130_fd_sc_hd__mux2_1 _4424_ (.A0(\as1802.regs[11][2] ),
    .A1(_0548_),
    .S(_1600_),
    .X(_1603_));
 sky130_fd_sc_hd__clkbuf_1 _4425_ (.A(_1603_),
    .X(_0194_));
 sky130_fd_sc_hd__mux2_1 _4426_ (.A0(\as1802.regs[11][3] ),
    .A1(_0612_),
    .S(_1600_),
    .X(_1604_));
 sky130_fd_sc_hd__clkbuf_1 _4427_ (.A(_1604_),
    .X(_0195_));
 sky130_fd_sc_hd__mux2_1 _4428_ (.A0(\as1802.regs[11][4] ),
    .A1(_0682_),
    .S(_1600_),
    .X(_1605_));
 sky130_fd_sc_hd__clkbuf_1 _4429_ (.A(_1605_),
    .X(_0196_));
 sky130_fd_sc_hd__mux2_1 _4430_ (.A0(\as1802.regs[11][5] ),
    .A1(_0749_),
    .S(_1600_),
    .X(_1606_));
 sky130_fd_sc_hd__clkbuf_1 _4431_ (.A(_1606_),
    .X(_0197_));
 sky130_fd_sc_hd__mux2_1 _4432_ (.A0(\as1802.regs[11][6] ),
    .A1(_0805_),
    .S(_1600_),
    .X(_1607_));
 sky130_fd_sc_hd__clkbuf_1 _4433_ (.A(_1607_),
    .X(_0198_));
 sky130_fd_sc_hd__mux2_1 _4434_ (.A0(\as1802.regs[11][7] ),
    .A1(_0870_),
    .S(_1600_),
    .X(_1608_));
 sky130_fd_sc_hd__clkbuf_1 _4435_ (.A(_1608_),
    .X(_0199_));
 sky130_fd_sc_hd__and3_1 _4436_ (.A(_1430_),
    .B(_0941_),
    .C(_0943_),
    .X(_1609_));
 sky130_fd_sc_hd__buf_4 _4437_ (.A(_1609_),
    .X(_1610_));
 sky130_fd_sc_hd__mux2_1 _4438_ (.A0(\as1802.regs[10][0] ),
    .A1(_0394_),
    .S(_1610_),
    .X(_1611_));
 sky130_fd_sc_hd__clkbuf_1 _4439_ (.A(_1611_),
    .X(_0200_));
 sky130_fd_sc_hd__mux2_1 _4440_ (.A0(\as1802.regs[10][1] ),
    .A1(_0486_),
    .S(_1610_),
    .X(_1612_));
 sky130_fd_sc_hd__clkbuf_1 _4441_ (.A(_1612_),
    .X(_0201_));
 sky130_fd_sc_hd__mux2_1 _4442_ (.A0(\as1802.regs[10][2] ),
    .A1(_0548_),
    .S(_1610_),
    .X(_1613_));
 sky130_fd_sc_hd__clkbuf_1 _4443_ (.A(_1613_),
    .X(_0202_));
 sky130_fd_sc_hd__mux2_1 _4444_ (.A0(\as1802.regs[10][3] ),
    .A1(_0612_),
    .S(_1610_),
    .X(_1614_));
 sky130_fd_sc_hd__clkbuf_1 _4445_ (.A(_1614_),
    .X(_0203_));
 sky130_fd_sc_hd__mux2_1 _4446_ (.A0(\as1802.regs[10][4] ),
    .A1(_0682_),
    .S(_1610_),
    .X(_1615_));
 sky130_fd_sc_hd__clkbuf_1 _4447_ (.A(_1615_),
    .X(_0204_));
 sky130_fd_sc_hd__mux2_1 _4448_ (.A0(\as1802.regs[10][5] ),
    .A1(_0749_),
    .S(_1610_),
    .X(_1616_));
 sky130_fd_sc_hd__clkbuf_1 _4449_ (.A(_1616_),
    .X(_0205_));
 sky130_fd_sc_hd__mux2_1 _4450_ (.A0(\as1802.regs[10][6] ),
    .A1(_0805_),
    .S(_1610_),
    .X(_1617_));
 sky130_fd_sc_hd__clkbuf_1 _4451_ (.A(_1617_),
    .X(_0206_));
 sky130_fd_sc_hd__mux2_1 _4452_ (.A0(\as1802.regs[10][7] ),
    .A1(_0870_),
    .S(_1610_),
    .X(_1618_));
 sky130_fd_sc_hd__clkbuf_1 _4453_ (.A(_1618_),
    .X(_0207_));
 sky130_fd_sc_hd__and3_1 _4454_ (.A(_1430_),
    .B(_1355_),
    .C(_1357_),
    .X(_1619_));
 sky130_fd_sc_hd__buf_4 _4455_ (.A(_1619_),
    .X(_1620_));
 sky130_fd_sc_hd__mux2_1 _4456_ (.A0(\as1802.regs[0][0] ),
    .A1(_0394_),
    .S(_1620_),
    .X(_1621_));
 sky130_fd_sc_hd__clkbuf_1 _4457_ (.A(_1621_),
    .X(_0208_));
 sky130_fd_sc_hd__mux2_1 _4458_ (.A0(\as1802.regs[0][1] ),
    .A1(_0486_),
    .S(_1620_),
    .X(_1622_));
 sky130_fd_sc_hd__clkbuf_1 _4459_ (.A(_1622_),
    .X(_0209_));
 sky130_fd_sc_hd__mux2_1 _4460_ (.A0(\as1802.regs[0][2] ),
    .A1(_0548_),
    .S(_1620_),
    .X(_1623_));
 sky130_fd_sc_hd__clkbuf_1 _4461_ (.A(_1623_),
    .X(_0210_));
 sky130_fd_sc_hd__mux2_1 _4462_ (.A0(\as1802.regs[0][3] ),
    .A1(_0612_),
    .S(_1620_),
    .X(_1624_));
 sky130_fd_sc_hd__clkbuf_1 _4463_ (.A(_1624_),
    .X(_0211_));
 sky130_fd_sc_hd__mux2_1 _4464_ (.A0(\as1802.regs[0][4] ),
    .A1(_0682_),
    .S(_1620_),
    .X(_1625_));
 sky130_fd_sc_hd__clkbuf_1 _4465_ (.A(_1625_),
    .X(_0212_));
 sky130_fd_sc_hd__mux2_1 _4466_ (.A0(\as1802.regs[0][5] ),
    .A1(_0749_),
    .S(_1620_),
    .X(_1626_));
 sky130_fd_sc_hd__clkbuf_1 _4467_ (.A(_1626_),
    .X(_0213_));
 sky130_fd_sc_hd__mux2_1 _4468_ (.A0(\as1802.regs[0][6] ),
    .A1(_0805_),
    .S(_1620_),
    .X(_1627_));
 sky130_fd_sc_hd__clkbuf_1 _4469_ (.A(_1627_),
    .X(_0214_));
 sky130_fd_sc_hd__mux2_1 _4470_ (.A0(\as1802.regs[0][7] ),
    .A1(_0870_),
    .S(_1620_),
    .X(_1628_));
 sky130_fd_sc_hd__clkbuf_1 _4471_ (.A(_1628_),
    .X(_0215_));
 sky130_fd_sc_hd__and3_1 _4472_ (.A(_0409_),
    .B(_0941_),
    .C(_0945_),
    .X(_1629_));
 sky130_fd_sc_hd__buf_4 _4473_ (.A(_1629_),
    .X(_1630_));
 sky130_fd_sc_hd__mux2_1 _4474_ (.A0(\as1802.regs[14][8] ),
    .A1(_0939_),
    .S(_1630_),
    .X(_1631_));
 sky130_fd_sc_hd__clkbuf_1 _4475_ (.A(_1631_),
    .X(_0216_));
 sky130_fd_sc_hd__mux2_1 _4476_ (.A0(\as1802.regs[14][9] ),
    .A1(_1007_),
    .S(_1630_),
    .X(_1632_));
 sky130_fd_sc_hd__clkbuf_1 _4477_ (.A(_1632_),
    .X(_0217_));
 sky130_fd_sc_hd__mux2_1 _4478_ (.A0(\as1802.regs[14][10] ),
    .A1(_1068_),
    .S(_1630_),
    .X(_1633_));
 sky130_fd_sc_hd__clkbuf_1 _4479_ (.A(_1633_),
    .X(_0218_));
 sky130_fd_sc_hd__mux2_1 _4480_ (.A0(\as1802.regs[14][11] ),
    .A1(_1134_),
    .S(_1630_),
    .X(_1634_));
 sky130_fd_sc_hd__clkbuf_1 _4481_ (.A(_1634_),
    .X(_0219_));
 sky130_fd_sc_hd__mux2_1 _4482_ (.A0(\as1802.regs[14][12] ),
    .A1(_1188_),
    .S(_1630_),
    .X(_1635_));
 sky130_fd_sc_hd__clkbuf_1 _4483_ (.A(_1635_),
    .X(_0220_));
 sky130_fd_sc_hd__mux2_1 _4484_ (.A0(\as1802.regs[14][13] ),
    .A1(_1246_),
    .S(_1630_),
    .X(_1636_));
 sky130_fd_sc_hd__clkbuf_1 _4485_ (.A(_1636_),
    .X(_0221_));
 sky130_fd_sc_hd__mux2_1 _4486_ (.A0(\as1802.regs[14][14] ),
    .A1(_1298_),
    .S(_1630_),
    .X(_1637_));
 sky130_fd_sc_hd__clkbuf_1 _4487_ (.A(_1637_),
    .X(_0222_));
 sky130_fd_sc_hd__mux2_1 _4488_ (.A0(\as1802.regs[14][15] ),
    .A1(_1351_),
    .S(_1630_),
    .X(_1638_));
 sky130_fd_sc_hd__clkbuf_1 _4489_ (.A(_1638_),
    .X(_0223_));
 sky130_fd_sc_hd__and3_1 _4490_ (.A(_0409_),
    .B(_1354_),
    .C(_1389_),
    .X(_1639_));
 sky130_fd_sc_hd__buf_4 _4491_ (.A(_1639_),
    .X(_1640_));
 sky130_fd_sc_hd__mux2_1 _4492_ (.A0(\as1802.regs[13][8] ),
    .A1(_0939_),
    .S(_1640_),
    .X(_1641_));
 sky130_fd_sc_hd__clkbuf_1 _4493_ (.A(_1641_),
    .X(_0224_));
 sky130_fd_sc_hd__mux2_1 _4494_ (.A0(\as1802.regs[13][9] ),
    .A1(_1007_),
    .S(_1640_),
    .X(_1642_));
 sky130_fd_sc_hd__clkbuf_1 _4495_ (.A(_1642_),
    .X(_0225_));
 sky130_fd_sc_hd__mux2_1 _4496_ (.A0(\as1802.regs[13][10] ),
    .A1(_1068_),
    .S(_1640_),
    .X(_1643_));
 sky130_fd_sc_hd__clkbuf_1 _4497_ (.A(_1643_),
    .X(_0226_));
 sky130_fd_sc_hd__mux2_1 _4498_ (.A0(\as1802.regs[13][11] ),
    .A1(_1134_),
    .S(_1640_),
    .X(_1644_));
 sky130_fd_sc_hd__clkbuf_1 _4499_ (.A(_1644_),
    .X(_0227_));
 sky130_fd_sc_hd__mux2_1 _4500_ (.A0(\as1802.regs[13][12] ),
    .A1(_1188_),
    .S(_1640_),
    .X(_1645_));
 sky130_fd_sc_hd__clkbuf_1 _4501_ (.A(_1645_),
    .X(_0228_));
 sky130_fd_sc_hd__mux2_1 _4502_ (.A0(\as1802.regs[13][13] ),
    .A1(_1246_),
    .S(_1640_),
    .X(_1646_));
 sky130_fd_sc_hd__clkbuf_1 _4503_ (.A(_1646_),
    .X(_0229_));
 sky130_fd_sc_hd__mux2_1 _4504_ (.A0(\as1802.regs[13][14] ),
    .A1(_1298_),
    .S(_1640_),
    .X(_1647_));
 sky130_fd_sc_hd__clkbuf_1 _4505_ (.A(_1647_),
    .X(_0230_));
 sky130_fd_sc_hd__mux2_1 _4506_ (.A0(\as1802.regs[13][15] ),
    .A1(_1351_),
    .S(_1640_),
    .X(_1648_));
 sky130_fd_sc_hd__clkbuf_1 _4507_ (.A(_1648_),
    .X(_0231_));
 sky130_fd_sc_hd__and3_1 _4508_ (.A(_0409_),
    .B(_0411_),
    .C(_1355_),
    .X(_1649_));
 sky130_fd_sc_hd__buf_4 _4509_ (.A(_1649_),
    .X(_1650_));
 sky130_fd_sc_hd__mux2_1 _4510_ (.A0(\as1802.regs[12][0] ),
    .A1(_0394_),
    .S(_1650_),
    .X(_1651_));
 sky130_fd_sc_hd__clkbuf_1 _4511_ (.A(_1651_),
    .X(_0232_));
 sky130_fd_sc_hd__mux2_1 _4512_ (.A0(\as1802.regs[12][1] ),
    .A1(_0486_),
    .S(_1650_),
    .X(_1652_));
 sky130_fd_sc_hd__clkbuf_1 _4513_ (.A(_1652_),
    .X(_0233_));
 sky130_fd_sc_hd__mux2_1 _4514_ (.A0(\as1802.regs[12][2] ),
    .A1(_0548_),
    .S(_1650_),
    .X(_1653_));
 sky130_fd_sc_hd__clkbuf_1 _4515_ (.A(_1653_),
    .X(_0234_));
 sky130_fd_sc_hd__mux2_1 _4516_ (.A0(\as1802.regs[12][3] ),
    .A1(_0612_),
    .S(_1650_),
    .X(_1654_));
 sky130_fd_sc_hd__clkbuf_1 _4517_ (.A(_1654_),
    .X(_0235_));
 sky130_fd_sc_hd__mux2_1 _4518_ (.A0(\as1802.regs[12][4] ),
    .A1(_0682_),
    .S(_1650_),
    .X(_1655_));
 sky130_fd_sc_hd__clkbuf_1 _4519_ (.A(_1655_),
    .X(_0236_));
 sky130_fd_sc_hd__mux2_1 _4520_ (.A0(\as1802.regs[12][5] ),
    .A1(_0749_),
    .S(_1650_),
    .X(_1656_));
 sky130_fd_sc_hd__clkbuf_1 _4521_ (.A(_1656_),
    .X(_0237_));
 sky130_fd_sc_hd__mux2_1 _4522_ (.A0(\as1802.regs[12][6] ),
    .A1(_0805_),
    .S(_1650_),
    .X(_1657_));
 sky130_fd_sc_hd__clkbuf_1 _4523_ (.A(_1657_),
    .X(_0238_));
 sky130_fd_sc_hd__mux2_1 _4524_ (.A0(\as1802.regs[12][7] ),
    .A1(_0870_),
    .S(_1650_),
    .X(_1658_));
 sky130_fd_sc_hd__clkbuf_1 _4525_ (.A(_1658_),
    .X(_0239_));
 sky130_fd_sc_hd__and3_1 _4526_ (.A(_0402_),
    .B(_0943_),
    .C(_0945_),
    .X(_1659_));
 sky130_fd_sc_hd__buf_4 _4527_ (.A(_1659_),
    .X(_1660_));
 sky130_fd_sc_hd__mux2_1 _4528_ (.A0(\as1802.regs[11][8] ),
    .A1(_0939_),
    .S(_1660_),
    .X(_1661_));
 sky130_fd_sc_hd__clkbuf_1 _4529_ (.A(_1661_),
    .X(_0240_));
 sky130_fd_sc_hd__mux2_1 _4530_ (.A0(\as1802.regs[11][9] ),
    .A1(_1007_),
    .S(_1660_),
    .X(_1662_));
 sky130_fd_sc_hd__clkbuf_1 _4531_ (.A(_1662_),
    .X(_0241_));
 sky130_fd_sc_hd__mux2_1 _4532_ (.A0(\as1802.regs[11][10] ),
    .A1(_1068_),
    .S(_1660_),
    .X(_1663_));
 sky130_fd_sc_hd__clkbuf_1 _4533_ (.A(_1663_),
    .X(_0242_));
 sky130_fd_sc_hd__mux2_1 _4534_ (.A0(\as1802.regs[11][11] ),
    .A1(_1134_),
    .S(_1660_),
    .X(_1664_));
 sky130_fd_sc_hd__clkbuf_1 _4535_ (.A(_1664_),
    .X(_0243_));
 sky130_fd_sc_hd__mux2_1 _4536_ (.A0(\as1802.regs[11][12] ),
    .A1(_1188_),
    .S(_1660_),
    .X(_1665_));
 sky130_fd_sc_hd__clkbuf_1 _4537_ (.A(_1665_),
    .X(_0244_));
 sky130_fd_sc_hd__mux2_1 _4538_ (.A0(\as1802.regs[11][13] ),
    .A1(_1246_),
    .S(_1660_),
    .X(_1666_));
 sky130_fd_sc_hd__clkbuf_1 _4539_ (.A(_1666_),
    .X(_0245_));
 sky130_fd_sc_hd__mux2_1 _4540_ (.A0(\as1802.regs[11][14] ),
    .A1(_1298_),
    .S(_1660_),
    .X(_1667_));
 sky130_fd_sc_hd__clkbuf_1 _4541_ (.A(_1667_),
    .X(_0246_));
 sky130_fd_sc_hd__mux2_1 _4542_ (.A0(\as1802.regs[11][15] ),
    .A1(_1351_),
    .S(_1660_),
    .X(_1668_));
 sky130_fd_sc_hd__clkbuf_1 _4543_ (.A(_1668_),
    .X(_0247_));
 sky130_fd_sc_hd__inv_2 _4544_ (.A(\as1802.mem_write ),
    .Y(_1669_));
 sky130_fd_sc_hd__inv_2 _4545_ (.A(\as1802.addr_buff[15] ),
    .Y(_1670_));
 sky130_fd_sc_hd__inv_2 _4546_ (.A(\as1802.last_hi_addr[5] ),
    .Y(_1671_));
 sky130_fd_sc_hd__xnor2_1 _4547_ (.A(\as1802.last_hi_addr[1] ),
    .B(\as1802.addr_buff[9] ),
    .Y(_1672_));
 sky130_fd_sc_hd__o221a_1 _4548_ (.A1(\as1802.last_hi_addr[7] ),
    .A2(_1670_),
    .B1(_1671_),
    .B2(\as1802.addr_buff[13] ),
    .C1(_1672_),
    .X(_1673_));
 sky130_fd_sc_hd__inv_2 _4549_ (.A(\as1802.addr_buff[13] ),
    .Y(_1674_));
 sky130_fd_sc_hd__inv_2 _4550_ (.A(\as1802.last_hi_addr[0] ),
    .Y(_1675_));
 sky130_fd_sc_hd__xnor2_1 _4551_ (.A(\as1802.last_hi_addr[3] ),
    .B(\as1802.addr_buff[11] ),
    .Y(_1676_));
 sky130_fd_sc_hd__o221a_1 _4552_ (.A1(\as1802.last_hi_addr[5] ),
    .A2(_1674_),
    .B1(_1675_),
    .B2(\as1802.addr_buff[8] ),
    .C1(_1676_),
    .X(_1677_));
 sky130_fd_sc_hd__xnor2_1 _4553_ (.A(\as1802.last_hi_addr[6] ),
    .B(\as1802.addr_buff[14] ),
    .Y(_1678_));
 sky130_fd_sc_hd__inv_2 _4554_ (.A(\as1802.last_hi_addr[7] ),
    .Y(_1679_));
 sky130_fd_sc_hd__inv_2 _4555_ (.A(\as1802.addr_buff[8] ),
    .Y(_1680_));
 sky130_fd_sc_hd__xnor2_1 _4556_ (.A(\as1802.last_hi_addr[4] ),
    .B(\as1802.addr_buff[12] ),
    .Y(_1681_));
 sky130_fd_sc_hd__o221a_1 _4557_ (.A1(_1679_),
    .A2(\as1802.addr_buff[15] ),
    .B1(\as1802.last_hi_addr[0] ),
    .B2(_1680_),
    .C1(_1681_),
    .X(_1682_));
 sky130_fd_sc_hd__xnor2_1 _4558_ (.A(\as1802.last_hi_addr[2] ),
    .B(\as1802.addr_buff[10] ),
    .Y(_1683_));
 sky130_fd_sc_hd__and3_1 _4559_ (.A(_1678_),
    .B(_1682_),
    .C(_1683_),
    .X(_1684_));
 sky130_fd_sc_hd__a31o_1 _4560_ (.A1(_1673_),
    .A2(_1677_),
    .A3(_1684_),
    .B1(\as1802.mem_cycle[1] ),
    .X(_1685_));
 sky130_fd_sc_hd__clkbuf_4 _4561_ (.A(_1685_),
    .X(_1686_));
 sky130_fd_sc_hd__inv_2 _4562_ (.A(\as1802.mem_cycle[0] ),
    .Y(_1687_));
 sky130_fd_sc_hd__nor2_1 _4563_ (.A(\as1802.mem_cycle[2] ),
    .B(_1687_),
    .Y(_1688_));
 sky130_fd_sc_hd__clkbuf_2 _4564_ (.A(_1688_),
    .X(_1689_));
 sky130_fd_sc_hd__and4b_1 _4565_ (.A_N(\as1802.will_interrupt ),
    .B(_2580_),
    .C(_2547_),
    .D(_2489_),
    .X(_1690_));
 sky130_fd_sc_hd__nor2_1 _4566_ (.A(_2580_),
    .B(_2460_),
    .Y(_1691_));
 sky130_fd_sc_hd__and3_1 _4567_ (.A(_2474_),
    .B(_2523_),
    .C(_1691_),
    .X(_1692_));
 sky130_fd_sc_hd__nor2_1 _4568_ (.A(_2460_),
    .B(_1476_),
    .Y(_1693_));
 sky130_fd_sc_hd__or2_1 _4569_ (.A(_2456_),
    .B(_1693_),
    .X(_1694_));
 sky130_fd_sc_hd__clkbuf_4 _4570_ (.A(_2611_),
    .X(_1695_));
 sky130_fd_sc_hd__o21a_1 _4571_ (.A1(_2610_),
    .A2(_1695_),
    .B1(_2613_),
    .X(_1696_));
 sky130_fd_sc_hd__or4b_1 _4572_ (.A(_1690_),
    .B(_1692_),
    .C(_1694_),
    .D_N(_1696_),
    .X(_1697_));
 sky130_fd_sc_hd__and2b_1 _4573_ (.A_N(_2477_),
    .B(_1474_),
    .X(_1698_));
 sky130_fd_sc_hd__nand2_1 _4574_ (.A(_1698_),
    .B(_0449_),
    .Y(_1699_));
 sky130_fd_sc_hd__or2_1 _4575_ (.A(_2463_),
    .B(_2478_),
    .X(_1700_));
 sky130_fd_sc_hd__a21o_1 _4576_ (.A1(_0383_),
    .A2(_1700_),
    .B1(_2610_),
    .X(_1701_));
 sky130_fd_sc_hd__nand2_1 _4577_ (.A(_2711_),
    .B(_2712_),
    .Y(_1702_));
 sky130_fd_sc_hd__and3_1 _4578_ (.A(_2542_),
    .B(_2565_),
    .C(_2544_),
    .X(_1703_));
 sky130_fd_sc_hd__a22oi_2 _4579_ (.A1(_2558_),
    .A2(_2711_),
    .B1(_1484_),
    .B2(_1703_),
    .Y(_1704_));
 sky130_fd_sc_hd__a221o_1 _4580_ (.A1(_2549_),
    .A2(_2521_),
    .B1(_1702_),
    .B2(_1704_),
    .C1(_2460_),
    .X(_1705_));
 sky130_fd_sc_hd__nand4_1 _4581_ (.A(_2486_),
    .B(_2482_),
    .C(_2520_),
    .D(_2551_),
    .Y(_1706_));
 sky130_fd_sc_hd__nor2_1 _4582_ (.A(_2555_),
    .B(_2600_),
    .Y(_1707_));
 sky130_fd_sc_hd__o21ai_1 _4583_ (.A1(_2555_),
    .A2(_2511_),
    .B1(_2593_),
    .Y(_1708_));
 sky130_fd_sc_hd__o31ai_1 _4584_ (.A1(_1707_),
    .A2(_1482_),
    .A3(_1708_),
    .B1(_2709_),
    .Y(_1709_));
 sky130_fd_sc_hd__nand2_1 _4585_ (.A(_2717_),
    .B(_2721_),
    .Y(_1710_));
 sky130_fd_sc_hd__or2_1 _4586_ (.A(_1709_),
    .B(_1710_),
    .X(_1711_));
 sky130_fd_sc_hd__inv_2 _4587_ (.A(_1711_),
    .Y(_1712_));
 sky130_fd_sc_hd__a31o_1 _4588_ (.A1(_0443_),
    .A2(_1706_),
    .A3(_1712_),
    .B1(_2460_),
    .X(_1713_));
 sky130_fd_sc_hd__o2111a_1 _4589_ (.A1(_2461_),
    .A2(_1699_),
    .B1(_1701_),
    .C1(_1705_),
    .D1(_1713_),
    .X(_1714_));
 sky130_fd_sc_hd__and3b_1 _4590_ (.A_N(_1697_),
    .B(_1714_),
    .C(_0385_),
    .X(_1715_));
 sky130_fd_sc_hd__nand2_1 _4591_ (.A(\as1802.mem_cycle[0] ),
    .B(_1715_),
    .Y(_1716_));
 sky130_fd_sc_hd__or2_1 _4592_ (.A(\as1802.mem_cycle[0] ),
    .B(_1715_),
    .X(_1717_));
 sky130_fd_sc_hd__a32o_1 _4593_ (.A1(_1669_),
    .A2(_1686_),
    .A3(_1689_),
    .B1(_1716_),
    .B2(_1717_),
    .X(_0248_));
 sky130_fd_sc_hd__inv_2 _4594_ (.A(_1685_),
    .Y(_1718_));
 sky130_fd_sc_hd__a32o_1 _4595_ (.A1(_1715_),
    .A2(_1718_),
    .A3(_1689_),
    .B1(_1716_),
    .B2(\as1802.mem_cycle[1] ),
    .X(_0249_));
 sky130_fd_sc_hd__a32o_1 _4596_ (.A1(_1715_),
    .A2(_1686_),
    .A3(_1689_),
    .B1(_1716_),
    .B2(\as1802.mem_cycle[2] ),
    .X(_0250_));
 sky130_fd_sc_hd__nand2_1 _4597_ (.A(_1702_),
    .B(_1706_),
    .Y(_1719_));
 sky130_fd_sc_hd__or2_1 _4598_ (.A(_2568_),
    .B(_2525_),
    .X(_1720_));
 sky130_fd_sc_hd__o211a_1 _4599_ (.A1(\as1802.will_interrupt ),
    .A2(_2487_),
    .B1(_2488_),
    .C1(_2580_),
    .X(_1721_));
 sky130_fd_sc_hd__and4_1 _4600_ (.A(_2486_),
    .B(_2464_),
    .C(_2561_),
    .D(_1700_),
    .X(_1722_));
 sky130_fd_sc_hd__o221a_1 _4601_ (.A1(_2580_),
    .A2(_1720_),
    .B1(_1721_),
    .B2(_1722_),
    .C1(_2467_),
    .X(_1723_));
 sky130_fd_sc_hd__nand4_1 _4602_ (.A(_1476_),
    .B(_1704_),
    .C(_1699_),
    .D(_1723_),
    .Y(_1724_));
 sky130_fd_sc_hd__or3_1 _4603_ (.A(_1711_),
    .B(_1719_),
    .C(_1724_),
    .X(_1725_));
 sky130_fd_sc_hd__clkbuf_4 _4604_ (.A(_1725_),
    .X(_1726_));
 sky130_fd_sc_hd__clkbuf_4 _4605_ (.A(_1726_),
    .X(_1727_));
 sky130_fd_sc_hd__buf_2 _4606_ (.A(_1727_),
    .X(_1728_));
 sky130_fd_sc_hd__nor2_4 _4607_ (.A(_2580_),
    .B(_2551_),
    .Y(_1729_));
 sky130_fd_sc_hd__clkbuf_4 _4608_ (.A(_1729_),
    .X(_1730_));
 sky130_fd_sc_hd__nor2_2 _4609_ (.A(_1698_),
    .B(_2563_),
    .Y(_1731_));
 sky130_fd_sc_hd__clkbuf_4 _4610_ (.A(_2704_),
    .X(_1732_));
 sky130_fd_sc_hd__buf_4 _4611_ (.A(_1288_),
    .X(_1733_));
 sky130_fd_sc_hd__o21a_1 _4612_ (.A1(_1733_),
    .A2(_2665_),
    .B1(_2695_),
    .X(_1734_));
 sky130_fd_sc_hd__nor2_1 _4613_ (.A(_1732_),
    .B(_2696_),
    .Y(_1735_));
 sky130_fd_sc_hd__a211o_1 _4614_ (.A1(_1732_),
    .A2(_1734_),
    .B1(_1735_),
    .C1(_1491_),
    .X(_1736_));
 sky130_fd_sc_hd__nor2_1 _4615_ (.A(_2513_),
    .B(_2593_),
    .Y(_1737_));
 sky130_fd_sc_hd__clkbuf_4 _4616_ (.A(_1737_),
    .X(_1738_));
 sky130_fd_sc_hd__a221o_1 _4617_ (.A1(_2590_),
    .A2(_1738_),
    .B1(_1734_),
    .B2(_2571_),
    .C1(_1495_),
    .X(_1739_));
 sky130_fd_sc_hd__buf_2 _4618_ (.A(_2570_),
    .X(_1740_));
 sky130_fd_sc_hd__clkbuf_4 _4619_ (.A(_2594_),
    .X(_1741_));
 sky130_fd_sc_hd__a31o_4 _4620_ (.A1(_1490_),
    .A2(_1740_),
    .A3(_1741_),
    .B1(_2563_),
    .X(_1742_));
 sky130_fd_sc_hd__a32o_1 _4621_ (.A1(_1731_),
    .A2(_1736_),
    .A3(_1739_),
    .B1(_2665_),
    .B2(_1742_),
    .X(_1743_));
 sky130_fd_sc_hd__nor2_1 _4622_ (.A(_2581_),
    .B(_2466_),
    .Y(_1744_));
 sky130_fd_sc_hd__buf_2 _4623_ (.A(_1744_),
    .X(_1745_));
 sky130_fd_sc_hd__buf_2 _4624_ (.A(_1475_),
    .X(_1746_));
 sky130_fd_sc_hd__a221o_1 _4625_ (.A1(_1745_),
    .A2(_2665_),
    .B1(_2720_),
    .B2(_1746_),
    .C1(_1726_),
    .X(_1747_));
 sky130_fd_sc_hd__a21oi_1 _4626_ (.A1(_1730_),
    .A2(_1743_),
    .B1(_1747_),
    .Y(_1748_));
 sky130_fd_sc_hd__a21o_1 _4627_ (.A1(\as1802.addr_buff[0] ),
    .A2(_1728_),
    .B1(_1748_),
    .X(_0251_));
 sky130_fd_sc_hd__or2_1 _4628_ (.A(_1698_),
    .B(_2563_),
    .X(_1749_));
 sky130_fd_sc_hd__buf_2 _4629_ (.A(_1749_),
    .X(_1750_));
 sky130_fd_sc_hd__inv_2 _4630_ (.A(_2572_),
    .Y(_1751_));
 sky130_fd_sc_hd__clkbuf_4 _4631_ (.A(_1741_),
    .X(_1752_));
 sky130_fd_sc_hd__or2_1 _4632_ (.A(_2553_),
    .B(_2570_),
    .X(_1753_));
 sky130_fd_sc_hd__nand2_1 _4633_ (.A(_2556_),
    .B(_0469_),
    .Y(_1754_));
 sky130_fd_sc_hd__o21ai_1 _4634_ (.A1(_1288_),
    .A2(_0439_),
    .B1(_1754_),
    .Y(_1755_));
 sky130_fd_sc_hd__mux2_1 _4635_ (.A0(_0469_),
    .A1(_1755_),
    .S(_2704_),
    .X(_1756_));
 sky130_fd_sc_hd__o22a_1 _4636_ (.A1(_1753_),
    .A2(_1755_),
    .B1(_1756_),
    .B2(_1490_),
    .X(_1757_));
 sky130_fd_sc_hd__o31a_1 _4637_ (.A1(\as1802.regs[2][1] ),
    .A2(_1751_),
    .A3(_1752_),
    .B1(_1757_),
    .X(_1758_));
 sky130_fd_sc_hd__a2bb2o_1 _4638_ (.A1_N(_1750_),
    .A2_N(_1758_),
    .B1(_1742_),
    .B2(_0439_),
    .X(_1759_));
 sky130_fd_sc_hd__a2bb2o_1 _4639_ (.A1_N(_0469_),
    .A2_N(_1729_),
    .B1(_1744_),
    .B2(_0439_),
    .X(_1760_));
 sky130_fd_sc_hd__a211o_1 _4640_ (.A1(_1730_),
    .A2(_1759_),
    .B1(_1760_),
    .C1(_1727_),
    .X(_1761_));
 sky130_fd_sc_hd__a21bo_1 _4641_ (.A1(\as1802.addr_buff[1] ),
    .A2(_1728_),
    .B1_N(_1761_),
    .X(_0252_));
 sky130_fd_sc_hd__mux2_1 _4642_ (.A0(_0507_),
    .A1(_0523_),
    .S(_1733_),
    .X(_1762_));
 sky130_fd_sc_hd__mux2_1 _4643_ (.A0(_0523_),
    .A1(_1762_),
    .S(_1732_),
    .X(_1763_));
 sky130_fd_sc_hd__buf_2 _4644_ (.A(_1740_),
    .X(_1764_));
 sky130_fd_sc_hd__o21ai_1 _4645_ (.A1(\as1802.regs[2][2] ),
    .A2(_1752_),
    .B1(_1740_),
    .Y(_1765_));
 sky130_fd_sc_hd__clkbuf_4 _4646_ (.A(_1490_),
    .X(_1766_));
 sky130_fd_sc_hd__o211a_1 _4647_ (.A1(_1764_),
    .A2(_1762_),
    .B1(_1765_),
    .C1(_1766_),
    .X(_1767_));
 sky130_fd_sc_hd__a21o_1 _4648_ (.A1(_1496_),
    .A2(_1763_),
    .B1(_1767_),
    .X(_1768_));
 sky130_fd_sc_hd__a22o_1 _4649_ (.A1(_0507_),
    .A2(_1742_),
    .B1(_1768_),
    .B2(_1731_),
    .X(_1769_));
 sky130_fd_sc_hd__a221o_1 _4650_ (.A1(_1745_),
    .A2(_0507_),
    .B1(_0523_),
    .B2(_1746_),
    .C1(_1726_),
    .X(_1770_));
 sky130_fd_sc_hd__a21oi_1 _4651_ (.A1(_1730_),
    .A2(_1769_),
    .B1(_1770_),
    .Y(_1771_));
 sky130_fd_sc_hd__a21o_1 _4652_ (.A1(\as1802.addr_buff[2] ),
    .A2(_1728_),
    .B1(_1771_),
    .X(_0253_));
 sky130_fd_sc_hd__nor2_1 _4653_ (.A(_2493_),
    .B(_0593_),
    .Y(_1772_));
 sky130_fd_sc_hd__a21o_1 _4654_ (.A1(_2493_),
    .A2(_0570_),
    .B1(_1772_),
    .X(_1773_));
 sky130_fd_sc_hd__or2_1 _4655_ (.A(_2479_),
    .B(_1773_),
    .X(_1774_));
 sky130_fd_sc_hd__nand2_1 _4656_ (.A(_2480_),
    .B(_0593_),
    .Y(_1775_));
 sky130_fd_sc_hd__o21ai_1 _4657_ (.A1(\as1802.regs[2][3] ),
    .A2(_2594_),
    .B1(_2570_),
    .Y(_1776_));
 sky130_fd_sc_hd__o211a_1 _4658_ (.A1(_2570_),
    .A2(_1773_),
    .B1(_1776_),
    .C1(_2526_),
    .X(_1777_));
 sky130_fd_sc_hd__a31o_1 _4659_ (.A1(_2554_),
    .A2(_1774_),
    .A3(_1775_),
    .B1(_1777_),
    .X(_1778_));
 sky130_fd_sc_hd__a22o_1 _4660_ (.A1(_0570_),
    .A2(_1742_),
    .B1(_1778_),
    .B2(_1731_),
    .X(_1779_));
 sky130_fd_sc_hd__a22o_1 _4661_ (.A1(_1744_),
    .A2(_0570_),
    .B1(_1729_),
    .B2(_1779_),
    .X(_1780_));
 sky130_fd_sc_hd__o21ba_1 _4662_ (.A1(_0593_),
    .A2(_1729_),
    .B1_N(_1780_),
    .X(_1781_));
 sky130_fd_sc_hd__mux2_1 _4663_ (.A0(_1781_),
    .A1(\as1802.addr_buff[3] ),
    .S(_1727_),
    .X(_1782_));
 sky130_fd_sc_hd__clkbuf_1 _4664_ (.A(_1782_),
    .X(_0254_));
 sky130_fd_sc_hd__a21oi_4 _4665_ (.A1(_2572_),
    .A2(_1741_),
    .B1(_2563_),
    .Y(_1783_));
 sky130_fd_sc_hd__nor2_1 _4666_ (.A(_2494_),
    .B(_0663_),
    .Y(_1784_));
 sky130_fd_sc_hd__a21o_1 _4667_ (.A1(_2494_),
    .A2(_0642_),
    .B1(_1784_),
    .X(_1785_));
 sky130_fd_sc_hd__o21ai_1 _4668_ (.A1(\as1802.regs[2][4] ),
    .A2(_1741_),
    .B1(_2570_),
    .Y(_1786_));
 sky130_fd_sc_hd__o211a_1 _4669_ (.A1(_2570_),
    .A2(_1785_),
    .B1(_1786_),
    .C1(_1490_),
    .X(_1787_));
 sky130_fd_sc_hd__nand2_1 _4670_ (.A(_2480_),
    .B(_0663_),
    .Y(_1788_));
 sky130_fd_sc_hd__o211a_1 _4671_ (.A1(_2480_),
    .A2(_1785_),
    .B1(_1788_),
    .C1(_2554_),
    .X(_1789_));
 sky130_fd_sc_hd__nor2_1 _4672_ (.A(_1787_),
    .B(_1789_),
    .Y(_1790_));
 sky130_fd_sc_hd__o22a_1 _4673_ (.A1(_0649_),
    .A2(_1783_),
    .B1(_1790_),
    .B2(_1750_),
    .X(_1791_));
 sky130_fd_sc_hd__o22a_1 _4674_ (.A1(_2466_),
    .A2(_0649_),
    .B1(_1791_),
    .B2(_2551_),
    .X(_1792_));
 sky130_fd_sc_hd__o22a_1 _4675_ (.A1(_0663_),
    .A2(_1729_),
    .B1(_1792_),
    .B2(_1489_),
    .X(_1793_));
 sky130_fd_sc_hd__mux2_1 _4676_ (.A0(_1793_),
    .A1(\as1802.addr_buff[4] ),
    .S(_1727_),
    .X(_1794_));
 sky130_fd_sc_hd__clkbuf_1 _4677_ (.A(_1794_),
    .X(_0255_));
 sky130_fd_sc_hd__nand2_1 _4678_ (.A(_1288_),
    .B(_0729_),
    .Y(_1795_));
 sky130_fd_sc_hd__o21a_1 _4679_ (.A1(_1288_),
    .A2(_0710_),
    .B1(_1795_),
    .X(_1796_));
 sky130_fd_sc_hd__or2_1 _4680_ (.A(_2480_),
    .B(_1796_),
    .X(_1797_));
 sky130_fd_sc_hd__nand2_1 _4681_ (.A(_2480_),
    .B(_0729_),
    .Y(_1798_));
 sky130_fd_sc_hd__o21ai_1 _4682_ (.A1(\as1802.regs[2][5] ),
    .A2(_1741_),
    .B1(_1740_),
    .Y(_1799_));
 sky130_fd_sc_hd__o211a_1 _4683_ (.A1(_1740_),
    .A2(_1796_),
    .B1(_1799_),
    .C1(_1490_),
    .X(_1800_));
 sky130_fd_sc_hd__a31o_1 _4684_ (.A1(_1495_),
    .A2(_1797_),
    .A3(_1798_),
    .B1(_1800_),
    .X(_1801_));
 sky130_fd_sc_hd__a22o_1 _4685_ (.A1(_0710_),
    .A2(_1742_),
    .B1(_1801_),
    .B2(_1731_),
    .X(_1802_));
 sky130_fd_sc_hd__o21bai_1 _4686_ (.A1(_0729_),
    .A2(_1730_),
    .B1_N(_1726_),
    .Y(_1803_));
 sky130_fd_sc_hd__a221o_1 _4687_ (.A1(_1745_),
    .A2(_0710_),
    .B1(_1730_),
    .B2(_1802_),
    .C1(_1803_),
    .X(_1804_));
 sky130_fd_sc_hd__a21bo_1 _4688_ (.A1(\as1802.addr_buff[5] ),
    .A2(_1727_),
    .B1_N(_1804_),
    .X(_0256_));
 sky130_fd_sc_hd__or2_1 _4689_ (.A(_2493_),
    .B(_0761_),
    .X(_1805_));
 sky130_fd_sc_hd__o211a_1 _4690_ (.A1(_2556_),
    .A2(_0792_),
    .B1(_1805_),
    .C1(_2571_),
    .X(_1806_));
 sky130_fd_sc_hd__o31a_1 _4691_ (.A1(\as1802.regs[2][6] ),
    .A2(_2553_),
    .A3(_1741_),
    .B1(_1753_),
    .X(_1807_));
 sky130_fd_sc_hd__o211a_1 _4692_ (.A1(_1288_),
    .A2(_0792_),
    .B1(_1805_),
    .C1(_2704_),
    .X(_1808_));
 sky130_fd_sc_hd__a21o_1 _4693_ (.A1(_2480_),
    .A2(_0761_),
    .B1(_1490_),
    .X(_1809_));
 sky130_fd_sc_hd__o22a_1 _4694_ (.A1(_1806_),
    .A2(_1807_),
    .B1(_1808_),
    .B2(_1809_),
    .X(_1810_));
 sky130_fd_sc_hd__o22a_1 _4695_ (.A1(_0792_),
    .A2(_1783_),
    .B1(_1810_),
    .B2(_1750_),
    .X(_1811_));
 sky130_fd_sc_hd__o22a_1 _4696_ (.A1(_2466_),
    .A2(_0792_),
    .B1(_1811_),
    .B2(_2551_),
    .X(_1812_));
 sky130_fd_sc_hd__o22a_1 _4697_ (.A1(_0761_),
    .A2(_1729_),
    .B1(_1812_),
    .B2(_1489_),
    .X(_1813_));
 sky130_fd_sc_hd__mux2_1 _4698_ (.A0(_1813_),
    .A1(\as1802.addr_buff[6] ),
    .S(_1727_),
    .X(_1814_));
 sky130_fd_sc_hd__clkbuf_1 _4699_ (.A(_1814_),
    .X(_0257_));
 sky130_fd_sc_hd__mux2_1 _4700_ (.A0(_0832_),
    .A1(_0853_),
    .S(_2556_),
    .X(_1815_));
 sky130_fd_sc_hd__or3_1 _4701_ (.A(\as1802.regs[2][7] ),
    .B(_2553_),
    .C(_2594_),
    .X(_1816_));
 sky130_fd_sc_hd__a22o_1 _4702_ (.A1(_2571_),
    .A2(_1815_),
    .B1(_1816_),
    .B2(_1753_),
    .X(_1817_));
 sky130_fd_sc_hd__a21o_1 _4703_ (.A1(_2479_),
    .A2(_0853_),
    .B1(_2526_),
    .X(_1818_));
 sky130_fd_sc_hd__a21o_1 _4704_ (.A1(_2704_),
    .A2(_1815_),
    .B1(_1818_),
    .X(_1819_));
 sky130_fd_sc_hd__a21oi_1 _4705_ (.A1(_1817_),
    .A2(_1819_),
    .B1(_1750_),
    .Y(_1820_));
 sky130_fd_sc_hd__a21oi_1 _4706_ (.A1(_0831_),
    .A2(_1742_),
    .B1(_1820_),
    .Y(_1821_));
 sky130_fd_sc_hd__o22a_1 _4707_ (.A1(_2466_),
    .A2(_0832_),
    .B1(_1821_),
    .B2(_2551_),
    .X(_1822_));
 sky130_fd_sc_hd__o22a_1 _4708_ (.A1(_0853_),
    .A2(_1729_),
    .B1(_1822_),
    .B2(_1489_),
    .X(_1823_));
 sky130_fd_sc_hd__mux2_1 _4709_ (.A0(_1823_),
    .A1(\as1802.addr_buff[7] ),
    .S(_1727_),
    .X(_1824_));
 sky130_fd_sc_hd__clkbuf_1 _4710_ (.A(_1824_),
    .X(_0258_));
 sky130_fd_sc_hd__mux2_1 _4711_ (.A0(_0904_),
    .A1(_0919_),
    .S(_1733_),
    .X(_1825_));
 sky130_fd_sc_hd__mux2_1 _4712_ (.A0(_0919_),
    .A1(_1825_),
    .S(_1732_),
    .X(_1826_));
 sky130_fd_sc_hd__o21ai_1 _4713_ (.A1(\as1802.regs[2][8] ),
    .A2(_1752_),
    .B1(_1740_),
    .Y(_1827_));
 sky130_fd_sc_hd__o211a_1 _4714_ (.A1(_1764_),
    .A2(_1825_),
    .B1(_1827_),
    .C1(_1766_),
    .X(_1828_));
 sky130_fd_sc_hd__a21o_1 _4715_ (.A1(_1496_),
    .A2(_1826_),
    .B1(_1828_),
    .X(_1829_));
 sky130_fd_sc_hd__a22o_1 _4716_ (.A1(_0904_),
    .A2(_1742_),
    .B1(_1829_),
    .B2(_1731_),
    .X(_1830_));
 sky130_fd_sc_hd__a221o_1 _4717_ (.A1(_1745_),
    .A2(_0904_),
    .B1(_0919_),
    .B2(_1746_),
    .C1(_1726_),
    .X(_1831_));
 sky130_fd_sc_hd__a21oi_1 _4718_ (.A1(_1730_),
    .A2(_1830_),
    .B1(_1831_),
    .Y(_1832_));
 sky130_fd_sc_hd__a21o_1 _4719_ (.A1(\as1802.addr_buff[8] ),
    .A2(_1728_),
    .B1(_1832_),
    .X(_0259_));
 sky130_fd_sc_hd__mux2_1 _4720_ (.A0(_0969_),
    .A1(_0998_),
    .S(_1288_),
    .X(_1833_));
 sky130_fd_sc_hd__mux2_1 _4721_ (.A0(_0998_),
    .A1(_1833_),
    .S(_1732_),
    .X(_1834_));
 sky130_fd_sc_hd__o21ai_1 _4722_ (.A1(\as1802.regs[2][9] ),
    .A2(_1752_),
    .B1(_1740_),
    .Y(_1835_));
 sky130_fd_sc_hd__o211a_1 _4723_ (.A1(_1764_),
    .A2(_1833_),
    .B1(_1835_),
    .C1(_1766_),
    .X(_1836_));
 sky130_fd_sc_hd__a21oi_1 _4724_ (.A1(_1496_),
    .A2(_1834_),
    .B1(_1836_),
    .Y(_1837_));
 sky130_fd_sc_hd__o22a_1 _4725_ (.A1(_1034_),
    .A2(_1783_),
    .B1(_1837_),
    .B2(_1750_),
    .X(_1838_));
 sky130_fd_sc_hd__a221o_1 _4726_ (.A1(_1745_),
    .A2(_0969_),
    .B1(_0998_),
    .B2(_1475_),
    .C1(_1726_),
    .X(_1839_));
 sky130_fd_sc_hd__o21ba_1 _4727_ (.A1(_1746_),
    .A2(_1838_),
    .B1_N(_1839_),
    .X(_1840_));
 sky130_fd_sc_hd__a21o_1 _4728_ (.A1(\as1802.addr_buff[9] ),
    .A2(_1728_),
    .B1(_1840_),
    .X(_0260_));
 sky130_fd_sc_hd__nand2_1 _4729_ (.A(_2556_),
    .B(_1050_),
    .Y(_1841_));
 sky130_fd_sc_hd__o211a_1 _4730_ (.A1(_2556_),
    .A2(_1032_),
    .B1(_1841_),
    .C1(_2704_),
    .X(_1842_));
 sky130_fd_sc_hd__nor2_1 _4731_ (.A(_2704_),
    .B(_1050_),
    .Y(_1843_));
 sky130_fd_sc_hd__o211a_1 _4732_ (.A1(_1288_),
    .A2(_1032_),
    .B1(_1841_),
    .C1(_2571_),
    .X(_1844_));
 sky130_fd_sc_hd__o31a_1 _4733_ (.A1(\as1802.regs[2][10] ),
    .A2(_2553_),
    .A3(_1741_),
    .B1(_1753_),
    .X(_1845_));
 sky130_fd_sc_hd__o32a_1 _4734_ (.A1(_1490_),
    .A2(_1842_),
    .A3(_1843_),
    .B1(_1844_),
    .B2(_1845_),
    .X(_1846_));
 sky130_fd_sc_hd__o22a_1 _4735_ (.A1(_1032_),
    .A2(_1783_),
    .B1(_1846_),
    .B2(_1750_),
    .X(_1847_));
 sky130_fd_sc_hd__o22a_1 _4736_ (.A1(_2466_),
    .A2(_1032_),
    .B1(_1847_),
    .B2(_2551_),
    .X(_1848_));
 sky130_fd_sc_hd__o22a_1 _4737_ (.A1(_1052_),
    .A2(_1729_),
    .B1(_1848_),
    .B2(_1489_),
    .X(_1849_));
 sky130_fd_sc_hd__mux2_1 _4738_ (.A0(_1849_),
    .A1(\as1802.addr_buff[10] ),
    .S(_1727_),
    .X(_1850_));
 sky130_fd_sc_hd__clkbuf_1 _4739_ (.A(_1850_),
    .X(_0261_));
 sky130_fd_sc_hd__mux2_1 _4740_ (.A0(_1115_),
    .A1(_1099_),
    .S(_2494_),
    .X(_1851_));
 sky130_fd_sc_hd__mux2_1 _4741_ (.A0(_1115_),
    .A1(_1851_),
    .S(_1732_),
    .X(_1852_));
 sky130_fd_sc_hd__o21ai_1 _4742_ (.A1(\as1802.regs[2][11] ),
    .A2(_1752_),
    .B1(_1764_),
    .Y(_1853_));
 sky130_fd_sc_hd__o211a_1 _4743_ (.A1(_1764_),
    .A2(_1851_),
    .B1(_1853_),
    .C1(_1491_),
    .X(_1854_));
 sky130_fd_sc_hd__a21oi_1 _4744_ (.A1(_1496_),
    .A2(_1852_),
    .B1(_1854_),
    .Y(_1855_));
 sky130_fd_sc_hd__o22a_1 _4745_ (.A1(_1093_),
    .A2(_1783_),
    .B1(_1855_),
    .B2(_1750_),
    .X(_1856_));
 sky130_fd_sc_hd__nor2_1 _4746_ (.A(_1746_),
    .B(_1856_),
    .Y(_1857_));
 sky130_fd_sc_hd__a221o_1 _4747_ (.A1(_1745_),
    .A2(_1099_),
    .B1(_1746_),
    .B2(_1115_),
    .C1(_1727_),
    .X(_1858_));
 sky130_fd_sc_hd__a2bb2o_1 _4748_ (.A1_N(_1857_),
    .A2_N(_1858_),
    .B1(\as1802.addr_buff[11] ),
    .B2(_1728_),
    .X(_0262_));
 sky130_fd_sc_hd__mux2_1 _4749_ (.A0(_1155_),
    .A1(_1171_),
    .S(_1733_),
    .X(_1859_));
 sky130_fd_sc_hd__mux2_1 _4750_ (.A0(_1171_),
    .A1(_1859_),
    .S(_1732_),
    .X(_1860_));
 sky130_fd_sc_hd__o21ai_1 _4751_ (.A1(\as1802.regs[2][12] ),
    .A2(_1752_),
    .B1(_1740_),
    .Y(_1861_));
 sky130_fd_sc_hd__o211a_1 _4752_ (.A1(_1764_),
    .A2(_1859_),
    .B1(_1861_),
    .C1(_1766_),
    .X(_1862_));
 sky130_fd_sc_hd__a21oi_1 _4753_ (.A1(_1496_),
    .A2(_1860_),
    .B1(_1862_),
    .Y(_1863_));
 sky130_fd_sc_hd__a2bb2o_1 _4754_ (.A1_N(_1750_),
    .A2_N(_1863_),
    .B1(_1742_),
    .B2(_1155_),
    .X(_1864_));
 sky130_fd_sc_hd__a221o_1 _4755_ (.A1(_1745_),
    .A2(_1155_),
    .B1(_1171_),
    .B2(_1746_),
    .C1(_1726_),
    .X(_1865_));
 sky130_fd_sc_hd__a21oi_1 _4756_ (.A1(_1730_),
    .A2(_1864_),
    .B1(_1865_),
    .Y(_1866_));
 sky130_fd_sc_hd__a21o_1 _4757_ (.A1(\as1802.addr_buff[12] ),
    .A2(_1728_),
    .B1(_1866_),
    .X(_0263_));
 sky130_fd_sc_hd__mux2_1 _4758_ (.A0(_1211_),
    .A1(_1233_),
    .S(_1733_),
    .X(_1867_));
 sky130_fd_sc_hd__mux2_1 _4759_ (.A0(_1233_),
    .A1(_1867_),
    .S(_1732_),
    .X(_1868_));
 sky130_fd_sc_hd__o21ai_1 _4760_ (.A1(\as1802.regs[2][13] ),
    .A2(_1741_),
    .B1(_1740_),
    .Y(_1869_));
 sky130_fd_sc_hd__o211a_1 _4761_ (.A1(_1764_),
    .A2(_1867_),
    .B1(_1869_),
    .C1(_1766_),
    .X(_1870_));
 sky130_fd_sc_hd__a21o_1 _4762_ (.A1(_1496_),
    .A2(_1868_),
    .B1(_1870_),
    .X(_1871_));
 sky130_fd_sc_hd__a22o_1 _4763_ (.A1(_1211_),
    .A2(_1742_),
    .B1(_1871_),
    .B2(_1731_),
    .X(_1872_));
 sky130_fd_sc_hd__a221o_1 _4764_ (.A1(_1745_),
    .A2(_1211_),
    .B1(_1233_),
    .B2(_1746_),
    .C1(_1726_),
    .X(_1873_));
 sky130_fd_sc_hd__a21oi_1 _4765_ (.A1(_1730_),
    .A2(_1872_),
    .B1(_1873_),
    .Y(_1874_));
 sky130_fd_sc_hd__a21o_1 _4766_ (.A1(\as1802.addr_buff[13] ),
    .A2(_1728_),
    .B1(_1874_),
    .X(_0264_));
 sky130_fd_sc_hd__mux2_1 _4767_ (.A0(_1265_),
    .A1(_1281_),
    .S(_1733_),
    .X(_1875_));
 sky130_fd_sc_hd__mux2_1 _4768_ (.A0(_1281_),
    .A1(_1875_),
    .S(_1732_),
    .X(_1876_));
 sky130_fd_sc_hd__o21ai_1 _4769_ (.A1(\as1802.regs[2][14] ),
    .A2(_1741_),
    .B1(_1740_),
    .Y(_1877_));
 sky130_fd_sc_hd__o211a_1 _4770_ (.A1(_1764_),
    .A2(_1875_),
    .B1(_1877_),
    .C1(_1766_),
    .X(_1878_));
 sky130_fd_sc_hd__a21o_1 _4771_ (.A1(_1495_),
    .A2(_1876_),
    .B1(_1878_),
    .X(_1879_));
 sky130_fd_sc_hd__a22o_1 _4772_ (.A1(_1265_),
    .A2(_1742_),
    .B1(_1879_),
    .B2(_1731_),
    .X(_1880_));
 sky130_fd_sc_hd__a221o_1 _4773_ (.A1(_1745_),
    .A2(_1265_),
    .B1(_1281_),
    .B2(_1475_),
    .C1(_1726_),
    .X(_1881_));
 sky130_fd_sc_hd__a21oi_1 _4774_ (.A1(_1730_),
    .A2(_1880_),
    .B1(_1881_),
    .Y(_1882_));
 sky130_fd_sc_hd__a21o_1 _4775_ (.A1(\as1802.addr_buff[14] ),
    .A2(_1728_),
    .B1(_1882_),
    .X(_0265_));
 sky130_fd_sc_hd__mux2_1 _4776_ (.A0(_1316_),
    .A1(_1334_),
    .S(_1733_),
    .X(_1883_));
 sky130_fd_sc_hd__o21ai_1 _4777_ (.A1(\as1802.regs[2][15] ),
    .A2(_1752_),
    .B1(_1764_),
    .Y(_1884_));
 sky130_fd_sc_hd__o211a_1 _4778_ (.A1(_1764_),
    .A2(_1883_),
    .B1(_1884_),
    .C1(_1766_),
    .X(_1885_));
 sky130_fd_sc_hd__nand2_1 _4779_ (.A(_2480_),
    .B(_1333_),
    .Y(_1886_));
 sky130_fd_sc_hd__o211a_1 _4780_ (.A1(_2480_),
    .A2(_1883_),
    .B1(_1886_),
    .C1(_1495_),
    .X(_1887_));
 sky130_fd_sc_hd__nor2_1 _4781_ (.A(_1885_),
    .B(_1887_),
    .Y(_1888_));
 sky130_fd_sc_hd__o22a_1 _4782_ (.A1(_1317_),
    .A2(_1783_),
    .B1(_1888_),
    .B2(_1750_),
    .X(_1889_));
 sky130_fd_sc_hd__nor2_1 _4783_ (.A(_1746_),
    .B(_1889_),
    .Y(_1890_));
 sky130_fd_sc_hd__a221o_1 _4784_ (.A1(_1745_),
    .A2(_1316_),
    .B1(_1334_),
    .B2(_1746_),
    .C1(_1727_),
    .X(_1891_));
 sky130_fd_sc_hd__a2bb2o_1 _4785_ (.A1_N(_1890_),
    .A2_N(_1891_),
    .B1(\as1802.addr_buff[15] ),
    .B2(_1728_),
    .X(_0266_));
 sky130_fd_sc_hd__inv_2 _4786_ (.A(\as1802.mem_cycle[2] ),
    .Y(_1892_));
 sky130_fd_sc_hd__nand2_2 _4787_ (.A(_1892_),
    .B(\as1802.mem_cycle[0] ),
    .Y(_1893_));
 sky130_fd_sc_hd__mux2_1 _4788_ (.A0(\as1802.addr_buff[8] ),
    .A1(\as1802.addr_buff[0] ),
    .S(_1686_),
    .X(_1894_));
 sky130_fd_sc_hd__or2_1 _4789_ (.A(io_out[13]),
    .B(_1689_),
    .X(_1895_));
 sky130_fd_sc_hd__o211a_1 _4790_ (.A1(_1893_),
    .A2(_1894_),
    .B1(_1895_),
    .C1(_1494_),
    .X(_0267_));
 sky130_fd_sc_hd__mux2_1 _4791_ (.A0(\as1802.addr_buff[9] ),
    .A1(\as1802.addr_buff[1] ),
    .S(_1686_),
    .X(_1896_));
 sky130_fd_sc_hd__or2_1 _4792_ (.A(io_out[14]),
    .B(_1689_),
    .X(_1897_));
 sky130_fd_sc_hd__o211a_1 _4793_ (.A1(_1893_),
    .A2(_1896_),
    .B1(_1897_),
    .C1(_1494_),
    .X(_0268_));
 sky130_fd_sc_hd__mux2_1 _4794_ (.A0(\as1802.addr_buff[10] ),
    .A1(\as1802.addr_buff[2] ),
    .S(_1686_),
    .X(_1898_));
 sky130_fd_sc_hd__or2_1 _4795_ (.A(io_out[15]),
    .B(_1689_),
    .X(_1899_));
 sky130_fd_sc_hd__o211a_1 _4796_ (.A1(_1893_),
    .A2(_1898_),
    .B1(_1899_),
    .C1(_1494_),
    .X(_0269_));
 sky130_fd_sc_hd__mux2_1 _4797_ (.A0(\as1802.addr_buff[11] ),
    .A1(\as1802.addr_buff[3] ),
    .S(_1686_),
    .X(_1900_));
 sky130_fd_sc_hd__or2_1 _4798_ (.A(io_out[16]),
    .B(_1689_),
    .X(_1901_));
 sky130_fd_sc_hd__o211a_1 _4799_ (.A1(_1893_),
    .A2(_1900_),
    .B1(_1901_),
    .C1(_1494_),
    .X(_0270_));
 sky130_fd_sc_hd__mux2_1 _4800_ (.A0(\as1802.addr_buff[12] ),
    .A1(\as1802.addr_buff[4] ),
    .S(_1686_),
    .X(_1902_));
 sky130_fd_sc_hd__or2_1 _4801_ (.A(io_out[17]),
    .B(_1689_),
    .X(_1903_));
 sky130_fd_sc_hd__o211a_1 _4802_ (.A1(_1893_),
    .A2(_1902_),
    .B1(_1903_),
    .C1(_1494_),
    .X(_0271_));
 sky130_fd_sc_hd__mux2_1 _4803_ (.A0(\as1802.addr_buff[13] ),
    .A1(\as1802.addr_buff[5] ),
    .S(_1686_),
    .X(_1904_));
 sky130_fd_sc_hd__or2_1 _4804_ (.A(io_out[18]),
    .B(_1689_),
    .X(_1905_));
 sky130_fd_sc_hd__o211a_1 _4805_ (.A1(_1893_),
    .A2(_1904_),
    .B1(_1905_),
    .C1(_2458_),
    .X(_0272_));
 sky130_fd_sc_hd__mux2_1 _4806_ (.A0(\as1802.addr_buff[14] ),
    .A1(\as1802.addr_buff[6] ),
    .S(_1686_),
    .X(_1906_));
 sky130_fd_sc_hd__or2_1 _4807_ (.A(io_out[19]),
    .B(_1689_),
    .X(_1907_));
 sky130_fd_sc_hd__o211a_1 _4808_ (.A1(_1893_),
    .A2(_1906_),
    .B1(_1907_),
    .C1(_2458_),
    .X(_0273_));
 sky130_fd_sc_hd__mux2_1 _4809_ (.A0(\as1802.addr_buff[15] ),
    .A1(\as1802.addr_buff[7] ),
    .S(_1685_),
    .X(_1908_));
 sky130_fd_sc_hd__or2_1 _4810_ (.A(io_out[20]),
    .B(_1688_),
    .X(_1909_));
 sky130_fd_sc_hd__o211a_1 _4811_ (.A1(_1893_),
    .A2(_1908_),
    .B1(_1909_),
    .C1(_2458_),
    .X(_0274_));
 sky130_fd_sc_hd__or2_1 _4812_ (.A(\as1802.mem_cycle[1] ),
    .B(_1687_),
    .X(_1910_));
 sky130_fd_sc_hd__or2_2 _4813_ (.A(_1892_),
    .B(_1910_),
    .X(_1911_));
 sky130_fd_sc_hd__or3b_1 _4814_ (.A(\as1802.mem_write ),
    .B(_1911_),
    .C_N(_2482_),
    .X(_1912_));
 sky130_fd_sc_hd__nor2_4 _4815_ (.A(_2456_),
    .B(_1912_),
    .Y(_1913_));
 sky130_fd_sc_hd__mux2_1 _4816_ (.A0(_2469_),
    .A1(net1),
    .S(_1913_),
    .X(_1914_));
 sky130_fd_sc_hd__clkbuf_1 _4817_ (.A(_1914_),
    .X(_0275_));
 sky130_fd_sc_hd__mux2_1 _4818_ (.A0(_2504_),
    .A1(net5),
    .S(_1913_),
    .X(_1915_));
 sky130_fd_sc_hd__clkbuf_1 _4819_ (.A(_1915_),
    .X(_0276_));
 sky130_fd_sc_hd__mux2_1 _4820_ (.A0(_2496_),
    .A1(net6),
    .S(_1913_),
    .X(_1916_));
 sky130_fd_sc_hd__clkbuf_1 _4821_ (.A(_1916_),
    .X(_0277_));
 sky130_fd_sc_hd__mux2_1 _4822_ (.A0(_1733_),
    .A1(net7),
    .S(_1913_),
    .X(_1917_));
 sky130_fd_sc_hd__clkbuf_1 _4823_ (.A(_1917_),
    .X(_0278_));
 sky130_fd_sc_hd__mux2_1 _4824_ (.A0(_2474_),
    .A1(net8),
    .S(_1913_),
    .X(_1918_));
 sky130_fd_sc_hd__clkbuf_1 _4825_ (.A(_1918_),
    .X(_0279_));
 sky130_fd_sc_hd__mux2_1 _4826_ (.A0(_2473_),
    .A1(net9),
    .S(_1913_),
    .X(_1919_));
 sky130_fd_sc_hd__clkbuf_1 _4827_ (.A(_1919_),
    .X(_0280_));
 sky130_fd_sc_hd__mux2_1 _4828_ (.A0(_2477_),
    .A1(net10),
    .S(_1913_),
    .X(_1920_));
 sky130_fd_sc_hd__clkbuf_1 _4829_ (.A(_1920_),
    .X(_0281_));
 sky130_fd_sc_hd__mux2_1 _4830_ (.A0(_2476_),
    .A1(net11),
    .S(_1913_),
    .X(_1921_));
 sky130_fd_sc_hd__clkbuf_1 _4831_ (.A(_1921_),
    .X(_0282_));
 sky130_fd_sc_hd__nor2_4 _4832_ (.A(\as1802.mem_cycle[2] ),
    .B(_1910_),
    .Y(_1922_));
 sky130_fd_sc_hd__mux2_1 _4833_ (.A0(_1675_),
    .A1(_1680_),
    .S(_1922_),
    .X(_1923_));
 sky130_fd_sc_hd__nand2_1 _4834_ (.A(_1494_),
    .B(_1923_),
    .Y(_0283_));
 sky130_fd_sc_hd__mux2_1 _4835_ (.A0(\as1802.last_hi_addr[1] ),
    .A1(\as1802.addr_buff[9] ),
    .S(_1922_),
    .X(_1924_));
 sky130_fd_sc_hd__or2_1 _4836_ (.A(_1499_),
    .B(_1924_),
    .X(_1925_));
 sky130_fd_sc_hd__clkbuf_1 _4837_ (.A(_1925_),
    .X(_0284_));
 sky130_fd_sc_hd__mux2_1 _4838_ (.A0(\as1802.last_hi_addr[2] ),
    .A1(\as1802.addr_buff[10] ),
    .S(_1922_),
    .X(_1926_));
 sky130_fd_sc_hd__or2_1 _4839_ (.A(_1499_),
    .B(_1926_),
    .X(_1927_));
 sky130_fd_sc_hd__clkbuf_1 _4840_ (.A(_1927_),
    .X(_0285_));
 sky130_fd_sc_hd__mux2_1 _4841_ (.A0(\as1802.last_hi_addr[3] ),
    .A1(\as1802.addr_buff[11] ),
    .S(_1922_),
    .X(_1928_));
 sky130_fd_sc_hd__or2_1 _4842_ (.A(_1499_),
    .B(_1928_),
    .X(_1929_));
 sky130_fd_sc_hd__clkbuf_1 _4843_ (.A(_1929_),
    .X(_0286_));
 sky130_fd_sc_hd__mux2_1 _4844_ (.A0(\as1802.last_hi_addr[4] ),
    .A1(\as1802.addr_buff[12] ),
    .S(_1922_),
    .X(_1930_));
 sky130_fd_sc_hd__or2_1 _4845_ (.A(_1499_),
    .B(_1930_),
    .X(_1931_));
 sky130_fd_sc_hd__clkbuf_1 _4846_ (.A(_1931_),
    .X(_0287_));
 sky130_fd_sc_hd__mux2_1 _4847_ (.A0(_1671_),
    .A1(_1674_),
    .S(_1922_),
    .X(_1932_));
 sky130_fd_sc_hd__nand2_1 _4848_ (.A(_1494_),
    .B(_1932_),
    .Y(_0288_));
 sky130_fd_sc_hd__mux2_1 _4849_ (.A0(\as1802.last_hi_addr[6] ),
    .A1(\as1802.addr_buff[14] ),
    .S(_1922_),
    .X(_1933_));
 sky130_fd_sc_hd__or2_1 _4850_ (.A(_2456_),
    .B(_1933_),
    .X(_1934_));
 sky130_fd_sc_hd__clkbuf_1 _4851_ (.A(_1934_),
    .X(_0289_));
 sky130_fd_sc_hd__mux2_1 _4852_ (.A0(_1679_),
    .A1(_1670_),
    .S(_1922_),
    .X(_1935_));
 sky130_fd_sc_hd__nand2_1 _4853_ (.A(_1494_),
    .B(_1935_),
    .Y(_0290_));
 sky130_fd_sc_hd__a41o_1 _4854_ (.A1(_1489_),
    .A2(\as1802.IE ),
    .A3(net12),
    .A4(_2548_),
    .B1(\as1802.will_interrupt ),
    .X(_1936_));
 sky130_fd_sc_hd__and2b_1 _4855_ (.A_N(_1694_),
    .B(_1936_),
    .X(_1937_));
 sky130_fd_sc_hd__clkbuf_1 _4856_ (.A(_1937_),
    .X(_0291_));
 sky130_fd_sc_hd__a31o_1 _4857_ (.A1(_2464_),
    .A2(_2525_),
    .A3(_1729_),
    .B1(_1477_),
    .X(_1938_));
 sky130_fd_sc_hd__nor2_1 _4858_ (.A(_1473_),
    .B(_1938_),
    .Y(_1939_));
 sky130_fd_sc_hd__a21boi_1 _4859_ (.A1(_1483_),
    .A2(_1939_),
    .B1_N(\as1802.IE ),
    .Y(_1940_));
 sky130_fd_sc_hd__a311o_1 _4860_ (.A1(_0449_),
    .A2(_1483_),
    .A3(_1939_),
    .B1(_1940_),
    .C1(_1499_),
    .X(_0292_));
 sky130_fd_sc_hd__nand2_1 _4861_ (.A(_1476_),
    .B(_1699_),
    .Y(_1941_));
 sky130_fd_sc_hd__and3_1 _4862_ (.A(_2547_),
    .B(_1479_),
    .C(_1941_),
    .X(_1942_));
 sky130_fd_sc_hd__mux2_1 _4863_ (.A0(_2487_),
    .A1(_1489_),
    .S(_1942_),
    .X(_1943_));
 sky130_fd_sc_hd__nor2_1 _4864_ (.A(_1499_),
    .B(_1943_),
    .Y(_0293_));
 sky130_fd_sc_hd__or3_1 _4865_ (.A(_1892_),
    .B(\as1802.mem_cycle[1] ),
    .C(\as1802.mem_cycle[0] ),
    .X(_1944_));
 sky130_fd_sc_hd__nor2_1 _4866_ (.A(_1892_),
    .B(\as1802.mem_cycle[1] ),
    .Y(_1945_));
 sky130_fd_sc_hd__o22a_1 _4867_ (.A1(_1669_),
    .A2(_1944_),
    .B1(_1945_),
    .B2(io_oeb),
    .X(_1946_));
 sky130_fd_sc_hd__or2_1 _4868_ (.A(_2456_),
    .B(_1946_),
    .X(_1947_));
 sky130_fd_sc_hd__clkbuf_1 _4869_ (.A(_1947_),
    .X(_0294_));
 sky130_fd_sc_hd__a21oi_1 _4870_ (.A1(io_out[22]),
    .A2(_1910_),
    .B1(_1499_),
    .Y(_1948_));
 sky130_fd_sc_hd__nand2_1 _4871_ (.A(_1911_),
    .B(_1948_),
    .Y(_0295_));
 sky130_fd_sc_hd__o21a_1 _4872_ (.A1(\as1802.mem_cycle[1] ),
    .A2(\as1802.mem_cycle[0] ),
    .B1(_1892_),
    .X(_1949_));
 sky130_fd_sc_hd__o21ai_1 _4873_ (.A1(_1687_),
    .A2(_1718_),
    .B1(_1949_),
    .Y(_1950_));
 sky130_fd_sc_hd__o2bb2a_1 _4874_ (.A1_N(io_out[24]),
    .A2_N(_1950_),
    .B1(_1893_),
    .B2(_1686_),
    .X(_1951_));
 sky130_fd_sc_hd__nor2_1 _4875_ (.A(_1499_),
    .B(_1951_),
    .Y(_0296_));
 sky130_fd_sc_hd__and3_1 _4876_ (.A(_2504_),
    .B(_2503_),
    .C(_1733_),
    .X(_1952_));
 sky130_fd_sc_hd__and3_1 _4877_ (.A(_1491_),
    .B(_1691_),
    .C(_1952_),
    .X(_1953_));
 sky130_fd_sc_hd__mux2_1 _4878_ (.A0(_2501_),
    .A1(_2513_),
    .S(_1953_),
    .X(_1954_));
 sky130_fd_sc_hd__nor2_1 _4879_ (.A(_1499_),
    .B(_1954_),
    .Y(_0297_));
 sky130_fd_sc_hd__and3_1 _4880_ (.A(_1732_),
    .B(_1495_),
    .C(_2516_),
    .X(_1955_));
 sky130_fd_sc_hd__o31a_1 _4881_ (.A1(_1474_),
    .A2(_2572_),
    .A3(_1955_),
    .B1(_1730_),
    .X(_1956_));
 sky130_fd_sc_hd__nor2_1 _4882_ (.A(_1707_),
    .B(_1482_),
    .Y(_1957_));
 sky130_fd_sc_hd__nand2_2 _4883_ (.A(_2474_),
    .B(_2563_),
    .Y(_1958_));
 sky130_fd_sc_hd__nor2_1 _4884_ (.A(_2581_),
    .B(_1958_),
    .Y(_1959_));
 sky130_fd_sc_hd__or4_1 _4885_ (.A(_2708_),
    .B(_1957_),
    .C(_1724_),
    .D(_1959_),
    .X(_1960_));
 sky130_fd_sc_hd__or3_1 _4886_ (.A(_1710_),
    .B(_1719_),
    .C(_1960_),
    .X(_1961_));
 sky130_fd_sc_hd__mux2_1 _4887_ (.A0(_1956_),
    .A1(\as1802.lda ),
    .S(_1961_),
    .X(_1962_));
 sky130_fd_sc_hd__clkbuf_1 _4888_ (.A(_1962_),
    .X(_0298_));
 sky130_fd_sc_hd__inv_2 _4889_ (.A(\as1802.DF ),
    .Y(_1963_));
 sky130_fd_sc_hd__nand2_1 _4890_ (.A(_2477_),
    .B(_2496_),
    .Y(_1964_));
 sky130_fd_sc_hd__a2111o_1 _4891_ (.A1(_2482_),
    .A2(_2497_),
    .B1(_2610_),
    .C1(_1964_),
    .D1(_2521_),
    .X(_1965_));
 sky130_fd_sc_hd__o21a_1 _4892_ (.A1(_1288_),
    .A2(_2500_),
    .B1(_2496_),
    .X(_1966_));
 sky130_fd_sc_hd__or2_1 _4893_ (.A(_0840_),
    .B(io_out[7]),
    .X(_1967_));
 sky130_fd_sc_hd__nor2b_2 _4894_ (.A(_0797_),
    .B_N(io_out[6]),
    .Y(_1968_));
 sky130_fd_sc_hd__and2_1 _4895_ (.A(_0840_),
    .B(io_out[7]),
    .X(_1969_));
 sky130_fd_sc_hd__a21oi_1 _4896_ (.A1(_1967_),
    .A2(_1968_),
    .B1(_1969_),
    .Y(_1970_));
 sky130_fd_sc_hd__nor2_1 _4897_ (.A(_0840_),
    .B(io_out[7]),
    .Y(_1971_));
 sky130_fd_sc_hd__nor2_2 _4898_ (.A(_1971_),
    .B(_1969_),
    .Y(_1972_));
 sky130_fd_sc_hd__nand2_1 _4899_ (.A(_1968_),
    .B(_1972_),
    .Y(_1973_));
 sky130_fd_sc_hd__or2_1 _4900_ (.A(_1968_),
    .B(_1972_),
    .X(_1974_));
 sky130_fd_sc_hd__nand2b_2 _4901_ (.A_N(_0716_),
    .B(io_out[5]),
    .Y(_1975_));
 sky130_fd_sc_hd__nor2b_2 _4902_ (.A(io_out[6]),
    .B_N(\as1802.D[6] ),
    .Y(_1976_));
 sky130_fd_sc_hd__or2_1 _4903_ (.A(_1976_),
    .B(_1968_),
    .X(_1977_));
 sky130_fd_sc_hd__buf_2 _4904_ (.A(_1977_),
    .X(_1978_));
 sky130_fd_sc_hd__nor2_1 _4905_ (.A(_1975_),
    .B(_1978_),
    .Y(_1979_));
 sky130_fd_sc_hd__nand2b_2 _4906_ (.A_N(io_out[5]),
    .B(_0716_),
    .Y(_1980_));
 sky130_fd_sc_hd__and2_1 _4907_ (.A(_1975_),
    .B(_1980_),
    .X(_1981_));
 sky130_fd_sc_hd__buf_2 _4908_ (.A(_1981_),
    .X(_1982_));
 sky130_fd_sc_hd__nor2b_2 _4909_ (.A(_0646_),
    .B_N(io_out[4]),
    .Y(_1983_));
 sky130_fd_sc_hd__nand2_1 _4910_ (.A(_1982_),
    .B(_1983_),
    .Y(_1984_));
 sky130_fd_sc_hd__and2b_1 _4911_ (.A_N(io_out[4]),
    .B(\as1802.D[4] ),
    .X(_1985_));
 sky130_fd_sc_hd__clkbuf_2 _4912_ (.A(_1985_),
    .X(_1986_));
 sky130_fd_sc_hd__or2_1 _4913_ (.A(_1983_),
    .B(_1986_),
    .X(_1987_));
 sky130_fd_sc_hd__buf_2 _4914_ (.A(_1987_),
    .X(_1988_));
 sky130_fd_sc_hd__nand2b_2 _4915_ (.A_N(_0579_),
    .B(io_out[3]),
    .Y(_1989_));
 sky130_fd_sc_hd__nor2_1 _4916_ (.A(_1988_),
    .B(_1989_),
    .Y(_1990_));
 sky130_fd_sc_hd__nand2b_2 _4917_ (.A_N(io_out[3]),
    .B(_0579_),
    .Y(_1991_));
 sky130_fd_sc_hd__nand2_1 _4918_ (.A(_1989_),
    .B(_1991_),
    .Y(_1992_));
 sky130_fd_sc_hd__buf_2 _4919_ (.A(_1992_),
    .X(_1993_));
 sky130_fd_sc_hd__or2_2 _4920_ (.A(_0539_),
    .B(_0527_),
    .X(_1994_));
 sky130_fd_sc_hd__nor2_1 _4921_ (.A(_1993_),
    .B(_1994_),
    .Y(_1995_));
 sky130_fd_sc_hd__nand2_2 _4922_ (.A(_0539_),
    .B(_0527_),
    .Y(_1996_));
 sky130_fd_sc_hd__nand2_4 _4923_ (.A(_1994_),
    .B(_1996_),
    .Y(_1997_));
 sky130_fd_sc_hd__or2_1 _4924_ (.A(_0452_),
    .B(_1997_),
    .X(_1998_));
 sky130_fd_sc_hd__or2b_1 _4925_ (.A(\as1802.DF ),
    .B_N(\as1802.D[0] ),
    .X(_1999_));
 sky130_fd_sc_hd__and2b_1 _4926_ (.A_N(\as1802.D[0] ),
    .B(\as1802.DF ),
    .X(_2000_));
 sky130_fd_sc_hd__a21o_1 _4927_ (.A1(_2702_),
    .A2(_1999_),
    .B1(_2000_),
    .X(_2001_));
 sky130_fd_sc_hd__xor2_1 _4928_ (.A(\as1802.D[1] ),
    .B(_2001_),
    .X(_2002_));
 sky130_fd_sc_hd__and2_1 _4929_ (.A(_0474_),
    .B(_2002_),
    .X(_2003_));
 sky130_fd_sc_hd__a21o_1 _4930_ (.A1(_0452_),
    .A2(_2001_),
    .B1(_2003_),
    .X(_2004_));
 sky130_fd_sc_hd__nand2_1 _4931_ (.A(_0452_),
    .B(_1997_),
    .Y(_2005_));
 sky130_fd_sc_hd__and2_1 _4932_ (.A(_1998_),
    .B(_2005_),
    .X(_2006_));
 sky130_fd_sc_hd__nand2_1 _4933_ (.A(_2004_),
    .B(_2006_),
    .Y(_2007_));
 sky130_fd_sc_hd__and2_1 _4934_ (.A(_1993_),
    .B(_1994_),
    .X(_2008_));
 sky130_fd_sc_hd__a211oi_2 _4935_ (.A1(_1998_),
    .A2(_2007_),
    .B1(_1995_),
    .C1(_2008_),
    .Y(_2009_));
 sky130_fd_sc_hd__and2_1 _4936_ (.A(_1988_),
    .B(_1989_),
    .X(_2010_));
 sky130_fd_sc_hd__or2_1 _4937_ (.A(_1990_),
    .B(_2010_),
    .X(_2011_));
 sky130_fd_sc_hd__o21ba_1 _4938_ (.A1(_1995_),
    .A2(_2009_),
    .B1_N(_2011_),
    .X(_2012_));
 sky130_fd_sc_hd__or2_1 _4939_ (.A(_1981_),
    .B(_1983_),
    .X(_2013_));
 sky130_fd_sc_hd__o211ai_2 _4940_ (.A1(_1990_),
    .A2(_2012_),
    .B1(_2013_),
    .C1(_1984_),
    .Y(_2014_));
 sky130_fd_sc_hd__and2_1 _4941_ (.A(_1975_),
    .B(_1978_),
    .X(_2015_));
 sky130_fd_sc_hd__a211oi_1 _4942_ (.A1(_1984_),
    .A2(_2014_),
    .B1(_1979_),
    .C1(_2015_),
    .Y(_2016_));
 sky130_fd_sc_hd__or2_1 _4943_ (.A(_1979_),
    .B(_2016_),
    .X(_2017_));
 sky130_fd_sc_hd__and3_1 _4944_ (.A(_1973_),
    .B(_1974_),
    .C(_2017_),
    .X(_2018_));
 sky130_fd_sc_hd__mux2_1 _4945_ (.A0(_1970_),
    .A1(_1969_),
    .S(_2018_),
    .X(_2019_));
 sky130_fd_sc_hd__or2_2 _4946_ (.A(_2503_),
    .B(_2505_),
    .X(_2020_));
 sky130_fd_sc_hd__or2b_1 _4947_ (.A(\as1802.D[1] ),
    .B_N(io_out[1]),
    .X(_2021_));
 sky130_fd_sc_hd__nand2b_2 _4948_ (.A_N(io_out[1]),
    .B(\as1802.D[1] ),
    .Y(_2022_));
 sky130_fd_sc_hd__nand2_1 _4949_ (.A(_2021_),
    .B(_2022_),
    .Y(_2023_));
 sky130_fd_sc_hd__inv_2 _4950_ (.A(io_out[0]),
    .Y(_2024_));
 sky130_fd_sc_hd__nor2_1 _4951_ (.A(_0382_),
    .B(_2024_),
    .Y(_2025_));
 sky130_fd_sc_hd__or2_1 _4952_ (.A(_2023_),
    .B(_2025_),
    .X(_2026_));
 sky130_fd_sc_hd__or2_2 _4953_ (.A(_1971_),
    .B(_1969_),
    .X(_2027_));
 sky130_fd_sc_hd__nand2_1 _4954_ (.A(_1975_),
    .B(_1980_),
    .Y(_2028_));
 sky130_fd_sc_hd__and2b_1 _4955_ (.A_N(_2702_),
    .B(_0382_),
    .X(_2029_));
 sky130_fd_sc_hd__or4_1 _4956_ (.A(_2028_),
    .B(_1988_),
    .C(_1993_),
    .D(_2029_),
    .X(_2030_));
 sky130_fd_sc_hd__or4_1 _4957_ (.A(_1997_),
    .B(_1978_),
    .C(_2027_),
    .D(_2030_),
    .X(_2031_));
 sky130_fd_sc_hd__inv_2 _4958_ (.A(_1976_),
    .Y(_2032_));
 sky130_fd_sc_hd__or2_1 _4959_ (.A(_2029_),
    .B(_2023_),
    .X(_2033_));
 sky130_fd_sc_hd__a21o_1 _4960_ (.A1(_2021_),
    .A2(_2033_),
    .B1(_1997_),
    .X(_2034_));
 sky130_fd_sc_hd__a21o_1 _4961_ (.A1(_1994_),
    .A2(_2034_),
    .B1(_1993_),
    .X(_2035_));
 sky130_fd_sc_hd__a21oi_1 _4962_ (.A1(_1989_),
    .A2(_2035_),
    .B1(_1988_),
    .Y(_2036_));
 sky130_fd_sc_hd__o21ai_1 _4963_ (.A1(_1983_),
    .A2(_2036_),
    .B1(_1981_),
    .Y(_2037_));
 sky130_fd_sc_hd__nand2_1 _4964_ (.A(_1975_),
    .B(_2037_),
    .Y(_2038_));
 sky130_fd_sc_hd__a21o_1 _4965_ (.A1(_2032_),
    .A2(_2038_),
    .B1(_1968_),
    .X(_2039_));
 sky130_fd_sc_hd__a21o_1 _4966_ (.A1(_1967_),
    .A2(_2039_),
    .B1(_1969_),
    .X(_2040_));
 sky130_fd_sc_hd__o21a_1 _4967_ (.A1(_2026_),
    .A2(_2031_),
    .B1(_2040_),
    .X(_2041_));
 sky130_fd_sc_hd__a2bb2o_1 _4968_ (.A1_N(_2020_),
    .A2_N(_2041_),
    .B1(_2040_),
    .B2(_2508_),
    .X(_2042_));
 sky130_fd_sc_hd__nand2_1 _4969_ (.A(\as1802.D[7] ),
    .B(io_out[7]),
    .Y(_2043_));
 sky130_fd_sc_hd__nand2_1 _4970_ (.A(_0797_),
    .B(io_out[6]),
    .Y(_2044_));
 sky130_fd_sc_hd__nand2_1 _4971_ (.A(_0716_),
    .B(io_out[5]),
    .Y(_2045_));
 sky130_fd_sc_hd__nand2_1 _4972_ (.A(_0646_),
    .B(io_out[4]),
    .Y(_2046_));
 sky130_fd_sc_hd__nand2_1 _4973_ (.A(_0579_),
    .B(io_out[3]),
    .Y(_2047_));
 sky130_fd_sc_hd__nand2_1 _4974_ (.A(_0539_),
    .B(io_out[2]),
    .Y(_2048_));
 sky130_fd_sc_hd__nand2_1 _4975_ (.A(\as1802.D[1] ),
    .B(_0474_),
    .Y(_2049_));
 sky130_fd_sc_hd__and2_1 _4976_ (.A(_2021_),
    .B(_2022_),
    .X(_2050_));
 sky130_fd_sc_hd__nand2_1 _4977_ (.A(_0382_),
    .B(_2702_),
    .Y(_2051_));
 sky130_fd_sc_hd__or2_1 _4978_ (.A(_2050_),
    .B(_2051_),
    .X(_2052_));
 sky130_fd_sc_hd__or2_1 _4979_ (.A(_0382_),
    .B(_2702_),
    .X(_2053_));
 sky130_fd_sc_hd__and2_1 _4980_ (.A(\as1802.DF ),
    .B(_2053_),
    .X(_2054_));
 sky130_fd_sc_hd__nand2_1 _4981_ (.A(_2023_),
    .B(_2054_),
    .Y(_2055_));
 sky130_fd_sc_hd__and2_1 _4982_ (.A(_1994_),
    .B(_1996_),
    .X(_2056_));
 sky130_fd_sc_hd__clkbuf_2 _4983_ (.A(_2056_),
    .X(_2057_));
 sky130_fd_sc_hd__a31o_1 _4984_ (.A1(_2049_),
    .A2(_2052_),
    .A3(_2055_),
    .B1(_2057_),
    .X(_2058_));
 sky130_fd_sc_hd__and2_1 _4985_ (.A(_1989_),
    .B(_1991_),
    .X(_2059_));
 sky130_fd_sc_hd__a21o_1 _4986_ (.A1(_2048_),
    .A2(_2058_),
    .B1(_2059_),
    .X(_2060_));
 sky130_fd_sc_hd__nor2_1 _4987_ (.A(_1983_),
    .B(_1986_),
    .Y(_2061_));
 sky130_fd_sc_hd__a21o_1 _4988_ (.A1(_2047_),
    .A2(_2060_),
    .B1(_2061_),
    .X(_2062_));
 sky130_fd_sc_hd__a21o_1 _4989_ (.A1(_2046_),
    .A2(_2062_),
    .B1(_1982_),
    .X(_2063_));
 sky130_fd_sc_hd__nor2_1 _4990_ (.A(_1976_),
    .B(_1968_),
    .Y(_2064_));
 sky130_fd_sc_hd__a21o_1 _4991_ (.A1(_2045_),
    .A2(_2063_),
    .B1(_2064_),
    .X(_2065_));
 sky130_fd_sc_hd__a21o_1 _4992_ (.A1(_2044_),
    .A2(_2065_),
    .B1(_1972_),
    .X(_2066_));
 sky130_fd_sc_hd__a21oi_1 _4993_ (.A1(_2043_),
    .A2(_2066_),
    .B1(_2557_),
    .Y(_2067_));
 sky130_fd_sc_hd__nand2_1 _4994_ (.A(_1976_),
    .B(_1972_),
    .Y(_2068_));
 sky130_fd_sc_hd__nor2_2 _4995_ (.A(_0453_),
    .B(_2020_),
    .Y(_2069_));
 sky130_fd_sc_hd__nor2_1 _4996_ (.A(_1980_),
    .B(_1978_),
    .Y(_2070_));
 sky130_fd_sc_hd__nand2_1 _4997_ (.A(_1982_),
    .B(_1986_),
    .Y(_2071_));
 sky130_fd_sc_hd__nor2_1 _4998_ (.A(_1988_),
    .B(_1991_),
    .Y(_2072_));
 sky130_fd_sc_hd__nor2_1 _4999_ (.A(_1993_),
    .B(_1996_),
    .Y(_2073_));
 sky130_fd_sc_hd__nor2_1 _5000_ (.A(_0474_),
    .B(_1997_),
    .Y(_2074_));
 sky130_fd_sc_hd__xnor2_1 _5001_ (.A(_0474_),
    .B(_2057_),
    .Y(_2075_));
 sky130_fd_sc_hd__nor2_1 _5002_ (.A(\as1802.D[1] ),
    .B(io_out[1]),
    .Y(_2076_));
 sky130_fd_sc_hd__nor2_1 _5003_ (.A(\as1802.DF ),
    .B(_2029_),
    .Y(_2077_));
 sky130_fd_sc_hd__or2_1 _5004_ (.A(_2025_),
    .B(_2077_),
    .X(_2078_));
 sky130_fd_sc_hd__o21ai_1 _5005_ (.A1(_2076_),
    .A2(_2078_),
    .B1(_2049_),
    .Y(_2079_));
 sky130_fd_sc_hd__and2_1 _5006_ (.A(_2075_),
    .B(_2079_),
    .X(_2080_));
 sky130_fd_sc_hd__and2_1 _5007_ (.A(_1992_),
    .B(_1996_),
    .X(_2081_));
 sky130_fd_sc_hd__nor2_1 _5008_ (.A(_2073_),
    .B(_2081_),
    .Y(_2082_));
 sky130_fd_sc_hd__o21a_1 _5009_ (.A1(_2074_),
    .A2(_2080_),
    .B1(_2082_),
    .X(_2083_));
 sky130_fd_sc_hd__inv_2 _5010_ (.A(_2072_),
    .Y(_2084_));
 sky130_fd_sc_hd__nand2_1 _5011_ (.A(_1988_),
    .B(_1991_),
    .Y(_2085_));
 sky130_fd_sc_hd__o211a_1 _5012_ (.A1(_2073_),
    .A2(_2083_),
    .B1(_2084_),
    .C1(_2085_),
    .X(_2086_));
 sky130_fd_sc_hd__xnor2_1 _5013_ (.A(_2028_),
    .B(_1986_),
    .Y(_2087_));
 sky130_fd_sc_hd__o21ai_2 _5014_ (.A1(_2072_),
    .A2(_2086_),
    .B1(_2087_),
    .Y(_2088_));
 sky130_fd_sc_hd__and2_1 _5015_ (.A(_1980_),
    .B(_1978_),
    .X(_2089_));
 sky130_fd_sc_hd__a211oi_2 _5016_ (.A1(_2071_),
    .A2(_2088_),
    .B1(_2070_),
    .C1(_2089_),
    .Y(_2090_));
 sky130_fd_sc_hd__nand2_1 _5017_ (.A(_2032_),
    .B(_2027_),
    .Y(_2091_));
 sky130_fd_sc_hd__o211a_1 _5018_ (.A1(_2070_),
    .A2(_2090_),
    .B1(_2068_),
    .C1(_2091_),
    .X(_2092_));
 sky130_fd_sc_hd__xnor2_1 _5019_ (.A(_1971_),
    .B(_2092_),
    .Y(_2093_));
 sky130_fd_sc_hd__nor2_4 _5020_ (.A(_2533_),
    .B(_2543_),
    .Y(_2094_));
 sky130_fd_sc_hd__nor2_4 _5021_ (.A(_2493_),
    .B(_2543_),
    .Y(_2095_));
 sky130_fd_sc_hd__a22o_1 _5022_ (.A1(_0382_),
    .A2(_2094_),
    .B1(_2095_),
    .B2(\as1802.D[7] ),
    .X(_2096_));
 sky130_fd_sc_hd__o21ai_4 _5023_ (.A1(_0453_),
    .A2(_2500_),
    .B1(_2496_),
    .Y(_2097_));
 sky130_fd_sc_hd__or2_1 _5024_ (.A(_2096_),
    .B(_2097_),
    .X(_2098_));
 sky130_fd_sc_hd__a31o_1 _5025_ (.A1(_2068_),
    .A2(_2069_),
    .A3(_2093_),
    .B1(_2098_),
    .X(_2099_));
 sky130_fd_sc_hd__a211o_1 _5026_ (.A1(_1733_),
    .A2(_2042_),
    .B1(_2067_),
    .C1(_2099_),
    .X(_2100_));
 sky130_fd_sc_hd__o211a_1 _5027_ (.A1(_1966_),
    .A2(_2019_),
    .B1(_2100_),
    .C1(_1491_),
    .X(_2101_));
 sky130_fd_sc_hd__inv_2 _5028_ (.A(_2048_),
    .Y(_2102_));
 sky130_fd_sc_hd__a21oi_1 _5029_ (.A1(_2049_),
    .A2(_2052_),
    .B1(_2057_),
    .Y(_2103_));
 sky130_fd_sc_hd__o21ai_1 _5030_ (.A1(_2102_),
    .A2(_2103_),
    .B1(_1993_),
    .Y(_2104_));
 sky130_fd_sc_hd__a21o_1 _5031_ (.A1(_2047_),
    .A2(_2104_),
    .B1(_2061_),
    .X(_2105_));
 sky130_fd_sc_hd__a21o_1 _5032_ (.A1(_2046_),
    .A2(_2105_),
    .B1(_1982_),
    .X(_2106_));
 sky130_fd_sc_hd__a21o_1 _5033_ (.A1(_2045_),
    .A2(_2106_),
    .B1(_2064_),
    .X(_2107_));
 sky130_fd_sc_hd__a21oi_1 _5034_ (.A1(_2044_),
    .A2(_2107_),
    .B1(_1972_),
    .Y(_2108_));
 sky130_fd_sc_hd__o21ai_1 _5035_ (.A1(_2503_),
    .A2(_2470_),
    .B1(_2043_),
    .Y(_2109_));
 sky130_fd_sc_hd__or4_1 _5036_ (.A(_2503_),
    .B(_2470_),
    .C(_2042_),
    .D(_2096_),
    .X(_2110_));
 sky130_fd_sc_hd__o211a_1 _5037_ (.A1(_2108_),
    .A2(_2109_),
    .B1(_1496_),
    .C1(_2110_),
    .X(_2111_));
 sky130_fd_sc_hd__o31a_1 _5038_ (.A1(_2101_),
    .A2(_2111_),
    .A3(_1965_),
    .B1(_2457_),
    .X(_2112_));
 sky130_fd_sc_hd__a21boi_1 _5039_ (.A1(_1963_),
    .A2(_1965_),
    .B1_N(_2112_),
    .Y(_0299_));
 sky130_fd_sc_hd__o32a_1 _5040_ (.A1(_2581_),
    .A2(_2567_),
    .A3(_2478_),
    .B1(_1737_),
    .B2(_1483_),
    .X(_2113_));
 sky130_fd_sc_hd__and2_1 _5041_ (.A(_1480_),
    .B(_2113_),
    .X(_2114_));
 sky130_fd_sc_hd__clkbuf_2 _5042_ (.A(_2114_),
    .X(_2115_));
 sky130_fd_sc_hd__mux2_1 _5043_ (.A0(\as1802.P[0] ),
    .A1(io_out[4]),
    .S(_1752_),
    .X(_2116_));
 sky130_fd_sc_hd__mux2_1 _5044_ (.A0(_2469_),
    .A1(_2116_),
    .S(_1491_),
    .X(_2117_));
 sky130_fd_sc_hd__a21bo_1 _5045_ (.A1(_2486_),
    .A2(_2117_),
    .B1_N(_2115_),
    .X(_2118_));
 sky130_fd_sc_hd__o211a_1 _5046_ (.A1(\as1802.X[0] ),
    .A2(_2115_),
    .B1(_2118_),
    .C1(_2458_),
    .X(_0300_));
 sky130_fd_sc_hd__mux2_1 _5047_ (.A0(\as1802.P[1] ),
    .A1(io_out[5]),
    .S(_1752_),
    .X(_2119_));
 sky130_fd_sc_hd__nand2_1 _5048_ (.A(_1491_),
    .B(_2119_),
    .Y(_2120_));
 sky130_fd_sc_hd__nand4_1 _5049_ (.A(_2486_),
    .B(_1497_),
    .C(_2115_),
    .D(_2120_),
    .Y(_2121_));
 sky130_fd_sc_hd__o211a_1 _5050_ (.A1(\as1802.X[1] ),
    .A2(_2115_),
    .B1(_2121_),
    .C1(_2458_),
    .X(_0301_));
 sky130_fd_sc_hd__mux2_1 _5051_ (.A0(\as1802.P[2] ),
    .A1(io_out[6]),
    .S(_1752_),
    .X(_2122_));
 sky130_fd_sc_hd__nor2_1 _5052_ (.A(_1496_),
    .B(_2122_),
    .Y(_2123_));
 sky130_fd_sc_hd__o31ai_1 _5053_ (.A1(_1489_),
    .A2(_1502_),
    .A3(_2123_),
    .B1(_2115_),
    .Y(_2124_));
 sky130_fd_sc_hd__o211a_1 _5054_ (.A1(\as1802.X[2] ),
    .A2(_2115_),
    .B1(_2124_),
    .C1(_2458_),
    .X(_0302_));
 sky130_fd_sc_hd__mux2_1 _5055_ (.A0(\as1802.P[3] ),
    .A1(io_out[7]),
    .S(_1741_),
    .X(_2125_));
 sky130_fd_sc_hd__o21a_1 _5056_ (.A1(_1495_),
    .A2(_2125_),
    .B1(_1505_),
    .X(_2126_));
 sky130_fd_sc_hd__mux2_1 _5057_ (.A0(\as1802.X[3] ),
    .A1(_2126_),
    .S(_2115_),
    .X(_2127_));
 sky130_fd_sc_hd__and2_1 _5058_ (.A(_1504_),
    .B(_2127_),
    .X(_2128_));
 sky130_fd_sc_hd__clkbuf_1 _5059_ (.A(_2128_),
    .X(_0303_));
 sky130_fd_sc_hd__o211a_4 _5060_ (.A1(_1738_),
    .A2(_1482_),
    .B1(_1939_),
    .C1(_1479_),
    .X(_2129_));
 sky130_fd_sc_hd__mux2_1 _5061_ (.A0(\as1802.T[0] ),
    .A1(\as1802.P[0] ),
    .S(_2129_),
    .X(_2130_));
 sky130_fd_sc_hd__and2_1 _5062_ (.A(_1504_),
    .B(_2130_),
    .X(_2131_));
 sky130_fd_sc_hd__clkbuf_1 _5063_ (.A(_2131_),
    .X(_0304_));
 sky130_fd_sc_hd__mux2_1 _5064_ (.A0(\as1802.T[1] ),
    .A1(\as1802.P[1] ),
    .S(_2129_),
    .X(_2132_));
 sky130_fd_sc_hd__and2_1 _5065_ (.A(_1504_),
    .B(_2132_),
    .X(_2133_));
 sky130_fd_sc_hd__clkbuf_1 _5066_ (.A(_2133_),
    .X(_0305_));
 sky130_fd_sc_hd__mux2_1 _5067_ (.A0(\as1802.T[2] ),
    .A1(\as1802.P[2] ),
    .S(_2129_),
    .X(_2134_));
 sky130_fd_sc_hd__and2_1 _5068_ (.A(_1504_),
    .B(_2134_),
    .X(_2135_));
 sky130_fd_sc_hd__clkbuf_1 _5069_ (.A(_2135_),
    .X(_0306_));
 sky130_fd_sc_hd__mux2_1 _5070_ (.A0(\as1802.T[3] ),
    .A1(\as1802.P[3] ),
    .S(_2129_),
    .X(_2136_));
 sky130_fd_sc_hd__and2_1 _5071_ (.A(_1504_),
    .B(_2136_),
    .X(_2137_));
 sky130_fd_sc_hd__clkbuf_1 _5072_ (.A(_2137_),
    .X(_0307_));
 sky130_fd_sc_hd__mux2_1 _5073_ (.A0(\as1802.T[4] ),
    .A1(\as1802.X[0] ),
    .S(_2129_),
    .X(_2138_));
 sky130_fd_sc_hd__and2_1 _5074_ (.A(_1504_),
    .B(_2138_),
    .X(_2139_));
 sky130_fd_sc_hd__clkbuf_1 _5075_ (.A(_2139_),
    .X(_0308_));
 sky130_fd_sc_hd__mux2_1 _5076_ (.A0(\as1802.T[5] ),
    .A1(\as1802.X[1] ),
    .S(_2129_),
    .X(_2140_));
 sky130_fd_sc_hd__and2_1 _5077_ (.A(_1504_),
    .B(_2140_),
    .X(_2141_));
 sky130_fd_sc_hd__clkbuf_1 _5078_ (.A(_2141_),
    .X(_0309_));
 sky130_fd_sc_hd__o21ai_1 _5079_ (.A1(\as1802.T[6] ),
    .A2(_2129_),
    .B1(_1504_),
    .Y(_2142_));
 sky130_fd_sc_hd__a21oi_1 _5080_ (.A1(_2634_),
    .A2(_2129_),
    .B1(_2142_),
    .Y(_0310_));
 sky130_fd_sc_hd__o21ai_1 _5081_ (.A1(\as1802.T[7] ),
    .A2(_2129_),
    .B1(_1504_),
    .Y(_2143_));
 sky130_fd_sc_hd__a21oi_1 _5082_ (.A1(_0436_),
    .A2(_2129_),
    .B1(_2143_),
    .Y(_0311_));
 sky130_fd_sc_hd__clkbuf_4 _5083_ (.A(_2612_),
    .X(_2144_));
 sky130_fd_sc_hd__nor3_4 _5084_ (.A(_2473_),
    .B(_2567_),
    .C(_2561_),
    .Y(_2145_));
 sky130_fd_sc_hd__nand2_1 _5085_ (.A(_0452_),
    .B(_2094_),
    .Y(_2146_));
 sky130_fd_sc_hd__nor2_1 _5086_ (.A(_2504_),
    .B(_2496_),
    .Y(_2147_));
 sky130_fd_sc_hd__o211a_1 _5087_ (.A1(_2051_),
    .A2(_2147_),
    .B1(_2053_),
    .C1(_2497_),
    .X(_2148_));
 sky130_fd_sc_hd__nor2_1 _5088_ (.A(_2145_),
    .B(_2148_),
    .Y(_2149_));
 sky130_fd_sc_hd__o211a_1 _5089_ (.A1(_2600_),
    .A2(_2051_),
    .B1(_2146_),
    .C1(_2149_),
    .X(_2150_));
 sky130_fd_sc_hd__a211o_1 _5090_ (.A1(_2145_),
    .A2(_0904_),
    .B1(_2150_),
    .C1(_2562_),
    .X(_2151_));
 sky130_fd_sc_hd__o211a_1 _5091_ (.A1(_2144_),
    .A2(_2665_),
    .B1(_2151_),
    .C1(_1495_),
    .X(_2152_));
 sky130_fd_sc_hd__a221o_1 _5092_ (.A1(_0452_),
    .A2(_2094_),
    .B1(_2095_),
    .B2(\as1802.DF ),
    .C1(_2554_),
    .X(_2153_));
 sky130_fd_sc_hd__clkbuf_4 _5093_ (.A(_2515_),
    .X(_2154_));
 sky130_fd_sc_hd__nand2_1 _5094_ (.A(_2702_),
    .B(_1999_),
    .Y(_2155_));
 sky130_fd_sc_hd__o22ai_1 _5095_ (.A1(_2077_),
    .A2(_2054_),
    .B1(_2000_),
    .B2(_2155_),
    .Y(_2156_));
 sky130_fd_sc_hd__mux2_1 _5096_ (.A0(_2514_),
    .A1(_2154_),
    .S(_2156_),
    .X(_2157_));
 sky130_fd_sc_hd__nor2_4 _5097_ (.A(_2461_),
    .B(_2569_),
    .Y(_2158_));
 sky130_fd_sc_hd__o21ai_1 _5098_ (.A1(_2153_),
    .A2(_2157_),
    .B1(_2158_),
    .Y(_2159_));
 sky130_fd_sc_hd__a2bb2o_1 _5099_ (.A1_N(_2152_),
    .A2_N(_2159_),
    .B1(net1),
    .B2(_2462_),
    .X(_2160_));
 sky130_fd_sc_hd__o311a_1 _5100_ (.A1(_2581_),
    .A2(_1720_),
    .A3(_0448_),
    .B1(_1472_),
    .C1(_2705_),
    .X(_2161_));
 sky130_fd_sc_hd__a21oi_1 _5101_ (.A1(_2494_),
    .A2(_2466_),
    .B1(_2516_),
    .Y(_2162_));
 sky130_fd_sc_hd__or4_1 _5102_ (.A(_2580_),
    .B(_1720_),
    .C(_2602_),
    .D(_2162_),
    .X(_2163_));
 sky130_fd_sc_hd__a21oi_1 _5103_ (.A1(_2545_),
    .A2(_1484_),
    .B1(_1959_),
    .Y(_2164_));
 sky130_fd_sc_hd__o211a_1 _5104_ (.A1(_2496_),
    .A2(_1482_),
    .B1(_2163_),
    .C1(_2164_),
    .X(_2165_));
 sky130_fd_sc_hd__a31o_1 _5105_ (.A1(_0444_),
    .A2(_2161_),
    .A3(_2165_),
    .B1(_2461_),
    .X(_2166_));
 sky130_fd_sc_hd__or3_1 _5106_ (.A(_2482_),
    .B(\as1802.mem_write ),
    .C(_1911_),
    .X(_2167_));
 sky130_fd_sc_hd__a21o_1 _5107_ (.A1(_2486_),
    .A2(_2583_),
    .B1(_2460_),
    .X(_2168_));
 sky130_fd_sc_hd__and2_1 _5108_ (.A(_1912_),
    .B(_2168_),
    .X(_2169_));
 sky130_fd_sc_hd__o221a_1 _5109_ (.A1(_2524_),
    .A2(_2699_),
    .B1(_2167_),
    .B2(\as1802.lda ),
    .C1(_2169_),
    .X(_2170_));
 sky130_fd_sc_hd__a211o_1 _5110_ (.A1(\as1802.mem_cycle[0] ),
    .A2(\as1802.mem_write ),
    .B1(_2456_),
    .C1(\as1802.mem_cycle[1] ),
    .X(_2171_));
 sky130_fd_sc_hd__or3b_1 _5111_ (.A(_2171_),
    .B(_1949_),
    .C_N(_1944_),
    .X(_2172_));
 sky130_fd_sc_hd__a311oi_1 _5112_ (.A1(_2549_),
    .A2(_2463_),
    .A3(_1691_),
    .B1(_1692_),
    .C1(_2172_),
    .Y(_2173_));
 sky130_fd_sc_hd__and4_1 _5113_ (.A(_0385_),
    .B(_1701_),
    .C(_2170_),
    .D(_2173_),
    .X(_2174_));
 sky130_fd_sc_hd__nand2_4 _5114_ (.A(_2166_),
    .B(_2174_),
    .Y(_2175_));
 sky130_fd_sc_hd__mux2_1 _5115_ (.A0(_2160_),
    .A1(_0382_),
    .S(_2175_),
    .X(_2176_));
 sky130_fd_sc_hd__clkbuf_1 _5116_ (.A(_2176_),
    .X(_0312_));
 sky130_fd_sc_hd__a22o_1 _5117_ (.A1(_0539_),
    .A2(_2094_),
    .B1(_2095_),
    .B2(_0382_),
    .X(_2177_));
 sky130_fd_sc_hd__nand2_1 _5118_ (.A(_2050_),
    .B(_2051_),
    .Y(_2178_));
 sky130_fd_sc_hd__and3_1 _5119_ (.A(_2515_),
    .B(_2052_),
    .C(_2178_),
    .X(_2179_));
 sky130_fd_sc_hd__nand2_1 _5120_ (.A(_2023_),
    .B(_2025_),
    .Y(_2180_));
 sky130_fd_sc_hd__nand2_1 _5121_ (.A(_2029_),
    .B(_2023_),
    .Y(_2181_));
 sky130_fd_sc_hd__and3_1 _5122_ (.A(_2508_),
    .B(_2033_),
    .C(_2181_),
    .X(_2182_));
 sky130_fd_sc_hd__a31o_1 _5123_ (.A1(_2506_),
    .A2(_2026_),
    .A3(_2180_),
    .B1(_2182_),
    .X(_2183_));
 sky130_fd_sc_hd__or2_1 _5124_ (.A(_2504_),
    .B(_2495_),
    .X(_2184_));
 sky130_fd_sc_hd__clkbuf_4 _5125_ (.A(_2184_),
    .X(_2185_));
 sky130_fd_sc_hd__or2_1 _5126_ (.A(_2600_),
    .B(_2049_),
    .X(_2186_));
 sky130_fd_sc_hd__o221a_1 _5127_ (.A1(_2511_),
    .A2(_2050_),
    .B1(_2076_),
    .B2(_2185_),
    .C1(_2186_),
    .X(_2187_));
 sky130_fd_sc_hd__or4b_1 _5128_ (.A(_2177_),
    .B(_2179_),
    .C(_2183_),
    .D_N(_2187_),
    .X(_2188_));
 sky130_fd_sc_hd__mux2_1 _5129_ (.A0(_1034_),
    .A1(_2188_),
    .S(_1695_),
    .X(_2189_));
 sky130_fd_sc_hd__nor2_1 _5130_ (.A(_2144_),
    .B(_0439_),
    .Y(_2190_));
 sky130_fd_sc_hd__a211o_1 _5131_ (.A1(_2144_),
    .A2(_2189_),
    .B1(_2190_),
    .C1(_1766_),
    .X(_2191_));
 sky130_fd_sc_hd__nor2_1 _5132_ (.A(_0474_),
    .B(_2002_),
    .Y(_2192_));
 sky130_fd_sc_hd__or2_1 _5133_ (.A(_2003_),
    .B(_2192_),
    .X(_2193_));
 sky130_fd_sc_hd__inv_2 _5134_ (.A(_2508_),
    .Y(_2194_));
 sky130_fd_sc_hd__nor2_2 _5135_ (.A(_2494_),
    .B(_2194_),
    .Y(_2195_));
 sky130_fd_sc_hd__nor2_4 _5136_ (.A(_2493_),
    .B(_2020_),
    .Y(_2196_));
 sky130_fd_sc_hd__or2_1 _5137_ (.A(_2023_),
    .B(_2078_),
    .X(_2197_));
 sky130_fd_sc_hd__nand2_1 _5138_ (.A(_2023_),
    .B(_2078_),
    .Y(_2198_));
 sky130_fd_sc_hd__and2_1 _5139_ (.A(_2197_),
    .B(_2198_),
    .X(_2199_));
 sky130_fd_sc_hd__mux2_1 _5140_ (.A0(_2069_),
    .A1(_2196_),
    .S(_2199_),
    .X(_2200_));
 sky130_fd_sc_hd__and3_1 _5141_ (.A(_2154_),
    .B(_2052_),
    .C(_2055_),
    .X(_2201_));
 sky130_fd_sc_hd__o21a_1 _5142_ (.A1(_2054_),
    .A2(_2178_),
    .B1(_2201_),
    .X(_2202_));
 sky130_fd_sc_hd__or4_1 _5143_ (.A(_2554_),
    .B(_2177_),
    .C(_2200_),
    .D(_2202_),
    .X(_2203_));
 sky130_fd_sc_hd__nor2_1 _5144_ (.A(_1966_),
    .B(_2193_),
    .Y(_2204_));
 sky130_fd_sc_hd__a211o_1 _5145_ (.A1(_2193_),
    .A2(_2195_),
    .B1(_2203_),
    .C1(_2204_),
    .X(_2205_));
 sky130_fd_sc_hd__a32o_1 _5146_ (.A1(_2158_),
    .A2(_2191_),
    .A3(_2205_),
    .B1(_2462_),
    .B2(net5),
    .X(_2206_));
 sky130_fd_sc_hd__mux2_1 _5147_ (.A0(_2206_),
    .A1(_0452_),
    .S(_2175_),
    .X(_2207_));
 sky130_fd_sc_hd__clkbuf_1 _5148_ (.A(_2207_),
    .X(_0313_));
 sky130_fd_sc_hd__a21o_1 _5149_ (.A1(_2022_),
    .A2(_2026_),
    .B1(_1997_),
    .X(_2208_));
 sky130_fd_sc_hd__nand2_1 _5150_ (.A(_2506_),
    .B(_2208_),
    .Y(_2209_));
 sky130_fd_sc_hd__a31o_1 _5151_ (.A1(_1997_),
    .A2(_2022_),
    .A3(_2026_),
    .B1(_2209_),
    .X(_2210_));
 sky130_fd_sc_hd__a22o_1 _5152_ (.A1(_0579_),
    .A2(_2094_),
    .B1(_2095_),
    .B2(_0452_),
    .X(_2211_));
 sky130_fd_sc_hd__o221a_1 _5153_ (.A1(_2511_),
    .A2(_2057_),
    .B1(_2048_),
    .B2(_2600_),
    .C1(_2185_),
    .X(_2212_));
 sky130_fd_sc_hd__nand2_1 _5154_ (.A(_2508_),
    .B(_2034_),
    .Y(_2213_));
 sky130_fd_sc_hd__a31o_1 _5155_ (.A1(_1997_),
    .A2(_2021_),
    .A3(_2033_),
    .B1(_2213_),
    .X(_2214_));
 sky130_fd_sc_hd__and3_1 _5156_ (.A(_2057_),
    .B(_2049_),
    .C(_2052_),
    .X(_2215_));
 sky130_fd_sc_hd__or3_1 _5157_ (.A(_2557_),
    .B(_2103_),
    .C(_2215_),
    .X(_2216_));
 sky130_fd_sc_hd__and4b_1 _5158_ (.A_N(_2211_),
    .B(_2212_),
    .C(_2214_),
    .D(_2216_),
    .X(_2217_));
 sky130_fd_sc_hd__nand2_1 _5159_ (.A(_2210_),
    .B(_2217_),
    .Y(_2218_));
 sky130_fd_sc_hd__o311a_1 _5160_ (.A1(_0539_),
    .A2(io_out[2]),
    .A3(_2185_),
    .B1(_2218_),
    .C1(_1695_),
    .X(_2219_));
 sky130_fd_sc_hd__a21oi_1 _5161_ (.A1(_2145_),
    .A2(_1032_),
    .B1(_2219_),
    .Y(_2220_));
 sky130_fd_sc_hd__o21a_1 _5162_ (.A1(_2144_),
    .A2(_0507_),
    .B1(_1495_),
    .X(_2221_));
 sky130_fd_sc_hd__o21ai_1 _5163_ (.A1(_2562_),
    .A2(_2220_),
    .B1(_2221_),
    .Y(_2222_));
 sky130_fd_sc_hd__a21bo_1 _5164_ (.A1(_2022_),
    .A2(_2001_),
    .B1_N(_2021_),
    .X(_2223_));
 sky130_fd_sc_hd__or2_1 _5165_ (.A(_2057_),
    .B(_2223_),
    .X(_2224_));
 sky130_fd_sc_hd__nand2_1 _5166_ (.A(_2057_),
    .B(_2223_),
    .Y(_2225_));
 sky130_fd_sc_hd__or2_1 _5167_ (.A(_2004_),
    .B(_2006_),
    .X(_2226_));
 sky130_fd_sc_hd__o21ai_1 _5168_ (.A1(_2075_),
    .A2(_2079_),
    .B1(_2069_),
    .Y(_2227_));
 sky130_fd_sc_hd__nor2_1 _5169_ (.A(_2080_),
    .B(_2227_),
    .Y(_2228_));
 sky130_fd_sc_hd__nand2_1 _5170_ (.A(_2055_),
    .B(_2215_),
    .Y(_2229_));
 sky130_fd_sc_hd__nand3_1 _5171_ (.A(_1997_),
    .B(_2022_),
    .C(_2197_),
    .Y(_2230_));
 sky130_fd_sc_hd__a21o_1 _5172_ (.A1(_2022_),
    .A2(_2197_),
    .B1(_1997_),
    .X(_2231_));
 sky130_fd_sc_hd__and3_1 _5173_ (.A(_2196_),
    .B(_2230_),
    .C(_2231_),
    .X(_2232_));
 sky130_fd_sc_hd__a31o_1 _5174_ (.A1(_2154_),
    .A2(_2058_),
    .A3(_2229_),
    .B1(_2232_),
    .X(_2233_));
 sky130_fd_sc_hd__or4_1 _5175_ (.A(_2553_),
    .B(_2211_),
    .C(_2228_),
    .D(_2233_),
    .X(_2234_));
 sky130_fd_sc_hd__a31o_1 _5176_ (.A1(_2097_),
    .A2(_2007_),
    .A3(_2226_),
    .B1(_2234_),
    .X(_2235_));
 sky130_fd_sc_hd__a31o_1 _5177_ (.A1(_2195_),
    .A2(_2224_),
    .A3(_2225_),
    .B1(_2235_),
    .X(_2236_));
 sky130_fd_sc_hd__a32o_1 _5178_ (.A1(_2158_),
    .A2(_2222_),
    .A3(_2236_),
    .B1(_2462_),
    .B2(net6),
    .X(_2237_));
 sky130_fd_sc_hd__mux2_1 _5179_ (.A0(_2237_),
    .A1(_0539_),
    .S(_2175_),
    .X(_2238_));
 sky130_fd_sc_hd__clkbuf_1 _5180_ (.A(_2238_),
    .X(_0314_));
 sky130_fd_sc_hd__or3b_1 _5181_ (.A(_1993_),
    .B(_2102_),
    .C_N(_2058_),
    .X(_2239_));
 sky130_fd_sc_hd__nand2_1 _5182_ (.A(_2494_),
    .B(_2506_),
    .Y(_2240_));
 sky130_fd_sc_hd__nor3_1 _5183_ (.A(_2082_),
    .B(_2074_),
    .C(_2080_),
    .Y(_2241_));
 sky130_fd_sc_hd__a21o_1 _5184_ (.A1(_1994_),
    .A2(_2225_),
    .B1(_1993_),
    .X(_2242_));
 sky130_fd_sc_hd__nand2_1 _5185_ (.A(_0453_),
    .B(_2508_),
    .Y(_2243_));
 sky130_fd_sc_hd__a21oi_1 _5186_ (.A1(_2008_),
    .A2(_2225_),
    .B1(_2243_),
    .Y(_2244_));
 sky130_fd_sc_hd__a21o_1 _5187_ (.A1(_1996_),
    .A2(_2231_),
    .B1(_1993_),
    .X(_2245_));
 sky130_fd_sc_hd__nand2_1 _5188_ (.A(_2081_),
    .B(_2231_),
    .Y(_2246_));
 sky130_fd_sc_hd__a22o_1 _5189_ (.A1(_0646_),
    .A2(_2094_),
    .B1(_2095_),
    .B2(_0539_),
    .X(_2247_));
 sky130_fd_sc_hd__a311o_1 _5190_ (.A1(_2196_),
    .A2(_2245_),
    .A3(_2246_),
    .B1(_2247_),
    .C1(_2097_),
    .X(_2248_));
 sky130_fd_sc_hd__a21oi_1 _5191_ (.A1(_2242_),
    .A2(_2244_),
    .B1(_2248_),
    .Y(_2249_));
 sky130_fd_sc_hd__o31ai_1 _5192_ (.A1(_2083_),
    .A2(_2240_),
    .A3(_2241_),
    .B1(_2249_),
    .Y(_2250_));
 sky130_fd_sc_hd__a31o_1 _5193_ (.A1(_2154_),
    .A2(_2060_),
    .A3(_2239_),
    .B1(_2250_),
    .X(_2251_));
 sky130_fd_sc_hd__o211a_1 _5194_ (.A1(_1995_),
    .A2(_2008_),
    .B1(_1998_),
    .C1(_2007_),
    .X(_2252_));
 sky130_fd_sc_hd__o21ai_1 _5195_ (.A1(_2009_),
    .A2(_2252_),
    .B1(_2097_),
    .Y(_2253_));
 sky130_fd_sc_hd__nand2_1 _5196_ (.A(_2034_),
    .B(_2008_),
    .Y(_2254_));
 sky130_fd_sc_hd__a21o_1 _5197_ (.A1(_1996_),
    .A2(_2208_),
    .B1(_1992_),
    .X(_2255_));
 sky130_fd_sc_hd__inv_2 _5198_ (.A(_2255_),
    .Y(_2256_));
 sky130_fd_sc_hd__a211oi_1 _5199_ (.A1(_2081_),
    .A2(_2208_),
    .B1(_2256_),
    .C1(_2020_),
    .Y(_2257_));
 sky130_fd_sc_hd__or3_1 _5200_ (.A(_1993_),
    .B(_2102_),
    .C(_2103_),
    .X(_2258_));
 sky130_fd_sc_hd__and3_1 _5201_ (.A(_2515_),
    .B(_2104_),
    .C(_2258_),
    .X(_2259_));
 sky130_fd_sc_hd__o221a_1 _5202_ (.A1(_2511_),
    .A2(_2059_),
    .B1(_2047_),
    .B2(_2600_),
    .C1(_2184_),
    .X(_2260_));
 sky130_fd_sc_hd__or4b_1 _5203_ (.A(_2257_),
    .B(_2259_),
    .C(_2247_),
    .D_N(_2260_),
    .X(_2261_));
 sky130_fd_sc_hd__a31o_1 _5204_ (.A1(_2508_),
    .A2(_2035_),
    .A3(_2254_),
    .B1(_2261_),
    .X(_2262_));
 sky130_fd_sc_hd__o311a_1 _5205_ (.A1(_0579_),
    .A2(io_out[3]),
    .A3(_2185_),
    .B1(_2262_),
    .C1(_1695_),
    .X(_2263_));
 sky130_fd_sc_hd__a21oi_1 _5206_ (.A1(_2145_),
    .A2(_1093_),
    .B1(_2263_),
    .Y(_2264_));
 sky130_fd_sc_hd__mux2_1 _5207_ (.A0(_0570_),
    .A1(_2264_),
    .S(_2144_),
    .X(_2265_));
 sky130_fd_sc_hd__nor2_1 _5208_ (.A(_1490_),
    .B(_2265_),
    .Y(_2266_));
 sky130_fd_sc_hd__a31o_1 _5209_ (.A1(_1491_),
    .A2(_2251_),
    .A3(_2253_),
    .B1(_2266_),
    .X(_2267_));
 sky130_fd_sc_hd__a22o_1 _5210_ (.A1(net7),
    .A2(_2462_),
    .B1(_2158_),
    .B2(_2267_),
    .X(_2268_));
 sky130_fd_sc_hd__mux2_1 _5211_ (.A0(_2268_),
    .A1(_0579_),
    .S(_2175_),
    .X(_2269_));
 sky130_fd_sc_hd__clkbuf_1 _5212_ (.A(_2269_),
    .X(_0315_));
 sky130_fd_sc_hd__a211o_1 _5213_ (.A1(_2035_),
    .A2(_2010_),
    .B1(_2036_),
    .C1(_2194_),
    .X(_2270_));
 sky130_fd_sc_hd__a21o_1 _5214_ (.A1(_1991_),
    .A2(_2255_),
    .B1(_1988_),
    .X(_2271_));
 sky130_fd_sc_hd__o211a_1 _5215_ (.A1(_2085_),
    .A2(_2256_),
    .B1(_2271_),
    .C1(_2506_),
    .X(_2272_));
 sky130_fd_sc_hd__a22o_1 _5216_ (.A1(_0716_),
    .A2(_2094_),
    .B1(_2095_),
    .B2(_0579_),
    .X(_2273_));
 sky130_fd_sc_hd__o221a_1 _5217_ (.A1(_2511_),
    .A2(_2061_),
    .B1(_2046_),
    .B2(_2600_),
    .C1(_2185_),
    .X(_2274_));
 sky130_fd_sc_hd__nand2_1 _5218_ (.A(_2515_),
    .B(_2105_),
    .Y(_2275_));
 sky130_fd_sc_hd__a31o_1 _5219_ (.A1(_2061_),
    .A2(_2047_),
    .A3(_2104_),
    .B1(_2275_),
    .X(_2276_));
 sky130_fd_sc_hd__and4bb_1 _5220_ (.A_N(_2272_),
    .B_N(_2273_),
    .C(_2274_),
    .D(_2276_),
    .X(_2277_));
 sky130_fd_sc_hd__o31a_1 _5221_ (.A1(_0646_),
    .A2(io_out[4]),
    .A3(_2185_),
    .B1(_1695_),
    .X(_2278_));
 sky130_fd_sc_hd__a21bo_1 _5222_ (.A1(_2270_),
    .A2(_2277_),
    .B1_N(_2278_),
    .X(_2279_));
 sky130_fd_sc_hd__o211a_1 _5223_ (.A1(_1695_),
    .A2(_1155_),
    .B1(_2279_),
    .C1(_2144_),
    .X(_2280_));
 sky130_fd_sc_hd__a211o_1 _5224_ (.A1(_2562_),
    .A2(_0642_),
    .B1(_2280_),
    .C1(_1490_),
    .X(_2281_));
 sky130_fd_sc_hd__nor2_1 _5225_ (.A(_1995_),
    .B(_2009_),
    .Y(_2282_));
 sky130_fd_sc_hd__xnor2_1 _5226_ (.A(_2011_),
    .B(_2282_),
    .Y(_2283_));
 sky130_fd_sc_hd__a21oi_1 _5227_ (.A1(_1989_),
    .A2(_2242_),
    .B1(_1988_),
    .Y(_2284_));
 sky130_fd_sc_hd__a211o_1 _5228_ (.A1(_2010_),
    .A2(_2242_),
    .B1(_2284_),
    .C1(_2243_),
    .X(_2285_));
 sky130_fd_sc_hd__a21oi_1 _5229_ (.A1(_1991_),
    .A2(_2245_),
    .B1(_1988_),
    .Y(_2286_));
 sky130_fd_sc_hd__inv_2 _5230_ (.A(_2196_),
    .Y(_2287_));
 sky130_fd_sc_hd__a311o_1 _5231_ (.A1(_1988_),
    .A2(_1991_),
    .A3(_2245_),
    .B1(_2286_),
    .C1(_2287_),
    .X(_2288_));
 sky130_fd_sc_hd__and4bb_1 _5232_ (.A_N(_2097_),
    .B_N(_2273_),
    .C(_2285_),
    .D(_2288_),
    .X(_2289_));
 sky130_fd_sc_hd__nand2_1 _5233_ (.A(_2154_),
    .B(_2062_),
    .Y(_2290_));
 sky130_fd_sc_hd__a31o_1 _5234_ (.A1(_2061_),
    .A2(_2047_),
    .A3(_2060_),
    .B1(_2290_),
    .X(_2291_));
 sky130_fd_sc_hd__a211oi_1 _5235_ (.A1(_2084_),
    .A2(_2085_),
    .B1(_2073_),
    .C1(_2083_),
    .Y(_2292_));
 sky130_fd_sc_hd__or3_1 _5236_ (.A(_2086_),
    .B(_2240_),
    .C(_2292_),
    .X(_2293_));
 sky130_fd_sc_hd__a31o_1 _5237_ (.A1(_2289_),
    .A2(_2291_),
    .A3(_2293_),
    .B1(_2554_),
    .X(_2294_));
 sky130_fd_sc_hd__a21o_1 _5238_ (.A1(_2097_),
    .A2(_2283_),
    .B1(_2294_),
    .X(_2295_));
 sky130_fd_sc_hd__nand2_1 _5239_ (.A(_2281_),
    .B(_2295_),
    .Y(_2296_));
 sky130_fd_sc_hd__a22o_1 _5240_ (.A1(net8),
    .A2(_2462_),
    .B1(_2158_),
    .B2(_2296_),
    .X(_2297_));
 sky130_fd_sc_hd__mux2_1 _5241_ (.A0(_2297_),
    .A1(_0646_),
    .S(_2175_),
    .X(_2298_));
 sky130_fd_sc_hd__clkbuf_1 _5242_ (.A(_2298_),
    .X(_0316_));
 sky130_fd_sc_hd__a22o_1 _5243_ (.A1(_0797_),
    .A2(_2094_),
    .B1(_2095_),
    .B2(_0646_),
    .X(_2299_));
 sky130_fd_sc_hd__o22a_1 _5244_ (.A1(_2511_),
    .A2(_1982_),
    .B1(_2045_),
    .B2(_2600_),
    .X(_2300_));
 sky130_fd_sc_hd__or3b_1 _5245_ (.A(_2147_),
    .B(_2299_),
    .C_N(_2300_),
    .X(_2301_));
 sky130_fd_sc_hd__nand3_1 _5246_ (.A(_1982_),
    .B(_2046_),
    .C(_2105_),
    .Y(_2302_));
 sky130_fd_sc_hd__or2b_1 _5247_ (.A(io_out[4]),
    .B_N(_0646_),
    .X(_2303_));
 sky130_fd_sc_hd__a21o_1 _5248_ (.A1(_2303_),
    .A2(_2271_),
    .B1(_2028_),
    .X(_2304_));
 sky130_fd_sc_hd__or3b_1 _5249_ (.A(_1981_),
    .B(_1986_),
    .C_N(_2271_),
    .X(_2305_));
 sky130_fd_sc_hd__o211a_1 _5250_ (.A1(_2036_),
    .A2(_2013_),
    .B1(_2037_),
    .C1(_2508_),
    .X(_2306_));
 sky130_fd_sc_hd__a31o_1 _5251_ (.A1(_2506_),
    .A2(_2304_),
    .A3(_2305_),
    .B1(_2306_),
    .X(_2307_));
 sky130_fd_sc_hd__a31o_1 _5252_ (.A1(_2154_),
    .A2(_2106_),
    .A3(_2302_),
    .B1(_2307_),
    .X(_2308_));
 sky130_fd_sc_hd__o32a_1 _5253_ (.A1(_0716_),
    .A2(io_out[5]),
    .A3(_2185_),
    .B1(_2301_),
    .B2(_2308_),
    .X(_2309_));
 sky130_fd_sc_hd__nand2_1 _5254_ (.A(_2145_),
    .B(_1211_),
    .Y(_2310_));
 sky130_fd_sc_hd__o211a_1 _5255_ (.A1(_2145_),
    .A2(_2309_),
    .B1(_2310_),
    .C1(_2144_),
    .X(_2311_));
 sky130_fd_sc_hd__a211o_1 _5256_ (.A1(_2562_),
    .A2(_0709_),
    .B1(_2311_),
    .C1(_1766_),
    .X(_2312_));
 sky130_fd_sc_hd__o31a_1 _5257_ (.A1(_2087_),
    .A2(_2072_),
    .A3(_2086_),
    .B1(_2069_),
    .X(_2313_));
 sky130_fd_sc_hd__o21ai_1 _5258_ (.A1(_1986_),
    .A2(_2286_),
    .B1(_1982_),
    .Y(_2314_));
 sky130_fd_sc_hd__o311a_1 _5259_ (.A1(_1982_),
    .A2(_1986_),
    .A3(_2286_),
    .B1(_2314_),
    .C1(_2196_),
    .X(_2315_));
 sky130_fd_sc_hd__a211o_1 _5260_ (.A1(_2088_),
    .A2(_2313_),
    .B1(_2315_),
    .C1(_2299_),
    .X(_2316_));
 sky130_fd_sc_hd__a211o_1 _5261_ (.A1(_1984_),
    .A2(_2013_),
    .B1(_2012_),
    .C1(_1990_),
    .X(_2317_));
 sky130_fd_sc_hd__a31o_1 _5262_ (.A1(_2097_),
    .A2(_2014_),
    .A3(_2317_),
    .B1(_2554_),
    .X(_2318_));
 sky130_fd_sc_hd__nand3_1 _5263_ (.A(_1982_),
    .B(_2046_),
    .C(_2062_),
    .Y(_2319_));
 sky130_fd_sc_hd__o21ai_1 _5264_ (.A1(_1983_),
    .A2(_2284_),
    .B1(_1982_),
    .Y(_2320_));
 sky130_fd_sc_hd__o211a_1 _5265_ (.A1(_2013_),
    .A2(_2284_),
    .B1(_2320_),
    .C1(_2195_),
    .X(_2321_));
 sky130_fd_sc_hd__a31o_1 _5266_ (.A1(_2154_),
    .A2(_2063_),
    .A3(_2319_),
    .B1(_2321_),
    .X(_2322_));
 sky130_fd_sc_hd__or3_1 _5267_ (.A(_2316_),
    .B(_2318_),
    .C(_2322_),
    .X(_2323_));
 sky130_fd_sc_hd__a32o_1 _5268_ (.A1(_2158_),
    .A2(_2312_),
    .A3(_2323_),
    .B1(_2462_),
    .B2(net9),
    .X(_2324_));
 sky130_fd_sc_hd__mux2_1 _5269_ (.A0(_2324_),
    .A1(_0716_),
    .S(_2175_),
    .X(_2325_));
 sky130_fd_sc_hd__clkbuf_1 _5270_ (.A(_2325_),
    .X(_0317_));
 sky130_fd_sc_hd__o211a_1 _5271_ (.A1(_1979_),
    .A2(_2015_),
    .B1(_1984_),
    .C1(_2014_),
    .X(_2326_));
 sky130_fd_sc_hd__o211a_1 _5272_ (.A1(_2070_),
    .A2(_2089_),
    .B1(_2071_),
    .C1(_2088_),
    .X(_2327_));
 sky130_fd_sc_hd__nand2_1 _5273_ (.A(_2154_),
    .B(_2065_),
    .Y(_2328_));
 sky130_fd_sc_hd__a31o_1 _5274_ (.A1(_2064_),
    .A2(_2045_),
    .A3(_2063_),
    .B1(_2328_),
    .X(_2329_));
 sky130_fd_sc_hd__a21o_1 _5275_ (.A1(_1980_),
    .A2(_2314_),
    .B1(_1978_),
    .X(_2330_));
 sky130_fd_sc_hd__nand2_1 _5276_ (.A(_2089_),
    .B(_2314_),
    .Y(_2331_));
 sky130_fd_sc_hd__a22o_1 _5277_ (.A1(\as1802.D[7] ),
    .A2(_2094_),
    .B1(_2095_),
    .B2(_0716_),
    .X(_2332_));
 sky130_fd_sc_hd__a311oi_1 _5278_ (.A1(_2196_),
    .A2(_2330_),
    .A3(_2331_),
    .B1(_2332_),
    .C1(_2553_),
    .Y(_2333_));
 sky130_fd_sc_hd__o311a_1 _5279_ (.A1(_2090_),
    .A2(_2240_),
    .A3(_2327_),
    .B1(_2329_),
    .C1(_2333_),
    .X(_2334_));
 sky130_fd_sc_hd__o31a_1 _5280_ (.A1(_1966_),
    .A2(_2016_),
    .A3(_2326_),
    .B1(_2334_),
    .X(_2335_));
 sky130_fd_sc_hd__a21oi_1 _5281_ (.A1(_1975_),
    .A2(_2320_),
    .B1(_1978_),
    .Y(_2336_));
 sky130_fd_sc_hd__a211o_1 _5282_ (.A1(_2015_),
    .A2(_2320_),
    .B1(_2336_),
    .C1(_2243_),
    .X(_2337_));
 sky130_fd_sc_hd__nand3_1 _5283_ (.A(_2064_),
    .B(_2045_),
    .C(_2106_),
    .Y(_2338_));
 sky130_fd_sc_hd__nand2_1 _5284_ (.A(_2038_),
    .B(_2064_),
    .Y(_2339_));
 sky130_fd_sc_hd__nand2_1 _5285_ (.A(_2037_),
    .B(_2015_),
    .Y(_2340_));
 sky130_fd_sc_hd__a21oi_1 _5286_ (.A1(_1980_),
    .A2(_2304_),
    .B1(_1978_),
    .Y(_2341_));
 sky130_fd_sc_hd__a211oi_1 _5287_ (.A1(_2089_),
    .A2(_2304_),
    .B1(_2341_),
    .C1(_2020_),
    .Y(_2342_));
 sky130_fd_sc_hd__o21ai_1 _5288_ (.A1(_2600_),
    .A2(_2044_),
    .B1(_2184_),
    .Y(_2343_));
 sky130_fd_sc_hd__a211o_1 _5289_ (.A1(_2512_),
    .A2(_1978_),
    .B1(_2332_),
    .C1(_2343_),
    .X(_2344_));
 sky130_fd_sc_hd__a311o_1 _5290_ (.A1(_2508_),
    .A2(_2339_),
    .A3(_2340_),
    .B1(_2342_),
    .C1(_2344_),
    .X(_2345_));
 sky130_fd_sc_hd__a31o_1 _5291_ (.A1(_2154_),
    .A2(_2107_),
    .A3(_2338_),
    .B1(_2345_),
    .X(_2346_));
 sky130_fd_sc_hd__o31a_1 _5292_ (.A1(_0797_),
    .A2(io_out[6]),
    .A3(_2185_),
    .B1(_1695_),
    .X(_2347_));
 sky130_fd_sc_hd__a2bb2o_1 _5293_ (.A1_N(_1695_),
    .A2_N(_1265_),
    .B1(_2346_),
    .B2(_2347_),
    .X(_2348_));
 sky130_fd_sc_hd__mux2_1 _5294_ (.A0(_0792_),
    .A1(_2348_),
    .S(_2144_),
    .X(_2349_));
 sky130_fd_sc_hd__o2bb2a_1 _5295_ (.A1_N(_2335_),
    .A2_N(_2337_),
    .B1(_2349_),
    .B2(_1766_),
    .X(_2350_));
 sky130_fd_sc_hd__a22o_1 _5296_ (.A1(net10),
    .A2(_2461_),
    .B1(_2158_),
    .B2(_2350_),
    .X(_2351_));
 sky130_fd_sc_hd__mux2_1 _5297_ (.A0(_2351_),
    .A1(_0797_),
    .S(_2175_),
    .X(_2352_));
 sky130_fd_sc_hd__clkbuf_1 _5298_ (.A(_2352_),
    .X(_0318_));
 sky130_fd_sc_hd__xnor2_1 _5299_ (.A(_2039_),
    .B(_2027_),
    .Y(_2353_));
 sky130_fd_sc_hd__o21ai_1 _5300_ (.A1(_1976_),
    .A2(_2341_),
    .B1(_1972_),
    .Y(_2354_));
 sky130_fd_sc_hd__o211a_1 _5301_ (.A1(_2091_),
    .A2(_2341_),
    .B1(_2354_),
    .C1(_2506_),
    .X(_2355_));
 sky130_fd_sc_hd__o221ai_1 _5302_ (.A1(_2511_),
    .A2(_1972_),
    .B1(_2043_),
    .B2(_2600_),
    .C1(_2185_),
    .Y(_2356_));
 sky130_fd_sc_hd__a211o_1 _5303_ (.A1(_0797_),
    .A2(_2095_),
    .B1(_2355_),
    .C1(_2356_),
    .X(_2357_));
 sky130_fd_sc_hd__and3_1 _5304_ (.A(_1972_),
    .B(_2044_),
    .C(_2107_),
    .X(_2358_));
 sky130_fd_sc_hd__nor3_1 _5305_ (.A(_2557_),
    .B(_2108_),
    .C(_2358_),
    .Y(_2359_));
 sky130_fd_sc_hd__a211o_1 _5306_ (.A1(_2508_),
    .A2(_2353_),
    .B1(_2357_),
    .C1(_2359_),
    .X(_2360_));
 sky130_fd_sc_hd__o311a_1 _5307_ (.A1(\as1802.D[7] ),
    .A2(io_out[7]),
    .A3(_2185_),
    .B1(_2360_),
    .C1(_1695_),
    .X(_2361_));
 sky130_fd_sc_hd__nor2_1 _5308_ (.A(_1695_),
    .B(_1316_),
    .Y(_2362_));
 sky130_fd_sc_hd__o21a_1 _5309_ (.A1(_2361_),
    .A2(_2362_),
    .B1(_2144_),
    .X(_2363_));
 sky130_fd_sc_hd__nor2_1 _5310_ (.A(_2144_),
    .B(_0831_),
    .Y(_2364_));
 sky130_fd_sc_hd__nand3_1 _5311_ (.A(_1972_),
    .B(_2044_),
    .C(_2065_),
    .Y(_2365_));
 sky130_fd_sc_hd__a211o_1 _5312_ (.A1(_2068_),
    .A2(_2091_),
    .B1(_2070_),
    .C1(_2090_),
    .X(_2366_));
 sky130_fd_sc_hd__and3b_1 _5313_ (.A_N(_2092_),
    .B(_2069_),
    .C(_2366_),
    .X(_2367_));
 sky130_fd_sc_hd__a31o_1 _5314_ (.A1(_2154_),
    .A2(_2066_),
    .A3(_2365_),
    .B1(_2367_),
    .X(_2368_));
 sky130_fd_sc_hd__mux2_1 _5315_ (.A0(_2027_),
    .A1(_2091_),
    .S(_2330_),
    .X(_2369_));
 sky130_fd_sc_hd__mux2_1 _5316_ (.A0(_1974_),
    .A1(_2027_),
    .S(_2336_),
    .X(_2370_));
 sky130_fd_sc_hd__a221o_1 _5317_ (.A1(\as1802.DF ),
    .A2(_2094_),
    .B1(_2095_),
    .B2(_0797_),
    .C1(_2554_),
    .X(_2371_));
 sky130_fd_sc_hd__a31o_1 _5318_ (.A1(_1973_),
    .A2(_2195_),
    .A3(_2370_),
    .B1(_2371_),
    .X(_2372_));
 sky130_fd_sc_hd__a31o_1 _5319_ (.A1(_2068_),
    .A2(_2196_),
    .A3(_2369_),
    .B1(_2372_),
    .X(_2373_));
 sky130_fd_sc_hd__a21o_1 _5320_ (.A1(_1973_),
    .A2(_1974_),
    .B1(_2017_),
    .X(_2374_));
 sky130_fd_sc_hd__or3b_1 _5321_ (.A(_1966_),
    .B(_2018_),
    .C_N(_2374_),
    .X(_2375_));
 sky130_fd_sc_hd__or3b_1 _5322_ (.A(_2368_),
    .B(_2373_),
    .C_N(_2375_),
    .X(_2376_));
 sky130_fd_sc_hd__o311a_1 _5323_ (.A1(_1491_),
    .A2(_2363_),
    .A3(_2364_),
    .B1(_2376_),
    .C1(_2158_),
    .X(_2377_));
 sky130_fd_sc_hd__a21o_1 _5324_ (.A1(net11),
    .A2(_2462_),
    .B1(_2175_),
    .X(_2378_));
 sky130_fd_sc_hd__o2bb2a_1 _5325_ (.A1_N(_0840_),
    .A2_N(_2175_),
    .B1(_2377_),
    .B2(_2378_),
    .X(_0319_));
 sky130_fd_sc_hd__o211a_1 _5326_ (.A1(\as1802.P[0] ),
    .A2(_1488_),
    .B1(_1493_),
    .C1(_2458_),
    .X(_0320_));
 sky130_fd_sc_hd__o21a_1 _5327_ (.A1(\as1802.P[1] ),
    .A2(_1488_),
    .B1(_1500_),
    .X(_0321_));
 sky130_fd_sc_hd__o211a_1 _5328_ (.A1(\as1802.P[2] ),
    .A2(_1488_),
    .B1(_1503_),
    .C1(_2458_),
    .X(_0322_));
 sky130_fd_sc_hd__and2_1 _5329_ (.A(_2457_),
    .B(_1507_),
    .X(_2379_));
 sky130_fd_sc_hd__clkbuf_1 _5330_ (.A(_2379_),
    .X(_0323_));
 sky130_fd_sc_hd__nor2_4 _5331_ (.A(_2494_),
    .B(_2542_),
    .Y(_2380_));
 sky130_fd_sc_hd__a22o_1 _5332_ (.A1(\as1802.P[0] ),
    .A2(_1738_),
    .B1(_2380_),
    .B2(\as1802.T[0] ),
    .X(_2381_));
 sky130_fd_sc_hd__a21o_2 _5333_ (.A1(_2474_),
    .A2(_2563_),
    .B1(_2593_),
    .X(_2382_));
 sky130_fd_sc_hd__a22o_1 _5334_ (.A1(_1958_),
    .A2(_2381_),
    .B1(_2382_),
    .B2(_0382_),
    .X(_2383_));
 sky130_fd_sc_hd__mux2_1 _5335_ (.A0(net1),
    .A1(_2383_),
    .S(_2548_),
    .X(_2384_));
 sky130_fd_sc_hd__or3b_1 _5336_ (.A(_2460_),
    .B(_2581_),
    .C_N(_2476_),
    .X(_2385_));
 sky130_fd_sc_hd__inv_2 _5337_ (.A(\as1802.lda ),
    .Y(_2386_));
 sky130_fd_sc_hd__o221a_1 _5338_ (.A1(_2461_),
    .A2(_0443_),
    .B1(_2167_),
    .B2(_2386_),
    .C1(_2169_),
    .X(_2387_));
 sky130_fd_sc_hd__o32a_1 _5339_ (.A1(_2584_),
    .A2(_1482_),
    .A3(_1708_),
    .B1(_1472_),
    .B2(_2524_),
    .X(_2388_));
 sky130_fd_sc_hd__and4_1 _5340_ (.A(_2173_),
    .B(_2385_),
    .C(_2387_),
    .D(_2388_),
    .X(_2389_));
 sky130_fd_sc_hd__buf_2 _5341_ (.A(_2389_),
    .X(_2390_));
 sky130_fd_sc_hd__mux2_1 _5342_ (.A0(_2702_),
    .A1(_2384_),
    .S(_2390_),
    .X(_2391_));
 sky130_fd_sc_hd__clkbuf_1 _5343_ (.A(_2391_),
    .X(_0324_));
 sky130_fd_sc_hd__a22o_1 _5344_ (.A1(\as1802.P[1] ),
    .A2(_1738_),
    .B1(_2380_),
    .B2(\as1802.T[1] ),
    .X(_2392_));
 sky130_fd_sc_hd__a22o_1 _5345_ (.A1(_0452_),
    .A2(_2382_),
    .B1(_2392_),
    .B2(_1958_),
    .X(_2393_));
 sky130_fd_sc_hd__mux2_1 _5346_ (.A0(net5),
    .A1(_2393_),
    .S(_2548_),
    .X(_2394_));
 sky130_fd_sc_hd__mux2_1 _5347_ (.A0(_0474_),
    .A1(_2394_),
    .S(_2390_),
    .X(_2395_));
 sky130_fd_sc_hd__clkbuf_1 _5348_ (.A(_2395_),
    .X(_0325_));
 sky130_fd_sc_hd__a22o_1 _5349_ (.A1(\as1802.P[2] ),
    .A2(_1738_),
    .B1(_2380_),
    .B2(\as1802.T[2] ),
    .X(_2396_));
 sky130_fd_sc_hd__a22o_1 _5350_ (.A1(_0539_),
    .A2(_2382_),
    .B1(_2396_),
    .B2(_1958_),
    .X(_2397_));
 sky130_fd_sc_hd__mux2_1 _5351_ (.A0(net6),
    .A1(_2397_),
    .S(_2548_),
    .X(_2398_));
 sky130_fd_sc_hd__mux2_1 _5352_ (.A0(io_out[2]),
    .A1(_2398_),
    .S(_2390_),
    .X(_2399_));
 sky130_fd_sc_hd__clkbuf_1 _5353_ (.A(_2399_),
    .X(_0326_));
 sky130_fd_sc_hd__a22o_1 _5354_ (.A1(\as1802.P[3] ),
    .A2(_1738_),
    .B1(_2380_),
    .B2(\as1802.T[3] ),
    .X(_2400_));
 sky130_fd_sc_hd__a22o_1 _5355_ (.A1(_0579_),
    .A2(_2382_),
    .B1(_2400_),
    .B2(_1958_),
    .X(_2401_));
 sky130_fd_sc_hd__mux2_1 _5356_ (.A0(net7),
    .A1(_2401_),
    .S(_2548_),
    .X(_2402_));
 sky130_fd_sc_hd__mux2_1 _5357_ (.A0(io_out[3]),
    .A1(_2402_),
    .S(_2390_),
    .X(_2403_));
 sky130_fd_sc_hd__clkbuf_1 _5358_ (.A(_2403_),
    .X(_0327_));
 sky130_fd_sc_hd__a22o_1 _5359_ (.A1(\as1802.X[0] ),
    .A2(_1738_),
    .B1(_2380_),
    .B2(\as1802.T[4] ),
    .X(_2404_));
 sky130_fd_sc_hd__a22o_1 _5360_ (.A1(_0646_),
    .A2(_2382_),
    .B1(_2404_),
    .B2(_1958_),
    .X(_2405_));
 sky130_fd_sc_hd__mux2_1 _5361_ (.A0(net8),
    .A1(_2405_),
    .S(_2548_),
    .X(_2406_));
 sky130_fd_sc_hd__mux2_1 _5362_ (.A0(io_out[4]),
    .A1(_2406_),
    .S(_2390_),
    .X(_2407_));
 sky130_fd_sc_hd__clkbuf_1 _5363_ (.A(_2407_),
    .X(_0328_));
 sky130_fd_sc_hd__a22o_1 _5364_ (.A1(\as1802.X[1] ),
    .A2(_1738_),
    .B1(_2380_),
    .B2(\as1802.T[5] ),
    .X(_2408_));
 sky130_fd_sc_hd__a22o_1 _5365_ (.A1(_0716_),
    .A2(_2382_),
    .B1(_2408_),
    .B2(_1958_),
    .X(_2409_));
 sky130_fd_sc_hd__mux2_1 _5366_ (.A0(net9),
    .A1(_2409_),
    .S(_2548_),
    .X(_2410_));
 sky130_fd_sc_hd__mux2_1 _5367_ (.A0(io_out[5]),
    .A1(_2410_),
    .S(_2390_),
    .X(_2411_));
 sky130_fd_sc_hd__clkbuf_1 _5368_ (.A(_2411_),
    .X(_0329_));
 sky130_fd_sc_hd__a22o_1 _5369_ (.A1(\as1802.X[2] ),
    .A2(_1738_),
    .B1(_2380_),
    .B2(\as1802.T[6] ),
    .X(_2412_));
 sky130_fd_sc_hd__a22o_1 _5370_ (.A1(_0797_),
    .A2(_2382_),
    .B1(_2412_),
    .B2(_1958_),
    .X(_2413_));
 sky130_fd_sc_hd__mux2_1 _5371_ (.A0(net10),
    .A1(_2413_),
    .S(_2548_),
    .X(_2414_));
 sky130_fd_sc_hd__mux2_1 _5372_ (.A0(io_out[6]),
    .A1(_2414_),
    .S(_2390_),
    .X(_2415_));
 sky130_fd_sc_hd__clkbuf_1 _5373_ (.A(_2415_),
    .X(_0330_));
 sky130_fd_sc_hd__a22o_1 _5374_ (.A1(\as1802.X[3] ),
    .A2(_1738_),
    .B1(_2380_),
    .B2(\as1802.T[7] ),
    .X(_2416_));
 sky130_fd_sc_hd__a22o_1 _5375_ (.A1(\as1802.D[7] ),
    .A2(_2382_),
    .B1(_2416_),
    .B2(_1958_),
    .X(_2417_));
 sky130_fd_sc_hd__mux2_1 _5376_ (.A0(net11),
    .A1(_2417_),
    .S(_2547_),
    .X(_2418_));
 sky130_fd_sc_hd__mux2_1 _5377_ (.A0(io_out[7]),
    .A1(_2418_),
    .S(_2390_),
    .X(_2419_));
 sky130_fd_sc_hd__clkbuf_1 _5378_ (.A(_2419_),
    .X(_0331_));
 sky130_fd_sc_hd__and3_1 _5379_ (.A(_0943_),
    .B(_0945_),
    .C(_1389_),
    .X(_2420_));
 sky130_fd_sc_hd__buf_4 _5380_ (.A(_2420_),
    .X(_2421_));
 sky130_fd_sc_hd__mux2_1 _5381_ (.A0(\as1802.regs[9][8] ),
    .A1(_0939_),
    .S(_2421_),
    .X(_2422_));
 sky130_fd_sc_hd__clkbuf_1 _5382_ (.A(_2422_),
    .X(_0332_));
 sky130_fd_sc_hd__mux2_1 _5383_ (.A0(\as1802.regs[9][9] ),
    .A1(_1007_),
    .S(_2421_),
    .X(_2423_));
 sky130_fd_sc_hd__clkbuf_1 _5384_ (.A(_2423_),
    .X(_0333_));
 sky130_fd_sc_hd__mux2_1 _5385_ (.A0(\as1802.regs[9][10] ),
    .A1(_1068_),
    .S(_2421_),
    .X(_2424_));
 sky130_fd_sc_hd__clkbuf_1 _5386_ (.A(_2424_),
    .X(_0334_));
 sky130_fd_sc_hd__mux2_1 _5387_ (.A0(\as1802.regs[9][11] ),
    .A1(_1134_),
    .S(_2421_),
    .X(_2425_));
 sky130_fd_sc_hd__clkbuf_1 _5388_ (.A(_2425_),
    .X(_0335_));
 sky130_fd_sc_hd__mux2_1 _5389_ (.A0(\as1802.regs[9][12] ),
    .A1(_1188_),
    .S(_2421_),
    .X(_2426_));
 sky130_fd_sc_hd__clkbuf_1 _5390_ (.A(_2426_),
    .X(_0336_));
 sky130_fd_sc_hd__mux2_1 _5391_ (.A0(\as1802.regs[9][13] ),
    .A1(_1246_),
    .S(_2421_),
    .X(_2427_));
 sky130_fd_sc_hd__clkbuf_1 _5392_ (.A(_2427_),
    .X(_0337_));
 sky130_fd_sc_hd__mux2_1 _5393_ (.A0(\as1802.regs[9][14] ),
    .A1(_1298_),
    .S(_2421_),
    .X(_2428_));
 sky130_fd_sc_hd__clkbuf_1 _5394_ (.A(_2428_),
    .X(_0338_));
 sky130_fd_sc_hd__mux2_1 _5395_ (.A0(\as1802.regs[9][15] ),
    .A1(_1351_),
    .S(_2421_),
    .X(_2429_));
 sky130_fd_sc_hd__clkbuf_1 _5396_ (.A(_2429_),
    .X(_0339_));
 sky130_fd_sc_hd__and3_1 _5397_ (.A(_0941_),
    .B(_0945_),
    .C(_1357_),
    .X(_2430_));
 sky130_fd_sc_hd__clkbuf_4 _5398_ (.A(_2430_),
    .X(_2431_));
 sky130_fd_sc_hd__mux2_1 _5399_ (.A0(\as1802.regs[2][8] ),
    .A1(_0939_),
    .S(_2431_),
    .X(_2432_));
 sky130_fd_sc_hd__clkbuf_1 _5400_ (.A(_2432_),
    .X(_0340_));
 sky130_fd_sc_hd__mux2_1 _5401_ (.A0(\as1802.regs[2][9] ),
    .A1(_1007_),
    .S(_2431_),
    .X(_2433_));
 sky130_fd_sc_hd__clkbuf_1 _5402_ (.A(_2433_),
    .X(_0341_));
 sky130_fd_sc_hd__mux2_1 _5403_ (.A0(\as1802.regs[2][10] ),
    .A1(_1068_),
    .S(_2431_),
    .X(_2434_));
 sky130_fd_sc_hd__clkbuf_1 _5404_ (.A(_2434_),
    .X(_0342_));
 sky130_fd_sc_hd__mux2_1 _5405_ (.A0(\as1802.regs[2][11] ),
    .A1(_1134_),
    .S(_2431_),
    .X(_2435_));
 sky130_fd_sc_hd__clkbuf_1 _5406_ (.A(_2435_),
    .X(_0343_));
 sky130_fd_sc_hd__mux2_1 _5407_ (.A0(\as1802.regs[2][12] ),
    .A1(_1188_),
    .S(_2431_),
    .X(_2436_));
 sky130_fd_sc_hd__clkbuf_1 _5408_ (.A(_2436_),
    .X(_0344_));
 sky130_fd_sc_hd__mux2_1 _5409_ (.A0(\as1802.regs[2][13] ),
    .A1(_1246_),
    .S(_2431_),
    .X(_2437_));
 sky130_fd_sc_hd__clkbuf_1 _5410_ (.A(_2437_),
    .X(_0345_));
 sky130_fd_sc_hd__mux2_1 _5411_ (.A0(\as1802.regs[2][14] ),
    .A1(_1298_),
    .S(_2431_),
    .X(_2438_));
 sky130_fd_sc_hd__clkbuf_1 _5412_ (.A(_2438_),
    .X(_0346_));
 sky130_fd_sc_hd__mux2_1 _5413_ (.A0(\as1802.regs[2][15] ),
    .A1(_1351_),
    .S(_2431_),
    .X(_2439_));
 sky130_fd_sc_hd__clkbuf_1 _5414_ (.A(_2439_),
    .X(_0347_));
 sky130_fd_sc_hd__a21o_1 _5415_ (.A1(_1481_),
    .A2(_1708_),
    .B1(_1959_),
    .X(_2440_));
 sky130_fd_sc_hd__mux2_1 _5416_ (.A0(_2440_),
    .A1(\as1802.mem_write ),
    .S(_1726_),
    .X(_2441_));
 sky130_fd_sc_hd__clkbuf_1 _5417_ (.A(_2441_),
    .X(_0348_));
 sky130_fd_sc_hd__and3_1 _5418_ (.A(_1354_),
    .B(_1357_),
    .C(_1389_),
    .X(_2442_));
 sky130_fd_sc_hd__buf_4 _5419_ (.A(_2442_),
    .X(_2443_));
 sky130_fd_sc_hd__mux2_1 _5420_ (.A0(\as1802.regs[1][8] ),
    .A1(_0939_),
    .S(_2443_),
    .X(_2444_));
 sky130_fd_sc_hd__clkbuf_1 _5421_ (.A(_2444_),
    .X(_0349_));
 sky130_fd_sc_hd__mux2_1 _5422_ (.A0(\as1802.regs[1][9] ),
    .A1(_1007_),
    .S(_2443_),
    .X(_2445_));
 sky130_fd_sc_hd__clkbuf_1 _5423_ (.A(_2445_),
    .X(_0350_));
 sky130_fd_sc_hd__mux2_1 _5424_ (.A0(\as1802.regs[1][10] ),
    .A1(_1068_),
    .S(_2443_),
    .X(_2446_));
 sky130_fd_sc_hd__clkbuf_1 _5425_ (.A(_2446_),
    .X(_0351_));
 sky130_fd_sc_hd__mux2_1 _5426_ (.A0(\as1802.regs[1][11] ),
    .A1(_1134_),
    .S(_2443_),
    .X(_2447_));
 sky130_fd_sc_hd__clkbuf_1 _5427_ (.A(_2447_),
    .X(_0352_));
 sky130_fd_sc_hd__mux2_1 _5428_ (.A0(\as1802.regs[1][12] ),
    .A1(_1188_),
    .S(_2443_),
    .X(_2448_));
 sky130_fd_sc_hd__clkbuf_1 _5429_ (.A(_2448_),
    .X(_0353_));
 sky130_fd_sc_hd__mux2_1 _5430_ (.A0(\as1802.regs[1][13] ),
    .A1(_1246_),
    .S(_2443_),
    .X(_2449_));
 sky130_fd_sc_hd__clkbuf_1 _5431_ (.A(_2449_),
    .X(_0354_));
 sky130_fd_sc_hd__mux2_1 _5432_ (.A0(\as1802.regs[1][14] ),
    .A1(_1298_),
    .S(_2443_),
    .X(_2450_));
 sky130_fd_sc_hd__clkbuf_1 _5433_ (.A(_2450_),
    .X(_0355_));
 sky130_fd_sc_hd__mux2_1 _5434_ (.A0(\as1802.regs[1][15] ),
    .A1(_1351_),
    .S(_2443_),
    .X(_2451_));
 sky130_fd_sc_hd__clkbuf_1 _5435_ (.A(_2451_),
    .X(_0356_));
 sky130_fd_sc_hd__a21oi_1 _5436_ (.A1(_2581_),
    .A2(_1479_),
    .B1(_2461_),
    .Y(_2452_));
 sky130_fd_sc_hd__or4b_1 _5437_ (.A(_1690_),
    .B(_2172_),
    .C(_2452_),
    .D_N(_2167_),
    .X(_2453_));
 sky130_fd_sc_hd__mux2_1 _5438_ (.A0(_2578_),
    .A1(io_out[25]),
    .S(_2453_),
    .X(_2454_));
 sky130_fd_sc_hd__clkbuf_1 _5439_ (.A(_2454_),
    .X(_0357_));
 sky130_fd_sc_hd__mux2_1 _5440_ (.A0(_1693_),
    .A1(io_out[26]),
    .S(_2453_),
    .X(_2455_));
 sky130_fd_sc_hd__clkbuf_1 _5441_ (.A(_2455_),
    .X(_0358_));
 sky130_fd_sc_hd__dfxtp_1 _5442_ (.CLK(clknet_leaf_30_clk),
    .D(_0012_),
    .Q(\as1802.regs[15][0] ));
 sky130_fd_sc_hd__dfxtp_1 _5443_ (.CLK(clknet_leaf_35_clk),
    .D(_0013_),
    .Q(\as1802.regs[15][1] ));
 sky130_fd_sc_hd__dfxtp_1 _5444_ (.CLK(clknet_leaf_42_clk),
    .D(_0014_),
    .Q(\as1802.regs[15][2] ));
 sky130_fd_sc_hd__dfxtp_1 _5445_ (.CLK(clknet_leaf_33_clk),
    .D(_0015_),
    .Q(\as1802.regs[15][3] ));
 sky130_fd_sc_hd__dfxtp_1 _5446_ (.CLK(clknet_leaf_33_clk),
    .D(_0016_),
    .Q(\as1802.regs[15][4] ));
 sky130_fd_sc_hd__dfxtp_1 _5447_ (.CLK(clknet_leaf_16_clk),
    .D(_0017_),
    .Q(\as1802.regs[15][5] ));
 sky130_fd_sc_hd__dfxtp_1 _5448_ (.CLK(clknet_leaf_22_clk),
    .D(_0018_),
    .Q(\as1802.regs[15][6] ));
 sky130_fd_sc_hd__dfxtp_1 _5449_ (.CLK(clknet_leaf_17_clk),
    .D(_0019_),
    .Q(\as1802.regs[15][7] ));
 sky130_fd_sc_hd__dfxtp_1 _5450_ (.CLK(clknet_leaf_19_clk),
    .D(_0020_),
    .Q(\as1802.regs[10][8] ));
 sky130_fd_sc_hd__dfxtp_1 _5451_ (.CLK(clknet_leaf_12_clk),
    .D(_0021_),
    .Q(\as1802.regs[10][9] ));
 sky130_fd_sc_hd__dfxtp_1 _5452_ (.CLK(clknet_leaf_13_clk),
    .D(_0022_),
    .Q(\as1802.regs[10][10] ));
 sky130_fd_sc_hd__dfxtp_1 _5453_ (.CLK(clknet_leaf_14_clk),
    .D(_0023_),
    .Q(\as1802.regs[10][11] ));
 sky130_fd_sc_hd__dfxtp_1 _5454_ (.CLK(clknet_leaf_11_clk),
    .D(_0024_),
    .Q(\as1802.regs[10][12] ));
 sky130_fd_sc_hd__dfxtp_1 _5455_ (.CLK(clknet_leaf_9_clk),
    .D(_0025_),
    .Q(\as1802.regs[10][13] ));
 sky130_fd_sc_hd__dfxtp_1 _5456_ (.CLK(clknet_leaf_6_clk),
    .D(_0026_),
    .Q(\as1802.regs[10][14] ));
 sky130_fd_sc_hd__dfxtp_1 _5457_ (.CLK(clknet_leaf_4_clk),
    .D(_0027_),
    .Q(\as1802.regs[10][15] ));
 sky130_fd_sc_hd__dfxtp_1 _5458_ (.CLK(clknet_leaf_17_clk),
    .D(_0028_),
    .Q(\as1802.regs[0][8] ));
 sky130_fd_sc_hd__dfxtp_1 _5459_ (.CLK(clknet_leaf_12_clk),
    .D(_0029_),
    .Q(\as1802.regs[0][9] ));
 sky130_fd_sc_hd__dfxtp_1 _5460_ (.CLK(clknet_leaf_13_clk),
    .D(_0030_),
    .Q(\as1802.regs[0][10] ));
 sky130_fd_sc_hd__dfxtp_1 _5461_ (.CLK(clknet_leaf_13_clk),
    .D(_0031_),
    .Q(\as1802.regs[0][11] ));
 sky130_fd_sc_hd__dfxtp_1 _5462_ (.CLK(clknet_leaf_10_clk),
    .D(_0032_),
    .Q(\as1802.regs[0][12] ));
 sky130_fd_sc_hd__dfxtp_1 _5463_ (.CLK(clknet_leaf_9_clk),
    .D(_0033_),
    .Q(\as1802.regs[0][13] ));
 sky130_fd_sc_hd__dfxtp_1 _5464_ (.CLK(clknet_leaf_6_clk),
    .D(_0034_),
    .Q(\as1802.regs[0][14] ));
 sky130_fd_sc_hd__dfxtp_1 _5465_ (.CLK(clknet_leaf_4_clk),
    .D(_0035_),
    .Q(\as1802.regs[0][15] ));
 sky130_fd_sc_hd__dfxtp_1 _5466_ (.CLK(clknet_leaf_19_clk),
    .D(_0036_),
    .Q(\as1802.regs[8][8] ));
 sky130_fd_sc_hd__dfxtp_1 _5467_ (.CLK(clknet_leaf_12_clk),
    .D(_0037_),
    .Q(\as1802.regs[8][9] ));
 sky130_fd_sc_hd__dfxtp_1 _5468_ (.CLK(clknet_leaf_15_clk),
    .D(_0038_),
    .Q(\as1802.regs[8][10] ));
 sky130_fd_sc_hd__dfxtp_1 _5469_ (.CLK(clknet_leaf_10_clk),
    .D(_0039_),
    .Q(\as1802.regs[8][11] ));
 sky130_fd_sc_hd__dfxtp_1 _5470_ (.CLK(clknet_leaf_11_clk),
    .D(_0040_),
    .Q(\as1802.regs[8][12] ));
 sky130_fd_sc_hd__dfxtp_1 _5471_ (.CLK(clknet_leaf_8_clk),
    .D(_0041_),
    .Q(\as1802.regs[8][13] ));
 sky130_fd_sc_hd__dfxtp_1 _5472_ (.CLK(clknet_leaf_6_clk),
    .D(_0042_),
    .Q(\as1802.regs[8][14] ));
 sky130_fd_sc_hd__dfxtp_1 _5473_ (.CLK(clknet_leaf_4_clk),
    .D(_0043_),
    .Q(\as1802.regs[8][15] ));
 sky130_fd_sc_hd__dfxtp_1 _5474_ (.CLK(clknet_leaf_20_clk),
    .D(_0044_),
    .Q(\as1802.regs[4][8] ));
 sky130_fd_sc_hd__dfxtp_1 _5475_ (.CLK(clknet_leaf_20_clk),
    .D(_0045_),
    .Q(\as1802.regs[4][9] ));
 sky130_fd_sc_hd__dfxtp_1 _5476_ (.CLK(clknet_leaf_18_clk),
    .D(_0046_),
    .Q(\as1802.regs[4][10] ));
 sky130_fd_sc_hd__dfxtp_1 _5477_ (.CLK(clknet_leaf_11_clk),
    .D(_0047_),
    .Q(\as1802.regs[4][11] ));
 sky130_fd_sc_hd__dfxtp_1 _5478_ (.CLK(clknet_leaf_12_clk),
    .D(_0048_),
    .Q(\as1802.regs[4][12] ));
 sky130_fd_sc_hd__dfxtp_1 _5479_ (.CLK(clknet_leaf_8_clk),
    .D(_0049_),
    .Q(\as1802.regs[4][13] ));
 sky130_fd_sc_hd__dfxtp_1 _5480_ (.CLK(clknet_leaf_7_clk),
    .D(_0050_),
    .Q(\as1802.regs[4][14] ));
 sky130_fd_sc_hd__dfxtp_1 _5481_ (.CLK(clknet_leaf_4_clk),
    .D(_0051_),
    .Q(\as1802.regs[4][15] ));
 sky130_fd_sc_hd__dfxtp_1 _5482_ (.CLK(clknet_leaf_17_clk),
    .D(_0052_),
    .Q(\as1802.regs[5][8] ));
 sky130_fd_sc_hd__dfxtp_1 _5483_ (.CLK(clknet_leaf_20_clk),
    .D(_0053_),
    .Q(\as1802.regs[5][9] ));
 sky130_fd_sc_hd__dfxtp_1 _5484_ (.CLK(clknet_leaf_18_clk),
    .D(_0054_),
    .Q(\as1802.regs[5][10] ));
 sky130_fd_sc_hd__dfxtp_1 _5485_ (.CLK(clknet_leaf_11_clk),
    .D(_0055_),
    .Q(\as1802.regs[5][11] ));
 sky130_fd_sc_hd__dfxtp_1 _5486_ (.CLK(clknet_leaf_11_clk),
    .D(_0056_),
    .Q(\as1802.regs[5][12] ));
 sky130_fd_sc_hd__dfxtp_1 _5487_ (.CLK(clknet_leaf_8_clk),
    .D(_0057_),
    .Q(\as1802.regs[5][13] ));
 sky130_fd_sc_hd__dfxtp_1 _5488_ (.CLK(clknet_leaf_7_clk),
    .D(_0058_),
    .Q(\as1802.regs[5][14] ));
 sky130_fd_sc_hd__dfxtp_1 _5489_ (.CLK(clknet_leaf_4_clk),
    .D(_0059_),
    .Q(\as1802.regs[5][15] ));
 sky130_fd_sc_hd__dfxtp_1 _5490_ (.CLK(clknet_leaf_19_clk),
    .D(_0060_),
    .Q(\as1802.regs[7][8] ));
 sky130_fd_sc_hd__dfxtp_1 _5491_ (.CLK(clknet_leaf_19_clk),
    .D(_0061_),
    .Q(\as1802.regs[7][9] ));
 sky130_fd_sc_hd__dfxtp_1 _5492_ (.CLK(clknet_leaf_15_clk),
    .D(_0062_),
    .Q(\as1802.regs[7][10] ));
 sky130_fd_sc_hd__dfxtp_1 _5493_ (.CLK(clknet_leaf_11_clk),
    .D(_0063_),
    .Q(\as1802.regs[7][11] ));
 sky130_fd_sc_hd__dfxtp_1 _5494_ (.CLK(clknet_leaf_11_clk),
    .D(_0064_),
    .Q(\as1802.regs[7][12] ));
 sky130_fd_sc_hd__dfxtp_1 _5495_ (.CLK(clknet_leaf_7_clk),
    .D(_0065_),
    .Q(\as1802.regs[7][13] ));
 sky130_fd_sc_hd__dfxtp_1 _5496_ (.CLK(clknet_leaf_6_clk),
    .D(_0066_),
    .Q(\as1802.regs[7][14] ));
 sky130_fd_sc_hd__dfxtp_1 _5497_ (.CLK(clknet_leaf_4_clk),
    .D(_0067_),
    .Q(\as1802.regs[7][15] ));
 sky130_fd_sc_hd__dfxtp_1 _5498_ (.CLK(clknet_leaf_19_clk),
    .D(_0068_),
    .Q(\as1802.regs[6][8] ));
 sky130_fd_sc_hd__dfxtp_1 _5499_ (.CLK(clknet_leaf_20_clk),
    .D(_0069_),
    .Q(\as1802.regs[6][9] ));
 sky130_fd_sc_hd__dfxtp_1 _5500_ (.CLK(clknet_leaf_13_clk),
    .D(_0070_),
    .Q(\as1802.regs[6][10] ));
 sky130_fd_sc_hd__dfxtp_1 _5501_ (.CLK(clknet_leaf_11_clk),
    .D(_0071_),
    .Q(\as1802.regs[6][11] ));
 sky130_fd_sc_hd__dfxtp_1 _5502_ (.CLK(clknet_leaf_11_clk),
    .D(_0072_),
    .Q(\as1802.regs[6][12] ));
 sky130_fd_sc_hd__dfxtp_1 _5503_ (.CLK(clknet_leaf_7_clk),
    .D(_0073_),
    .Q(\as1802.regs[6][13] ));
 sky130_fd_sc_hd__dfxtp_1 _5504_ (.CLK(clknet_leaf_6_clk),
    .D(_0074_),
    .Q(\as1802.regs[6][14] ));
 sky130_fd_sc_hd__dfxtp_1 _5505_ (.CLK(clknet_leaf_4_clk),
    .D(_0075_),
    .Q(\as1802.regs[6][15] ));
 sky130_fd_sc_hd__dfxtp_1 _5506_ (.CLK(clknet_leaf_18_clk),
    .D(_0076_),
    .Q(\as1802.regs[3][8] ));
 sky130_fd_sc_hd__dfxtp_1 _5507_ (.CLK(clknet_leaf_12_clk),
    .D(_0077_),
    .Q(\as1802.regs[3][9] ));
 sky130_fd_sc_hd__dfxtp_1 _5508_ (.CLK(clknet_leaf_13_clk),
    .D(_0078_),
    .Q(\as1802.regs[3][10] ));
 sky130_fd_sc_hd__dfxtp_1 _5509_ (.CLK(clknet_leaf_13_clk),
    .D(_0079_),
    .Q(\as1802.regs[3][11] ));
 sky130_fd_sc_hd__dfxtp_1 _5510_ (.CLK(clknet_leaf_10_clk),
    .D(_0080_),
    .Q(\as1802.regs[3][12] ));
 sky130_fd_sc_hd__dfxtp_1 _5511_ (.CLK(clknet_leaf_9_clk),
    .D(_0081_),
    .Q(\as1802.regs[3][13] ));
 sky130_fd_sc_hd__dfxtp_1 _5512_ (.CLK(clknet_leaf_5_clk),
    .D(_0082_),
    .Q(\as1802.regs[3][14] ));
 sky130_fd_sc_hd__dfxtp_1 _5513_ (.CLK(clknet_leaf_4_clk),
    .D(_0083_),
    .Q(\as1802.regs[3][15] ));
 sky130_fd_sc_hd__dfxtp_1 _5514_ (.CLK(clknet_leaf_28_clk),
    .D(_0084_),
    .Q(\as1802.regs[9][0] ));
 sky130_fd_sc_hd__dfxtp_1 _5515_ (.CLK(clknet_leaf_34_clk),
    .D(_0085_),
    .Q(\as1802.regs[9][1] ));
 sky130_fd_sc_hd__dfxtp_1 _5516_ (.CLK(clknet_leaf_34_clk),
    .D(_0086_),
    .Q(\as1802.regs[9][2] ));
 sky130_fd_sc_hd__dfxtp_1 _5517_ (.CLK(clknet_leaf_33_clk),
    .D(_0087_),
    .Q(\as1802.regs[9][3] ));
 sky130_fd_sc_hd__dfxtp_1 _5518_ (.CLK(clknet_leaf_25_clk),
    .D(_0088_),
    .Q(\as1802.regs[9][4] ));
 sky130_fd_sc_hd__dfxtp_1 _5519_ (.CLK(clknet_leaf_27_clk),
    .D(_0089_),
    .Q(\as1802.regs[9][5] ));
 sky130_fd_sc_hd__dfxtp_1 _5520_ (.CLK(clknet_leaf_22_clk),
    .D(_0090_),
    .Q(\as1802.regs[9][6] ));
 sky130_fd_sc_hd__dfxtp_1 _5521_ (.CLK(clknet_leaf_21_clk),
    .D(_0091_),
    .Q(\as1802.regs[9][7] ));
 sky130_fd_sc_hd__dfxtp_1 _5522_ (.CLK(clknet_leaf_28_clk),
    .D(_0092_),
    .Q(\as1802.regs[8][0] ));
 sky130_fd_sc_hd__dfxtp_1 _5523_ (.CLK(clknet_leaf_34_clk),
    .D(_0093_),
    .Q(\as1802.regs[8][1] ));
 sky130_fd_sc_hd__dfxtp_1 _5524_ (.CLK(clknet_leaf_34_clk),
    .D(_0094_),
    .Q(\as1802.regs[8][2] ));
 sky130_fd_sc_hd__dfxtp_1 _5525_ (.CLK(clknet_leaf_33_clk),
    .D(_0095_),
    .Q(\as1802.regs[8][3] ));
 sky130_fd_sc_hd__dfxtp_1 _5526_ (.CLK(clknet_leaf_25_clk),
    .D(_0096_),
    .Q(\as1802.regs[8][4] ));
 sky130_fd_sc_hd__dfxtp_1 _5527_ (.CLK(clknet_leaf_27_clk),
    .D(_0097_),
    .Q(\as1802.regs[8][5] ));
 sky130_fd_sc_hd__dfxtp_1 _5528_ (.CLK(clknet_leaf_22_clk),
    .D(_0098_),
    .Q(\as1802.regs[8][6] ));
 sky130_fd_sc_hd__dfxtp_1 _5529_ (.CLK(clknet_leaf_20_clk),
    .D(_0099_),
    .Q(\as1802.regs[8][7] ));
 sky130_fd_sc_hd__dfxtp_1 _5530_ (.CLK(clknet_leaf_30_clk),
    .D(_0100_),
    .Q(\as1802.regs[7][0] ));
 sky130_fd_sc_hd__dfxtp_1 _5531_ (.CLK(clknet_leaf_36_clk),
    .D(_0101_),
    .Q(\as1802.regs[7][1] ));
 sky130_fd_sc_hd__dfxtp_1 _5532_ (.CLK(clknet_leaf_34_clk),
    .D(_0102_),
    .Q(\as1802.regs[7][2] ));
 sky130_fd_sc_hd__dfxtp_1 _5533_ (.CLK(clknet_leaf_34_clk),
    .D(_0103_),
    .Q(\as1802.regs[7][3] ));
 sky130_fd_sc_hd__dfxtp_1 _5534_ (.CLK(clknet_leaf_25_clk),
    .D(_0104_),
    .Q(\as1802.regs[7][4] ));
 sky130_fd_sc_hd__dfxtp_1 _5535_ (.CLK(clknet_leaf_25_clk),
    .D(_0105_),
    .Q(\as1802.regs[7][5] ));
 sky130_fd_sc_hd__dfxtp_1 _5536_ (.CLK(clknet_leaf_24_clk),
    .D(_0106_),
    .Q(\as1802.regs[7][6] ));
 sky130_fd_sc_hd__dfxtp_1 _5537_ (.CLK(clknet_leaf_24_clk),
    .D(_0107_),
    .Q(\as1802.regs[7][7] ));
 sky130_fd_sc_hd__dfxtp_1 _5538_ (.CLK(clknet_leaf_30_clk),
    .D(_0108_),
    .Q(\as1802.regs[6][0] ));
 sky130_fd_sc_hd__dfxtp_1 _5539_ (.CLK(clknet_leaf_36_clk),
    .D(_0109_),
    .Q(\as1802.regs[6][1] ));
 sky130_fd_sc_hd__dfxtp_1 _5540_ (.CLK(clknet_leaf_35_clk),
    .D(_0110_),
    .Q(\as1802.regs[6][2] ));
 sky130_fd_sc_hd__dfxtp_1 _5541_ (.CLK(clknet_leaf_34_clk),
    .D(_0111_),
    .Q(\as1802.regs[6][3] ));
 sky130_fd_sc_hd__dfxtp_1 _5542_ (.CLK(clknet_leaf_25_clk),
    .D(_0112_),
    .Q(\as1802.regs[6][4] ));
 sky130_fd_sc_hd__dfxtp_1 _5543_ (.CLK(clknet_leaf_25_clk),
    .D(_0113_),
    .Q(\as1802.regs[6][5] ));
 sky130_fd_sc_hd__dfxtp_1 _5544_ (.CLK(clknet_leaf_24_clk),
    .D(_0114_),
    .Q(\as1802.regs[6][6] ));
 sky130_fd_sc_hd__dfxtp_1 _5545_ (.CLK(clknet_leaf_22_clk),
    .D(_0115_),
    .Q(\as1802.regs[6][7] ));
 sky130_fd_sc_hd__dfxtp_2 _5546_ (.CLK(clknet_leaf_46_clk),
    .D(_0004_),
    .Q(\as1802.instr_cycle[0] ));
 sky130_fd_sc_hd__dfxtp_2 _5547_ (.CLK(clknet_leaf_47_clk),
    .D(_0005_),
    .Q(\as1802.instr_cycle[1] ));
 sky130_fd_sc_hd__dfxtp_2 _5548_ (.CLK(clknet_leaf_0_clk),
    .D(_0006_),
    .Q(\as1802.instr_cycle[2] ));
 sky130_fd_sc_hd__dfxtp_1 _5549_ (.CLK(clknet_2_0__leaf_clk),
    .D(_0007_),
    .Q(\as1802.instr_cycle[3] ));
 sky130_fd_sc_hd__dfxtp_2 _5550_ (.CLK(clknet_leaf_37_clk),
    .D(_0116_),
    .Q(_0000_));
 sky130_fd_sc_hd__dfxtp_2 _5551_ (.CLK(clknet_leaf_37_clk),
    .D(_0117_),
    .Q(_0001_));
 sky130_fd_sc_hd__dfxtp_1 _5552_ (.CLK(clknet_leaf_38_clk),
    .D(_0118_),
    .Q(_0002_));
 sky130_fd_sc_hd__dfxtp_4 _5553_ (.CLK(clknet_leaf_38_clk),
    .D(_0119_),
    .Q(_0003_));
 sky130_fd_sc_hd__dfxtp_1 _5554_ (.CLK(clknet_leaf_32_clk),
    .D(_0120_),
    .Q(\as1802.regs[5][0] ));
 sky130_fd_sc_hd__dfxtp_1 _5555_ (.CLK(clknet_leaf_34_clk),
    .D(_0121_),
    .Q(\as1802.regs[5][1] ));
 sky130_fd_sc_hd__dfxtp_1 _5556_ (.CLK(clknet_leaf_34_clk),
    .D(_0122_),
    .Q(\as1802.regs[5][2] ));
 sky130_fd_sc_hd__dfxtp_1 _5557_ (.CLK(clknet_leaf_34_clk),
    .D(_0123_),
    .Q(\as1802.regs[5][3] ));
 sky130_fd_sc_hd__dfxtp_1 _5558_ (.CLK(clknet_leaf_33_clk),
    .D(_0124_),
    .Q(\as1802.regs[5][4] ));
 sky130_fd_sc_hd__dfxtp_1 _5559_ (.CLK(clknet_leaf_25_clk),
    .D(_0125_),
    .Q(\as1802.regs[5][5] ));
 sky130_fd_sc_hd__dfxtp_1 _5560_ (.CLK(clknet_leaf_24_clk),
    .D(_0126_),
    .Q(\as1802.regs[5][6] ));
 sky130_fd_sc_hd__dfxtp_1 _5561_ (.CLK(clknet_leaf_24_clk),
    .D(_0127_),
    .Q(\as1802.regs[5][7] ));
 sky130_fd_sc_hd__dfxtp_1 _5562_ (.CLK(clknet_leaf_28_clk),
    .D(_0128_),
    .Q(\as1802.regs[4][0] ));
 sky130_fd_sc_hd__dfxtp_1 _5563_ (.CLK(clknet_leaf_34_clk),
    .D(_0129_),
    .Q(\as1802.regs[4][1] ));
 sky130_fd_sc_hd__dfxtp_1 _5564_ (.CLK(clknet_leaf_34_clk),
    .D(_0130_),
    .Q(\as1802.regs[4][2] ));
 sky130_fd_sc_hd__dfxtp_1 _5565_ (.CLK(clknet_leaf_34_clk),
    .D(_0131_),
    .Q(\as1802.regs[4][3] ));
 sky130_fd_sc_hd__dfxtp_1 _5566_ (.CLK(clknet_leaf_25_clk),
    .D(_0132_),
    .Q(\as1802.regs[4][4] ));
 sky130_fd_sc_hd__dfxtp_1 _5567_ (.CLK(clknet_leaf_25_clk),
    .D(_0133_),
    .Q(\as1802.regs[4][5] ));
 sky130_fd_sc_hd__dfxtp_1 _5568_ (.CLK(clknet_leaf_24_clk),
    .D(_0134_),
    .Q(\as1802.regs[4][6] ));
 sky130_fd_sc_hd__dfxtp_1 _5569_ (.CLK(clknet_leaf_24_clk),
    .D(_0135_),
    .Q(\as1802.regs[4][7] ));
 sky130_fd_sc_hd__dfxtp_1 _5570_ (.CLK(clknet_leaf_30_clk),
    .D(_0136_),
    .Q(\as1802.regs[3][0] ));
 sky130_fd_sc_hd__dfxtp_1 _5571_ (.CLK(clknet_leaf_38_clk),
    .D(_0137_),
    .Q(\as1802.regs[3][1] ));
 sky130_fd_sc_hd__dfxtp_1 _5572_ (.CLK(clknet_leaf_38_clk),
    .D(_0138_),
    .Q(\as1802.regs[3][2] ));
 sky130_fd_sc_hd__dfxtp_1 _5573_ (.CLK(clknet_leaf_33_clk),
    .D(_0139_),
    .Q(\as1802.regs[3][3] ));
 sky130_fd_sc_hd__dfxtp_1 _5574_ (.CLK(clknet_leaf_25_clk),
    .D(_0140_),
    .Q(\as1802.regs[3][4] ));
 sky130_fd_sc_hd__dfxtp_1 _5575_ (.CLK(clknet_leaf_26_clk),
    .D(_0141_),
    .Q(\as1802.regs[3][5] ));
 sky130_fd_sc_hd__dfxtp_1 _5576_ (.CLK(clknet_leaf_24_clk),
    .D(_0142_),
    .Q(\as1802.regs[3][6] ));
 sky130_fd_sc_hd__dfxtp_1 _5577_ (.CLK(clknet_leaf_27_clk),
    .D(_0143_),
    .Q(\as1802.regs[3][7] ));
 sky130_fd_sc_hd__dfxtp_2 _5578_ (.CLK(clknet_leaf_30_clk),
    .D(_0144_),
    .Q(\as1802.regs[2][0] ));
 sky130_fd_sc_hd__dfxtp_2 _5579_ (.CLK(clknet_leaf_35_clk),
    .D(_0145_),
    .Q(\as1802.regs[2][1] ));
 sky130_fd_sc_hd__dfxtp_1 _5580_ (.CLK(clknet_leaf_42_clk),
    .D(_0146_),
    .Q(\as1802.regs[2][2] ));
 sky130_fd_sc_hd__dfxtp_2 _5581_ (.CLK(clknet_leaf_33_clk),
    .D(_0147_),
    .Q(\as1802.regs[2][3] ));
 sky130_fd_sc_hd__dfxtp_2 _5582_ (.CLK(clknet_leaf_33_clk),
    .D(_0148_),
    .Q(\as1802.regs[2][4] ));
 sky130_fd_sc_hd__dfxtp_1 _5583_ (.CLK(clknet_leaf_28_clk),
    .D(_0149_),
    .Q(\as1802.regs[2][5] ));
 sky130_fd_sc_hd__dfxtp_2 _5584_ (.CLK(clknet_leaf_24_clk),
    .D(_0150_),
    .Q(\as1802.regs[2][6] ));
 sky130_fd_sc_hd__dfxtp_2 _5585_ (.CLK(clknet_leaf_27_clk),
    .D(_0151_),
    .Q(\as1802.regs[2][7] ));
 sky130_fd_sc_hd__dfxtp_1 _5586_ (.CLK(clknet_leaf_30_clk),
    .D(_0152_),
    .Q(\as1802.regs[1][0] ));
 sky130_fd_sc_hd__dfxtp_1 _5587_ (.CLK(clknet_leaf_38_clk),
    .D(_0153_),
    .Q(\as1802.regs[1][1] ));
 sky130_fd_sc_hd__dfxtp_1 _5588_ (.CLK(clknet_leaf_38_clk),
    .D(_0154_),
    .Q(\as1802.regs[1][2] ));
 sky130_fd_sc_hd__dfxtp_1 _5589_ (.CLK(clknet_leaf_33_clk),
    .D(_0155_),
    .Q(\as1802.regs[1][3] ));
 sky130_fd_sc_hd__dfxtp_1 _5590_ (.CLK(clknet_leaf_33_clk),
    .D(_0156_),
    .Q(\as1802.regs[1][4] ));
 sky130_fd_sc_hd__dfxtp_1 _5591_ (.CLK(clknet_leaf_25_clk),
    .D(_0157_),
    .Q(\as1802.regs[1][5] ));
 sky130_fd_sc_hd__dfxtp_1 _5592_ (.CLK(clknet_leaf_24_clk),
    .D(_0158_),
    .Q(\as1802.regs[1][6] ));
 sky130_fd_sc_hd__dfxtp_1 _5593_ (.CLK(clknet_leaf_27_clk),
    .D(_0159_),
    .Q(\as1802.regs[1][7] ));
 sky130_fd_sc_hd__dfxtp_1 _5594_ (.CLK(clknet_leaf_19_clk),
    .D(_0160_),
    .Q(\as1802.regs[15][8] ));
 sky130_fd_sc_hd__dfxtp_1 _5595_ (.CLK(clknet_leaf_19_clk),
    .D(_0161_),
    .Q(\as1802.regs[15][9] ));
 sky130_fd_sc_hd__dfxtp_1 _5596_ (.CLK(clknet_leaf_16_clk),
    .D(_0162_),
    .Q(\as1802.regs[15][10] ));
 sky130_fd_sc_hd__dfxtp_1 _5597_ (.CLK(clknet_leaf_1_clk),
    .D(_0163_),
    .Q(\as1802.regs[15][11] ));
 sky130_fd_sc_hd__dfxtp_1 _5598_ (.CLK(clknet_leaf_12_clk),
    .D(_0164_),
    .Q(\as1802.regs[15][12] ));
 sky130_fd_sc_hd__dfxtp_1 _5599_ (.CLK(clknet_leaf_8_clk),
    .D(_0165_),
    .Q(\as1802.regs[15][13] ));
 sky130_fd_sc_hd__dfxtp_1 _5600_ (.CLK(clknet_leaf_6_clk),
    .D(_0166_),
    .Q(\as1802.regs[15][14] ));
 sky130_fd_sc_hd__dfxtp_1 _5601_ (.CLK(clknet_leaf_4_clk),
    .D(_0167_),
    .Q(\as1802.regs[15][15] ));
 sky130_fd_sc_hd__dfxtp_1 _5602_ (.CLK(clknet_leaf_28_clk),
    .D(_0168_),
    .Q(\as1802.regs[14][0] ));
 sky130_fd_sc_hd__dfxtp_1 _5603_ (.CLK(clknet_leaf_35_clk),
    .D(_0169_),
    .Q(\as1802.regs[14][1] ));
 sky130_fd_sc_hd__dfxtp_1 _5604_ (.CLK(clknet_leaf_31_clk),
    .D(_0170_),
    .Q(\as1802.regs[14][2] ));
 sky130_fd_sc_hd__dfxtp_1 _5605_ (.CLK(clknet_leaf_32_clk),
    .D(_0171_),
    .Q(\as1802.regs[14][3] ));
 sky130_fd_sc_hd__dfxtp_1 _5606_ (.CLK(clknet_leaf_32_clk),
    .D(_0172_),
    .Q(\as1802.regs[14][4] ));
 sky130_fd_sc_hd__dfxtp_1 _5607_ (.CLK(clknet_leaf_16_clk),
    .D(_0173_),
    .Q(\as1802.regs[14][5] ));
 sky130_fd_sc_hd__dfxtp_1 _5608_ (.CLK(clknet_leaf_23_clk),
    .D(_0174_),
    .Q(\as1802.regs[14][6] ));
 sky130_fd_sc_hd__dfxtp_1 _5609_ (.CLK(clknet_leaf_17_clk),
    .D(_0175_),
    .Q(\as1802.regs[14][7] ));
 sky130_fd_sc_hd__dfxtp_1 _5610_ (.CLK(clknet_leaf_16_clk),
    .D(_0176_),
    .Q(\as1802.regs[13][0] ));
 sky130_fd_sc_hd__dfxtp_1 _5611_ (.CLK(clknet_leaf_35_clk),
    .D(_0177_),
    .Q(\as1802.regs[13][1] ));
 sky130_fd_sc_hd__dfxtp_1 _5612_ (.CLK(clknet_leaf_42_clk),
    .D(_0178_),
    .Q(\as1802.regs[13][2] ));
 sky130_fd_sc_hd__dfxtp_1 _5613_ (.CLK(clknet_leaf_32_clk),
    .D(_0179_),
    .Q(\as1802.regs[13][3] ));
 sky130_fd_sc_hd__dfxtp_1 _5614_ (.CLK(clknet_leaf_32_clk),
    .D(_0180_),
    .Q(\as1802.regs[13][4] ));
 sky130_fd_sc_hd__dfxtp_1 _5615_ (.CLK(clknet_leaf_16_clk),
    .D(_0181_),
    .Q(\as1802.regs[13][5] ));
 sky130_fd_sc_hd__dfxtp_1 _5616_ (.CLK(clknet_leaf_22_clk),
    .D(_0182_),
    .Q(\as1802.regs[13][6] ));
 sky130_fd_sc_hd__dfxtp_1 _5617_ (.CLK(clknet_leaf_16_clk),
    .D(_0183_),
    .Q(\as1802.regs[13][7] ));
 sky130_fd_sc_hd__dfxtp_1 _5618_ (.CLK(clknet_leaf_20_clk),
    .D(_0184_),
    .Q(\as1802.regs[12][8] ));
 sky130_fd_sc_hd__dfxtp_1 _5619_ (.CLK(clknet_leaf_19_clk),
    .D(_0185_),
    .Q(\as1802.regs[12][9] ));
 sky130_fd_sc_hd__dfxtp_1 _5620_ (.CLK(clknet_leaf_18_clk),
    .D(_0186_),
    .Q(\as1802.regs[12][10] ));
 sky130_fd_sc_hd__dfxtp_1 _5621_ (.CLK(clknet_leaf_14_clk),
    .D(_0187_),
    .Q(\as1802.regs[12][11] ));
 sky130_fd_sc_hd__dfxtp_1 _5622_ (.CLK(clknet_leaf_12_clk),
    .D(_0188_),
    .Q(\as1802.regs[12][12] ));
 sky130_fd_sc_hd__dfxtp_1 _5623_ (.CLK(clknet_leaf_8_clk),
    .D(_0189_),
    .Q(\as1802.regs[12][13] ));
 sky130_fd_sc_hd__dfxtp_1 _5624_ (.CLK(clknet_leaf_6_clk),
    .D(_0190_),
    .Q(\as1802.regs[12][14] ));
 sky130_fd_sc_hd__dfxtp_1 _5625_ (.CLK(clknet_leaf_4_clk),
    .D(_0191_),
    .Q(\as1802.regs[12][15] ));
 sky130_fd_sc_hd__dfxtp_1 _5626_ (.CLK(clknet_leaf_28_clk),
    .D(_0192_),
    .Q(\as1802.regs[11][0] ));
 sky130_fd_sc_hd__dfxtp_1 _5627_ (.CLK(clknet_leaf_31_clk),
    .D(_0193_),
    .Q(\as1802.regs[11][1] ));
 sky130_fd_sc_hd__dfxtp_1 _5628_ (.CLK(clknet_leaf_31_clk),
    .D(_0194_),
    .Q(\as1802.regs[11][2] ));
 sky130_fd_sc_hd__dfxtp_1 _5629_ (.CLK(clknet_leaf_32_clk),
    .D(_0195_),
    .Q(\as1802.regs[11][3] ));
 sky130_fd_sc_hd__dfxtp_1 _5630_ (.CLK(clknet_leaf_26_clk),
    .D(_0196_),
    .Q(\as1802.regs[11][4] ));
 sky130_fd_sc_hd__dfxtp_1 _5631_ (.CLK(clknet_leaf_28_clk),
    .D(_0197_),
    .Q(\as1802.regs[11][5] ));
 sky130_fd_sc_hd__dfxtp_1 _5632_ (.CLK(clknet_leaf_21_clk),
    .D(_0198_),
    .Q(\as1802.regs[11][6] ));
 sky130_fd_sc_hd__dfxtp_1 _5633_ (.CLK(clknet_leaf_21_clk),
    .D(_0199_),
    .Q(\as1802.regs[11][7] ));
 sky130_fd_sc_hd__dfxtp_1 _5634_ (.CLK(clknet_leaf_28_clk),
    .D(_0200_),
    .Q(\as1802.regs[10][0] ));
 sky130_fd_sc_hd__dfxtp_1 _5635_ (.CLK(clknet_leaf_31_clk),
    .D(_0201_),
    .Q(\as1802.regs[10][1] ));
 sky130_fd_sc_hd__dfxtp_1 _5636_ (.CLK(clknet_leaf_31_clk),
    .D(_0202_),
    .Q(\as1802.regs[10][2] ));
 sky130_fd_sc_hd__dfxtp_1 _5637_ (.CLK(clknet_leaf_31_clk),
    .D(_0203_),
    .Q(\as1802.regs[10][3] ));
 sky130_fd_sc_hd__dfxtp_1 _5638_ (.CLK(clknet_leaf_26_clk),
    .D(_0204_),
    .Q(\as1802.regs[10][4] ));
 sky130_fd_sc_hd__dfxtp_1 _5639_ (.CLK(clknet_leaf_27_clk),
    .D(_0205_),
    .Q(\as1802.regs[10][5] ));
 sky130_fd_sc_hd__dfxtp_1 _5640_ (.CLK(clknet_leaf_17_clk),
    .D(_0206_),
    .Q(\as1802.regs[10][6] ));
 sky130_fd_sc_hd__dfxtp_1 _5641_ (.CLK(clknet_leaf_17_clk),
    .D(_0207_),
    .Q(\as1802.regs[10][7] ));
 sky130_fd_sc_hd__dfxtp_1 _5642_ (.CLK(clknet_leaf_30_clk),
    .D(_0208_),
    .Q(\as1802.regs[0][0] ));
 sky130_fd_sc_hd__dfxtp_1 _5643_ (.CLK(clknet_leaf_35_clk),
    .D(_0209_),
    .Q(\as1802.regs[0][1] ));
 sky130_fd_sc_hd__dfxtp_1 _5644_ (.CLK(clknet_leaf_42_clk),
    .D(_0210_),
    .Q(\as1802.regs[0][2] ));
 sky130_fd_sc_hd__dfxtp_1 _5645_ (.CLK(clknet_leaf_32_clk),
    .D(_0211_),
    .Q(\as1802.regs[0][3] ));
 sky130_fd_sc_hd__dfxtp_1 _5646_ (.CLK(clknet_leaf_25_clk),
    .D(_0212_),
    .Q(\as1802.regs[0][4] ));
 sky130_fd_sc_hd__dfxtp_1 _5647_ (.CLK(clknet_leaf_27_clk),
    .D(_0213_),
    .Q(\as1802.regs[0][5] ));
 sky130_fd_sc_hd__dfxtp_1 _5648_ (.CLK(clknet_leaf_24_clk),
    .D(_0214_),
    .Q(\as1802.regs[0][6] ));
 sky130_fd_sc_hd__dfxtp_1 _5649_ (.CLK(clknet_leaf_23_clk),
    .D(_0215_),
    .Q(\as1802.regs[0][7] ));
 sky130_fd_sc_hd__dfxtp_1 _5650_ (.CLK(clknet_leaf_19_clk),
    .D(_0216_),
    .Q(\as1802.regs[14][8] ));
 sky130_fd_sc_hd__dfxtp_1 _5651_ (.CLK(clknet_leaf_12_clk),
    .D(_0217_),
    .Q(\as1802.regs[14][9] ));
 sky130_fd_sc_hd__dfxtp_1 _5652_ (.CLK(clknet_leaf_15_clk),
    .D(_0218_),
    .Q(\as1802.regs[14][10] ));
 sky130_fd_sc_hd__dfxtp_1 _5653_ (.CLK(clknet_leaf_1_clk),
    .D(_0219_),
    .Q(\as1802.regs[14][11] ));
 sky130_fd_sc_hd__dfxtp_1 _5654_ (.CLK(clknet_leaf_12_clk),
    .D(_0220_),
    .Q(\as1802.regs[14][12] ));
 sky130_fd_sc_hd__dfxtp_1 _5655_ (.CLK(clknet_leaf_8_clk),
    .D(_0221_),
    .Q(\as1802.regs[14][13] ));
 sky130_fd_sc_hd__dfxtp_1 _5656_ (.CLK(clknet_leaf_6_clk),
    .D(_0222_),
    .Q(\as1802.regs[14][14] ));
 sky130_fd_sc_hd__dfxtp_1 _5657_ (.CLK(clknet_leaf_2_clk),
    .D(_0223_),
    .Q(\as1802.regs[14][15] ));
 sky130_fd_sc_hd__dfxtp_1 _5658_ (.CLK(clknet_leaf_20_clk),
    .D(_0224_),
    .Q(\as1802.regs[13][8] ));
 sky130_fd_sc_hd__dfxtp_1 _5659_ (.CLK(clknet_leaf_19_clk),
    .D(_0225_),
    .Q(\as1802.regs[13][9] ));
 sky130_fd_sc_hd__dfxtp_1 _5660_ (.CLK(clknet_leaf_16_clk),
    .D(_0226_),
    .Q(\as1802.regs[13][10] ));
 sky130_fd_sc_hd__dfxtp_1 _5661_ (.CLK(clknet_leaf_14_clk),
    .D(_0227_),
    .Q(\as1802.regs[13][11] ));
 sky130_fd_sc_hd__dfxtp_1 _5662_ (.CLK(clknet_leaf_13_clk),
    .D(_0228_),
    .Q(\as1802.regs[13][12] ));
 sky130_fd_sc_hd__dfxtp_1 _5663_ (.CLK(clknet_leaf_9_clk),
    .D(_0229_),
    .Q(\as1802.regs[13][13] ));
 sky130_fd_sc_hd__dfxtp_1 _5664_ (.CLK(clknet_leaf_5_clk),
    .D(_0230_),
    .Q(\as1802.regs[13][14] ));
 sky130_fd_sc_hd__dfxtp_1 _5665_ (.CLK(clknet_leaf_1_clk),
    .D(_0231_),
    .Q(\as1802.regs[13][15] ));
 sky130_fd_sc_hd__dfxtp_1 _5666_ (.CLK(clknet_2_3__leaf_clk),
    .D(_0232_),
    .Q(\as1802.regs[12][0] ));
 sky130_fd_sc_hd__dfxtp_1 _5667_ (.CLK(clknet_leaf_35_clk),
    .D(_0233_),
    .Q(\as1802.regs[12][1] ));
 sky130_fd_sc_hd__dfxtp_1 _5668_ (.CLK(clknet_leaf_31_clk),
    .D(_0234_),
    .Q(\as1802.regs[12][2] ));
 sky130_fd_sc_hd__dfxtp_1 _5669_ (.CLK(clknet_leaf_33_clk),
    .D(_0235_),
    .Q(\as1802.regs[12][3] ));
 sky130_fd_sc_hd__dfxtp_1 _5670_ (.CLK(clknet_leaf_26_clk),
    .D(_0236_),
    .Q(\as1802.regs[12][4] ));
 sky130_fd_sc_hd__dfxtp_1 _5671_ (.CLK(clknet_leaf_27_clk),
    .D(_0237_),
    .Q(\as1802.regs[12][5] ));
 sky130_fd_sc_hd__dfxtp_1 _5672_ (.CLK(clknet_leaf_22_clk),
    .D(_0238_),
    .Q(\as1802.regs[12][6] ));
 sky130_fd_sc_hd__dfxtp_1 _5673_ (.CLK(clknet_leaf_16_clk),
    .D(_0239_),
    .Q(\as1802.regs[12][7] ));
 sky130_fd_sc_hd__dfxtp_1 _5674_ (.CLK(clknet_leaf_19_clk),
    .D(_0240_),
    .Q(\as1802.regs[11][8] ));
 sky130_fd_sc_hd__dfxtp_1 _5675_ (.CLK(clknet_leaf_12_clk),
    .D(_0241_),
    .Q(\as1802.regs[11][9] ));
 sky130_fd_sc_hd__dfxtp_1 _5676_ (.CLK(clknet_leaf_15_clk),
    .D(_0242_),
    .Q(\as1802.regs[11][10] ));
 sky130_fd_sc_hd__dfxtp_1 _5677_ (.CLK(clknet_leaf_10_clk),
    .D(_0243_),
    .Q(\as1802.regs[11][11] ));
 sky130_fd_sc_hd__dfxtp_1 _5678_ (.CLK(clknet_leaf_11_clk),
    .D(_0244_),
    .Q(\as1802.regs[11][12] ));
 sky130_fd_sc_hd__dfxtp_1 _5679_ (.CLK(clknet_leaf_11_clk),
    .D(_0245_),
    .Q(\as1802.regs[11][13] ));
 sky130_fd_sc_hd__dfxtp_1 _5680_ (.CLK(clknet_leaf_10_clk),
    .D(_0246_),
    .Q(\as1802.regs[11][14] ));
 sky130_fd_sc_hd__dfxtp_1 _5681_ (.CLK(clknet_leaf_1_clk),
    .D(_0247_),
    .Q(\as1802.regs[11][15] ));
 sky130_fd_sc_hd__dfxtp_4 _5682_ (.CLK(clknet_leaf_39_clk),
    .D(_0248_),
    .Q(\as1802.mem_cycle[0] ));
 sky130_fd_sc_hd__dfxtp_4 _5683_ (.CLK(clknet_leaf_39_clk),
    .D(_0249_),
    .Q(\as1802.mem_cycle[1] ));
 sky130_fd_sc_hd__dfxtp_4 _5684_ (.CLK(clknet_leaf_39_clk),
    .D(_0250_),
    .Q(\as1802.mem_cycle[2] ));
 sky130_fd_sc_hd__dfxtp_1 _5685_ (.CLK(clknet_leaf_41_clk),
    .D(_0251_),
    .Q(\as1802.addr_buff[0] ));
 sky130_fd_sc_hd__dfxtp_1 _5686_ (.CLK(clknet_leaf_39_clk),
    .D(_0252_),
    .Q(\as1802.addr_buff[1] ));
 sky130_fd_sc_hd__dfxtp_1 _5687_ (.CLK(clknet_leaf_39_clk),
    .D(_0253_),
    .Q(\as1802.addr_buff[2] ));
 sky130_fd_sc_hd__dfxtp_1 _5688_ (.CLK(clknet_leaf_41_clk),
    .D(_0254_),
    .Q(\as1802.addr_buff[3] ));
 sky130_fd_sc_hd__dfxtp_1 _5689_ (.CLK(clknet_leaf_41_clk),
    .D(_0255_),
    .Q(\as1802.addr_buff[4] ));
 sky130_fd_sc_hd__dfxtp_1 _5690_ (.CLK(clknet_leaf_42_clk),
    .D(_0256_),
    .Q(\as1802.addr_buff[5] ));
 sky130_fd_sc_hd__dfxtp_1 _5691_ (.CLK(clknet_leaf_39_clk),
    .D(_0257_),
    .Q(\as1802.addr_buff[6] ));
 sky130_fd_sc_hd__dfxtp_1 _5692_ (.CLK(clknet_leaf_38_clk),
    .D(_0258_),
    .Q(\as1802.addr_buff[7] ));
 sky130_fd_sc_hd__dfxtp_1 _5693_ (.CLK(clknet_leaf_41_clk),
    .D(_0259_),
    .Q(\as1802.addr_buff[8] ));
 sky130_fd_sc_hd__dfxtp_1 _5694_ (.CLK(clknet_leaf_40_clk),
    .D(_0260_),
    .Q(\as1802.addr_buff[9] ));
 sky130_fd_sc_hd__dfxtp_1 _5695_ (.CLK(clknet_leaf_41_clk),
    .D(_0261_),
    .Q(\as1802.addr_buff[10] ));
 sky130_fd_sc_hd__dfxtp_1 _5696_ (.CLK(clknet_leaf_31_clk),
    .D(_0262_),
    .Q(\as1802.addr_buff[11] ));
 sky130_fd_sc_hd__dfxtp_1 _5697_ (.CLK(clknet_leaf_42_clk),
    .D(_0263_),
    .Q(\as1802.addr_buff[12] ));
 sky130_fd_sc_hd__dfxtp_1 _5698_ (.CLK(clknet_leaf_41_clk),
    .D(_0264_),
    .Q(\as1802.addr_buff[13] ));
 sky130_fd_sc_hd__dfxtp_1 _5699_ (.CLK(clknet_leaf_42_clk),
    .D(_0265_),
    .Q(\as1802.addr_buff[14] ));
 sky130_fd_sc_hd__dfxtp_1 _5700_ (.CLK(clknet_leaf_31_clk),
    .D(_0266_),
    .Q(\as1802.addr_buff[15] ));
 sky130_fd_sc_hd__dfxtp_2 _5701_ (.CLK(clknet_leaf_40_clk),
    .D(_0267_),
    .Q(io_out[13]));
 sky130_fd_sc_hd__dfxtp_2 _5702_ (.CLK(clknet_leaf_40_clk),
    .D(_0268_),
    .Q(io_out[14]));
 sky130_fd_sc_hd__dfxtp_2 _5703_ (.CLK(clknet_leaf_39_clk),
    .D(_0269_),
    .Q(io_out[15]));
 sky130_fd_sc_hd__dfxtp_2 _5704_ (.CLK(clknet_leaf_39_clk),
    .D(_0270_),
    .Q(io_out[16]));
 sky130_fd_sc_hd__dfxtp_2 _5705_ (.CLK(clknet_leaf_39_clk),
    .D(_0271_),
    .Q(io_out[17]));
 sky130_fd_sc_hd__dfxtp_2 _5706_ (.CLK(clknet_leaf_39_clk),
    .D(_0272_),
    .Q(io_out[18]));
 sky130_fd_sc_hd__dfxtp_2 _5707_ (.CLK(clknet_leaf_37_clk),
    .D(_0273_),
    .Q(io_out[19]));
 sky130_fd_sc_hd__dfxtp_2 _5708_ (.CLK(clknet_leaf_37_clk),
    .D(_0274_),
    .Q(io_out[20]));
 sky130_fd_sc_hd__dfxtp_1 _5709_ (.CLK(clknet_leaf_48_clk),
    .D(_0275_),
    .Q(\as1802.instr_latch[0] ));
 sky130_fd_sc_hd__dfxtp_4 _5710_ (.CLK(clknet_leaf_48_clk),
    .D(_0276_),
    .Q(\as1802.instr_latch[1] ));
 sky130_fd_sc_hd__dfxtp_4 _5711_ (.CLK(clknet_leaf_47_clk),
    .D(_0277_),
    .Q(\as1802.instr_latch[2] ));
 sky130_fd_sc_hd__dfxtp_2 _5712_ (.CLK(clknet_leaf_47_clk),
    .D(_0278_),
    .Q(\as1802.cond_inv ));
 sky130_fd_sc_hd__dfxtp_1 _5713_ (.CLK(clknet_leaf_48_clk),
    .D(_0279_),
    .Q(\as1802.instr_latch[4] ));
 sky130_fd_sc_hd__dfxtp_2 _5714_ (.CLK(clknet_leaf_46_clk),
    .D(_0280_),
    .Q(\as1802.instr_latch[5] ));
 sky130_fd_sc_hd__dfxtp_1 _5715_ (.CLK(clknet_leaf_48_clk),
    .D(_0281_),
    .Q(\as1802.instr_latch[6] ));
 sky130_fd_sc_hd__dfxtp_2 _5716_ (.CLK(clknet_leaf_46_clk),
    .D(_0282_),
    .Q(\as1802.instr_latch[7] ));
 sky130_fd_sc_hd__dfxtp_1 _5717_ (.CLK(clknet_leaf_38_clk),
    .D(_0283_),
    .Q(\as1802.last_hi_addr[0] ));
 sky130_fd_sc_hd__dfxtp_1 _5718_ (.CLK(clknet_leaf_37_clk),
    .D(_0284_),
    .Q(\as1802.last_hi_addr[1] ));
 sky130_fd_sc_hd__dfxtp_1 _5719_ (.CLK(clknet_leaf_39_clk),
    .D(_0285_),
    .Q(\as1802.last_hi_addr[2] ));
 sky130_fd_sc_hd__dfxtp_1 _5720_ (.CLK(clknet_leaf_38_clk),
    .D(_0286_),
    .Q(\as1802.last_hi_addr[3] ));
 sky130_fd_sc_hd__dfxtp_1 _5721_ (.CLK(clknet_leaf_38_clk),
    .D(_0287_),
    .Q(\as1802.last_hi_addr[4] ));
 sky130_fd_sc_hd__dfxtp_1 _5722_ (.CLK(clknet_leaf_38_clk),
    .D(_0288_),
    .Q(\as1802.last_hi_addr[5] ));
 sky130_fd_sc_hd__dfxtp_1 _5723_ (.CLK(clknet_leaf_39_clk),
    .D(_0289_),
    .Q(\as1802.last_hi_addr[6] ));
 sky130_fd_sc_hd__dfxtp_1 _5724_ (.CLK(clknet_leaf_37_clk),
    .D(_0290_),
    .Q(\as1802.last_hi_addr[7] ));
 sky130_fd_sc_hd__dfxtp_1 _5725_ (.CLK(clknet_leaf_45_clk),
    .D(_0291_),
    .Q(\as1802.will_interrupt ));
 sky130_fd_sc_hd__dfxtp_2 _5726_ (.CLK(clknet_leaf_44_clk),
    .D(_0292_),
    .Q(\as1802.IE ));
 sky130_fd_sc_hd__dfxtp_1 _5727_ (.CLK(clknet_leaf_45_clk),
    .D(_0293_),
    .Q(\as1802.idle ));
 sky130_fd_sc_hd__dfxtp_2 _5728_ (.CLK(clknet_leaf_39_clk),
    .D(_0294_),
    .Q(io_oeb));
 sky130_fd_sc_hd__dfxtp_2 _5729_ (.CLK(clknet_leaf_37_clk),
    .D(_0295_),
    .Q(io_out[22]));
 sky130_fd_sc_hd__dfxtp_2 _5730_ (.CLK(clknet_leaf_37_clk),
    .D(_0296_),
    .Q(io_out[24]));
 sky130_fd_sc_hd__dfxtp_4 _5731_ (.CLK(clknet_leaf_45_clk),
    .D(_0297_),
    .Q(io_out[21]));
 sky130_fd_sc_hd__dfxtp_1 _5732_ (.CLK(clknet_leaf_3_clk),
    .D(_0008_),
    .Q(\as1802.EF_l[0] ));
 sky130_fd_sc_hd__dfxtp_1 _5733_ (.CLK(clknet_leaf_3_clk),
    .D(_0009_),
    .Q(\as1802.EF_l[1] ));
 sky130_fd_sc_hd__dfxtp_1 _5734_ (.CLK(clknet_leaf_3_clk),
    .D(_0010_),
    .Q(\as1802.EF_l[2] ));
 sky130_fd_sc_hd__dfxtp_1 _5735_ (.CLK(clknet_leaf_7_clk),
    .D(_0011_),
    .Q(\as1802.EF_l[3] ));
 sky130_fd_sc_hd__dfxtp_1 _5736_ (.CLK(clknet_leaf_44_clk),
    .D(_0298_),
    .Q(\as1802.lda ));
 sky130_fd_sc_hd__dfxtp_2 _5737_ (.CLK(clknet_leaf_47_clk),
    .D(_0299_),
    .Q(\as1802.DF ));
 sky130_fd_sc_hd__dfxtp_2 _5738_ (.CLK(clknet_leaf_40_clk),
    .D(_0300_),
    .Q(\as1802.X[0] ));
 sky130_fd_sc_hd__dfxtp_2 _5739_ (.CLK(clknet_leaf_40_clk),
    .D(_0301_),
    .Q(\as1802.X[1] ));
 sky130_fd_sc_hd__dfxtp_2 _5740_ (.CLK(clknet_leaf_41_clk),
    .D(_0302_),
    .Q(\as1802.X[2] ));
 sky130_fd_sc_hd__dfxtp_2 _5741_ (.CLK(clknet_leaf_41_clk),
    .D(_0303_),
    .Q(\as1802.X[3] ));
 sky130_fd_sc_hd__dfxtp_1 _5742_ (.CLK(clknet_leaf_40_clk),
    .D(_0304_),
    .Q(\as1802.T[0] ));
 sky130_fd_sc_hd__dfxtp_1 _5743_ (.CLK(clknet_leaf_40_clk),
    .D(_0305_),
    .Q(\as1802.T[1] ));
 sky130_fd_sc_hd__dfxtp_1 _5744_ (.CLK(clknet_leaf_40_clk),
    .D(_0306_),
    .Q(\as1802.T[2] ));
 sky130_fd_sc_hd__dfxtp_1 _5745_ (.CLK(clknet_leaf_45_clk),
    .D(_0307_),
    .Q(\as1802.T[3] ));
 sky130_fd_sc_hd__dfxtp_1 _5746_ (.CLK(clknet_leaf_40_clk),
    .D(_0308_),
    .Q(\as1802.T[4] ));
 sky130_fd_sc_hd__dfxtp_1 _5747_ (.CLK(clknet_leaf_45_clk),
    .D(_0309_),
    .Q(\as1802.T[5] ));
 sky130_fd_sc_hd__dfxtp_1 _5748_ (.CLK(clknet_leaf_41_clk),
    .D(_0310_),
    .Q(\as1802.T[6] ));
 sky130_fd_sc_hd__dfxtp_1 _5749_ (.CLK(clknet_leaf_41_clk),
    .D(_0311_),
    .Q(\as1802.T[7] ));
 sky130_fd_sc_hd__dfxtp_1 _5750_ (.CLK(clknet_leaf_49_clk),
    .D(_0312_),
    .Q(\as1802.D[0] ));
 sky130_fd_sc_hd__dfxtp_2 _5751_ (.CLK(clknet_leaf_49_clk),
    .D(_0313_),
    .Q(\as1802.D[1] ));
 sky130_fd_sc_hd__dfxtp_1 _5752_ (.CLK(clknet_leaf_49_clk),
    .D(_0314_),
    .Q(\as1802.D[2] ));
 sky130_fd_sc_hd__dfxtp_1 _5753_ (.CLK(clknet_leaf_49_clk),
    .D(_0315_),
    .Q(\as1802.D[3] ));
 sky130_fd_sc_hd__dfxtp_1 _5754_ (.CLK(clknet_leaf_50_clk),
    .D(_0316_),
    .Q(\as1802.D[4] ));
 sky130_fd_sc_hd__dfxtp_1 _5755_ (.CLK(clknet_leaf_2_clk),
    .D(_0317_),
    .Q(\as1802.D[5] ));
 sky130_fd_sc_hd__dfxtp_1 _5756_ (.CLK(clknet_leaf_50_clk),
    .D(_0318_),
    .Q(\as1802.D[6] ));
 sky130_fd_sc_hd__dfxtp_4 _5757_ (.CLK(clknet_leaf_0_clk),
    .D(_0319_),
    .Q(\as1802.D[7] ));
 sky130_fd_sc_hd__dfxtp_1 _5758_ (.CLK(clknet_leaf_40_clk),
    .D(_0320_),
    .Q(\as1802.P[0] ));
 sky130_fd_sc_hd__dfxtp_1 _5759_ (.CLK(clknet_leaf_44_clk),
    .D(_0321_),
    .Q(\as1802.P[1] ));
 sky130_fd_sc_hd__dfxtp_1 _5760_ (.CLK(clknet_leaf_41_clk),
    .D(_0322_),
    .Q(\as1802.P[2] ));
 sky130_fd_sc_hd__dfxtp_2 _5761_ (.CLK(clknet_leaf_44_clk),
    .D(_0323_),
    .Q(\as1802.P[3] ));
 sky130_fd_sc_hd__dfxtp_4 _5762_ (.CLK(clknet_leaf_49_clk),
    .D(_0324_),
    .Q(io_out[0]));
 sky130_fd_sc_hd__dfxtp_4 _5763_ (.CLK(clknet_leaf_49_clk),
    .D(_0325_),
    .Q(io_out[1]));
 sky130_fd_sc_hd__dfxtp_4 _5764_ (.CLK(clknet_leaf_49_clk),
    .D(_0326_),
    .Q(io_out[2]));
 sky130_fd_sc_hd__dfxtp_4 _5765_ (.CLK(clknet_leaf_48_clk),
    .D(_0327_),
    .Q(io_out[3]));
 sky130_fd_sc_hd__dfxtp_4 _5766_ (.CLK(clknet_leaf_48_clk),
    .D(_0328_),
    .Q(io_out[4]));
 sky130_fd_sc_hd__dfxtp_4 _5767_ (.CLK(clknet_leaf_48_clk),
    .D(_0329_),
    .Q(io_out[5]));
 sky130_fd_sc_hd__dfxtp_4 _5768_ (.CLK(clknet_leaf_48_clk),
    .D(_0330_),
    .Q(io_out[6]));
 sky130_fd_sc_hd__dfxtp_4 _5769_ (.CLK(clknet_leaf_48_clk),
    .D(_0331_),
    .Q(io_out[7]));
 sky130_fd_sc_hd__dfxtp_1 _5770_ (.CLK(clknet_leaf_19_clk),
    .D(_0332_),
    .Q(\as1802.regs[9][8] ));
 sky130_fd_sc_hd__dfxtp_1 _5771_ (.CLK(clknet_leaf_12_clk),
    .D(_0333_),
    .Q(\as1802.regs[9][9] ));
 sky130_fd_sc_hd__dfxtp_1 _5772_ (.CLK(clknet_leaf_15_clk),
    .D(_0334_),
    .Q(\as1802.regs[9][10] ));
 sky130_fd_sc_hd__dfxtp_1 _5773_ (.CLK(clknet_leaf_14_clk),
    .D(_0335_),
    .Q(\as1802.regs[9][11] ));
 sky130_fd_sc_hd__dfxtp_1 _5774_ (.CLK(clknet_leaf_12_clk),
    .D(_0336_),
    .Q(\as1802.regs[9][12] ));
 sky130_fd_sc_hd__dfxtp_1 _5775_ (.CLK(clknet_leaf_8_clk),
    .D(_0337_),
    .Q(\as1802.regs[9][13] ));
 sky130_fd_sc_hd__dfxtp_1 _5776_ (.CLK(clknet_leaf_10_clk),
    .D(_0338_),
    .Q(\as1802.regs[9][14] ));
 sky130_fd_sc_hd__dfxtp_1 _5777_ (.CLK(clknet_leaf_1_clk),
    .D(_0339_),
    .Q(\as1802.regs[9][15] ));
 sky130_fd_sc_hd__dfxtp_2 _5778_ (.CLK(clknet_leaf_15_clk),
    .D(_0340_),
    .Q(\as1802.regs[2][8] ));
 sky130_fd_sc_hd__dfxtp_2 _5779_ (.CLK(clknet_leaf_15_clk),
    .D(_0341_),
    .Q(\as1802.regs[2][9] ));
 sky130_fd_sc_hd__dfxtp_2 _5780_ (.CLK(clknet_leaf_15_clk),
    .D(_0342_),
    .Q(\as1802.regs[2][10] ));
 sky130_fd_sc_hd__dfxtp_2 _5781_ (.CLK(clknet_leaf_1_clk),
    .D(_0343_),
    .Q(\as1802.regs[2][11] ));
 sky130_fd_sc_hd__dfxtp_2 _5782_ (.CLK(clknet_leaf_14_clk),
    .D(_0344_),
    .Q(\as1802.regs[2][12] ));
 sky130_fd_sc_hd__dfxtp_2 _5783_ (.CLK(clknet_leaf_1_clk),
    .D(_0345_),
    .Q(\as1802.regs[2][13] ));
 sky130_fd_sc_hd__dfxtp_2 _5784_ (.CLK(clknet_leaf_2_clk),
    .D(_0346_),
    .Q(\as1802.regs[2][14] ));
 sky130_fd_sc_hd__dfxtp_2 _5785_ (.CLK(clknet_leaf_2_clk),
    .D(_0347_),
    .Q(\as1802.regs[2][15] ));
 sky130_fd_sc_hd__dfxtp_1 _5786_ (.CLK(clknet_leaf_44_clk),
    .D(_0348_),
    .Q(\as1802.mem_write ));
 sky130_fd_sc_hd__dfxtp_1 _5787_ (.CLK(clknet_leaf_16_clk),
    .D(_0349_),
    .Q(\as1802.regs[1][8] ));
 sky130_fd_sc_hd__dfxtp_1 _5788_ (.CLK(clknet_leaf_13_clk),
    .D(_0350_),
    .Q(\as1802.regs[1][9] ));
 sky130_fd_sc_hd__dfxtp_1 _5789_ (.CLK(clknet_leaf_15_clk),
    .D(_0351_),
    .Q(\as1802.regs[1][10] ));
 sky130_fd_sc_hd__dfxtp_1 _5790_ (.CLK(clknet_leaf_14_clk),
    .D(_0352_),
    .Q(\as1802.regs[1][11] ));
 sky130_fd_sc_hd__dfxtp_1 _5791_ (.CLK(clknet_leaf_13_clk),
    .D(_0353_),
    .Q(\as1802.regs[1][12] ));
 sky130_fd_sc_hd__dfxtp_1 _5792_ (.CLK(clknet_leaf_10_clk),
    .D(_0354_),
    .Q(\as1802.regs[1][13] ));
 sky130_fd_sc_hd__dfxtp_1 _5793_ (.CLK(clknet_leaf_5_clk),
    .D(_0355_),
    .Q(\as1802.regs[1][14] ));
 sky130_fd_sc_hd__dfxtp_1 _5794_ (.CLK(clknet_leaf_2_clk),
    .D(_0356_),
    .Q(\as1802.regs[1][15] ));
 sky130_fd_sc_hd__dfxtp_2 _5795_ (.CLK(clknet_leaf_46_clk),
    .D(_0357_),
    .Q(io_out[25]));
 sky130_fd_sc_hd__dfxtp_2 _5796_ (.CLK(clknet_leaf_45_clk),
    .D(_0358_),
    .Q(io_out[26]));
 sky130_fd_sc_hd__conb_1 wrapped_as1802_16 (.LO(net16));
 sky130_fd_sc_hd__conb_1 wrapped_as1802_17 (.LO(net17));
 sky130_fd_sc_hd__conb_1 wrapped_as1802_18 (.LO(net18));
 sky130_fd_sc_hd__conb_1 wrapped_as1802_19 (.LO(net19));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_0_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_0_clk));
 sky130_fd_sc_hd__buf_2 _5802_ (.A(io_oeb),
    .X(io_out[23]));
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__decap_3 PHY_166 ();
 sky130_fd_sc_hd__decap_3 PHY_167 ();
 sky130_fd_sc_hd__decap_3 PHY_168 ();
 sky130_fd_sc_hd__decap_3 PHY_169 ();
 sky130_fd_sc_hd__decap_3 PHY_170 ();
 sky130_fd_sc_hd__decap_3 PHY_171 ();
 sky130_fd_sc_hd__decap_3 PHY_172 ();
 sky130_fd_sc_hd__decap_3 PHY_173 ();
 sky130_fd_sc_hd__decap_3 PHY_174 ();
 sky130_fd_sc_hd__decap_3 PHY_175 ();
 sky130_fd_sc_hd__decap_3 PHY_176 ();
 sky130_fd_sc_hd__decap_3 PHY_177 ();
 sky130_fd_sc_hd__decap_3 PHY_178 ();
 sky130_fd_sc_hd__decap_3 PHY_179 ();
 sky130_fd_sc_hd__decap_3 PHY_180 ();
 sky130_fd_sc_hd__decap_3 PHY_181 ();
 sky130_fd_sc_hd__decap_3 PHY_182 ();
 sky130_fd_sc_hd__decap_3 PHY_183 ();
 sky130_fd_sc_hd__decap_3 PHY_184 ();
 sky130_fd_sc_hd__decap_3 PHY_185 ();
 sky130_fd_sc_hd__decap_3 PHY_186 ();
 sky130_fd_sc_hd__decap_3 PHY_187 ();
 sky130_fd_sc_hd__decap_3 PHY_188 ();
 sky130_fd_sc_hd__decap_3 PHY_189 ();
 sky130_fd_sc_hd__decap_3 PHY_190 ();
 sky130_fd_sc_hd__decap_3 PHY_191 ();
 sky130_fd_sc_hd__decap_3 PHY_192 ();
 sky130_fd_sc_hd__decap_3 PHY_193 ();
 sky130_fd_sc_hd__decap_3 PHY_194 ();
 sky130_fd_sc_hd__decap_3 PHY_195 ();
 sky130_fd_sc_hd__decap_3 PHY_196 ();
 sky130_fd_sc_hd__decap_3 PHY_197 ();
 sky130_fd_sc_hd__decap_3 PHY_198 ();
 sky130_fd_sc_hd__decap_3 PHY_199 ();
 sky130_fd_sc_hd__decap_3 PHY_200 ();
 sky130_fd_sc_hd__decap_3 PHY_201 ();
 sky130_fd_sc_hd__decap_3 PHY_202 ();
 sky130_fd_sc_hd__decap_3 PHY_203 ();
 sky130_fd_sc_hd__decap_3 PHY_204 ();
 sky130_fd_sc_hd__decap_3 PHY_205 ();
 sky130_fd_sc_hd__decap_3 PHY_206 ();
 sky130_fd_sc_hd__decap_3 PHY_207 ();
 sky130_fd_sc_hd__decap_3 PHY_208 ();
 sky130_fd_sc_hd__decap_3 PHY_209 ();
 sky130_fd_sc_hd__decap_3 PHY_210 ();
 sky130_fd_sc_hd__decap_3 PHY_211 ();
 sky130_fd_sc_hd__decap_3 PHY_212 ();
 sky130_fd_sc_hd__decap_3 PHY_213 ();
 sky130_fd_sc_hd__decap_3 PHY_214 ();
 sky130_fd_sc_hd__decap_3 PHY_215 ();
 sky130_fd_sc_hd__decap_3 PHY_216 ();
 sky130_fd_sc_hd__decap_3 PHY_217 ();
 sky130_fd_sc_hd__decap_3 PHY_218 ();
 sky130_fd_sc_hd__decap_3 PHY_219 ();
 sky130_fd_sc_hd__decap_3 PHY_220 ();
 sky130_fd_sc_hd__decap_3 PHY_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1577 ();
 sky130_fd_sc_hd__dlymetal6s2s_1 input1 (.A(io_in[0]),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(io_in[10]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(io_in[11]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(io_in[12]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(io_in[1]),
    .X(net5));
 sky130_fd_sc_hd__dlymetal6s2s_1 input6 (.A(io_in[2]),
    .X(net6));
 sky130_fd_sc_hd__dlymetal6s2s_1 input7 (.A(io_in[3]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_2 input8 (.A(io_in[4]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_2 input9 (.A(io_in[5]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_2 input10 (.A(io_in[6]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_2 input11 (.A(io_in[7]),
    .X(net11));
 sky130_fd_sc_hd__buf_2 input12 (.A(io_in[8]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_1 input13 (.A(io_in[9]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_4 input14 (.A(rst),
    .X(net14));
 sky130_fd_sc_hd__conb_1 wrapped_as1802_15 (.LO(net15));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_1_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_1_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_2_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_2_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_3_clk (.A(clknet_opt_1_0_clk),
    .X(clknet_leaf_3_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_4_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_4_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_5_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_5_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_6_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_6_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_7_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_7_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_8_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_8_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_9_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_9_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_10_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_10_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_11_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_11_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_12_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_12_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_13_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_13_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_14_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_14_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_15_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_15_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_16_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_16_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_17_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_17_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_18_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_18_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_19_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_19_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_20_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_20_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_21_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_21_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_22_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_22_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_23_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_23_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_24_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_24_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_25_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_25_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_26_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_26_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_27_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_27_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_28_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_28_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_30_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_30_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_31_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_31_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_32_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_32_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_33_clk (.A(clknet_opt_2_0_clk),
    .X(clknet_leaf_33_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_34_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_34_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_35_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_35_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_36_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_36_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_37_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_37_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_38_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_38_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_39_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_39_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_40_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_40_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_41_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_41_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_42_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_42_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_44_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_44_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_45_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_45_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_46_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_46_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_47_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_47_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_48_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_48_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_49_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_49_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_50_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_50_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_0__f_clk (.A(clknet_0_clk),
    .X(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_1__f_clk (.A(clknet_0_clk),
    .X(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_2__f_clk (.A(clknet_0_clk),
    .X(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_3__f_clk (.A(clknet_0_clk),
    .X(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_1_0_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_opt_1_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_2_0_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_opt_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__3304__S0 (.DIODE(_0000_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3303__S0 (.DIODE(_0000_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3233__S0 (.DIODE(_0000_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3232__S0 (.DIODE(_0000_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3098__A (.DIODE(_0000_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2943__A (.DIODE(_0000_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3304__S1 (.DIODE(_0001_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3303__S1 (.DIODE(_0001_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3298__B1_N (.DIODE(_0001_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3233__S1 (.DIODE(_0001_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3232__S1 (.DIODE(_0001_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3227__B1_N (.DIODE(_0001_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3106__S1 (.DIODE(_0001_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2946__A (.DIODE(_0001_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3499__B2 (.DIODE(_0003_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3406__B2 (.DIODE(_0003_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3373__B2 (.DIODE(_0003_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3306__B2 (.DIODE(_0003_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3235__B2 (.DIODE(_0003_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3160__A1 (.DIODE(_0003_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3159__B1 (.DIODE(_0003_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3108__B2 (.DIODE(_0003_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2966__A (.DIODE(_0003_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2941__A (.DIODE(_0003_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3994__B1 (.DIODE(_0366_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3940__B1 (.DIODE(_0366_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3834__A1 (.DIODE(_0366_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3775__A1 (.DIODE(_0366_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3513__A1 (.DIODE(_0366_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3417__A1 (.DIODE(_0366_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3387__A1 (.DIODE(_0366_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3321__A1 (.DIODE(_0366_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3247__A1 (.DIODE(_0366_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3006__C1 (.DIODE(_0366_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3649__A (.DIODE(_0379_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3123__C1 (.DIODE(_0379_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3045__A2 (.DIODE(_0379_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3043__A2 (.DIODE(_0379_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3039__A2 (.DIODE(_0379_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3019__A (.DIODE(_0379_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3947__A1 (.DIODE(_0380_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3777__A1 (.DIODE(_0380_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3713__A1 (.DIODE(_0380_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3578__C1 (.DIODE(_0380_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3514__B2 (.DIODE(_0380_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3445__A1 (.DIODE(_0380_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3389__A1 (.DIODE(_0380_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3249__A1 (.DIODE(_0380_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3038__A2 (.DIODE(_0380_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3020__C1 (.DIODE(_0380_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5334__B2 (.DIODE(_0382_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5117__B2 (.DIODE(_0382_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5115__A1 (.DIODE(_0382_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5022__A1 (.DIODE(_0382_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4979__A (.DIODE(_0382_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4977__A (.DIODE(_0382_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4955__B (.DIODE(_0382_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4951__A (.DIODE(_0382_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3585__A1 (.DIODE(_0382_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3031__A1 (.DIODE(_0382_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3488__A1 (.DIODE(_0384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3487__B (.DIODE(_0384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3362__A1 (.DIODE(_0384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3295__C1 (.DIODE(_0384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3224__C1 (.DIODE(_0384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3181__A2 (.DIODE(_0384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3124__A2 (.DIODE(_0384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3049__C (.DIODE(_0384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3035__A (.DIODE(_0384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3031__A2 (.DIODE(_0384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5113__A (.DIODE(_0385_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4590__C (.DIODE(_0385_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3581__B (.DIODE(_0385_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3025__B (.DIODE(_0385_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4000__A1 (.DIODE(_0390_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3999__B1 (.DIODE(_0390_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3896__C1 (.DIODE(_0390_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3716__A1 (.DIODE(_0390_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3030__B (.DIODE(_0390_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3871__B1 (.DIODE(_0397_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3488__C1 (.DIODE(_0397_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3443__B1 (.DIODE(_0397_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3290__A (.DIODE(_0397_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3225__B1 (.DIODE(_0397_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3045__B1 (.DIODE(_0397_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3043__B1 (.DIODE(_0397_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3039__B1 (.DIODE(_0397_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3037__A2 (.DIODE(_0397_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4068__A (.DIODE(_0399_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4010__B (.DIODE(_0399_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3588__A (.DIODE(_0399_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3041__A_N (.DIODE(_0399_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4068__B (.DIODE(_0401_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4010__A_N (.DIODE(_0401_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3588__B (.DIODE(_0401_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3041__B (.DIODE(_0401_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4508__B (.DIODE(_0411_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4418__B (.DIODE(_0411_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4382__B (.DIODE(_0411_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4364__B (.DIODE(_0411_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4292__B (.DIODE(_0411_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4141__A (.DIODE(_0411_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3051__C (.DIODE(_0411_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3518__S (.DIODE(_0413_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3452__S (.DIODE(_0413_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3395__S (.DIODE(_0413_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3327__S (.DIODE(_0413_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3256__S (.DIODE(_0413_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3191__S (.DIODE(_0413_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3128__S (.DIODE(_0413_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3053__S (.DIODE(_0413_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3895__A (.DIODE(_0415_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3579__C1 (.DIODE(_0415_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3056__A (.DIODE(_0415_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4001__D1 (.DIODE(_0416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3844__B1 (.DIODE(_0416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3838__B1 (.DIODE(_0416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3835__B1 (.DIODE(_0416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3597__B1 (.DIODE(_0416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3520__B1 (.DIODE(_0416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3455__B1 (.DIODE(_0416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3323__C1 (.DIODE(_0416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3253__B (.DIODE(_0416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3126__A1 (.DIODE(_0416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3436__B1 (.DIODE(_0437_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3352__A (.DIODE(_0437_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3341__B1 (.DIODE(_0437_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3284__B1 (.DIODE(_0437_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3211__B1 (.DIODE(_0437_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3148__A1 (.DIODE(_0437_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3078__B1 (.DIODE(_0437_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5130__B (.DIODE(_0439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4639__B2 (.DIODE(_0439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4638__B2 (.DIODE(_0439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4634__A2 (.DIODE(_0439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3219__A2 (.DIODE(_0439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3218__B (.DIODE(_0439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3214__A2 (.DIODE(_0439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3213__B (.DIODE(_0439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3081__B (.DIODE(_0439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3080__B (.DIODE(_0439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5105__A1 (.DIODE(_0444_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3095__B (.DIODE(_0444_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3085__B (.DIODE(_0444_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3976__A1 (.DIODE(_0447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3945__A1 (.DIODE(_0447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3944__B1 (.DIODE(_0447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3751__A1 (.DIODE(_0447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3688__A1 (.DIODE(_0447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3687__B1 (.DIODE(_0447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3584__A1 (.DIODE(_0447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3359__S (.DIODE(_0447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3295__A1 (.DIODE(_0447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3091__A2 (.DIODE(_0447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3651__A1 (.DIODE(_0450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3514__A1 (.DIODE(_0450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3446__B2 (.DIODE(_0450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3130__A (.DIODE(_0450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3091__B1 (.DIODE(_0450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5345__A1 (.DIODE(_0452_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5152__B2 (.DIODE(_0452_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5147__A1 (.DIODE(_0452_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5092__A1 (.DIODE(_0452_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5085__A (.DIODE(_0452_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4931__A (.DIODE(_0452_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4930__A1 (.DIODE(_0452_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4924__A (.DIODE(_0452_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3653__A (.DIODE(_0452_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3124__A1 (.DIODE(_0452_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5185__A (.DIODE(_0453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5023__A1 (.DIODE(_0453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4995__A (.DIODE(_0453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3941__A (.DIODE(_0453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3827__S (.DIODE(_0453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3710__A1 (.DIODE(_0453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3709__A (.DIODE(_0453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3648__A1 (.DIODE(_0453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3175__A (.DIODE(_0453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3094__A (.DIODE(_0453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3779__B1 (.DIODE(_0454_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3715__A (.DIODE(_0454_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3651__B2 (.DIODE(_0454_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3489__A (.DIODE(_0454_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3446__A1 (.DIODE(_0454_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3388__A1 (.DIODE(_0454_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3096__A (.DIODE(_0454_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3298__A1 (.DIODE(_0458_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3297__A_N (.DIODE(_0458_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3227__A1 (.DIODE(_0458_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3226__A_N (.DIODE(_0458_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3156__S0 (.DIODE(_0458_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3154__S (.DIODE(_0458_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3152__A_N (.DIODE(_0458_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3101__S (.DIODE(_0458_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3100__A1 (.DIODE(_0458_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3099__A_N (.DIODE(_0458_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4639__A1_N (.DIODE(_0469_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4635__A0 (.DIODE(_0469_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4633__B (.DIODE(_0469_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3236__A (.DIODE(_0469_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3165__A (.DIODE(_0469_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3162__A2 (.DIODE(_0469_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3118__B (.DIODE(_0469_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3115__B (.DIODE(_0469_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3111__B (.DIODE(_0469_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3110__B (.DIODE(_0469_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5347__A0 (.DIODE(_0474_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5132__A (.DIODE(_0474_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5001__A (.DIODE(_0474_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5000__A (.DIODE(_0474_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4975__B (.DIODE(_0474_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4929__A (.DIODE(_0474_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4242__A1_N (.DIODE(_0474_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3645__A1 (.DIODE(_0474_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3121__A (.DIODE(_0474_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3116__A0 (.DIODE(_0474_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4512__A1 (.DIODE(_0486_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4458__A1 (.DIODE(_0486_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4440__A1 (.DIODE(_0486_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4422__A1 (.DIODE(_0486_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4386__A1 (.DIODE(_0486_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4368__A1 (.DIODE(_0486_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3127__A (.DIODE(_0486_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5162__A2 (.DIODE(_0507_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4650__A2 (.DIODE(_0507_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4649__A1 (.DIODE(_0507_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4642__A0 (.DIODE(_0507_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3219__A3 (.DIODE(_0507_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3218__C (.DIODE(_0507_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3214__A3 (.DIODE(_0507_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3213__C (.DIODE(_0507_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3184__B (.DIODE(_0507_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3149__B (.DIODE(_0507_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3307__B (.DIODE(_0519_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3236__B (.DIODE(_0519_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3165__B (.DIODE(_0519_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3162__B1 (.DIODE(_0519_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3161__B (.DIODE(_0519_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4650__B1 (.DIODE(_0523_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4643__A0 (.DIODE(_0523_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4642__A1 (.DIODE(_0523_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3167__A0 (.DIODE(_0523_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4922__B (.DIODE(_0527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4920__B (.DIODE(_0527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3174__A1 (.DIODE(_0527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3169__A0 (.DIODE(_0527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5350__A1 (.DIODE(_0539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5189__B2 (.DIODE(_0539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5179__A1 (.DIODE(_0539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5160__A1 (.DIODE(_0539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5117__A1 (.DIODE(_0539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4974__A (.DIODE(_0539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4922__A (.DIODE(_0539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4920__A (.DIODE(_0539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3689__A (.DIODE(_0539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3181__A1 (.DIODE(_0539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4514__A1 (.DIODE(_0548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4460__A1 (.DIODE(_0548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4442__A1 (.DIODE(_0548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4424__A1 (.DIODE(_0548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4388__A1 (.DIODE(_0548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4370__A1 (.DIODE(_0548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3190__A (.DIODE(_0548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4334__A1 (.DIODE(_0549_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4316__A1 (.DIODE(_0549_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4298__A1 (.DIODE(_0549_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4280__A1 (.DIODE(_0549_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4262__A1 (.DIODE(_0549_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4202__A1 (.DIODE(_0549_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4184__A1 (.DIODE(_0549_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4166__A1 (.DIODE(_0549_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4148__A1 (.DIODE(_0549_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3191__A1 (.DIODE(_0549_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3473__C1 (.DIODE(_0560_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3459__C1 (.DIODE(_0560_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3435__C1 (.DIODE(_0560_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3423__C1 (.DIODE(_0560_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3340__A1 (.DIODE(_0560_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3335__C1 (.DIODE(_0560_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3332__C1 (.DIODE(_0560_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3281__A (.DIODE(_0560_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3260__A (.DIODE(_0560_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3206__A1 (.DIODE(_0560_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5207__A0 (.DIODE(_0570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4661__A2 (.DIODE(_0570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4660__A1 (.DIODE(_0570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4654__A2 (.DIODE(_0570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3219__B1 (.DIODE(_0570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3218__D (.DIODE(_0570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3214__B1 (.DIODE(_0570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3213__D (.DIODE(_0570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3923__A1 (.DIODE(_0575_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3780__A1 (.DIODE(_0575_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3580__A1 (.DIODE(_0575_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3388__B2 (.DIODE(_0575_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3324__A1 (.DIODE(_0575_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3250__A1 (.DIODE(_0575_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5355__A1 (.DIODE(_0579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5216__B2 (.DIODE(_0579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5211__A1 (.DIODE(_0579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5205__A1 (.DIODE(_0579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5152__A1 (.DIODE(_0579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4973__A (.DIODE(_0579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4917__B (.DIODE(_0579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4915__A_N (.DIODE(_0579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3753__A (.DIODE(_0579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3225__A1 (.DIODE(_0579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4662__A1 (.DIODE(_0593_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4656__B (.DIODE(_0593_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4653__B (.DIODE(_0593_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3307__C (.DIODE(_0593_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3240__B1 (.DIODE(_0593_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3239__A1 (.DIODE(_0593_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3237__B (.DIODE(_0593_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3236__C (.DIODE(_0593_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4516__A1 (.DIODE(_0612_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4462__A1 (.DIODE(_0612_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4444__A1 (.DIODE(_0612_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4426__A1 (.DIODE(_0612_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4390__A1 (.DIODE(_0612_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4372__A1 (.DIODE(_0612_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3255__A (.DIODE(_0612_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3604__C1 (.DIODE(_0617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3545__A (.DIODE(_0617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3523__A (.DIODE(_0617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3471__A1 (.DIODE(_0617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3464__A1 (.DIODE(_0617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3431__A1 (.DIODE(_0617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3421__A1 (.DIODE(_0617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3278__A1 (.DIODE(_0617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3273__A1 (.DIODE(_0617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3266__A1 (.DIODE(_0617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3466__A (.DIODE(_0618_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3418__S (.DIODE(_0618_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3347__A2 (.DIODE(_0618_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3345__A2 (.DIODE(_0618_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3343__A2 (.DIODE(_0618_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3332__A2 (.DIODE(_0618_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3330__S (.DIODE(_0618_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3275__A (.DIODE(_0618_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3267__S (.DIODE(_0618_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3262__S (.DIODE(_0618_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3475__C1 (.DIODE(_0628_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3470__C1 (.DIODE(_0628_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3463__C1 (.DIODE(_0628_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3433__C1 (.DIODE(_0628_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3429__C1 (.DIODE(_0628_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3425__C1 (.DIODE(_0628_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3420__C1 (.DIODE(_0628_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3283__A (.DIODE(_0628_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3277__C1 (.DIODE(_0628_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3272__C1 (.DIODE(_0628_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3537__A (.DIODE(_0632_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3524__A (.DIODE(_0632_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3475__A2 (.DIODE(_0632_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3465__S (.DIODE(_0632_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3463__A2 (.DIODE(_0632_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3459__A2 (.DIODE(_0632_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3435__A2 (.DIODE(_0632_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3433__A2 (.DIODE(_0632_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3429__A2 (.DIODE(_0632_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3277__A2 (.DIODE(_0632_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3861__B1 (.DIODE(_0636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3800__C1 (.DIODE(_0636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3611__C1 (.DIODE(_0636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3607__A1 (.DIODE(_0636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3543__A (.DIODE(_0636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3532__C1 (.DIODE(_0636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3476__A1 (.DIODE(_0636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3460__C1 (.DIODE(_0636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3436__A1 (.DIODE(_0636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3284__A1 (.DIODE(_0636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5224__A2 (.DIODE(_0642_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4667__A2 (.DIODE(_0642_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3621__B (.DIODE(_0642_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3482__B (.DIODE(_0642_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3480__B (.DIODE(_0642_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3439__B (.DIODE(_0642_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3356__A2 (.DIODE(_0642_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3355__B (.DIODE(_0642_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3287__B (.DIODE(_0642_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3286__B (.DIODE(_0642_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5360__A1 (.DIODE(_0646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5247__B_N (.DIODE(_0646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5243__B2 (.DIODE(_0646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5241__A1 (.DIODE(_0646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5221__A1 (.DIODE(_0646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5189__A1 (.DIODE(_0646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4972__A (.DIODE(_0646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4909__A (.DIODE(_0646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3810__A1 (.DIODE(_0646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3296__A1 (.DIODE(_0646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3970__A1 (.DIODE(_0648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3918__A1 (.DIODE(_0648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3854__B1 (.DIODE(_0648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3796__B1 (.DIODE(_0648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3749__A1 (.DIODE(_0648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3743__A1 (.DIODE(_0648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3670__B1 (.DIODE(_0648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3607__B1 (.DIODE(_0648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3549__B1 (.DIODE(_0648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3292__A1 (.DIODE(_0648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4674__A2 (.DIODE(_0649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4673__A1 (.DIODE(_0649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3456__A (.DIODE(_0649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3293__B (.DIODE(_0649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4675__A1 (.DIODE(_0663_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4670__B (.DIODE(_0663_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4666__B (.DIODE(_0663_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3312__B1 (.DIODE(_0663_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3311__A1 (.DIODE(_0663_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3309__B (.DIODE(_0663_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3307__D (.DIODE(_0663_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4518__A1 (.DIODE(_0682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4464__A1 (.DIODE(_0682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4446__A1 (.DIODE(_0682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4428__A1 (.DIODE(_0682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4392__A1 (.DIODE(_0682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4374__A1 (.DIODE(_0682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3326__A (.DIODE(_0682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3803__C1 (.DIODE(_0685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3799__C1 (.DIODE(_0685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3735__A (.DIODE(_0685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3613__C1 (.DIODE(_0685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3610__C1 (.DIODE(_0685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3606__C1 (.DIODE(_0685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3601__C1 (.DIODE(_0685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3530__A (.DIODE(_0685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3460__A1 (.DIODE(_0685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3333__A1 (.DIODE(_0685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3349__A2 (.DIODE(_0693_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3339__B (.DIODE(_0693_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3338__A2 (.DIODE(_0693_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3969__C1 (.DIODE(_0708_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3917__C1 (.DIODE(_0708_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3863__B2 (.DIODE(_0708_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3805__A (.DIODE(_0708_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3742__B1 (.DIODE(_0708_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3679__B1 (.DIODE(_0708_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3616__B1 (.DIODE(_0708_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3550__A1 (.DIODE(_0708_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3476__B1 (.DIODE(_0708_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3353__B2 (.DIODE(_0708_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5256__A2 (.DIODE(_0709_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3479__A (.DIODE(_0709_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3456__B (.DIODE(_0709_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3354__A (.DIODE(_0709_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4687__A2 (.DIODE(_0710_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4685__A1 (.DIODE(_0710_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4679__A2 (.DIODE(_0710_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3482__C (.DIODE(_0710_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3439__C (.DIODE(_0710_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3358__B (.DIODE(_0710_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3356__B1 (.DIODE(_0710_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3355__C (.DIODE(_0710_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5365__A1 (.DIODE(_0716_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5277__B2 (.DIODE(_0716_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5269__A1 (.DIODE(_0716_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5253__A1 (.DIODE(_0716_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5216__A1 (.DIODE(_0716_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4971__A (.DIODE(_0716_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4906__B (.DIODE(_0716_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4901__A_N (.DIODE(_0716_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3871__A1 (.DIODE(_0716_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3361__A1 (.DIODE(_0716_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4686__A1 (.DIODE(_0729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4681__B (.DIODE(_0729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4678__B (.DIODE(_0729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3505__A3 (.DIODE(_0729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3502__A2 (.DIODE(_0729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3500__B (.DIODE(_0729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3379__B1 (.DIODE(_0729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3377__A1 (.DIODE(_0729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3375__B (.DIODE(_0729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3374__B (.DIODE(_0729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4340__A1 (.DIODE(_0750_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4322__A1 (.DIODE(_0750_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4304__A1 (.DIODE(_0750_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4286__A1 (.DIODE(_0750_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4268__A1 (.DIODE(_0750_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4208__A1 (.DIODE(_0750_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4190__A1 (.DIODE(_0750_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4172__A1 (.DIODE(_0750_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4154__A1 (.DIODE(_0750_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3395__A1 (.DIODE(_0750_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4697__A1 (.DIODE(_0761_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4693__A2 (.DIODE(_0761_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4689__B (.DIODE(_0761_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3505__A4 (.DIODE(_0761_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3502__A3 (.DIODE(_0761_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3500__C (.DIODE(_0761_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3410__B (.DIODE(_0761_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3409__A1 (.DIODE(_0761_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3407__B (.DIODE(_0761_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3804__C1 (.DIODE(_0785_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3674__A (.DIODE(_0785_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3665__C1 (.DIODE(_0785_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3616__A1 (.DIODE(_0785_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3602__C1 (.DIODE(_0785_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3542__C1 (.DIODE(_0785_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3536__C1 (.DIODE(_0785_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3471__C1 (.DIODE(_0785_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3464__C1 (.DIODE(_0785_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3431__C1 (.DIODE(_0785_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5294__A0 (.DIODE(_0792_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4696__A2 (.DIODE(_0792_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4695__A1 (.DIODE(_0792_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4692__A2 (.DIODE(_0792_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4690__A2 (.DIODE(_0792_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3482__D_N (.DIODE(_0792_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3479__B (.DIODE(_0792_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3456__C (.DIODE(_0792_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3440__B (.DIODE(_0792_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3438__B (.DIODE(_0792_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5370__A1 (.DIODE(_0797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5317__B2 (.DIODE(_0797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5303__A1 (.DIODE(_0797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5297__A1 (.DIODE(_0797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5292__A1 (.DIODE(_0797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5243__A1 (.DIODE(_0797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4970__A (.DIODE(_0797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4894__A (.DIODE(_0797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3946__A1 (.DIODE(_0797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3443__A1 (.DIODE(_0797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4522__A1 (.DIODE(_0805_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4468__A1 (.DIODE(_0805_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4450__A1 (.DIODE(_0805_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4432__A1 (.DIODE(_0805_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4396__A1 (.DIODE(_0805_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4378__A1 (.DIODE(_0805_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3451__A (.DIODE(_0805_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3797__S (.DIODE(_0820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3740__S (.DIODE(_0820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3738__S (.DIODE(_0820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3677__S (.DIODE(_0820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3676__S (.DIODE(_0820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3599__S (.DIODE(_0820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3539__A (.DIODE(_0820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3526__A (.DIODE(_0820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3473__A2 (.DIODE(_0820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3470__A2 (.DIODE(_0820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3802__B (.DIODE(_0821_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3798__B (.DIODE(_0821_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3661__A (.DIODE(_0821_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3605__B (.DIODE(_0821_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3603__B (.DIODE(_0821_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3600__B (.DIODE(_0821_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3527__A (.DIODE(_0821_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3474__B (.DIODE(_0821_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3472__B (.DIODE(_0821_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3469__B (.DIODE(_0821_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3802__C (.DIODE(_0822_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3798__C (.DIODE(_0822_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3662__A (.DIODE(_0822_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3605__C (.DIODE(_0822_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3603__C (.DIODE(_0822_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3600__C (.DIODE(_0822_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3528__A (.DIODE(_0822_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3474__C (.DIODE(_0822_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3472__C (.DIODE(_0822_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3469__C (.DIODE(_0822_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5310__B (.DIODE(_0831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4706__A1 (.DIODE(_0831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3865__B (.DIODE(_0831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3846__B (.DIODE(_0831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3745__B (.DIODE(_0831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3619__B (.DIODE(_0831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3618__A2 (.DIODE(_0831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3522__B (.DIODE(_0831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3479__C_N (.DIODE(_0831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3478__A (.DIODE(_0831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4707__A2 (.DIODE(_0832_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4700__A0 (.DIODE(_0832_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3722__B (.DIODE(_0832_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3484__B (.DIODE(_0832_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3481__A2 (.DIODE(_0832_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5325__A1_N (.DIODE(_0840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4897__A (.DIODE(_0840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4895__A (.DIODE(_0840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4893__A (.DIODE(_0840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3487__A (.DIODE(_0840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4708__A1 (.DIODE(_0853_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4703__A2 (.DIODE(_0853_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4700__A1 (.DIODE(_0853_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3505__B1 (.DIODE(_0853_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3504__A1 (.DIODE(_0853_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3502__B1 (.DIODE(_0853_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3500__D (.DIODE(_0853_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4524__A1 (.DIODE(_0870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4470__A1 (.DIODE(_0870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4452__A1 (.DIODE(_0870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4434__A1 (.DIODE(_0870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4398__A1 (.DIODE(_0870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4380__A1 (.DIODE(_0870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3517__A (.DIODE(_0870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4344__A1 (.DIODE(_0871_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4326__A1 (.DIODE(_0871_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4308__A1 (.DIODE(_0871_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4290__A1 (.DIODE(_0871_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4272__A1 (.DIODE(_0871_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4212__A1 (.DIODE(_0871_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4194__A1 (.DIODE(_0871_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4176__A1 (.DIODE(_0871_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4158__A1 (.DIODE(_0871_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3518__A1 (.DIODE(_0871_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3861__A1 (.DIODE(_0876_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3804__A1 (.DIODE(_0876_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3731__A1 (.DIODE(_0876_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3727__A1 (.DIODE(_0876_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3675__A1 (.DIODE(_0876_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3665__A1 (.DIODE(_0876_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3611__A1 (.DIODE(_0876_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3542__A1 (.DIODE(_0876_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3536__A1 (.DIODE(_0876_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3532__A1 (.DIODE(_0876_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3856__S (.DIODE(_0877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3855__S (.DIODE(_0877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3852__S (.DIODE(_0877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3801__S (.DIODE(_0877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3794__S (.DIODE(_0877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3793__S (.DIODE(_0877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3724__A (.DIODE(_0877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3608__S (.DIODE(_0877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3533__S (.DIODE(_0877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3525__S (.DIODE(_0877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3730__C1 (.DIODE(_0883_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3726__C1 (.DIODE(_0883_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3678__S (.DIODE(_0883_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3673__C1 (.DIODE(_0883_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3667__C1 (.DIODE(_0883_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3664__C1 (.DIODE(_0883_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3548__C1 (.DIODE(_0883_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3541__C1 (.DIODE(_0883_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3535__C1 (.DIODE(_0883_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3531__C1 (.DIODE(_0883_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3966__S (.DIODE(_0890_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3860__S (.DIODE(_0890_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3858__S (.DIODE(_0890_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3851__S (.DIODE(_0890_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3803__A2 (.DIODE(_0890_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3799__A2 (.DIODE(_0890_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3606__A2 (.DIODE(_0890_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3604__A2 (.DIODE(_0890_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3601__A2 (.DIODE(_0890_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3538__S (.DIODE(_0890_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3959__S (.DIODE(_0892_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3956__S (.DIODE(_0892_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3733__S (.DIODE(_0892_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3728__S (.DIODE(_0892_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3723__S (.DIODE(_0892_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3673__A2 (.DIODE(_0892_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3669__A2 (.DIODE(_0892_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3667__A2 (.DIODE(_0892_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3664__A2 (.DIODE(_0892_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3541__A2 (.DIODE(_0892_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3968__C1 (.DIODE(_0896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3917__A1 (.DIODE(_0896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3905__C1 (.DIODE(_0896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3850__C1 (.DIODE(_0896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3796__A1 (.DIODE(_0896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3742__A1 (.DIODE(_0896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3727__C1 (.DIODE(_0896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3679__A1 (.DIODE(_0896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3670__A1 (.DIODE(_0896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3549__A1 (.DIODE(_0896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3857__S (.DIODE(_0898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3853__S (.DIODE(_0898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3800__A1 (.DIODE(_0898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3795__S (.DIODE(_0898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3739__A (.DIODE(_0898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3732__A (.DIODE(_0898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3669__C1 (.DIODE(_0898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3615__C1 (.DIODE(_0898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3602__A1 (.DIODE(_0898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3546__C1 (.DIODE(_0898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5090__A2 (.DIODE(_0904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4717__A2 (.DIODE(_0904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4716__A1 (.DIODE(_0904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4711__A0 (.DIODE(_0904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3745__C (.DIODE(_0904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3721__A (.DIODE(_0904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3619__C (.DIODE(_0904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3618__A3 (.DIODE(_0904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3553__B (.DIODE(_0904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3552__B (.DIODE(_0904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3819__S1 (.DIODE(_0911_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3818__S1 (.DIODE(_0911_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3813__B1_N (.DIODE(_0911_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3762__S1 (.DIODE(_0911_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3761__S1 (.DIODE(_0911_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3759__S1 (.DIODE(_0911_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3756__B1_N (.DIODE(_0911_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3693__B2 (.DIODE(_0911_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3632__S1 (.DIODE(_0911_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3560__B2 (.DIODE(_0911_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3986__S (.DIODE(_0912_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3981__C1 (.DIODE(_0912_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3932__C1 (.DIODE(_0912_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3883__C1 (.DIODE(_0912_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3815__C1 (.DIODE(_0912_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3763__S (.DIODE(_0912_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3758__C1 (.DIODE(_0912_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3693__C1 (.DIODE(_0912_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3630__C1 (.DIODE(_0912_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3560__C1 (.DIODE(_0912_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4717__B1 (.DIODE(_0919_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4712__A0 (.DIODE(_0919_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4711__A1 (.DIODE(_0919_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3575__B (.DIODE(_0919_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3571__B1 (.DIODE(_0919_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3567__A (.DIODE(_0919_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5420__A1 (.DIODE(_0939_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5399__A1 (.DIODE(_0939_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5381__A1 (.DIODE(_0939_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4528__A1 (.DIODE(_0939_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4492__A1 (.DIODE(_0939_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4474__A1 (.DIODE(_0939_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3587__A (.DIODE(_0939_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5379__A (.DIODE(_0943_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4526__B (.DIODE(_0943_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4436__C (.DIODE(_0943_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4418__C (.DIODE(_0943_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4160__B (.DIODE(_0943_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4142__B (.DIODE(_0943_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4031__A (.DIODE(_0943_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3593__B (.DIODE(_0943_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5397__B (.DIODE(_0945_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5379__B (.DIODE(_0945_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4526__C (.DIODE(_0945_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4472__C (.DIODE(_0945_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4346__C (.DIODE(_0945_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4009__A (.DIODE(_0945_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3593__C (.DIODE(_0945_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4007__S (.DIODE(_0947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3953__S (.DIODE(_0947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3900__S (.DIODE(_0947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3841__S (.DIODE(_0947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3786__S (.DIODE(_0947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3719__S (.DIODE(_0947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3657__S (.DIODE(_0947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3595__S (.DIODE(_0947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4726__A2 (.DIODE(_0969_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4720__A0 (.DIODE(_0969_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3721__B (.DIODE(_0969_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3686__A2 (.DIODE(_0969_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3683__A (.DIODE(_0969_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3623__B (.DIODE(_0969_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3619__D (.DIODE(_0969_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3618__B1 (.DIODE(_0969_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3877__A (.DIODE(_0977_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3816__S0 (.DIODE(_0977_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3814__S (.DIODE(_0977_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3812__A_N (.DIODE(_0977_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3759__S0 (.DIODE(_0977_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3757__S (.DIODE(_0977_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3754__A_N (.DIODE(_0977_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3628__S (.DIODE(_0977_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3627__A1 (.DIODE(_0977_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3626__A_N (.DIODE(_0977_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3930__B1_N (.DIODE(_0981_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3926__S1 (.DIODE(_0981_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3881__B1_N (.DIODE(_0981_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3878__A (.DIODE(_0981_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3875__S1 (.DIODE(_0981_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3874__S1 (.DIODE(_0981_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3816__S1 (.DIODE(_0981_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3815__B2 (.DIODE(_0981_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3758__B2 (.DIODE(_0981_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3630__B2 (.DIODE(_0981_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3983__A1 (.DIODE(_0983_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3933__A1 (.DIODE(_0983_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3927__S (.DIODE(_0983_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3884__A1 (.DIODE(_0983_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3876__S (.DIODE(_0983_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3820__S (.DIODE(_0983_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3817__A1 (.DIODE(_0983_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3760__A1 (.DIODE(_0983_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3636__S (.DIODE(_0983_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3633__A1 (.DIODE(_0983_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3702__C (.DIODE(_0989_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3646__A (.DIODE(_0989_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3643__B (.DIODE(_0989_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3642__A3 (.DIODE(_0989_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3639__D (.DIODE(_0989_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3638__B1 (.DIODE(_0989_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5422__A1 (.DIODE(_1007_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5401__A1 (.DIODE(_1007_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5383__A1 (.DIODE(_1007_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4530__A1 (.DIODE(_1007_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4494__A1 (.DIODE(_1007_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4476__A1 (.DIODE(_1007_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3656__A (.DIODE(_1007_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3914__B (.DIODE(_1012_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3907__B (.DIODE(_1012_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3903__B (.DIODE(_1012_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3848__B (.DIODE(_1012_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3790__B (.DIODE(_1012_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3734__B (.DIODE(_1012_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3729__B (.DIODE(_1012_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3725__B (.DIODE(_1012_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3672__B (.DIODE(_1012_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3663__B (.DIODE(_1012_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3914__C (.DIODE(_1013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3907__C (.DIODE(_1013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3903__C (.DIODE(_1013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3848__C (.DIODE(_1013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3790__C (.DIODE(_1013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3734__C (.DIODE(_1013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3729__C (.DIODE(_1013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3725__C (.DIODE(_1013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3672__C (.DIODE(_1013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3663__C (.DIODE(_1013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3969__A1 (.DIODE(_1025_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3961__S (.DIODE(_1025_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3916__C1 (.DIODE(_1025_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3909__C1 (.DIODE(_1025_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3862__A1 (.DIODE(_1025_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3854__A1 (.DIODE(_1025_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3792__C1 (.DIODE(_1025_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3737__C1 (.DIODE(_1025_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3731__C1 (.DIODE(_1025_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3675__C1 (.DIODE(_1025_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5161__A2 (.DIODE(_1032_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4736__A2 (.DIODE(_1032_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4735__A1 (.DIODE(_1032_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4732__A2 (.DIODE(_1032_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4730__A2 (.DIODE(_1032_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3747__B (.DIODE(_1032_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3722__D (.DIODE(_1032_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3686__B1_N (.DIODE(_1032_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3684__B (.DIODE(_1032_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3682__B (.DIODE(_1032_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5129__A0 (.DIODE(_1034_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4725__A1 (.DIODE(_1034_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3747__A (.DIODE(_1034_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3744__A (.DIODE(_1034_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3684__A (.DIODE(_1034_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4731__B (.DIODE(_1050_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4729__B (.DIODE(_1050_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3825__B (.DIODE(_1050_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3709__B (.DIODE(_1050_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3706__A2 (.DIODE(_1050_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3701__A (.DIODE(_1050_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3700__B (.DIODE(_1050_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3965__S (.DIODE(_1074_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3963__S (.DIODE(_1074_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3962__S (.DIODE(_1074_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3958__S (.DIODE(_1074_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3955__S (.DIODE(_1074_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3847__S (.DIODE(_1074_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3788__S (.DIODE(_1074_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3736__A2 (.DIODE(_1074_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3730__A2 (.DIODE(_1074_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3726__A2 (.DIODE(_1074_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3968__A1 (.DIODE(_1082_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3964__S (.DIODE(_1082_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3960__S (.DIODE(_1082_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3957__S (.DIODE(_1082_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3916__A1 (.DIODE(_1082_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3909__A1 (.DIODE(_1082_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3905__A1 (.DIODE(_1082_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3850__A1 (.DIODE(_1082_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3792__A1 (.DIODE(_1082_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3737__A1 (.DIODE(_1082_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3967__A (.DIODE(_1085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3915__C1 (.DIODE(_1085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3912__S (.DIODE(_1085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3908__C1 (.DIODE(_1085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3904__C1 (.DIODE(_1085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3859__A (.DIODE(_1085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3849__C1 (.DIODE(_1085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3791__C1 (.DIODE(_1085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3741__A (.DIODE(_1085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3736__C1 (.DIODE(_1085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5206__A2 (.DIODE(_1093_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4745__A1 (.DIODE(_1093_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3845__C (.DIODE(_1093_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3747__C (.DIODE(_1093_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3746__A2 (.DIODE(_1093_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3744__C (.DIODE(_1093_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4747__A2 (.DIODE(_1099_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4740__A1 (.DIODE(_1099_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3750__B1 (.DIODE(_1099_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3990__B (.DIODE(_1114_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3828__A3 (.DIODE(_1114_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3824__A (.DIODE(_1114_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3823__A3 (.DIODE(_1114_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3774__B (.DIODE(_1114_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3767__B (.DIODE(_1114_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3765__A (.DIODE(_1114_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4747__B2 (.DIODE(_1115_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4741__A0 (.DIODE(_1115_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4740__A0 (.DIODE(_1115_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3769__B (.DIODE(_1115_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3766__B (.DIODE(_1115_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4408__A1 (.DIODE(_1135_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4354__A1 (.DIODE(_1135_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4131__A1 (.DIODE(_1135_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4113__A1 (.DIODE(_1135_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4095__A1 (.DIODE(_1135_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4077__A1 (.DIODE(_1135_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4058__A1 (.DIODE(_1135_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4039__A1 (.DIODE(_1135_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4021__A1 (.DIODE(_1135_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3786__A1 (.DIODE(_1135_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3915__A2 (.DIODE(_1138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3913__S (.DIODE(_1138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3911__S (.DIODE(_1138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3910__S (.DIODE(_1138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3908__A2 (.DIODE(_1138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3906__S (.DIODE(_1138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3904__A2 (.DIODE(_1138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3902__S (.DIODE(_1138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3849__A2 (.DIODE(_1138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3791__A2 (.DIODE(_1138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5223__A2 (.DIODE(_1155_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4755__A2 (.DIODE(_1155_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4754__B2 (.DIODE(_1155_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4749__A0 (.DIODE(_1155_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3869__A3 (.DIODE(_1155_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3867__A (.DIODE(_1155_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3864__A (.DIODE(_1155_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3846__D (.DIODE(_1155_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3808__B (.DIODE(_1155_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3807__B (.DIODE(_1155_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3990__C (.DIODE(_1170_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3828__B1 (.DIODE(_1170_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3824__B (.DIODE(_1170_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3823__B1 (.DIODE(_1170_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3822__A (.DIODE(_1170_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4755__B1 (.DIODE(_1171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4750__A0 (.DIODE(_1171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4749__A1 (.DIODE(_1171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3827__A0 (.DIODE(_1171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5254__B (.DIODE(_1211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4764__A2 (.DIODE(_1211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4763__A1 (.DIODE(_1211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4758__A0 (.DIODE(_1211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3896__A2 (.DIODE(_1211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3869__B1 (.DIODE(_1211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3867__B (.DIODE(_1211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3866__A2 (.DIODE(_1211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3864__B (.DIODE(_1211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3985__S0 (.DIODE(_1225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3984__S0 (.DIODE(_1225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3982__S0 (.DIODE(_1225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3980__S (.DIODE(_1225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3979__A1 (.DIODE(_1225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3978__A_N (.DIODE(_1225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3930__A1 (.DIODE(_1225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3928__S0 (.DIODE(_1225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3925__S0 (.DIODE(_1225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3879__S0 (.DIODE(_1225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3985__S1 (.DIODE(_1226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3984__S1 (.DIODE(_1226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3982__S1 (.DIODE(_1226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3981__B2 (.DIODE(_1226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3979__B1_N (.DIODE(_1226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3932__B2 (.DIODE(_1226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3928__S1 (.DIODE(_1226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3925__S1 (.DIODE(_1226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3883__B2 (.DIODE(_1226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3879__S1 (.DIODE(_1226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4764__B1 (.DIODE(_1233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4759__A0 (.DIODE(_1233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4758__A1 (.DIODE(_1233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3989__A (.DIODE(_1233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3924__B (.DIODE(_1233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3889__C (.DIODE(_1233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3888__B1 (.DIODE(_1233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3887__A0 (.DIODE(_1233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3886__B (.DIODE(_1233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5430__A1 (.DIODE(_1246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5409__A1 (.DIODE(_1246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5391__A1 (.DIODE(_1246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4538__A1 (.DIODE(_1246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4502__A1 (.DIODE(_1246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4484__A1 (.DIODE(_1246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3899__A (.DIODE(_1246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5293__A2_N (.DIODE(_1265_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4773__A2 (.DIODE(_1265_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4772__A1 (.DIODE(_1265_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4767__A0 (.DIODE(_1265_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3973__C (.DIODE(_1265_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3972__A3 (.DIODE(_1265_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3921__B1 (.DIODE(_1265_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3920__D (.DIODE(_1265_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3919__B (.DIODE(_1265_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4773__B1 (.DIODE(_1281_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4768__A0 (.DIODE(_1281_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4767__A1 (.DIODE(_1281_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3989__B (.DIODE(_1281_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3942__B (.DIODE(_1281_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3937__B (.DIODE(_1281_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3936__B (.DIODE(_1281_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3935__B (.DIODE(_1281_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4892__A1 (.DIODE(_1288_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4732__A1 (.DIODE(_1288_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4720__S (.DIODE(_1288_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4692__A1 (.DIODE(_1288_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4679__A1 (.DIODE(_1288_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4678__A (.DIODE(_1288_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4634__A1 (.DIODE(_1288_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4611__A (.DIODE(_1288_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3943__A1 (.DIODE(_1288_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3942__A (.DIODE(_1288_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5432__A1 (.DIODE(_1298_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5411__A1 (.DIODE(_1298_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5393__A1 (.DIODE(_1298_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4540__A1 (.DIODE(_1298_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4504__A1 (.DIODE(_1298_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4486__A1 (.DIODE(_1298_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3952__A (.DIODE(_1298_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5308__B (.DIODE(_1316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4784__A2 (.DIODE(_1316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4776__A0 (.DIODE(_1316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3975__B (.DIODE(_1316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3971__A (.DIODE(_1316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4782__A1 (.DIODE(_1317_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3973__D (.DIODE(_1317_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3972__B1 (.DIODE(_1317_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4779__B (.DIODE(_1333_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3995__A0 (.DIODE(_1333_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3993__A0 (.DIODE(_1333_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3992__A0 (.DIODE(_1333_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3988__A (.DIODE(_1333_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4784__B1 (.DIODE(_1334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4776__A1 (.DIODE(_1334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3991__A (.DIODE(_1334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4029__S (.DIODE(_1359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4027__S (.DIODE(_1359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4025__S (.DIODE(_1359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4023__S (.DIODE(_1359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4021__S (.DIODE(_1359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4019__S (.DIODE(_1359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4017__S (.DIODE(_1359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4015__S (.DIODE(_1359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4047__S (.DIODE(_1369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4045__S (.DIODE(_1369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4043__S (.DIODE(_1369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4041__S (.DIODE(_1369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4039__S (.DIODE(_1369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4037__S (.DIODE(_1369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4035__S (.DIODE(_1369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4033__S (.DIODE(_1369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4066__S (.DIODE(_1380_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4064__S (.DIODE(_1380_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4062__S (.DIODE(_1380_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4060__S (.DIODE(_1380_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4058__S (.DIODE(_1380_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4056__S (.DIODE(_1380_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4054__S (.DIODE(_1380_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4052__S (.DIODE(_1380_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4085__S (.DIODE(_1391_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4083__S (.DIODE(_1391_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4081__S (.DIODE(_1391_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4079__S (.DIODE(_1391_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4077__S (.DIODE(_1391_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4075__S (.DIODE(_1391_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4073__S (.DIODE(_1391_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4071__S (.DIODE(_1391_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4103__S (.DIODE(_1401_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4101__S (.DIODE(_1401_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4099__S (.DIODE(_1401_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4097__S (.DIODE(_1401_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4095__S (.DIODE(_1401_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4093__S (.DIODE(_1401_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4091__S (.DIODE(_1401_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4089__S (.DIODE(_1401_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4121__S (.DIODE(_1411_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4119__S (.DIODE(_1411_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4117__S (.DIODE(_1411_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4115__S (.DIODE(_1411_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4113__S (.DIODE(_1411_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4111__S (.DIODE(_1411_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4109__S (.DIODE(_1411_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4107__S (.DIODE(_1411_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4139__S (.DIODE(_1421_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4137__S (.DIODE(_1421_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4135__S (.DIODE(_1421_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4133__S (.DIODE(_1421_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4131__S (.DIODE(_1421_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4129__S (.DIODE(_1421_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4127__S (.DIODE(_1421_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4125__S (.DIODE(_1421_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4158__S (.DIODE(_1432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4156__S (.DIODE(_1432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4154__S (.DIODE(_1432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4152__S (.DIODE(_1432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4150__S (.DIODE(_1432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4148__S (.DIODE(_1432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4146__S (.DIODE(_1432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4144__S (.DIODE(_1432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4176__S (.DIODE(_1442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4174__S (.DIODE(_1442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4172__S (.DIODE(_1442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4170__S (.DIODE(_1442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4168__S (.DIODE(_1442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4166__S (.DIODE(_1442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4164__S (.DIODE(_1442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4162__S (.DIODE(_1442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4194__S (.DIODE(_1452_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4192__S (.DIODE(_1452_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4190__S (.DIODE(_1452_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4188__S (.DIODE(_1452_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4186__S (.DIODE(_1452_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4184__S (.DIODE(_1452_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4182__S (.DIODE(_1452_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4180__S (.DIODE(_1452_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4212__S (.DIODE(_1462_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4210__S (.DIODE(_1462_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4208__S (.DIODE(_1462_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4206__S (.DIODE(_1462_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4204__S (.DIODE(_1462_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4202__S (.DIODE(_1462_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4200__S (.DIODE(_1462_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4198__S (.DIODE(_1462_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4773__B2 (.DIODE(_1475_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4726__B2 (.DIODE(_1475_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4624__A (.DIODE(_1475_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4220__A2 (.DIODE(_1475_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5053__A1 (.DIODE(_1489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4863__A1 (.DIODE(_1489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4854__A1 (.DIODE(_1489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4737__B2 (.DIODE(_1489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4708__B2 (.DIODE(_1489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4697__B2 (.DIODE(_1489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4675__B2 (.DIODE(_1489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4248__A1 (.DIODE(_1489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4242__B2 (.DIODE(_1489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4236__A (.DIODE(_1489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5224__C1 (.DIODE(_1490_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5208__A (.DIODE(_1490_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4734__A1 (.DIODE(_1490_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4693__B1 (.DIODE(_1490_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4683__C1 (.DIODE(_1490_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4669__C1 (.DIODE(_1490_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4646__A (.DIODE(_1490_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4636__B2 (.DIODE(_1490_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4620__A1 (.DIODE(_1490_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4234__A (.DIODE(_1490_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5323__A1 (.DIODE(_1491_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5209__A1 (.DIODE(_1491_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5048__A (.DIODE(_1491_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5044__S (.DIODE(_1491_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5027__C1 (.DIODE(_1491_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4877__A (.DIODE(_1491_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4743__C1 (.DIODE(_1491_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4614__C1 (.DIODE(_1491_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4247__B (.DIODE(_1491_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4235__S (.DIODE(_1491_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4853__A (.DIODE(_1494_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4848__A (.DIODE(_1494_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4834__A (.DIODE(_1494_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4802__C1 (.DIODE(_1494_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4799__C1 (.DIODE(_1494_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4796__C1 (.DIODE(_1494_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4793__C1 (.DIODE(_1494_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4790__C1 (.DIODE(_1494_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4249__C1 (.DIODE(_1494_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4238__C1 (.DIODE(_1494_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5162__B1 (.DIODE(_1495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5091__C1 (.DIODE(_1495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5056__A1 (.DIODE(_1495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4880__B (.DIODE(_1495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4780__C1 (.DIODE(_1495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4771__A1 (.DIODE(_1495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4684__A1 (.DIODE(_1495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4617__C1 (.DIODE(_1495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4252__A2 (.DIODE(_1495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4240__A (.DIODE(_1495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5052__A (.DIODE(_1496_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5037__B1 (.DIODE(_1496_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4762__A1 (.DIODE(_1496_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4753__A1 (.DIODE(_1496_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4744__A1 (.DIODE(_1496_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4724__A1 (.DIODE(_1496_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4715__A1 (.DIODE(_1496_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4648__A1 (.DIODE(_1496_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4246__B (.DIODE(_1496_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4241__B (.DIODE(_1496_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4879__A (.DIODE(_1499_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4875__A (.DIODE(_1499_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4870__B1 (.DIODE(_1499_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4864__A (.DIODE(_1499_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4860__C1 (.DIODE(_1499_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4845__A (.DIODE(_1499_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4842__A (.DIODE(_1499_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4839__A (.DIODE(_1499_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4836__A (.DIODE(_1499_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4244__B1 (.DIODE(_1499_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5081__B1 (.DIODE(_1504_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5079__B1 (.DIODE(_1504_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5077__A (.DIODE(_1504_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5074__A (.DIODE(_1504_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5071__A (.DIODE(_1504_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5068__A (.DIODE(_1504_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5065__A (.DIODE(_1504_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5062__A (.DIODE(_1504_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5058__A (.DIODE(_1504_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4254__A (.DIODE(_1504_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4272__S (.DIODE(_1510_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4270__S (.DIODE(_1510_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4268__S (.DIODE(_1510_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4266__S (.DIODE(_1510_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4264__S (.DIODE(_1510_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4262__S (.DIODE(_1510_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4260__S (.DIODE(_1510_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4258__S (.DIODE(_1510_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4290__S (.DIODE(_1520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4288__S (.DIODE(_1520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4286__S (.DIODE(_1520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4284__S (.DIODE(_1520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4282__S (.DIODE(_1520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4280__S (.DIODE(_1520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4278__S (.DIODE(_1520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4276__S (.DIODE(_1520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4308__S (.DIODE(_1530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4306__S (.DIODE(_1530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4304__S (.DIODE(_1530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4302__S (.DIODE(_1530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4300__S (.DIODE(_1530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4298__S (.DIODE(_1530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4296__S (.DIODE(_1530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4294__S (.DIODE(_1530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4326__S (.DIODE(_1540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4324__S (.DIODE(_1540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4322__S (.DIODE(_1540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4320__S (.DIODE(_1540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4318__S (.DIODE(_1540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4316__S (.DIODE(_1540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4314__S (.DIODE(_1540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4312__S (.DIODE(_1540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4344__S (.DIODE(_1550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4342__S (.DIODE(_1550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4340__S (.DIODE(_1550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4338__S (.DIODE(_1550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4336__S (.DIODE(_1550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4334__S (.DIODE(_1550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4332__S (.DIODE(_1550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4330__S (.DIODE(_1550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4362__S (.DIODE(_1560_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4360__S (.DIODE(_1560_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4358__S (.DIODE(_1560_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4356__S (.DIODE(_1560_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4354__S (.DIODE(_1560_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4352__S (.DIODE(_1560_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4350__S (.DIODE(_1560_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4348__S (.DIODE(_1560_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4380__S (.DIODE(_1570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4378__S (.DIODE(_1570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4376__S (.DIODE(_1570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4374__S (.DIODE(_1570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4372__S (.DIODE(_1570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4370__S (.DIODE(_1570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4368__S (.DIODE(_1570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4366__S (.DIODE(_1570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4398__S (.DIODE(_1580_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4396__S (.DIODE(_1580_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4394__S (.DIODE(_1580_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4392__S (.DIODE(_1580_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4390__S (.DIODE(_1580_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4388__S (.DIODE(_1580_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4386__S (.DIODE(_1580_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4384__S (.DIODE(_1580_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4416__S (.DIODE(_1590_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4414__S (.DIODE(_1590_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4412__S (.DIODE(_1590_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4410__S (.DIODE(_1590_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4408__S (.DIODE(_1590_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4406__S (.DIODE(_1590_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4404__S (.DIODE(_1590_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4402__S (.DIODE(_1590_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4434__S (.DIODE(_1600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4432__S (.DIODE(_1600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4430__S (.DIODE(_1600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4428__S (.DIODE(_1600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4426__S (.DIODE(_1600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4424__S (.DIODE(_1600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4422__S (.DIODE(_1600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4420__S (.DIODE(_1600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4452__S (.DIODE(_1610_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4450__S (.DIODE(_1610_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4448__S (.DIODE(_1610_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4446__S (.DIODE(_1610_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4444__S (.DIODE(_1610_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4442__S (.DIODE(_1610_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4440__S (.DIODE(_1610_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4438__S (.DIODE(_1610_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4470__S (.DIODE(_1620_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4468__S (.DIODE(_1620_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4466__S (.DIODE(_1620_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4464__S (.DIODE(_1620_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4462__S (.DIODE(_1620_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4460__S (.DIODE(_1620_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4458__S (.DIODE(_1620_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4456__S (.DIODE(_1620_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4488__S (.DIODE(_1630_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4486__S (.DIODE(_1630_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4484__S (.DIODE(_1630_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4482__S (.DIODE(_1630_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4480__S (.DIODE(_1630_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4478__S (.DIODE(_1630_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4476__S (.DIODE(_1630_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4474__S (.DIODE(_1630_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4506__S (.DIODE(_1640_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4504__S (.DIODE(_1640_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4502__S (.DIODE(_1640_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4500__S (.DIODE(_1640_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4498__S (.DIODE(_1640_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4496__S (.DIODE(_1640_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4494__S (.DIODE(_1640_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4492__S (.DIODE(_1640_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4524__S (.DIODE(_1650_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4522__S (.DIODE(_1650_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4520__S (.DIODE(_1650_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4518__S (.DIODE(_1650_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4516__S (.DIODE(_1650_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4514__S (.DIODE(_1650_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4512__S (.DIODE(_1650_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4510__S (.DIODE(_1650_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4542__S (.DIODE(_1660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4540__S (.DIODE(_1660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4538__S (.DIODE(_1660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4536__S (.DIODE(_1660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4534__S (.DIODE(_1660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4532__S (.DIODE(_1660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4530__S (.DIODE(_1660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4528__S (.DIODE(_1660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5308__A (.DIODE(_1695_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5307__C1 (.DIODE(_1695_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5293__A1_N (.DIODE(_1695_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5292__B1 (.DIODE(_1695_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5223__A1 (.DIODE(_1695_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5221__B1 (.DIODE(_1695_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5205__C1 (.DIODE(_1695_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5160__C1 (.DIODE(_1695_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5129__S (.DIODE(_1695_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4571__A2 (.DIODE(_1695_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5416__S (.DIODE(_1726_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4773__C1 (.DIODE(_1726_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4764__C1 (.DIODE(_1726_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4755__C1 (.DIODE(_1726_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4726__C1 (.DIODE(_1726_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4717__C1 (.DIODE(_1726_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4686__B1_N (.DIODE(_1726_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4650__C1 (.DIODE(_1726_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4625__C1 (.DIODE(_1726_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4605__A (.DIODE(_1726_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4784__C1 (.DIODE(_1727_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4747__C1 (.DIODE(_1727_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4738__S (.DIODE(_1727_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4709__S (.DIODE(_1727_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4698__S (.DIODE(_1727_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4688__A2 (.DIODE(_1727_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4676__S (.DIODE(_1727_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4663__S (.DIODE(_1727_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4640__C1 (.DIODE(_1727_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4606__A (.DIODE(_1727_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4785__B2 (.DIODE(_1728_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4775__A2 (.DIODE(_1728_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4766__A2 (.DIODE(_1728_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4757__A2 (.DIODE(_1728_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4748__B2 (.DIODE(_1728_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4728__A2 (.DIODE(_1728_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4719__A2 (.DIODE(_1728_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4652__A2 (.DIODE(_1728_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4641__A2 (.DIODE(_1728_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4627__A2 (.DIODE(_1728_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4881__B1 (.DIODE(_1730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4774__A1 (.DIODE(_1730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4765__A1 (.DIODE(_1730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4756__A1 (.DIODE(_1730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4718__A1 (.DIODE(_1730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4687__B1 (.DIODE(_1730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4686__A2 (.DIODE(_1730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4651__A1 (.DIODE(_1730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4640__A1 (.DIODE(_1730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4626__A1 (.DIODE(_1730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4880__A (.DIODE(_1732_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4768__S (.DIODE(_1732_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4759__S (.DIODE(_1732_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4750__S (.DIODE(_1732_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4741__S (.DIODE(_1732_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4721__S (.DIODE(_1732_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4712__S (.DIODE(_1732_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4643__S (.DIODE(_1732_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4614__A1 (.DIODE(_1732_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4613__A (.DIODE(_1732_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5026__A1 (.DIODE(_1733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4876__C (.DIODE(_1733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4822__A0 (.DIODE(_1733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4776__S (.DIODE(_1733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4767__S (.DIODE(_1733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4758__S (.DIODE(_1733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4749__S (.DIODE(_1733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4711__S (.DIODE(_1733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4642__S (.DIODE(_1733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4612__A1 (.DIODE(_1733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5374__A2 (.DIODE(_1738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5369__A2 (.DIODE(_1738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5364__A2 (.DIODE(_1738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5359__A2 (.DIODE(_1738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5354__A2 (.DIODE(_1738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5349__A2 (.DIODE(_1738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5344__A2 (.DIODE(_1738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5332__A2 (.DIODE(_1738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5060__A1 (.DIODE(_1738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4617__A2 (.DIODE(_1738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5055__S (.DIODE(_1741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4769__A2 (.DIODE(_1741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4760__A2 (.DIODE(_1741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4733__A3 (.DIODE(_1741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4691__A3 (.DIODE(_1741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4682__A2 (.DIODE(_1741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4668__A2 (.DIODE(_1741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4665__A2 (.DIODE(_1741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4631__A (.DIODE(_1741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4620__A3 (.DIODE(_1741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4782__B2 (.DIODE(_1750_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4754__A1_N (.DIODE(_1750_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4745__B2 (.DIODE(_1750_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4735__B2 (.DIODE(_1750_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4725__B2 (.DIODE(_1750_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4705__B1 (.DIODE(_1750_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4695__B2 (.DIODE(_1750_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4673__B2 (.DIODE(_1750_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4638__A1_N (.DIODE(_1750_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5051__S (.DIODE(_1752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5047__S (.DIODE(_1752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5043__S (.DIODE(_1752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4777__A2 (.DIODE(_1752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4751__A2 (.DIODE(_1752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4742__A2 (.DIODE(_1752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4722__A2 (.DIODE(_1752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4713__A2 (.DIODE(_1752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4645__A2 (.DIODE(_1752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4637__A3 (.DIODE(_1752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5295__B2 (.DIODE(_1766_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5256__C1 (.DIODE(_1766_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5131__C1 (.DIODE(_1766_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4778__C1 (.DIODE(_1766_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4770__C1 (.DIODE(_1766_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4761__C1 (.DIODE(_1766_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4752__C1 (.DIODE(_1766_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4723__C1 (.DIODE(_1766_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4714__C1 (.DIODE(_1766_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4647__C1 (.DIODE(_1766_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5106__C (.DIODE(_1911_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4871__A (.DIODE(_1911_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4814__B (.DIODE(_1911_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5321__A (.DIODE(_1966_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5280__A1 (.DIODE(_1966_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5144__A (.DIODE(_1966_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5027__A1 (.DIODE(_1966_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5313__B (.DIODE(_2069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5257__B1 (.DIODE(_2069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5168__B1 (.DIODE(_2069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5140__A0 (.DIODE(_2069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5025__A2 (.DIODE(_2069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5262__A1 (.DIODE(_2097_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5238__A1 (.DIODE(_2097_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5232__A_N (.DIODE(_2097_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5195__B1 (.DIODE(_2097_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5190__C1 (.DIODE(_2097_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5176__A1 (.DIODE(_2097_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5024__B (.DIODE(_2097_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5310__A (.DIODE(_2144_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5309__B1 (.DIODE(_2144_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5294__S (.DIODE(_2144_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5255__C1 (.DIODE(_2144_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5223__C1 (.DIODE(_2144_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5207__S (.DIODE(_2144_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5162__A1 (.DIODE(_2144_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5131__A1 (.DIODE(_2144_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5130__A (.DIODE(_2144_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5091__A1 (.DIODE(_2144_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5099__A1_N (.DIODE(_2152_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5323__C1 (.DIODE(_2158_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5296__B1 (.DIODE(_2158_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5268__A1 (.DIODE(_2158_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5240__B1 (.DIODE(_2158_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5210__B1 (.DIODE(_2158_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5178__A1 (.DIODE(_2158_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5146__A1 (.DIODE(_2158_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5098__B1 (.DIODE(_2158_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5437__B (.DIODE(_2172_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5112__C1 (.DIODE(_2172_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5325__A2_N (.DIODE(_2175_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5324__B1 (.DIODE(_2175_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5297__S (.DIODE(_2175_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5269__S (.DIODE(_2175_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5241__S (.DIODE(_2175_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5211__S (.DIODE(_2175_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5179__S (.DIODE(_2175_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5147__S (.DIODE(_2175_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5115__S (.DIODE(_2175_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5318__A2 (.DIODE(_2195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5265__C1 (.DIODE(_2195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5177__A1 (.DIODE(_2195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5145__A2 (.DIODE(_2195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5319__A2 (.DIODE(_2196_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5278__A1 (.DIODE(_2196_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5259__C1 (.DIODE(_2196_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5230__A (.DIODE(_2196_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5190__A1 (.DIODE(_2196_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5173__A (.DIODE(_2196_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5140__A1 (.DIODE(_2196_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5334__A2 (.DIODE(_2381_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5350__B1 (.DIODE(_2396_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5360__B1 (.DIODE(_2404_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5370__B1 (.DIODE(_2412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5375__B1 (.DIODE(_2416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5395__S (.DIODE(_2421_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5393__S (.DIODE(_2421_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5391__S (.DIODE(_2421_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5389__S (.DIODE(_2421_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5387__S (.DIODE(_2421_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5385__S (.DIODE(_2421_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5383__S (.DIODE(_2421_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5381__S (.DIODE(_2421_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5413__S (.DIODE(_2431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5411__S (.DIODE(_2431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5409__S (.DIODE(_2431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5407__S (.DIODE(_2431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5405__S (.DIODE(_2431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5403__S (.DIODE(_2431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5401__S (.DIODE(_2431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5399__S (.DIODE(_2431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5434__S (.DIODE(_2443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5432__S (.DIODE(_2443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5430__S (.DIODE(_2443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5428__S (.DIODE(_2443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5426__S (.DIODE(_2443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5424__S (.DIODE(_2443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5422__S (.DIODE(_2443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5420__S (.DIODE(_2443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5110__B1 (.DIODE(_2456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4868__A (.DIODE(_2456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4850__A (.DIODE(_2456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4815__A (.DIODE(_2456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4569__A (.DIODE(_2456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4243__A (.DIODE(_2456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3591__A (.DIODE(_2456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3049__A (.DIODE(_2456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2810__A1_N (.DIODE(_2456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2724__A (.DIODE(_2456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5328__C1 (.DIODE(_2458_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5326__C1 (.DIODE(_2458_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5054__C1 (.DIODE(_2458_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5050__C1 (.DIODE(_2458_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5046__C1 (.DIODE(_2458_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4811__C1 (.DIODE(_2458_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4808__C1 (.DIODE(_2458_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4805__C1 (.DIODE(_2458_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2760__A2 (.DIODE(_2458_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2749__A1 (.DIODE(_2458_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5436__B1 (.DIODE(_2461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5338__A1 (.DIODE(_2461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5296__A2 (.DIODE(_2461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5105__B1 (.DIODE(_2461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5097__A (.DIODE(_2461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4589__A1 (.DIODE(_2461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2857__A1 (.DIODE(_2461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2848__B (.DIODE(_2461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2799__A1 (.DIODE(_2461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2729__A (.DIODE(_2461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5324__A2 (.DIODE(_2462_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5268__B1 (.DIODE(_2462_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5240__A2 (.DIODE(_2462_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5210__A2 (.DIODE(_2462_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5178__B1 (.DIODE(_2462_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5146__B1 (.DIODE(_2462_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5099__B2 (.DIODE(_2462_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2815__A3 (.DIODE(_2462_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2760__A3 (.DIODE(_2462_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2749__A3 (.DIODE(_2462_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5101__A2 (.DIODE(_2466_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4736__A1 (.DIODE(_2466_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4707__A1 (.DIODE(_2466_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4696__A1 (.DIODE(_2466_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4674__A1 (.DIODE(_2466_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4622__B (.DIODE(_2466_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2890__A2 (.DIODE(_2466_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2735__B (.DIODE(_2466_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5044__A0 (.DIODE(_2469_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4816__A0 (.DIODE(_2469_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4235__A0 (.DIODE(_2469_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3039__B2 (.DIODE(_2469_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2785__B (.DIODE(_2469_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2776__A (.DIODE(_2469_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2774__B (.DIODE(_2469_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2769__B (.DIODE(_2469_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2766__A (.DIODE(_2469_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2737__B (.DIODE(_2469_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4780__A1 (.DIODE(_2480_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4779__A (.DIODE(_2480_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4693__A1 (.DIODE(_2480_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4681__A (.DIODE(_2480_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4680__A (.DIODE(_2480_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4671__A1 (.DIODE(_2480_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4670__A (.DIODE(_2480_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4656__A (.DIODE(_2480_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2844__A1 (.DIODE(_2480_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2748__C (.DIODE(_2480_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5106__A (.DIODE(_2482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4891__A1 (.DIODE(_2482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4814__C_N (.DIODE(_2482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4581__B (.DIODE(_2482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2860__A1 (.DIODE(_2482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2846__A (.DIODE(_2482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2845__A (.DIODE(_2482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2835__A (.DIODE(_2482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2816__A1 (.DIODE(_2482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2760__A1 (.DIODE(_2482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5107__A1 (.DIODE(_2486_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5049__A (.DIODE(_2486_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5045__A1 (.DIODE(_2486_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4600__A (.DIODE(_2486_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4581__A (.DIODE(_2486_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4227__C1 (.DIODE(_2486_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4218__A (.DIODE(_2486_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2990__A (.DIODE(_2486_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2885__A (.DIODE(_2486_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2758__B (.DIODE(_2486_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5136__A (.DIODE(_2493_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5021__A (.DIODE(_2493_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4689__A (.DIODE(_2493_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4654__A1 (.DIODE(_2493_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4653__A (.DIODE(_2493_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3624__A1 (.DIODE(_2493_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3569__A1 (.DIODE(_2493_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3088__A (.DIODE(_2493_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2868__C (.DIODE(_2493_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2763__A (.DIODE(_2493_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5331__A (.DIODE(_2494_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5182__A (.DIODE(_2494_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5135__A (.DIODE(_2494_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5101__A1 (.DIODE(_2494_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4740__S (.DIODE(_2494_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4667__A1 (.DIODE(_2494_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4666__A (.DIODE(_2494_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4251__A1 (.DIODE(_2494_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4226__A3 (.DIODE(_2494_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2789__A (.DIODE(_2494_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5104__A1 (.DIODE(_2496_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5086__B (.DIODE(_2496_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5023__B1 (.DIODE(_2496_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4892__B1 (.DIODE(_2496_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4890__B (.DIODE(_2496_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4820__A0 (.DIODE(_2496_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4247__A (.DIODE(_2496_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3045__B2 (.DIODE(_2496_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2827__A (.DIODE(_2496_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2788__A1 (.DIODE(_2496_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5036__A (.DIODE(_2503_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5035__A1 (.DIODE(_2503_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4946__A (.DIODE(_2503_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4876__B (.DIODE(_2503_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4226__A2 (.DIODE(_2503_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2911__A1 (.DIODE(_2503_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2875__A (.DIODE(_2503_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2811__A (.DIODE(_2503_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2777__A (.DIODE(_2503_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2775__A (.DIODE(_2503_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5124__A (.DIODE(_2504_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5086__A (.DIODE(_2504_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4876__A (.DIODE(_2504_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4818__A0 (.DIODE(_2504_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4241__A (.DIODE(_2504_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3037__A1 (.DIODE(_2504_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2868__A (.DIODE(_2504_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2784__A (.DIODE(_2504_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2776__B_N (.DIODE(_2504_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2774__A (.DIODE(_2504_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5301__C1 (.DIODE(_2506_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5251__A1 (.DIODE(_2506_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5215__C1 (.DIODE(_2506_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5182__B (.DIODE(_2506_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5150__A (.DIODE(_2506_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5123__A1 (.DIODE(_2506_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2787__A2 (.DIODE(_2506_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5306__A1 (.DIODE(_2508_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5290__A1 (.DIODE(_2508_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5250__C1 (.DIODE(_2508_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5204__A1 (.DIODE(_2508_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5185__B (.DIODE(_2508_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5154__A (.DIODE(_2508_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5134__A (.DIODE(_2508_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5122__A (.DIODE(_2508_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4968__B2 (.DIODE(_2508_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2778__B1 (.DIODE(_2508_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5302__A1 (.DIODE(_2511_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5244__A1 (.DIODE(_2511_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5217__A1 (.DIODE(_2511_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5202__A1 (.DIODE(_2511_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5153__A1 (.DIODE(_2511_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5127__A1 (.DIODE(_2511_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4583__A2 (.DIODE(_2511_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3094__B (.DIODE(_2511_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2880__B (.DIODE(_2511_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2781__A (.DIODE(_2511_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4878__A1 (.DIODE(_2513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4615__A (.DIODE(_2513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3337__B1 (.DIODE(_2513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2893__B1 (.DIODE(_2513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2869__A (.DIODE(_2513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2806__B (.DIODE(_2513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2783__A (.DIODE(_2513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5101__B1 (.DIODE(_2516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4880__C (.DIODE(_2516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3088__B (.DIODE(_2516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2836__A1 (.DIODE(_2516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2807__B1 (.DIODE(_2516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2786__C1 (.DIODE(_2516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4226__A1 (.DIODE(_2527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2900__B1 (.DIODE(_2527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2806__A (.DIODE(_2527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2797__A1 (.DIODE(_2527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4736__B2 (.DIODE(_2551_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4707__B2 (.DIODE(_2551_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4696__B2 (.DIODE(_2551_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4674__B2 (.DIODE(_2551_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4607__B (.DIODE(_2551_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4581__D (.DIODE(_2551_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2860__A4 (.DIODE(_2551_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5278__C1 (.DIODE(_2553_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5175__A (.DIODE(_2553_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4733__A2 (.DIODE(_2553_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4701__B (.DIODE(_2553_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4691__A2 (.DIODE(_2553_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4632__A (.DIODE(_2553_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4224__B (.DIODE(_2553_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2879__A1 (.DIODE(_2553_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2842__A (.DIODE(_2553_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2824__A (.DIODE(_2553_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5317__C1 (.DIODE(_2554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5262__B1 (.DIODE(_2554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5237__B1 (.DIODE(_2554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5143__A (.DIODE(_2554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5092__C1 (.DIODE(_2554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4671__C1 (.DIODE(_2554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4659__A1 (.DIODE(_2554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4251__A2 (.DIODE(_2554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4239__A (.DIODE(_2554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2829__A2 (.DIODE(_2554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4583__A1 (.DIODE(_2555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4582__A (.DIODE(_2555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3887__S (.DIODE(_2555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3774__A (.DIODE(_2555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3647__A (.DIODE(_2555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3576__A1 (.DIODE(_2555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3575__A (.DIODE(_2555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3093__A (.DIODE(_2555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2876__B2 (.DIODE(_2555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2826__A (.DIODE(_2555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4730__A1 (.DIODE(_2556_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4729__A (.DIODE(_2556_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4700__S (.DIODE(_2556_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4690__A1 (.DIODE(_2556_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4633__A (.DIODE(_2556_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3993__S (.DIODE(_2556_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3773__A (.DIODE(_2556_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3712__D_N (.DIODE(_2556_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3043__B2 (.DIODE(_2556_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2828__A (.DIODE(_2556_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5333__A2 (.DIODE(_2563_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4883__B (.DIODE(_2563_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4665__B1 (.DIODE(_2563_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4628__B (.DIODE(_2563_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4620__B1 (.DIODE(_2563_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4609__B (.DIODE(_2563_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2834__D1 (.DIODE(_2563_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4669__A1 (.DIODE(_2570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4668__B1 (.DIODE(_2570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4658__A1 (.DIODE(_2570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4657__B1 (.DIODE(_2570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4632__B (.DIODE(_2570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4618__A (.DIODE(_2570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4225__A (.DIODE(_2570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3170__A (.DIODE(_2570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2999__A (.DIODE(_2570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2841__A (.DIODE(_2570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5436__A1 (.DIODE(_2581_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5336__B (.DIODE(_2581_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5100__A1 (.DIODE(_2581_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5040__A1 (.DIODE(_2581_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4884__A (.DIODE(_2581_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4622__A (.DIODE(_2581_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4251__B1 (.DIODE(_2581_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4232__A (.DIODE(_2581_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4223__A1 (.DIODE(_2581_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2852__B1 (.DIODE(_2581_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3950__A (.DIODE(_2596_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3923__C1 (.DIODE(_2596_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3650__A (.DIODE(_2596_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3514__C1 (.DIODE(_2596_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3388__C1 (.DIODE(_2596_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3249__B1 (.DIODE(_2596_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3181__B1 (.DIODE(_2596_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3124__B1 (.DIODE(_2596_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3050__A (.DIODE(_2596_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2872__A (.DIODE(_2596_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4004__A (.DIODE(_2597_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3783__A (.DIODE(_2597_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3780__C1 (.DIODE(_2597_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3717__A1 (.DIODE(_2597_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3450__B2 (.DIODE(_2597_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3446__C1 (.DIODE(_2597_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3392__A (.DIODE(_2597_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3325__A1 (.DIODE(_2597_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3188__A (.DIODE(_2597_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3033__A2 (.DIODE(_2597_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5302__B2 (.DIODE(_2600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5288__A1 (.DIODE(_2600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5244__B2 (.DIODE(_2600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5217__B2 (.DIODE(_2600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5202__B2 (.DIODE(_2600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5153__B2 (.DIODE(_2600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5126__A (.DIODE(_2600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5089__A1 (.DIODE(_2600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4582__B (.DIODE(_2600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2876__B1 (.DIODE(_2600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5102__C (.DIODE(_2602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3217__A3 (.DIODE(_2602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2890__A3 (.DIODE(_2602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2878__B (.DIODE(_2602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4000__B1 (.DIODE(_2606_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3922__B1 (.DIODE(_2606_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3873__B1 (.DIODE(_2606_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3836__B2 (.DIODE(_2606_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3579__A1 (.DIODE(_2606_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3322__A (.DIODE(_2606_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3216__A (.DIODE(_2606_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3030__A (.DIODE(_2606_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2882__B1 (.DIODE(_2606_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4011__A2 (.DIODE(_2607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3589__A2 (.DIODE(_2607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3047__A2 (.DIODE(_2607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3044__A2 (.DIODE(_2607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3042__A (.DIODE(_2607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3040__S (.DIODE(_2607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3032__A1 (.DIODE(_2607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3337__A2 (.DIODE(_2616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3336__C (.DIODE(_2616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2910__B (.DIODE(_2616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2900__A2 (.DIODE(_2616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2899__C (.DIODE(_2616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2893__A2 (.DIODE(_2616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2892__C (.DIODE(_2616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3268__A (.DIODE(_2621_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3209__B (.DIODE(_2621_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3207__B (.DIODE(_2621_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3204__B (.DIODE(_2621_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2927__B (.DIODE(_2621_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2925__B (.DIODE(_2621_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2919__B (.DIODE(_2621_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2916__B (.DIODE(_2621_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2905__B (.DIODE(_2621_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2898__B (.DIODE(_2621_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3269__A (.DIODE(_2622_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3209__C (.DIODE(_2622_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3207__C (.DIODE(_2622_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3204__C (.DIODE(_2622_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2927__C (.DIODE(_2622_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2925__C (.DIODE(_2622_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2919__C (.DIODE(_2622_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2916__C (.DIODE(_2622_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2905__C (.DIODE(_2622_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2898__C (.DIODE(_2622_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3430__A (.DIODE(_2637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3421__C1 (.DIODE(_2637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3350__B1 (.DIODE(_2637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3278__C1 (.DIODE(_2637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3273__C1 (.DIODE(_2637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3211__A1 (.DIODE(_2637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3201__A1 (.DIODE(_2637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3071__C1 (.DIODE(_2637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2929__B1 (.DIODE(_2637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2913__B1 (.DIODE(_2637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3477__A1 (.DIODE(_2640_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3426__B1 (.DIODE(_2640_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3291__A (.DIODE(_2640_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3285__A1 (.DIODE(_2640_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3201__B1 (.DIODE(_2640_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3147__B1 (.DIODE(_2640_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3079__A1 (.DIODE(_2640_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2939__A2 (.DIODE(_2640_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2938__B1 (.DIODE(_2640_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3350__A1 (.DIODE(_2642_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3343__C1 (.DIODE(_2642_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3142__A1 (.DIODE(_2642_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3138__A1 (.DIODE(_2642_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3134__A1 (.DIODE(_2642_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3071__A1 (.DIODE(_2642_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3067__A1 (.DIODE(_2642_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2937__C1 (.DIODE(_2642_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2926__C1 (.DIODE(_2642_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2918__C1 (.DIODE(_2642_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3347__C1 (.DIODE(_2645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3345__C1 (.DIODE(_2645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3329__A (.DIODE(_2645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3271__A (.DIODE(_2645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3265__C1 (.DIODE(_2645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3196__A1 (.DIODE(_2645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3063__A1 (.DIODE(_2645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2935__C1 (.DIODE(_2645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2928__C1 (.DIODE(_2645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2921__C1 (.DIODE(_2645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3426__A1 (.DIODE(_2648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3351__A1 (.DIODE(_2648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3340__B1 (.DIODE(_2648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3333__C1 (.DIODE(_2648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3279__A (.DIODE(_2648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3266__C1 (.DIODE(_2648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3206__C1 (.DIODE(_2648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3196__C1 (.DIODE(_2648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2938__A1 (.DIODE(_2648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2924__B1 (.DIODE(_2648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3468__A (.DIODE(_2658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3348__C (.DIODE(_2658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3346__C (.DIODE(_2658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3344__C (.DIODE(_2658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3342__C (.DIODE(_2658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3334__C (.DIODE(_2658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3331__C (.DIODE(_2658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3264__C (.DIODE(_2658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2936__A2 (.DIODE(_2658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2934__A2 (.DIODE(_2658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5091__A2 (.DIODE(_2665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4625__A2 (.DIODE(_2665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4621__B1 (.DIODE(_2665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4612__A2 (.DIODE(_2665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3219__A1 (.DIODE(_2665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3214__A1 (.DIODE(_2665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3081__A (.DIODE(_2665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3080__A (.DIODE(_2665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3032__A2 (.DIODE(_2665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3031__B2 (.DIODE(_2665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3402__B1 (.DIODE(_2666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3369__B1 (.DIODE(_2666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3302__B1 (.DIODE(_2666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3231__B1 (.DIODE(_2666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3104__B1 (.DIODE(_2666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2942__A (.DIODE(_2666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3983__B1 (.DIODE(_2667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3933__C1 (.DIODE(_2667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3884__C1 (.DIODE(_2667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3817__B1 (.DIODE(_2667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3760__B1 (.DIODE(_2667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3695__B1 (.DIODE(_2667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3633__B1 (.DIODE(_2667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3562__B1 (.DIODE(_2667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3495__B1 (.DIODE(_2667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2968__A1 (.DIODE(_2667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3301__S0 (.DIODE(_2668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3299__S (.DIODE(_2668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3230__S0 (.DIODE(_2668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3228__S (.DIODE(_2668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3158__S0 (.DIODE(_2668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3150__S0 (.DIODE(_2668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3106__S0 (.DIODE(_2668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3105__S0 (.DIODE(_2668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3103__S0 (.DIODE(_2668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2944__A (.DIODE(_2668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3497__S0 (.DIODE(_2669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3496__S0 (.DIODE(_2669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3404__S0 (.DIODE(_2669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3403__S0 (.DIODE(_2669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3401__S0 (.DIODE(_2669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3371__S0 (.DIODE(_2669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3370__S0 (.DIODE(_2669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3363__A (.DIODE(_2669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3153__A1 (.DIODE(_2669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2945__A (.DIODE(_2669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3697__S0 (.DIODE(_2670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3696__S0 (.DIODE(_2670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3564__S0 (.DIODE(_2670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3491__A1 (.DIODE(_2670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2962__S (.DIODE(_2670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2958__A (.DIODE(_2670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2956__A (.DIODE(_2670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2955__S0 (.DIODE(_2670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2951__S0 (.DIODE(_2670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2950__S0 (.DIODE(_2670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3301__S1 (.DIODE(_2671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3230__S1 (.DIODE(_2671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3158__S1 (.DIODE(_2671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3156__S1 (.DIODE(_2671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3153__B1_N (.DIODE(_2671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3150__S1 (.DIODE(_2671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3105__S1 (.DIODE(_2671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3103__S1 (.DIODE(_2671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3100__B1_N (.DIODE(_2671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2947__A (.DIODE(_2671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3497__S1 (.DIODE(_2672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3404__S1 (.DIODE(_2672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3403__S1 (.DIODE(_2672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3371__S1 (.DIODE(_2672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3370__S1 (.DIODE(_2672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3300__B2 (.DIODE(_2672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3229__B2 (.DIODE(_2672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3155__B2 (.DIODE(_2672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3102__B2 (.DIODE(_2672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2948__A (.DIODE(_2672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3496__S1 (.DIODE(_2673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3494__S1 (.DIODE(_2673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3491__B1_N (.DIODE(_2673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3401__S1 (.DIODE(_2673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3398__B1_N (.DIODE(_2673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3368__S1 (.DIODE(_2673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3365__B1_N (.DIODE(_2673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2960__A (.DIODE(_2673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2951__S1 (.DIODE(_2673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2949__A (.DIODE(_2673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3697__S1 (.DIODE(_2674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3696__S1 (.DIODE(_2674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3691__B1_N (.DIODE(_2674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3564__S1 (.DIODE(_2674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3563__S1 (.DIODE(_2674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3493__B2 (.DIODE(_2674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3400__B2 (.DIODE(_2674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3367__B2 (.DIODE(_2674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2955__S1 (.DIODE(_2674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2950__S1 (.DIODE(_2674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3405__S (.DIODE(_2677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3305__S (.DIODE(_2677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3302__A1 (.DIODE(_2677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3234__S (.DIODE(_2677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3231__A1 (.DIODE(_2677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3159__A1 (.DIODE(_2677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3151__A (.DIODE(_2677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3107__S (.DIODE(_2677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3104__A1 (.DIODE(_2677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2953__A (.DIODE(_2677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3695__A1 (.DIODE(_2678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3631__A (.DIODE(_2678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3565__S (.DIODE(_2678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3562__A1 (.DIODE(_2678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3495__A1 (.DIODE(_2678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3402__A1 (.DIODE(_2678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3372__S (.DIODE(_2678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3369__A1 (.DIODE(_2678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2967__A1 (.DIODE(_2678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2954__S (.DIODE(_2678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3819__S0 (.DIODE(_2681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3818__S0 (.DIODE(_2681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3762__S0 (.DIODE(_2681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3761__S0 (.DIODE(_2681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3755__A (.DIODE(_2681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3635__S0 (.DIODE(_2681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3634__S0 (.DIODE(_2681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3632__S0 (.DIODE(_2681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3556__A1 (.DIODE(_2681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2961__A1 (.DIODE(_2681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3694__S0 (.DIODE(_2683_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3692__S (.DIODE(_2683_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3691__A1 (.DIODE(_2683_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3690__A_N (.DIODE(_2683_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3625__A (.DIODE(_2683_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3563__S0 (.DIODE(_2683_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3561__S0 (.DIODE(_2683_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3557__S (.DIODE(_2683_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3555__A_N (.DIODE(_2683_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2959__A (.DIODE(_2683_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3694__S1 (.DIODE(_2685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3635__S1 (.DIODE(_2685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3634__S1 (.DIODE(_2685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3629__A (.DIODE(_2685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3627__B1_N (.DIODE(_2685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3561__S1 (.DIODE(_2685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3558__A (.DIODE(_2685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3556__B1_N (.DIODE(_2685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2965__A1 (.DIODE(_2685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2961__C1 (.DIODE(_2685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3698__S (.DIODE(_2689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3559__A (.DIODE(_2689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3498__S (.DIODE(_2689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3493__C1 (.DIODE(_2689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3400__C1 (.DIODE(_2689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3367__C1 (.DIODE(_2689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3157__A (.DIODE(_2689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3155__C1 (.DIODE(_2689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3102__C1 (.DIODE(_2689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2965__B1 (.DIODE(_2689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3987__B2 (.DIODE(_2691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3934__A1 (.DIODE(_2691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3885__A1 (.DIODE(_2691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3821__B2 (.DIODE(_2691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3764__B2 (.DIODE(_2691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3699__B2 (.DIODE(_2691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3637__B2 (.DIODE(_2691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3566__B2 (.DIODE(_2691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3164__A1 (.DIODE(_2691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2967__C1 (.DIODE(_2691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3639__A (.DIODE(_2694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3506__A1 (.DIODE(_2694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3312__A1 (.DIODE(_2694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3240__A1 (.DIODE(_2694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3163__A1 (.DIODE(_2694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3162__A1 (.DIODE(_2694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3115__A (.DIODE(_2694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2995__A (.DIODE(_2694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2971__A (.DIODE(_2694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2970__B (.DIODE(_2694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4613__B (.DIODE(_2696_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3992__S (.DIODE(_2696_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3823__A1 (.DIODE(_2696_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3703__A (.DIODE(_2696_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3638__A1 (.DIODE(_2696_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3554__A (.DIODE(_2696_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3379__A1 (.DIODE(_2696_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3313__A1 (.DIODE(_2696_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3241__A1 (.DIODE(_2696_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2972__B (.DIODE(_2696_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5109__A2 (.DIODE(_2699_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3009__B1 (.DIODE(_2699_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3004__B (.DIODE(_2699_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2975__B (.DIODE(_2699_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3998__A1_N (.DIODE(_2701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3943__C1 (.DIODE(_2701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3772__B1 (.DIODE(_2701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3710__C1 (.DIODE(_2701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3416__B1 (.DIODE(_2701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3386__B1 (.DIODE(_2701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3320__B1 (.DIODE(_2701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3176__A1 (.DIODE(_2701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3123__A1 (.DIODE(_2701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3020__A2 (.DIODE(_2701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5342__A0 (.DIODE(_2702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5094__A (.DIODE(_2702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4979__B (.DIODE(_2702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4977__B (.DIODE(_2702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4955__A_N (.DIODE(_2702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4927__A1 (.DIODE(_2702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4235__A1 (.DIODE(_2702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3574__A1 (.DIODE(_2702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3006__A1 (.DIODE(_2702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2998__A0 (.DIODE(_2702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4731__A (.DIODE(_2704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4730__C1 (.DIODE(_2704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4704__A1 (.DIODE(_2704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4692__C1 (.DIODE(_2704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4635__S (.DIODE(_2704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4610__A (.DIODE(_2704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2991__B (.DIODE(_2704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2986__B (.DIODE(_2704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2983__D (.DIODE(_2704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2980__B (.DIODE(_2704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3995__S (.DIODE(_2719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3828__A1 (.DIODE(_2719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3706__B2 (.DIODE(_2719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3509__C1 (.DIODE(_2719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3413__C1 (.DIODE(_2719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3383__C1 (.DIODE(_2719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3316__C1 (.DIODE(_2719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3245__A1 (.DIODE(_2719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3173__A1 (.DIODE(_2719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3002__A (.DIODE(_2719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5375__A1 (.DIODE(\as1802.D[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5307__A1 (.DIODE(\as1802.D[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5277__A1 (.DIODE(\as1802.D[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5022__B2 (.DIODE(\as1802.D[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4969__A (.DIODE(\as1802.D[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3977__A1 (.DIODE(\as1802.D[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3486__A (.DIODE(\as1802.D[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2767__C (.DIODE(\as1802.D[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2786__B2 (.DIODE(\as1802.EF_l[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2778__B2 (.DIODE(\as1802.EF_l[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2778__A2 (.DIODE(\as1802.EF_l[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2787__A1 (.DIODE(\as1802.EF_l[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4859__B1_N (.DIODE(\as1802.IE ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4854__A2 (.DIODE(\as1802.IE ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4222__A (.DIODE(\as1802.IE ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2807__A1 (.DIODE(\as1802.IE ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2756__A (.DIODE(\as1802.IE ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5354__A1 (.DIODE(\as1802.P[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5070__A1 (.DIODE(\as1802.P[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5055__A0 (.DIODE(\as1802.P[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4253__A0 (.DIODE(\as1802.P[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3043__A1 (.DIODE(\as1802.P[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5359__A1 (.DIODE(\as1802.X[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5073__A1 (.DIODE(\as1802.X[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5046__A1 (.DIODE(\as1802.X[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3336__A (.DIODE(\as1802.X[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3040__A0 (.DIODE(\as1802.X[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2892__A (.DIODE(\as1802.X[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5364__A1 (.DIODE(\as1802.X[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5076__A1 (.DIODE(\as1802.X[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5050__A1 (.DIODE(\as1802.X[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3037__B2 (.DIODE(\as1802.X[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2899__A (.DIODE(\as1802.X[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5369__A1 (.DIODE(\as1802.X[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5054__A1 (.DIODE(\as1802.X[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3589__A1 (.DIODE(\as1802.X[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3047__A1 (.DIODE(\as1802.X[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2922__A0 (.DIODE(\as1802.X[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2909__A (.DIODE(\as1802.X[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5374__A1 (.DIODE(\as1802.X[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5057__A0 (.DIODE(\as1802.X[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4011__A1 (.DIODE(\as1802.X[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3076__A (.DIODE(\as1802.X[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3044__A1 (.DIODE(\as1802.X[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2914__A0 (.DIODE(\as1802.X[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4809__A0 (.DIODE(\as1802.addr_buff[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4785__B1 (.DIODE(\as1802.addr_buff[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4557__A2 (.DIODE(\as1802.addr_buff[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4545__A (.DIODE(\as1802.addr_buff[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2914__A1 (.DIODE(\as1802.cond_inv ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2877__D (.DIODE(\as1802.cond_inv ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2802__A (.DIODE(\as1802.cond_inv ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2761__A (.DIODE(\as1802.cond_inv ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2738__A1 (.DIODE(\as1802.cond_inv ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3641__A (.DIODE(\as1802.instr_cycle[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3120__A (.DIODE(\as1802.instr_cycle[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3017__A (.DIODE(\as1802.instr_cycle[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2984__A (.DIODE(\as1802.instr_cycle[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2982__A (.DIODE(\as1802.instr_cycle[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2847__A (.DIODE(\as1802.instr_cycle[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2845__B (.DIODE(\as1802.instr_cycle[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2815__A2 (.DIODE(\as1802.instr_cycle[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2749__B2 (.DIODE(\as1802.instr_cycle[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2922__A1 (.DIODE(\as1802.instr_latch[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2877__C (.DIODE(\as1802.instr_latch[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2803__A (.DIODE(\as1802.instr_latch[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2785__C (.DIODE(\as1802.instr_latch[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2772__A (.DIODE(\as1802.instr_latch[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2764__A (.DIODE(\as1802.instr_latch[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2738__B1 (.DIODE(\as1802.instr_latch[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5110__A1 (.DIODE(\as1802.mem_cycle[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4872__A2 (.DIODE(\as1802.mem_cycle[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4865__C (.DIODE(\as1802.mem_cycle[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4787__B (.DIODE(\as1802.mem_cycle[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4592__A (.DIODE(\as1802.mem_cycle[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4591__A (.DIODE(\as1802.mem_cycle[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4562__A (.DIODE(\as1802.mem_cycle[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2817__C (.DIODE(\as1802.mem_cycle[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2751__C (.DIODE(\as1802.mem_cycle[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2726__C (.DIODE(\as1802.mem_cycle[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5110__C1 (.DIODE(\as1802.mem_cycle[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4872__A1 (.DIODE(\as1802.mem_cycle[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4866__B (.DIODE(\as1802.mem_cycle[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4865__B (.DIODE(\as1802.mem_cycle[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4812__A (.DIODE(\as1802.mem_cycle[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4595__B2 (.DIODE(\as1802.mem_cycle[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4560__B1 (.DIODE(\as1802.mem_cycle[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2817__B (.DIODE(\as1802.mem_cycle[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2751__B (.DIODE(\as1802.mem_cycle[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2726__B (.DIODE(\as1802.mem_cycle[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4832__A (.DIODE(\as1802.mem_cycle[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4786__A (.DIODE(\as1802.mem_cycle[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4596__B2 (.DIODE(\as1802.mem_cycle[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4563__A (.DIODE(\as1802.mem_cycle[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2817__A (.DIODE(\as1802.mem_cycle[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2751__A (.DIODE(\as1802.mem_cycle[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2726__A (.DIODE(\as1802.mem_cycle[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5416__A1 (.DIODE(\as1802.mem_write ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5110__A2 (.DIODE(\as1802.mem_write ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5106__B (.DIODE(\as1802.mem_write ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4814__A (.DIODE(\as1802.mem_write ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4544__A (.DIODE(\as1802.mem_write ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5403__A0 (.DIODE(\as1802.regs[2][10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4733__A1 (.DIODE(\as1802.regs[2][10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3782__A1 (.DIODE(\as1802.regs[2][10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3781__A (.DIODE(\as1802.regs[2][10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3697__A2 (.DIODE(\as1802.regs[2][10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3663__A (.DIODE(\as1802.regs[2][10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3659__A (.DIODE(\as1802.regs[2][10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5405__A0 (.DIODE(\as1802.regs[2][11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4742__A1 (.DIODE(\as1802.regs[2][11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3782__B1 (.DIODE(\as1802.regs[2][11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3781__B (.DIODE(\as1802.regs[2][11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3762__A2 (.DIODE(\as1802.regs[2][11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3729__A (.DIODE(\as1802.regs[2][11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5407__A0 (.DIODE(\as1802.regs[2][12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4751__A1 (.DIODE(\as1802.regs[2][12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3838__A1 (.DIODE(\as1802.regs[2][12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3837__A (.DIODE(\as1802.regs[2][12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3818__A2 (.DIODE(\as1802.regs[2][12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3790__A (.DIODE(\as1802.regs[2][12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5409__A0 (.DIODE(\as1802.regs[2][13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4760__A1 (.DIODE(\as1802.regs[2][13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3874__A2 (.DIODE(\as1802.regs[2][13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3852__A0 (.DIODE(\as1802.regs[2][13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3844__A1 (.DIODE(\as1802.regs[2][13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3843__A (.DIODE(\as1802.regs[2][13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5411__A0 (.DIODE(\as1802.regs[2][14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4769__A1 (.DIODE(\as1802.regs[2][14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3949__A (.DIODE(\as1802.regs[2][14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3948__A (.DIODE(\as1802.regs[2][14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3925__A2 (.DIODE(\as1802.regs[2][14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3907__A (.DIODE(\as1802.regs[2][14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5413__A0 (.DIODE(\as1802.regs[2][15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4777__A1 (.DIODE(\as1802.regs[2][15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4003__A (.DIODE(\as1802.regs[2][15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4002__A (.DIODE(\as1802.regs[2][15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3985__A2 (.DIODE(\as1802.regs[2][15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3959__A0 (.DIODE(\as1802.regs[2][15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4637__A1 (.DIODE(\as1802.regs[2][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4314__A0 (.DIODE(\as1802.regs[2][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3187__B (.DIODE(\as1802.regs[2][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3186__A2 (.DIODE(\as1802.regs[2][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3105__A2 (.DIODE(\as1802.regs[2][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3065__A (.DIODE(\as1802.regs[2][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3058__B (.DIODE(\as1802.regs[2][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3057__B (.DIODE(\as1802.regs[2][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4645__A1 (.DIODE(\as1802.regs[2][2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4316__A0 (.DIODE(\as1802.regs[2][2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3187__C (.DIODE(\as1802.regs[2][2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3186__B1 (.DIODE(\as1802.regs[2][2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3156__A2 (.DIODE(\as1802.regs[2][2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3140__A (.DIODE(\as1802.regs[2][2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4657__A1 (.DIODE(\as1802.regs[2][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4318__A0 (.DIODE(\as1802.regs[2][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3252__A (.DIODE(\as1802.regs[2][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3251__A (.DIODE(\as1802.regs[2][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3232__A2 (.DIODE(\as1802.regs[2][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3199__A (.DIODE(\as1802.regs[2][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4668__A1 (.DIODE(\as1802.regs[2][4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4320__A0 (.DIODE(\as1802.regs[2][4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3303__A2 (.DIODE(\as1802.regs[2][4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3270__A (.DIODE(\as1802.regs[2][4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3259__A (.DIODE(\as1802.regs[2][4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3258__A (.DIODE(\as1802.regs[2][4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4682__A1 (.DIODE(\as1802.regs[2][5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4322__A0 (.DIODE(\as1802.regs[2][5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3391__A (.DIODE(\as1802.regs[2][5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3390__A (.DIODE(\as1802.regs[2][5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3370__A2 (.DIODE(\as1802.regs[2][5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3339__C_N (.DIODE(\as1802.regs[2][5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4691__A1 (.DIODE(\as1802.regs[2][6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4324__A0 (.DIODE(\as1802.regs[2][6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3448__A (.DIODE(\as1802.regs[2][6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3447__A (.DIODE(\as1802.regs[2][6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3419__A (.DIODE(\as1802.regs[2][6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3403__A2 (.DIODE(\as1802.regs[2][6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4701__A (.DIODE(\as1802.regs[2][7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4326__A0 (.DIODE(\as1802.regs[2][7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3497__A2 (.DIODE(\as1802.regs[2][7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3462__A (.DIODE(\as1802.regs[2][7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3455__A1 (.DIODE(\as1802.regs[2][7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3454__A (.DIODE(\as1802.regs[2][7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5399__A0 (.DIODE(\as1802.regs[2][8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4713__A1 (.DIODE(\as1802.regs[2][8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3563__A2 (.DIODE(\as1802.regs[2][8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3540__A (.DIODE(\as1802.regs[2][8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3521__A (.DIODE(\as1802.regs[2][8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3520__A1 (.DIODE(\as1802.regs[2][8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5401__A0 (.DIODE(\as1802.regs[2][9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4722__A1 (.DIODE(\as1802.regs[2][9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3634__A2 (.DIODE(\as1802.regs[2][9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3600__A (.DIODE(\as1802.regs[2][9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3598__A (.DIODE(\as1802.regs[2][9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3597__A1 (.DIODE(\as1802.regs[2][9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_clk_A (.DIODE(clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_A (.DIODE(io_in[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_A (.DIODE(io_in[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input3_A (.DIODE(io_in[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input4_A (.DIODE(io_in[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input5_A (.DIODE(io_in[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input6_A (.DIODE(io_in[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input7_A (.DIODE(io_in[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input8_A (.DIODE(io_in[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input9_A (.DIODE(io_in[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input10_A (.DIODE(io_in[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input11_A (.DIODE(io_in[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input12_A (.DIODE(io_in[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input13_A (.DIODE(io_in[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5802__A (.DIODE(io_oeb));
 sky130_fd_sc_hd__diode_2 ANTENNA__4867__B2 (.DIODE(io_oeb));
 sky130_fd_sc_hd__diode_2 ANTENNA__2801__A1 (.DIODE(io_out[21]));
 sky130_fd_sc_hd__diode_2 ANTENNA__2770__A (.DIODE(io_out[21]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5438__A1 (.DIODE(io_out[25]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5440__A1 (.DIODE(io_out[26]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5352__A0 (.DIODE(io_out[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5160__A2 (.DIODE(io_out[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA__4974__B (.DIODE(io_out[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA__4246__A (.DIODE(io_out[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3708__A1 (.DIODE(io_out[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3168__A (.DIODE(io_out[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5357__A0 (.DIODE(io_out[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5205__A2 (.DIODE(io_out[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA__4973__B (.DIODE(io_out[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA__4917__A_N (.DIODE(io_out[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA__4915__B (.DIODE(io_out[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA__4252__A1 (.DIODE(io_out[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3772__A1 (.DIODE(io_out[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3246__A1 (.DIODE(io_out[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3243__A1 (.DIODE(io_out[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5362__A0 (.DIODE(io_out[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5247__A (.DIODE(io_out[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5221__A2 (.DIODE(io_out[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5043__A1 (.DIODE(io_out[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA__4972__B (.DIODE(io_out[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA__4911__A_N (.DIODE(io_out[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA__4909__B_N (.DIODE(io_out[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3833__A1 (.DIODE(io_out[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3320__A1 (.DIODE(io_out[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3314__A (.DIODE(io_out[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5367__A0 (.DIODE(io_out[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5253__A2 (.DIODE(io_out[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5047__A1 (.DIODE(io_out[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA__4971__B (.DIODE(io_out[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA__4906__A_N (.DIODE(io_out[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA__4901__B (.DIODE(io_out[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3891__A1 (.DIODE(io_out[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3386__A1 (.DIODE(io_out[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3381__A (.DIODE(io_out[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5372__A0 (.DIODE(io_out[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5292__A2 (.DIODE(io_out[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5051__A1 (.DIODE(io_out[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA__4970__B (.DIODE(io_out[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA__4902__A (.DIODE(io_out[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA__4894__B_N (.DIODE(io_out[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3940__A1 (.DIODE(io_out[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3416__A1 (.DIODE(io_out[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3411__A (.DIODE(io_out[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5377__A0 (.DIODE(io_out[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5307__A2 (.DIODE(io_out[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5055__A1 (.DIODE(io_out[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA__4969__B (.DIODE(io_out[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA__4897__B (.DIODE(io_out[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA__4895__B (.DIODE(io_out[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA__4893__B (.DIODE(io_out[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3994__A1 (.DIODE(io_out[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3512__A1 (.DIODE(io_out[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3507__A (.DIODE(io_out[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input14_A (.DIODE(rst));
 sky130_fd_sc_hd__diode_2 ANTENNA__5356__A0 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__5210__A1 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__4822__A1 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__5361__A0 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__5240__A1 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__4824__A1 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__5366__A0 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__5268__B2 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__4826__A1 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__5371__A0 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__5296__A1 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__4828__A1 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__5376__A0 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__5324__A1 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__4830__A1 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__4854__A3 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__2756__B (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__3581__A (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__3025__A (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__2751__D (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__2734__A (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__2723__A (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_3__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_2__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_1__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_0__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_50_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_49_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_48_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_47_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_46_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_45_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_44_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__5549__CLK (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_2_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_0_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_18_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_15_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_14_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_13_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_12_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_11_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_10_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_9_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_8_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_7_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_6_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_5_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_4_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_opt_1_0_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_1_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_42_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_41_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_40_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_39_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_38_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_37_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_36_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_35_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_34_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_opt_2_0_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_32_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_31_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_30_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__5666__CLK (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_28_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_27_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_26_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_25_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_24_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_23_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_22_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_21_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_20_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_19_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_17_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_16_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__decap_3 FILLER_0_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_295 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_388 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_407 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_438 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_442 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_463 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_669 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_294 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_311 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_412 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_100 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_227 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_375 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_543 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_677 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_208 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_301 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_379 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_551 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_258 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_271 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_340 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_555 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_677 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_84 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_310 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_551 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_571 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_583 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_58 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_275 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_381 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_426 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_439 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_555 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_677 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_187 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_208 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_379 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_551 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_40 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_71 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_380 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_439 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_450 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_466 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_555 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_75 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_91 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_291 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_354 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_380 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_410 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_491 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_551 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_115 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_220 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_344 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_450 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_472 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_677 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_68 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_244 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_364 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_380 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_551 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_51 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_71 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_271 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_439 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_10 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_188 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_341 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_551 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_571 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_56 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_90 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_229 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_520 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_21 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_75 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_135 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_151 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_183 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_207 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_351 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_551 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_583 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_14 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_48 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_95 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_117 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_392 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_434 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_456 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_599 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_611 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_28 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_44 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_196 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_244 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_420 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_424 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_551 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_607 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_13 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_34 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_47 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_56 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_73 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_96 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_116 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_462 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_605 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_611 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_20 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_88 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_184 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_235 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_254 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_409 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_548 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_607 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_669 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_201 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_216 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_230 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_326 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_354 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_575 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_677 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_31 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_74 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_135 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_155 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_246 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_341 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_358 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_397 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_420 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_492 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_607 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_669 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_48 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_62 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_136 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_170 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_211 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_262 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_330 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_386 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_528 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_677 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_10 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_22 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_42 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_127 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_300 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_364 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_592 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_604 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_639 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_68 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_95 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_112 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_154 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_381 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_404 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_463 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_488 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_556 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_562 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_635 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_661 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_147 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_162 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_236 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_416 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_556 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_567 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_603 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_44 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_59 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_67 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_382 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_568 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_635 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_52 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_84 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_350 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_516 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_592 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_604 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_639 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_669 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_13 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_35 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_102 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_208 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_270 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_315 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_339 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_386 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_495 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_556 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_562 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_618 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_661 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_43 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_128 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_145 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_203 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_235 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_267 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_324 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_456 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_534 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_639 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_20 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_116 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_183 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_190 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_228 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_273 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_282 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_400 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_7 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_42 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_130 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_202 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_256 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_551 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_592 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_639 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_13 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_48 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_106 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_162 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_238 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_330 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_439 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_491 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_631 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_661 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_175 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_192 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_240 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_355 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_403 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_420 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_488 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_524 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_579 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_639 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_39 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_99 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_118 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_264 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_341 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_408 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_425 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_491 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_512 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_551 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_635 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_677 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_14 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_20 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_87 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_140 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_162 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_258 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_351 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_509 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_537 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_607 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_639 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_669 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_14 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_20 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_24 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_115 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_183 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_239 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_499 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_618 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_630 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_677 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_20 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_32 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_62 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_162 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_187 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_208 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_292 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_314 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_388 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_639 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_96 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_272 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_282 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_322 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_492 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_516 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_543 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_564 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_635 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_31 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_144 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_183 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_191 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_229 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_256 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_492 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_535 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_639 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_36 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_112 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_173 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_183 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_340 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_381 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_562 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_574 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_635 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_202 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_240 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_246 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_352 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_422 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_426 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_471 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_551 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_607 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_639 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_669 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_13 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_46 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_152 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_259 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_338 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_352 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_439 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_631 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_661 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_13 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_25 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_74 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_90 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_292 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_398 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_520 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_535 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_639 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_48 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_182 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_408 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_450 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_562 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_631 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_677 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_75 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_266 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_274 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_308 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_410 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_438 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_604 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_639 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_108 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_156 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_192 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_346 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_411 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_436 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_481 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_677 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_78 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_118 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_242 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_326 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_478 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_546 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_565 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_627 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_639 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_273 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_284 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_325 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_372 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_551 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_618 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_630 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_677 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_132 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_186 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_203 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_236 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_257 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_354 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_467 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_603 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_639 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_116 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_211 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_270 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_382 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_522 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_544 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_631 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_677 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_134 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_230 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_298 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_424 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_470 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_476 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_491 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_581 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_603 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_639 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_112 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_160 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_179 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_332 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_341 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_379 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_385 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_411 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_448 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_618 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_630 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_677 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_117 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_191 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_230 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_252 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_434 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_551 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_592 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_627 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_669 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_264 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_284 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_452 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_481 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_563 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_571 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_618 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_630 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_314 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_328 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_397 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_403 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_603 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_627 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_669 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_262 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_283 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_392 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_500 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_520 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_550 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_618 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_677 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_235 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_298 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_548 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_627 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_639 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_435 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_244 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_492 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_532 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_627 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_639 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_10 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_56 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_170 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_224 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_276 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_375 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_550 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_562 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_618 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_630 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_126 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_207 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_229 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_326 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_355 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_398 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_453 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_491 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_551 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_603 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_627 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_639 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_22 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_56 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_231 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_272 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_329 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_352 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_376 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_431 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_462 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_481 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_493 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_562 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_618 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_243 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_388 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_554 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_627 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_639 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_107 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_116 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_203 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_228 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_264 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_371 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_550 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_562 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_618 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_252 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_494 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_523 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_592 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_604 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_627 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_639 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_60 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_152 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_204 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_226 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_259 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_452 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_488 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_620 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_626 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_677 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_295 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_326 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_516 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_556 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_588 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_604 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_639 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_58 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_151 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_258 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_571 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_618 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_630 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_123 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_144 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_356 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_366 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_532 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_627 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_639 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_80 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_162 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_174 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_271 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_483 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_562 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_88 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_147 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_238 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_258 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_323 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_350 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_366 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_532 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_556 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_607 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_669 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_56 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_220 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_314 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_340 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_562 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_575 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_618 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_677 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_411 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_528 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_40 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_108 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_123 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_216 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_269 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_338 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_371 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_397 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_576 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_606 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_10 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_88 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_236 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_267 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_372 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_516 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_112 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_201 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_379 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_416 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_493 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_499 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_605 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_677 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_182 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_522 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_583 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_52 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_96 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_220 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_496 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_506 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_92 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_175 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_241 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_350 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_359 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_525 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_572 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_61 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_292 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_379 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_410 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_434 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_452 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_311 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_425 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_521 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_535 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_152 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_207 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_328 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_410 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_462 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_543 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_555 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_677 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_75 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_263 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_372 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_435 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_521 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_61 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_123 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_152 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_235 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_320 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_372 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_392 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_450 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_10 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_232 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_292 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_352 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_411 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_247 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_255 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_291 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_323 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_435 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_91 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_116 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_294 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_378 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_411 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_68 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_290 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_348 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_56 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_217 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_230 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_258 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_276 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_326 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_371 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_84 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_229 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_58 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_115 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_215 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_288 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_677 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_247 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_355 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_422 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_116 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_203 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_232 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_383 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_396 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_124 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_355 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_172 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_215 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_292 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_124 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_186 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_314 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_367 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_170 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_190 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_271 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_155 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_230 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_326 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_356 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_152 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_172 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_182 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_297 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_327 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_152 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_176 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_245 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_263 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_299 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_354 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_159 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_210 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_282 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_290 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_322 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_201 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_245 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_294 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_185 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_274 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_669 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_673 ();
 assign io_out[10] = net17;
 assign io_out[11] = net18;
 assign io_out[12] = net19;
 assign io_out[8] = net15;
 assign io_out[9] = net16;
endmodule

