VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO wrapped_as2650
  CLASS BLOCK ;
  FOREIGN wrapped_as2650 ;
  ORIGIN 0.000 0.000 ;
  SIZE 350.000 BY 350.000 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 297.250 0.000 297.530 4.000 ;
    END
  END clk
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.570 0.000 17.850 4.000 ;
    END
  END io_in[0]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.530 0.000 52.810 4.000 ;
    END
  END io_in[1]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.490 0.000 87.770 4.000 ;
    END
  END io_in[2]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.450 0.000 122.730 4.000 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.410 0.000 157.690 4.000 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 192.370 0.000 192.650 4.000 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 227.330 0.000 227.610 4.000 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 262.290 0.000 262.570 4.000 ;
    END
  END io_in[7]
  PIN io_oeb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 339.360 4.000 339.960 ;
    END
  END io_oeb
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 8.880 4.000 9.480 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 131.280 4.000 131.880 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 143.520 4.000 144.120 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 155.760 4.000 156.360 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 168.000 4.000 168.600 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 180.240 4.000 180.840 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 192.480 4.000 193.080 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 204.720 4.000 205.320 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 216.960 4.000 217.560 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 229.200 4.000 229.800 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 241.440 4.000 242.040 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 21.120 4.000 21.720 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 253.680 4.000 254.280 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 265.920 4.000 266.520 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 278.160 4.000 278.760 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 290.400 4.000 291.000 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 302.640 4.000 303.240 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 314.880 4.000 315.480 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 327.120 4.000 327.720 ;
    END
  END io_out[26]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 33.360 4.000 33.960 ;
    END
  END io_out[2]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 45.600 4.000 46.200 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.840 4.000 58.440 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 70.080 4.000 70.680 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 82.320 4.000 82.920 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 94.560 4.000 95.160 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 106.800 4.000 107.400 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 119.040 4.000 119.640 ;
    END
  END io_out[9]
  PIN rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 332.210 0.000 332.490 4.000 ;
    END
  END rst
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 337.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 337.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 337.520 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 337.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 337.520 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 344.080 337.365 ;
      LAYER met1 ;
        RECT 0.990 3.780 344.080 337.920 ;
      LAYER met2 ;
        RECT 1.010 4.280 340.760 339.845 ;
        RECT 1.010 3.750 17.290 4.280 ;
        RECT 18.130 3.750 52.250 4.280 ;
        RECT 53.090 3.750 87.210 4.280 ;
        RECT 88.050 3.750 122.170 4.280 ;
        RECT 123.010 3.750 157.130 4.280 ;
        RECT 157.970 3.750 192.090 4.280 ;
        RECT 192.930 3.750 227.050 4.280 ;
        RECT 227.890 3.750 262.010 4.280 ;
        RECT 262.850 3.750 296.970 4.280 ;
        RECT 297.810 3.750 331.930 4.280 ;
        RECT 332.770 3.750 340.760 4.280 ;
      LAYER met3 ;
        RECT 4.400 338.960 338.035 339.825 ;
        RECT 0.985 328.120 338.035 338.960 ;
        RECT 4.400 326.720 338.035 328.120 ;
        RECT 0.985 315.880 338.035 326.720 ;
        RECT 4.400 314.480 338.035 315.880 ;
        RECT 0.985 303.640 338.035 314.480 ;
        RECT 4.400 302.240 338.035 303.640 ;
        RECT 0.985 291.400 338.035 302.240 ;
        RECT 4.400 290.000 338.035 291.400 ;
        RECT 0.985 279.160 338.035 290.000 ;
        RECT 4.400 277.760 338.035 279.160 ;
        RECT 0.985 266.920 338.035 277.760 ;
        RECT 4.400 265.520 338.035 266.920 ;
        RECT 0.985 254.680 338.035 265.520 ;
        RECT 4.400 253.280 338.035 254.680 ;
        RECT 0.985 242.440 338.035 253.280 ;
        RECT 4.400 241.040 338.035 242.440 ;
        RECT 0.985 230.200 338.035 241.040 ;
        RECT 4.400 228.800 338.035 230.200 ;
        RECT 0.985 217.960 338.035 228.800 ;
        RECT 4.400 216.560 338.035 217.960 ;
        RECT 0.985 205.720 338.035 216.560 ;
        RECT 4.400 204.320 338.035 205.720 ;
        RECT 0.985 193.480 338.035 204.320 ;
        RECT 4.400 192.080 338.035 193.480 ;
        RECT 0.985 181.240 338.035 192.080 ;
        RECT 4.400 179.840 338.035 181.240 ;
        RECT 0.985 169.000 338.035 179.840 ;
        RECT 4.400 167.600 338.035 169.000 ;
        RECT 0.985 156.760 338.035 167.600 ;
        RECT 4.400 155.360 338.035 156.760 ;
        RECT 0.985 144.520 338.035 155.360 ;
        RECT 4.400 143.120 338.035 144.520 ;
        RECT 0.985 132.280 338.035 143.120 ;
        RECT 4.400 130.880 338.035 132.280 ;
        RECT 0.985 120.040 338.035 130.880 ;
        RECT 4.400 118.640 338.035 120.040 ;
        RECT 0.985 107.800 338.035 118.640 ;
        RECT 4.400 106.400 338.035 107.800 ;
        RECT 0.985 95.560 338.035 106.400 ;
        RECT 4.400 94.160 338.035 95.560 ;
        RECT 0.985 83.320 338.035 94.160 ;
        RECT 4.400 81.920 338.035 83.320 ;
        RECT 0.985 71.080 338.035 81.920 ;
        RECT 4.400 69.680 338.035 71.080 ;
        RECT 0.985 58.840 338.035 69.680 ;
        RECT 4.400 57.440 338.035 58.840 ;
        RECT 0.985 46.600 338.035 57.440 ;
        RECT 4.400 45.200 338.035 46.600 ;
        RECT 0.985 34.360 338.035 45.200 ;
        RECT 4.400 32.960 338.035 34.360 ;
        RECT 0.985 22.120 338.035 32.960 ;
        RECT 4.400 20.720 338.035 22.120 ;
        RECT 0.985 9.880 338.035 20.720 ;
        RECT 4.400 8.480 338.035 9.880 ;
        RECT 0.985 4.935 338.035 8.480 ;
      LAYER met4 ;
        RECT 3.055 10.240 20.640 331.665 ;
        RECT 23.040 10.240 97.440 331.665 ;
        RECT 99.840 10.240 174.240 331.665 ;
        RECT 176.640 10.240 251.040 331.665 ;
        RECT 253.440 10.240 297.785 331.665 ;
        RECT 3.055 4.935 297.785 10.240 ;
  END
END wrapped_as2650
END LIBRARY

