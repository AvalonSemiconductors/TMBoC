magic
tech sky130B
magscale 1 2
timestamp 1680173952
<< viali >>
rect 4905 33541 4939 33575
rect 7849 33541 7883 33575
rect 10793 33541 10827 33575
rect 14473 33541 14507 33575
rect 17049 33541 17083 33575
rect 19717 33541 19751 33575
rect 22661 33541 22695 33575
rect 25605 33541 25639 33575
rect 28549 33541 28583 33575
rect 31493 33541 31527 33575
rect 34253 33541 34287 33575
rect 8033 33337 8067 33371
rect 10977 33337 11011 33371
rect 14289 33337 14323 33371
rect 16865 33337 16899 33371
rect 19533 33337 19567 33371
rect 22477 33337 22511 33371
rect 25421 33337 25455 33371
rect 28365 33337 28399 33371
rect 31309 33337 31343 33371
rect 34069 33337 34103 33371
rect 4997 33269 5031 33303
rect 20637 32929 20671 32963
rect 10241 32861 10275 32895
rect 16313 32861 16347 32895
rect 16497 32861 16531 32895
rect 16589 32861 16623 32895
rect 20545 32861 20579 32895
rect 22477 32861 22511 32895
rect 15853 32793 15887 32827
rect 10149 32725 10183 32759
rect 20913 32725 20947 32759
rect 22385 32725 22419 32759
rect 12265 32521 12299 32555
rect 13461 32521 13495 32555
rect 17325 32521 17359 32555
rect 18061 32521 18095 32555
rect 13277 32453 13311 32487
rect 21189 32453 21223 32487
rect 22109 32453 22143 32487
rect 9873 32385 9907 32419
rect 10425 32385 10459 32419
rect 10517 32385 10551 32419
rect 12081 32385 12115 32419
rect 17233 32385 17267 32419
rect 18061 32385 18095 32419
rect 18245 32385 18279 32419
rect 21097 32385 21131 32419
rect 22017 32385 22051 32419
rect 22201 32385 22235 32419
rect 23121 32385 23155 32419
rect 23305 32385 23339 32419
rect 24501 32385 24535 32419
rect 24685 32385 24719 32419
rect 27721 32385 27755 32419
rect 28641 32385 28675 32419
rect 30481 32385 30515 32419
rect 33425 32385 33459 32419
rect 10701 32317 10735 32351
rect 12357 32317 12391 32351
rect 13553 32317 13587 32351
rect 17417 32317 17451 32351
rect 21281 32317 21315 32351
rect 16865 32249 16899 32283
rect 20729 32249 20763 32283
rect 23029 32249 23063 32283
rect 27169 32249 27203 32283
rect 9873 32181 9907 32215
rect 10609 32181 10643 32215
rect 11805 32181 11839 32215
rect 13001 32181 13035 32215
rect 24593 32181 24627 32215
rect 30297 32181 30331 32215
rect 33241 32181 33275 32215
rect 15761 31977 15795 32011
rect 18061 31977 18095 32011
rect 21281 31977 21315 32011
rect 23765 31977 23799 32011
rect 9321 31909 9355 31943
rect 11161 31909 11195 31943
rect 15945 31909 15979 31943
rect 18337 31909 18371 31943
rect 24593 31909 24627 31943
rect 8493 31841 8527 31875
rect 9781 31841 9815 31875
rect 9873 31841 9907 31875
rect 11621 31841 11655 31875
rect 12725 31841 12759 31875
rect 13553 31841 13587 31875
rect 14381 31841 14415 31875
rect 17141 31841 17175 31875
rect 19441 31841 19475 31875
rect 22109 31841 22143 31875
rect 22661 31841 22695 31875
rect 23121 31841 23155 31875
rect 25053 31841 25087 31875
rect 25145 31841 25179 31875
rect 8401 31773 8435 31807
rect 8585 31773 8619 31807
rect 9689 31773 9723 31807
rect 11713 31773 11747 31807
rect 13461 31773 13495 31807
rect 14289 31773 14323 31807
rect 14473 31773 14507 31807
rect 16405 31773 16439 31807
rect 16865 31773 16899 31807
rect 17325 31773 17359 31807
rect 18337 31773 18371 31807
rect 18521 31773 18555 31807
rect 20269 31773 20303 31807
rect 20453 31773 20487 31807
rect 21005 31773 21039 31807
rect 22937 31773 22971 31807
rect 23765 31773 23799 31807
rect 23949 31773 23983 31807
rect 26617 31773 26651 31807
rect 27353 31773 27387 31807
rect 15577 31705 15611 31739
rect 17233 31705 17267 31739
rect 21281 31705 21315 31739
rect 11621 31637 11655 31671
rect 15777 31637 15811 31671
rect 21097 31637 21131 31671
rect 23581 31637 23615 31671
rect 24961 31637 24995 31671
rect 9505 31433 9539 31467
rect 13553 31433 13587 31467
rect 16129 31433 16163 31467
rect 17049 31433 17083 31467
rect 17601 31433 17635 31467
rect 20846 31433 20880 31467
rect 24777 31433 24811 31467
rect 25881 31433 25915 31467
rect 28825 31433 28859 31467
rect 10701 31365 10735 31399
rect 16865 31365 16899 31399
rect 22201 31365 22235 31399
rect 9137 31297 9171 31331
rect 10241 31297 10275 31331
rect 10333 31297 10367 31331
rect 13185 31297 13219 31331
rect 14105 31297 14139 31331
rect 14841 31297 14875 31331
rect 14933 31297 14967 31331
rect 16129 31297 16163 31331
rect 16313 31297 16347 31331
rect 17141 31297 17175 31331
rect 17601 31297 17635 31331
rect 17785 31297 17819 31331
rect 20637 31297 20671 31331
rect 21097 31297 21131 31331
rect 22661 31297 22695 31331
rect 22753 31297 22787 31331
rect 23029 31297 23063 31331
rect 23305 31297 23339 31331
rect 23581 31297 23615 31331
rect 24225 31297 24259 31331
rect 24593 31297 24627 31331
rect 25237 31297 25271 31331
rect 25421 31297 25455 31331
rect 25697 31297 25731 31331
rect 27353 31297 27387 31331
rect 27629 31297 27663 31331
rect 28365 31297 28399 31331
rect 28641 31297 28675 31331
rect 9229 31229 9263 31263
rect 10425 31229 10459 31263
rect 13277 31229 13311 31263
rect 20545 31229 20579 31263
rect 25605 31229 25639 31263
rect 27169 31229 27203 31263
rect 10977 31161 11011 31195
rect 25513 31161 25547 31195
rect 28457 31161 28491 31195
rect 14289 31093 14323 31127
rect 16865 31093 16899 31127
rect 24593 31093 24627 31127
rect 9413 30889 9447 30923
rect 10057 30889 10091 30923
rect 10701 30889 10735 30923
rect 13553 30889 13587 30923
rect 17049 30889 17083 30923
rect 21005 30889 21039 30923
rect 22845 30889 22879 30923
rect 24961 30821 24995 30855
rect 13461 30753 13495 30787
rect 15761 30753 15795 30787
rect 20637 30753 20671 30787
rect 23213 30753 23247 30787
rect 27445 30753 27479 30787
rect 9321 30685 9355 30719
rect 9505 30685 9539 30719
rect 9965 30685 9999 30719
rect 10149 30685 10183 30719
rect 10609 30685 10643 30719
rect 10793 30685 10827 30719
rect 13645 30685 13679 30719
rect 13737 30685 13771 30719
rect 14565 30685 14599 30719
rect 14933 30685 14967 30719
rect 15485 30685 15519 30719
rect 15945 30685 15979 30719
rect 16129 30685 16163 30719
rect 16865 30685 16899 30719
rect 17049 30685 17083 30719
rect 20821 30685 20855 30719
rect 23029 30685 23063 30719
rect 23305 30685 23339 30719
rect 25145 30685 25179 30719
rect 25605 30685 25639 30719
rect 25789 30685 25823 30719
rect 26157 30685 26191 30719
rect 27629 30685 27663 30719
rect 28089 30685 28123 30719
rect 28457 30685 28491 30719
rect 28641 30685 28675 30719
rect 27445 30345 27479 30379
rect 28365 30345 28399 30379
rect 29561 30277 29595 30311
rect 30757 30277 30791 30311
rect 14289 30209 14323 30243
rect 14933 30209 14967 30243
rect 19165 30209 19199 30243
rect 19717 30209 19751 30243
rect 21005 30209 21039 30243
rect 24685 30209 24719 30243
rect 25237 30209 25271 30243
rect 25329 30209 25363 30243
rect 25697 30209 25731 30243
rect 25881 30209 25915 30243
rect 26065 30209 26099 30243
rect 27383 30209 27417 30243
rect 28549 30209 28583 30243
rect 28825 30209 28859 30243
rect 29009 30209 29043 30243
rect 29745 30209 29779 30243
rect 29929 30209 29963 30243
rect 30389 30209 30423 30243
rect 30573 30209 30607 30243
rect 27905 30141 27939 30175
rect 27261 30073 27295 30107
rect 27813 30073 27847 30107
rect 13461 30005 13495 30039
rect 20913 30005 20947 30039
rect 14841 29801 14875 29835
rect 25145 29801 25179 29835
rect 27353 29733 27387 29767
rect 20453 29665 20487 29699
rect 21557 29665 21591 29699
rect 27633 29665 27667 29699
rect 9597 29597 9631 29631
rect 9781 29597 9815 29631
rect 9873 29597 9907 29631
rect 10333 29597 10367 29631
rect 10425 29597 10459 29631
rect 13001 29597 13035 29631
rect 13185 29597 13219 29631
rect 14933 29597 14967 29631
rect 19625 29597 19659 29631
rect 20177 29597 20211 29631
rect 21005 29597 21039 29631
rect 21373 29597 21407 29631
rect 24777 29597 24811 29631
rect 24961 29597 24995 29631
rect 27537 29597 27571 29631
rect 27721 29597 27755 29631
rect 27813 29597 27847 29631
rect 28365 29597 28399 29631
rect 28549 29597 28583 29631
rect 28917 29597 28951 29631
rect 10609 29529 10643 29563
rect 15117 29529 15151 29563
rect 9413 29461 9447 29495
rect 10333 29461 10367 29495
rect 12817 29461 12851 29495
rect 19533 29461 19567 29495
rect 21373 29461 21407 29495
rect 28825 29461 28859 29495
rect 14565 29257 14599 29291
rect 20269 29257 20303 29291
rect 22109 29257 22143 29291
rect 27537 29257 27571 29291
rect 28289 29257 28323 29291
rect 28457 29257 28491 29291
rect 8309 29189 8343 29223
rect 15393 29189 15427 29223
rect 17785 29189 17819 29223
rect 23673 29189 23707 29223
rect 25237 29189 25271 29223
rect 28089 29189 28123 29223
rect 8125 29121 8159 29155
rect 8401 29121 8435 29155
rect 9045 29121 9079 29155
rect 9321 29121 9355 29155
rect 9505 29121 9539 29155
rect 11805 29121 11839 29155
rect 12541 29121 12575 29155
rect 12633 29121 12667 29155
rect 12909 29121 12943 29155
rect 13185 29121 13219 29155
rect 14749 29121 14783 29155
rect 15577 29121 15611 29155
rect 15761 29121 15795 29155
rect 19257 29121 19291 29155
rect 19441 29121 19475 29155
rect 20453 29121 20487 29155
rect 20545 29121 20579 29155
rect 20729 29121 20763 29155
rect 20821 29121 20855 29155
rect 21281 29121 21315 29155
rect 21465 29121 21499 29155
rect 22293 29121 22327 29155
rect 22569 29121 22603 29155
rect 22753 29121 22787 29155
rect 25329 29121 25363 29155
rect 25605 29121 25639 29155
rect 27445 29121 27479 29155
rect 27629 29121 27663 29155
rect 28917 29121 28951 29155
rect 29101 29121 29135 29155
rect 14933 29053 14967 29087
rect 22385 29053 22419 29087
rect 29193 29053 29227 29087
rect 21373 28985 21407 29019
rect 22477 28985 22511 29019
rect 23213 28985 23247 29019
rect 23397 28985 23431 29019
rect 7941 28917 7975 28951
rect 9413 28917 9447 28951
rect 11805 28917 11839 28951
rect 28273 28917 28307 28951
rect 21097 28713 21131 28747
rect 28917 28713 28951 28747
rect 10977 28645 11011 28679
rect 15209 28645 15243 28679
rect 11621 28577 11655 28611
rect 13185 28577 13219 28611
rect 13369 28577 13403 28611
rect 20085 28577 20119 28611
rect 26249 28577 26283 28611
rect 9137 28509 9171 28543
rect 9321 28509 9355 28543
rect 11253 28509 11287 28543
rect 12081 28509 12115 28543
rect 12357 28509 12391 28543
rect 13093 28509 13127 28543
rect 13277 28509 13311 28543
rect 14565 28509 14599 28543
rect 14933 28509 14967 28543
rect 15393 28509 15427 28543
rect 16313 28509 16347 28543
rect 19717 28509 19751 28543
rect 19901 28509 19935 28543
rect 20545 28509 20579 28543
rect 20637 28509 20671 28543
rect 20821 28509 20855 28543
rect 20913 28509 20947 28543
rect 22845 28509 22879 28543
rect 23397 28509 23431 28543
rect 29009 28509 29043 28543
rect 16681 28441 16715 28475
rect 9229 28373 9263 28407
rect 12909 28373 12943 28407
rect 27261 28373 27295 28407
rect 15393 28169 15427 28203
rect 22385 28169 22419 28203
rect 15945 28101 15979 28135
rect 19349 28101 19383 28135
rect 20637 28101 20671 28135
rect 22845 28101 22879 28135
rect 7757 28033 7791 28067
rect 7849 28033 7883 28067
rect 8033 28033 8067 28067
rect 8769 28033 8803 28067
rect 8861 28033 8895 28067
rect 9045 28033 9079 28067
rect 12173 28033 12207 28067
rect 12541 28033 12575 28067
rect 12909 28033 12943 28067
rect 13369 28033 13403 28067
rect 13829 28033 13863 28067
rect 14013 28033 14047 28067
rect 14197 28033 14231 28067
rect 15393 28033 15427 28067
rect 19257 28033 19291 28067
rect 19441 28033 19475 28067
rect 20269 28033 20303 28067
rect 20545 28033 20579 28067
rect 25053 28033 25087 28067
rect 25697 28033 25731 28067
rect 27261 28033 27295 28067
rect 27537 28033 27571 28067
rect 30113 28033 30147 28067
rect 30297 28033 30331 28067
rect 30389 28033 30423 28067
rect 8953 27965 8987 27999
rect 12449 27965 12483 27999
rect 15301 27965 15335 27999
rect 25789 27965 25823 27999
rect 27169 27965 27203 27999
rect 22569 27897 22603 27931
rect 24869 27897 24903 27931
rect 8217 27829 8251 27863
rect 9229 27829 9263 27863
rect 29929 27829 29963 27863
rect 16865 27557 16899 27591
rect 25237 27557 25271 27591
rect 27905 27557 27939 27591
rect 12817 27489 12851 27523
rect 14381 27489 14415 27523
rect 22385 27489 22419 27523
rect 28457 27489 28491 27523
rect 9321 27421 9355 27455
rect 9505 27421 9539 27455
rect 9689 27421 9723 27455
rect 13185 27421 13219 27455
rect 13369 27421 13403 27455
rect 14933 27421 14967 27455
rect 15945 27421 15979 27455
rect 16037 27421 16071 27455
rect 16221 27421 16255 27455
rect 18245 27421 18279 27455
rect 22109 27421 22143 27455
rect 25421 27421 25455 27455
rect 25697 27421 25731 27455
rect 26065 27421 26099 27455
rect 26341 27421 26375 27455
rect 26709 27421 26743 27455
rect 27445 27421 27479 27455
rect 27721 27421 27755 27455
rect 28365 27421 28399 27455
rect 28549 27421 28583 27455
rect 29745 27421 29779 27455
rect 10149 27353 10183 27387
rect 16405 27353 16439 27387
rect 17978 27353 18012 27387
rect 29990 27353 30024 27387
rect 27537 27285 27571 27319
rect 31125 27285 31159 27319
rect 8309 27081 8343 27115
rect 12081 27081 12115 27115
rect 19533 27081 19567 27115
rect 20821 27081 20855 27115
rect 31125 27081 31159 27115
rect 15485 27013 15519 27047
rect 27537 27013 27571 27047
rect 8217 26945 8251 26979
rect 8493 26945 8527 26979
rect 9229 26945 9263 26979
rect 9321 26945 9355 26979
rect 11897 26945 11931 26979
rect 12173 26945 12207 26979
rect 13645 26945 13679 26979
rect 15669 26945 15703 26979
rect 15761 26945 15795 26979
rect 18245 26945 18279 26979
rect 20729 26945 20763 26979
rect 21005 26945 21039 26979
rect 22109 26945 22143 26979
rect 24961 26945 24995 26979
rect 25145 26945 25179 26979
rect 25605 26945 25639 26979
rect 25697 26945 25731 26979
rect 25881 26945 25915 26979
rect 27261 26945 27295 26979
rect 27353 26945 27387 26979
rect 30021 26945 30055 26979
rect 9045 26877 9079 26911
rect 9137 26877 9171 26911
rect 13737 26877 13771 26911
rect 22661 26877 22695 26911
rect 26433 26877 26467 26911
rect 29745 26877 29779 26911
rect 8493 26809 8527 26843
rect 9505 26741 9539 26775
rect 11713 26741 11747 26775
rect 21189 26741 21223 26775
rect 12357 26537 12391 26571
rect 13461 26537 13495 26571
rect 25237 26537 25271 26571
rect 27077 26537 27111 26571
rect 29193 26537 29227 26571
rect 9413 26469 9447 26503
rect 13277 26469 13311 26503
rect 25605 26469 25639 26503
rect 31309 26469 31343 26503
rect 11161 26401 11195 26435
rect 11713 26401 11747 26435
rect 12725 26401 12759 26435
rect 17969 26401 18003 26435
rect 11345 26333 11379 26367
rect 12633 26333 12667 26367
rect 15669 26333 15703 26367
rect 15945 26333 15979 26367
rect 18613 26333 18647 26367
rect 18889 26333 18923 26367
rect 25421 26333 25455 26367
rect 25513 26333 25547 26367
rect 25696 26333 25730 26367
rect 25881 26333 25915 26367
rect 26525 26333 26559 26367
rect 26617 26333 26651 26367
rect 26801 26333 26835 26367
rect 26893 26333 26927 26367
rect 27537 26333 27571 26367
rect 28733 26333 28767 26367
rect 28825 26333 28859 26367
rect 29009 26333 29043 26367
rect 9137 26265 9171 26299
rect 11621 26265 11655 26299
rect 13429 26265 13463 26299
rect 13645 26265 13679 26299
rect 16129 26265 16163 26299
rect 17702 26265 17736 26299
rect 18429 26265 18463 26299
rect 18797 26265 18831 26299
rect 22569 26265 22603 26299
rect 27813 26265 27847 26299
rect 30021 26265 30055 26299
rect 9597 26197 9631 26231
rect 15761 26197 15795 26231
rect 16589 26197 16623 26231
rect 21097 26197 21131 26231
rect 10602 25993 10636 26027
rect 12265 25993 12299 26027
rect 21373 25993 21407 26027
rect 23581 25993 23615 26027
rect 25605 25993 25639 26027
rect 27169 25993 27203 26027
rect 29929 25993 29963 26027
rect 10517 25925 10551 25959
rect 12449 25925 12483 25959
rect 13093 25925 13127 25959
rect 13369 25925 13403 25959
rect 24593 25925 24627 25959
rect 25145 25925 25179 25959
rect 28641 25925 28675 25959
rect 9505 25857 9539 25891
rect 9781 25857 9815 25891
rect 10425 25857 10459 25891
rect 10701 25857 10735 25891
rect 12357 25857 12391 25891
rect 13277 25857 13311 25891
rect 13466 25857 13500 25891
rect 16957 25857 16991 25891
rect 19625 25857 19659 25891
rect 21189 25857 21223 25891
rect 21465 25857 21499 25891
rect 22293 25857 22327 25891
rect 24501 25857 24535 25891
rect 24685 25857 24719 25891
rect 26525 25857 26559 25891
rect 27629 25857 27663 25891
rect 32321 25857 32355 25891
rect 32413 25857 32447 25891
rect 32597 25857 32631 25891
rect 9597 25789 9631 25823
rect 12081 25789 12115 25823
rect 22017 25789 22051 25823
rect 26617 25789 26651 25823
rect 27353 25789 27387 25823
rect 27445 25789 27479 25823
rect 27537 25789 27571 25823
rect 25421 25721 25455 25755
rect 9965 25653 9999 25687
rect 12633 25653 12667 25687
rect 13093 25653 13127 25687
rect 17233 25653 17267 25687
rect 18337 25653 18371 25687
rect 21005 25653 21039 25687
rect 32781 25653 32815 25687
rect 15393 25449 15427 25483
rect 19809 25449 19843 25483
rect 26065 25449 26099 25483
rect 26249 25449 26283 25483
rect 28273 25449 28307 25483
rect 31493 25449 31527 25483
rect 16313 25381 16347 25415
rect 3985 25313 4019 25347
rect 21189 25313 21223 25347
rect 24777 25313 24811 25347
rect 26617 25313 26651 25347
rect 4169 25245 4203 25279
rect 4261 25245 4295 25279
rect 6745 25245 6779 25279
rect 6929 25245 6963 25279
rect 12265 25245 12299 25279
rect 12541 25245 12575 25279
rect 12725 25245 12759 25279
rect 16037 25245 16071 25279
rect 16313 25245 16347 25279
rect 20922 25245 20956 25279
rect 24593 25245 24627 25279
rect 27291 25245 27325 25279
rect 27438 25245 27472 25279
rect 28365 25245 28399 25279
rect 30113 25245 30147 25279
rect 30380 25245 30414 25279
rect 15577 25177 15611 25211
rect 21649 25177 21683 25211
rect 26249 25177 26283 25211
rect 3985 25109 4019 25143
rect 6745 25109 6779 25143
rect 12081 25109 12115 25143
rect 15209 25109 15243 25143
rect 15377 25109 15411 25143
rect 16129 25109 16163 25143
rect 22937 25109 22971 25143
rect 27077 25109 27111 25143
rect 5273 24837 5307 24871
rect 21465 24837 21499 24871
rect 23673 24837 23707 24871
rect 25053 24837 25087 24871
rect 28641 24837 28675 24871
rect 28825 24837 28859 24871
rect 6929 24769 6963 24803
rect 14841 24769 14875 24803
rect 15117 24769 15151 24803
rect 15209 24769 15243 24803
rect 15393 24769 15427 24803
rect 15945 24769 15979 24803
rect 16129 24769 16163 24803
rect 18153 24769 18187 24803
rect 21005 24769 21039 24803
rect 21097 24769 21131 24803
rect 21281 24769 21315 24803
rect 25145 24769 25179 24803
rect 25329 24769 25363 24803
rect 26157 24769 26191 24803
rect 29101 24769 29135 24803
rect 30380 24769 30414 24803
rect 3709 24701 3743 24735
rect 3985 24701 4019 24735
rect 4721 24701 4755 24735
rect 7941 24701 7975 24735
rect 15301 24701 15335 24735
rect 17877 24701 17911 24735
rect 19349 24701 19383 24735
rect 22017 24701 22051 24735
rect 22293 24701 22327 24735
rect 26433 24701 26467 24735
rect 30113 24701 30147 24735
rect 2605 24565 2639 24599
rect 16129 24565 16163 24599
rect 25973 24565 26007 24599
rect 26341 24565 26375 24599
rect 28825 24565 28859 24599
rect 31493 24565 31527 24599
rect 3341 24361 3375 24395
rect 4629 24361 4663 24395
rect 6837 24361 6871 24395
rect 30481 24361 30515 24395
rect 2605 24293 2639 24327
rect 22753 24293 22787 24327
rect 3985 24225 4019 24259
rect 4077 24225 4111 24259
rect 5089 24225 5123 24259
rect 5457 24225 5491 24259
rect 20913 24225 20947 24259
rect 2329 24157 2363 24191
rect 3249 24157 3283 24191
rect 3433 24157 3467 24191
rect 4353 24157 4387 24191
rect 4445 24157 4479 24191
rect 5273 24157 5307 24191
rect 5365 24157 5399 24191
rect 5549 24157 5583 24191
rect 7573 24157 7607 24191
rect 8493 24157 8527 24191
rect 11989 24157 12023 24191
rect 12173 24157 12207 24191
rect 14473 24157 14507 24191
rect 14565 24157 14599 24191
rect 14749 24157 14783 24191
rect 14841 24157 14875 24191
rect 15761 24157 15795 24191
rect 15945 24157 15979 24191
rect 17049 24157 17083 24191
rect 17233 24157 17267 24191
rect 17877 24157 17911 24191
rect 18153 24157 18187 24191
rect 20545 24157 20579 24191
rect 20729 24157 20763 24191
rect 21373 24157 21407 24191
rect 23397 24157 23431 24191
rect 23673 24157 23707 24191
rect 25237 24157 25271 24191
rect 25421 24157 25455 24191
rect 30665 24157 30699 24191
rect 30951 24157 30985 24191
rect 2605 24089 2639 24123
rect 18061 24089 18095 24123
rect 21640 24089 21674 24123
rect 23213 24089 23247 24123
rect 2421 24021 2455 24055
rect 12173 24021 12207 24055
rect 14289 24021 14323 24055
rect 15577 24021 15611 24055
rect 17141 24021 17175 24055
rect 17693 24021 17727 24055
rect 23581 24021 23615 24055
rect 25237 24021 25271 24055
rect 30849 24021 30883 24055
rect 5089 23817 5123 23851
rect 8401 23817 8435 23851
rect 15117 23817 15151 23851
rect 15945 23817 15979 23851
rect 30113 23817 30147 23851
rect 4629 23749 4663 23783
rect 14933 23749 14967 23783
rect 19993 23749 20027 23783
rect 22293 23749 22327 23783
rect 28641 23749 28675 23783
rect 3341 23681 3375 23715
rect 4077 23681 4111 23715
rect 5273 23681 5307 23715
rect 5549 23681 5583 23715
rect 9229 23681 9263 23715
rect 9873 23681 9907 23715
rect 10057 23681 10091 23715
rect 12909 23681 12943 23715
rect 13277 23681 13311 23715
rect 14381 23681 14415 23715
rect 16129 23681 16163 23715
rect 16313 23681 16347 23715
rect 20545 23681 20579 23715
rect 20729 23681 20763 23715
rect 22661 23681 22695 23715
rect 5365 23613 5399 23647
rect 5457 23613 5491 23647
rect 6837 23613 6871 23647
rect 7113 23613 7147 23647
rect 9045 23613 9079 23647
rect 9413 23613 9447 23647
rect 12265 23613 12299 23647
rect 13001 23613 13035 23647
rect 13185 23613 13219 23647
rect 14841 23613 14875 23647
rect 15209 23613 15243 23647
rect 15301 23613 15335 23647
rect 20821 23613 20855 23647
rect 9965 23545 9999 23579
rect 14289 23545 14323 23579
rect 15485 23545 15519 23579
rect 18705 23545 18739 23579
rect 3341 23273 3375 23307
rect 6929 23273 6963 23307
rect 18705 23273 18739 23307
rect 21925 23273 21959 23307
rect 4629 23205 4663 23239
rect 9137 23205 9171 23239
rect 15669 23205 15703 23239
rect 16221 23205 16255 23239
rect 19717 23205 19751 23239
rect 4169 23137 4203 23171
rect 4721 23137 4755 23171
rect 8217 23137 8251 23171
rect 8309 23137 8343 23171
rect 8401 23137 8435 23171
rect 15301 23137 15335 23171
rect 15393 23137 15427 23171
rect 16589 23137 16623 23171
rect 17325 23137 17359 23171
rect 25237 23137 25271 23171
rect 28733 23137 28767 23171
rect 31033 23137 31067 23171
rect 32689 23137 32723 23171
rect 33149 23137 33183 23171
rect 3433 23069 3467 23103
rect 4353 23069 4387 23103
rect 7113 23069 7147 23103
rect 7297 23069 7331 23103
rect 7573 23069 7607 23103
rect 8125 23069 8159 23103
rect 9413 23069 9447 23103
rect 12081 23069 12115 23103
rect 15209 23069 15243 23103
rect 15485 23069 15519 23103
rect 17592 23069 17626 23103
rect 19441 23069 19475 23103
rect 19717 23069 19751 23103
rect 20637 23069 20671 23103
rect 24777 23069 24811 23103
rect 24869 23069 24903 23103
rect 25789 23069 25823 23103
rect 25881 23069 25915 23103
rect 27537 23069 27571 23103
rect 27997 23069 28031 23103
rect 28273 23069 28307 23103
rect 28917 23069 28951 23103
rect 31769 23069 31803 23103
rect 32045 23069 32079 23103
rect 32781 23069 32815 23103
rect 33609 23069 33643 23103
rect 33793 23069 33827 23103
rect 7205 23001 7239 23035
rect 7435 23001 7469 23035
rect 9137 23001 9171 23035
rect 11805 23001 11839 23035
rect 12541 23001 12575 23035
rect 13277 23001 13311 23035
rect 24593 23001 24627 23035
rect 27813 23001 27847 23035
rect 29101 23001 29135 23035
rect 8585 22933 8619 22967
rect 9321 22933 9355 22967
rect 10333 22933 10367 22967
rect 16129 22933 16163 22967
rect 24961 22933 24995 22967
rect 25145 22933 25179 22967
rect 33701 22933 33735 22967
rect 3785 22729 3819 22763
rect 7205 22729 7239 22763
rect 32413 22729 32447 22763
rect 3985 22661 4019 22695
rect 8125 22661 8159 22695
rect 8309 22661 8343 22695
rect 8493 22661 8527 22695
rect 9689 22661 9723 22695
rect 12541 22661 12575 22695
rect 14473 22661 14507 22695
rect 15577 22661 15611 22695
rect 18705 22661 18739 22695
rect 23673 22661 23707 22695
rect 25237 22661 25271 22695
rect 33057 22661 33091 22695
rect 33517 22661 33551 22695
rect 4905 22593 4939 22627
rect 7389 22593 7423 22627
rect 7573 22593 7607 22627
rect 7665 22593 7699 22627
rect 9413 22593 9447 22627
rect 9505 22593 9539 22627
rect 10333 22593 10367 22627
rect 11713 22593 11747 22627
rect 11897 22593 11931 22627
rect 12909 22593 12943 22627
rect 13185 22593 13219 22627
rect 13369 22593 13403 22627
rect 13645 22593 13679 22627
rect 13921 22593 13955 22627
rect 14749 22593 14783 22627
rect 15393 22593 15427 22627
rect 15669 22593 15703 22627
rect 17417 22593 17451 22627
rect 17601 22593 17635 22627
rect 18337 22593 18371 22627
rect 20085 22593 20119 22627
rect 20177 22593 20211 22627
rect 20361 22593 20395 22627
rect 20453 22593 20487 22627
rect 22017 22593 22051 22627
rect 22201 22593 22235 22627
rect 23581 22593 23615 22627
rect 24869 22593 24903 22627
rect 27997 22593 28031 22627
rect 28825 22593 28859 22627
rect 31033 22593 31067 22627
rect 31217 22593 31251 22627
rect 32689 22593 32723 22627
rect 33701 22593 33735 22627
rect 10977 22525 11011 22559
rect 14473 22525 14507 22559
rect 18245 22525 18279 22559
rect 24777 22525 24811 22559
rect 25145 22525 25179 22559
rect 31125 22525 31159 22559
rect 31309 22525 31343 22559
rect 32551 22525 32585 22559
rect 32965 22525 32999 22559
rect 17509 22457 17543 22491
rect 22017 22457 22051 22491
rect 3617 22389 3651 22423
rect 3801 22389 3835 22423
rect 4537 22389 4571 22423
rect 11805 22389 11839 22423
rect 14657 22389 14691 22423
rect 15209 22389 15243 22423
rect 18061 22389 18095 22423
rect 19901 22389 19935 22423
rect 24593 22389 24627 22423
rect 27353 22389 27387 22423
rect 30849 22389 30883 22423
rect 33793 22389 33827 22423
rect 11817 22185 11851 22219
rect 23029 22185 23063 22219
rect 23213 22185 23247 22219
rect 33517 22185 33551 22219
rect 12913 22117 12947 22151
rect 13001 22117 13035 22151
rect 18107 22049 18141 22083
rect 24869 22049 24903 22083
rect 24961 22049 24995 22083
rect 26985 22049 27019 22083
rect 30021 22049 30055 22083
rect 33149 22049 33183 22083
rect 7205 21981 7239 22015
rect 9321 21981 9355 22015
rect 12081 21981 12115 22015
rect 12817 21981 12851 22015
rect 13093 21981 13127 22015
rect 17969 21981 18003 22015
rect 18337 21981 18371 22015
rect 19625 21981 19659 22015
rect 19901 21981 19935 22015
rect 20821 21981 20855 22015
rect 23213 21981 23247 22015
rect 23397 21981 23431 22015
rect 24777 21981 24811 22015
rect 25053 21981 25087 22015
rect 26065 21981 26099 22015
rect 26249 21981 26283 22015
rect 27077 21981 27111 22015
rect 27813 21981 27847 22015
rect 28641 21981 28675 22015
rect 30113 21981 30147 22015
rect 31033 21981 31067 22015
rect 31401 21981 31435 22015
rect 31585 21981 31619 22015
rect 32045 21981 32079 22015
rect 32413 21981 32447 22015
rect 32597 21981 32631 22015
rect 33333 21981 33367 22015
rect 18245 21913 18279 21947
rect 28273 21913 28307 21947
rect 28457 21913 28491 21947
rect 31125 21913 31159 21947
rect 32137 21913 32171 21947
rect 7205 21845 7239 21879
rect 9229 21845 9263 21879
rect 10333 21845 10367 21879
rect 12633 21845 12667 21879
rect 19441 21845 19475 21879
rect 19809 21845 19843 21879
rect 22293 21845 22327 21879
rect 25237 21845 25271 21879
rect 26157 21845 26191 21879
rect 27721 21845 27755 21879
rect 29745 21845 29779 21879
rect 27169 21641 27203 21675
rect 30389 21641 30423 21675
rect 31677 21641 31711 21675
rect 11713 21573 11747 21607
rect 30573 21573 30607 21607
rect 2881 21505 2915 21539
rect 3801 21505 3835 21539
rect 4077 21505 4111 21539
rect 11805 21505 11839 21539
rect 11989 21505 12023 21539
rect 14473 21505 14507 21539
rect 15301 21505 15335 21539
rect 15485 21505 15519 21539
rect 19625 21505 19659 21539
rect 19901 21505 19935 21539
rect 20545 21505 20579 21539
rect 20637 21505 20671 21539
rect 22017 21505 22051 21539
rect 22293 21505 22327 21539
rect 27537 21505 27571 21539
rect 28181 21505 28215 21539
rect 28365 21505 28399 21539
rect 30297 21505 30331 21539
rect 31493 21505 31527 21539
rect 31677 21505 31711 21539
rect 3157 21437 3191 21471
rect 3893 21437 3927 21471
rect 22385 21437 22419 21471
rect 23213 21437 23247 21471
rect 23489 21437 23523 21471
rect 24593 21437 24627 21471
rect 27445 21437 27479 21471
rect 2973 21369 3007 21403
rect 3985 21369 4019 21403
rect 3065 21301 3099 21335
rect 3617 21301 3651 21335
rect 14565 21301 14599 21335
rect 15485 21301 15519 21335
rect 19441 21301 19475 21335
rect 28365 21301 28399 21335
rect 30573 21301 30607 21335
rect 13461 21097 13495 21131
rect 14657 21097 14691 21131
rect 16129 21097 16163 21131
rect 18797 21097 18831 21131
rect 21281 21097 21315 21131
rect 23581 21097 23615 21131
rect 31493 21097 31527 21131
rect 32413 21097 32447 21131
rect 7389 20961 7423 20995
rect 20177 20961 20211 20995
rect 20269 20961 20303 20995
rect 33057 20961 33091 20995
rect 3249 20893 3283 20927
rect 3433 20893 3467 20927
rect 7573 20893 7607 20927
rect 7665 20893 7699 20927
rect 10425 20893 10459 20927
rect 10701 20893 10735 20927
rect 13553 20893 13587 20927
rect 14473 20893 14507 20927
rect 14657 20893 14691 20927
rect 17417 20893 17451 20927
rect 19809 20893 19843 20927
rect 19901 20893 19935 20927
rect 22569 20893 22603 20927
rect 23765 20893 23799 20927
rect 23949 20893 23983 20927
rect 24041 20893 24075 20927
rect 24777 20893 24811 20927
rect 25053 20893 25087 20927
rect 31584 20893 31618 20927
rect 31677 20893 31711 20927
rect 32229 20893 32263 20927
rect 32413 20893 32447 20927
rect 32965 20893 32999 20927
rect 33149 20893 33183 20927
rect 10609 20825 10643 20859
rect 18521 20825 18555 20859
rect 24593 20825 24627 20859
rect 3341 20757 3375 20791
rect 7389 20757 7423 20791
rect 10241 20757 10275 20791
rect 14289 20757 14323 20791
rect 19625 20757 19659 20791
rect 24961 20757 24995 20791
rect 7849 20553 7883 20587
rect 8401 20553 8435 20587
rect 21005 20553 21039 20587
rect 22201 20553 22235 20587
rect 31585 20553 31619 20587
rect 32597 20553 32631 20587
rect 3617 20485 3651 20519
rect 7481 20485 7515 20519
rect 20637 20485 20671 20519
rect 20729 20485 20763 20519
rect 23213 20485 23247 20519
rect 3157 20417 3191 20451
rect 3249 20417 3283 20451
rect 4445 20417 4479 20451
rect 7389 20417 7423 20451
rect 7665 20417 7699 20451
rect 8309 20417 8343 20451
rect 8493 20417 8527 20451
rect 8585 20417 8619 20451
rect 11069 20417 11103 20451
rect 13461 20417 13495 20451
rect 13829 20417 13863 20451
rect 14013 20417 14047 20451
rect 15117 20417 15151 20451
rect 15669 20417 15703 20451
rect 15853 20417 15887 20451
rect 19993 20417 20027 20451
rect 20453 20417 20487 20451
rect 20821 20417 20855 20451
rect 22109 20417 22143 20451
rect 27997 20417 28031 20451
rect 31585 20417 31619 20451
rect 31769 20417 31803 20451
rect 32781 20417 32815 20451
rect 33057 20417 33091 20451
rect 3525 20349 3559 20383
rect 4077 20349 4111 20383
rect 4353 20349 4387 20383
rect 10425 20349 10459 20383
rect 12817 20349 12851 20383
rect 13553 20349 13587 20383
rect 14749 20349 14783 20383
rect 16037 20349 16071 20383
rect 27905 20349 27939 20383
rect 24501 20281 24535 20315
rect 32965 20281 32999 20315
rect 2973 20213 3007 20247
rect 18705 20213 18739 20247
rect 27629 20213 27663 20247
rect 27997 20213 28031 20247
rect 3985 20009 4019 20043
rect 5089 20009 5123 20043
rect 7573 20009 7607 20043
rect 14565 20009 14599 20043
rect 20085 20009 20119 20043
rect 7113 19941 7147 19975
rect 7757 19941 7791 19975
rect 9137 19941 9171 19975
rect 32321 19941 32355 19975
rect 2421 19873 2455 19907
rect 10517 19873 10551 19907
rect 11897 19873 11931 19907
rect 13737 19873 13771 19907
rect 17417 19873 17451 19907
rect 22569 19873 22603 19907
rect 1685 19805 1719 19839
rect 1869 19805 1903 19839
rect 2881 19805 2915 19839
rect 3157 19805 3191 19839
rect 4169 19805 4203 19839
rect 4537 19805 4571 19839
rect 4629 19805 4663 19839
rect 5273 19805 5307 19839
rect 5457 19805 5491 19839
rect 6837 19805 6871 19839
rect 6929 19805 6963 19839
rect 7113 19805 7147 19839
rect 8033 19805 8067 19839
rect 9413 19805 9447 19839
rect 10425 19805 10459 19839
rect 10793 19805 10827 19839
rect 10885 19805 10919 19839
rect 11713 19805 11747 19839
rect 13369 19805 13403 19839
rect 13553 19805 13587 19839
rect 14473 19805 14507 19839
rect 15393 19805 15427 19839
rect 15669 19805 15703 19839
rect 16221 19805 16255 19839
rect 17969 19805 18003 19839
rect 19441 19805 19475 19839
rect 19534 19805 19568 19839
rect 19809 19805 19843 19839
rect 19906 19805 19940 19839
rect 28549 19805 28583 19839
rect 28825 19805 28859 19839
rect 29009 19805 29043 19839
rect 31953 19805 31987 19839
rect 32229 19805 32263 19839
rect 32413 19805 32447 19839
rect 32597 19805 32631 19839
rect 4261 19737 4295 19771
rect 4353 19737 4387 19771
rect 9137 19737 9171 19771
rect 9321 19737 9355 19771
rect 16773 19737 16807 19771
rect 19717 19737 19751 19771
rect 20821 19737 20855 19771
rect 1869 19669 1903 19703
rect 11529 19669 11563 19703
rect 15209 19669 15243 19703
rect 15577 19669 15611 19703
rect 28365 19669 28399 19703
rect 16313 19465 16347 19499
rect 17233 19465 17267 19499
rect 20821 19465 20855 19499
rect 22109 19465 22143 19499
rect 32689 19465 32723 19499
rect 32873 19465 32907 19499
rect 24777 19397 24811 19431
rect 32321 19397 32355 19431
rect 32505 19397 32539 19431
rect 2513 19329 2547 19363
rect 2789 19329 2823 19363
rect 4629 19329 4663 19363
rect 4813 19329 4847 19363
rect 4905 19329 4939 19363
rect 7113 19329 7147 19363
rect 7380 19329 7414 19363
rect 9045 19329 9079 19363
rect 9229 19329 9263 19363
rect 10793 19329 10827 19363
rect 12449 19329 12483 19363
rect 12725 19329 12759 19363
rect 15200 19329 15234 19363
rect 16865 19329 16899 19363
rect 17049 19329 17083 19363
rect 17325 19329 17359 19363
rect 19441 19329 19475 19363
rect 19708 19329 19742 19363
rect 22017 19329 22051 19363
rect 22293 19329 22327 19363
rect 23121 19329 23155 19363
rect 27261 19329 27295 19363
rect 27445 19329 27479 19363
rect 28825 19329 28859 19363
rect 29101 19329 29135 19363
rect 29377 19329 29411 19363
rect 29745 19329 29779 19363
rect 31217 19329 31251 19363
rect 31309 19329 31343 19363
rect 32597 19329 32631 19363
rect 10517 19261 10551 19295
rect 14933 19261 14967 19295
rect 22477 19261 22511 19295
rect 23397 19261 23431 19295
rect 28733 19261 28767 19295
rect 31493 19261 31527 19295
rect 4629 19193 4663 19227
rect 4077 19125 4111 19159
rect 8493 19125 8527 19159
rect 9137 19125 9171 19159
rect 10241 19125 10275 19159
rect 10701 19125 10735 19159
rect 27353 19125 27387 19159
rect 7665 18921 7699 18955
rect 16589 18921 16623 18955
rect 18613 18921 18647 18955
rect 25881 18921 25915 18955
rect 28273 18921 28307 18955
rect 33149 18921 33183 18955
rect 3157 18853 3191 18887
rect 7849 18785 7883 18819
rect 7941 18785 7975 18819
rect 8217 18785 8251 18819
rect 26065 18785 26099 18819
rect 26157 18785 26191 18819
rect 28733 18785 28767 18819
rect 28917 18785 28951 18819
rect 31861 18785 31895 18819
rect 32781 18785 32815 18819
rect 3341 18717 3375 18751
rect 3433 18717 3467 18751
rect 8309 18717 8343 18751
rect 10425 18717 10459 18751
rect 10517 18717 10551 18751
rect 11989 18717 12023 18751
rect 12265 18717 12299 18751
rect 15209 18717 15243 18751
rect 15465 18717 15499 18751
rect 18889 18717 18923 18751
rect 19441 18717 19475 18751
rect 23765 18717 23799 18751
rect 24041 18717 24075 18751
rect 24777 18717 24811 18751
rect 25053 18717 25087 18751
rect 26249 18717 26283 18751
rect 26342 18717 26376 18751
rect 27353 18717 27387 18751
rect 27537 18717 27571 18751
rect 28641 18717 28675 18751
rect 29009 18717 29043 18751
rect 29745 18717 29779 18751
rect 29837 18717 29871 18751
rect 30021 18717 30055 18751
rect 32045 18717 32079 18751
rect 32229 18717 32263 18751
rect 32689 18717 32723 18751
rect 32965 18717 32999 18751
rect 3157 18649 3191 18683
rect 12357 18649 12391 18683
rect 18429 18649 18463 18683
rect 8033 18581 8067 18615
rect 18613 18581 18647 18615
rect 20729 18581 20763 18615
rect 23581 18581 23615 18615
rect 23949 18581 23983 18615
rect 24593 18581 24627 18615
rect 24961 18581 24995 18615
rect 27261 18581 27295 18615
rect 8217 18377 8251 18411
rect 17141 18377 17175 18411
rect 20085 18377 20119 18411
rect 20913 18377 20947 18411
rect 25697 18377 25731 18411
rect 28825 18377 28859 18411
rect 32781 18377 32815 18411
rect 6837 18309 6871 18343
rect 14749 18309 14783 18343
rect 16221 18309 16255 18343
rect 17325 18309 17359 18343
rect 18972 18309 19006 18343
rect 24869 18309 24903 18343
rect 8033 18241 8067 18275
rect 8217 18241 8251 18275
rect 10333 18241 10367 18275
rect 12357 18241 12391 18275
rect 12449 18241 12483 18275
rect 13001 18241 13035 18275
rect 16037 18241 16071 18275
rect 16313 18241 16347 18275
rect 18705 18241 18739 18275
rect 20729 18241 20763 18275
rect 21005 18241 21039 18275
rect 23489 18241 23523 18275
rect 25329 18241 25363 18275
rect 28181 18241 28215 18275
rect 29009 18241 29043 18275
rect 29193 18241 29227 18275
rect 29285 18241 29319 18275
rect 32505 18241 32539 18275
rect 6745 18173 6779 18207
rect 6929 18173 6963 18207
rect 12173 18173 12207 18207
rect 23213 18173 23247 18207
rect 25421 18173 25455 18207
rect 27813 18173 27847 18207
rect 28273 18173 28307 18207
rect 32321 18173 32355 18207
rect 32873 18173 32907 18207
rect 34345 18173 34379 18207
rect 7297 18105 7331 18139
rect 10241 18037 10275 18071
rect 15853 18037 15887 18071
rect 16957 18037 16991 18071
rect 17141 18037 17175 18071
rect 20545 18037 20579 18071
rect 25329 18037 25363 18071
rect 6469 17833 6503 17867
rect 27997 17833 28031 17867
rect 30757 17833 30791 17867
rect 32689 17833 32723 17867
rect 3433 17765 3467 17799
rect 28549 17765 28583 17799
rect 27629 17697 27663 17731
rect 27813 17697 27847 17731
rect 33609 17697 33643 17731
rect 3249 17629 3283 17663
rect 6377 17629 6411 17663
rect 6561 17629 6595 17663
rect 13093 17629 13127 17663
rect 16957 17629 16991 17663
rect 19441 17629 19475 17663
rect 19708 17629 19742 17663
rect 25237 17629 25271 17663
rect 27537 17629 27571 17663
rect 27721 17629 27755 17663
rect 28549 17629 28583 17663
rect 28825 17629 28859 17663
rect 30941 17629 30975 17663
rect 31769 17629 31803 17663
rect 31953 17629 31987 17663
rect 32597 17629 32631 17663
rect 33241 17629 33275 17663
rect 33425 17629 33459 17663
rect 2881 17561 2915 17595
rect 12817 17561 12851 17595
rect 15209 17561 15243 17595
rect 24961 17561 24995 17595
rect 28641 17561 28675 17595
rect 31125 17561 31159 17595
rect 31861 17561 31895 17595
rect 32413 17561 32447 17595
rect 3065 17493 3099 17527
rect 3157 17493 3191 17527
rect 11345 17493 11379 17527
rect 20821 17493 20855 17527
rect 4445 17289 4479 17323
rect 24501 17289 24535 17323
rect 25697 17289 25731 17323
rect 29837 17289 29871 17323
rect 30757 17289 30791 17323
rect 30941 17289 30975 17323
rect 32521 17289 32555 17323
rect 32689 17289 32723 17323
rect 33241 17289 33275 17323
rect 2973 17221 3007 17255
rect 9597 17221 9631 17255
rect 13277 17221 13311 17255
rect 20821 17221 20855 17255
rect 21189 17221 21223 17255
rect 23388 17221 23422 17255
rect 25329 17221 25363 17255
rect 25421 17221 25455 17255
rect 30849 17221 30883 17255
rect 31493 17221 31527 17255
rect 32321 17221 32355 17255
rect 6745 17153 6779 17187
rect 7113 17153 7147 17187
rect 7573 17153 7607 17187
rect 8033 17153 8067 17187
rect 8217 17153 8251 17187
rect 9873 17153 9907 17187
rect 13553 17153 13587 17187
rect 16221 17153 16255 17187
rect 19156 17153 19190 17187
rect 25053 17153 25087 17187
rect 25146 17153 25180 17187
rect 25518 17153 25552 17187
rect 29745 17153 29779 17187
rect 29929 17153 29963 17187
rect 30481 17153 30515 17187
rect 30625 17153 30659 17187
rect 31677 17153 31711 17187
rect 31769 17153 31803 17187
rect 33149 17153 33183 17187
rect 33333 17153 33367 17187
rect 2697 17085 2731 17119
rect 6653 17085 6687 17119
rect 9781 17085 9815 17119
rect 15945 17085 15979 17119
rect 18889 17085 18923 17119
rect 23121 17085 23155 17119
rect 31493 17017 31527 17051
rect 8217 16949 8251 16983
rect 9689 16949 9723 16983
rect 10057 16949 10091 16983
rect 11805 16949 11839 16983
rect 20269 16949 20303 16983
rect 32505 16949 32539 16983
rect 3065 16745 3099 16779
rect 3249 16745 3283 16779
rect 4261 16745 4295 16779
rect 7343 16745 7377 16779
rect 9781 16745 9815 16779
rect 12265 16745 12299 16779
rect 19441 16745 19475 16779
rect 22109 16745 22143 16779
rect 31217 16745 31251 16779
rect 32229 16745 32263 16779
rect 5917 16677 5951 16711
rect 7205 16677 7239 16711
rect 14841 16677 14875 16711
rect 6745 16609 6779 16643
rect 7113 16609 7147 16643
rect 15301 16609 15335 16643
rect 20729 16609 20763 16643
rect 32597 16609 32631 16643
rect 4077 16541 4111 16575
rect 4353 16541 4387 16575
rect 9689 16541 9723 16575
rect 9905 16541 9939 16575
rect 10057 16541 10091 16575
rect 12173 16541 12207 16575
rect 12449 16541 12483 16575
rect 14381 16541 14415 16575
rect 14657 16541 14691 16575
rect 15568 16541 15602 16575
rect 17233 16541 17267 16575
rect 19625 16541 19659 16575
rect 19809 16541 19843 16575
rect 19901 16541 19935 16575
rect 24593 16541 24627 16575
rect 26433 16541 26467 16575
rect 30021 16541 30055 16575
rect 31401 16541 31435 16575
rect 31493 16541 31527 16575
rect 31621 16541 31655 16575
rect 32413 16541 32447 16575
rect 3433 16473 3467 16507
rect 5549 16473 5583 16507
rect 7481 16473 7515 16507
rect 17601 16473 17635 16507
rect 20996 16473 21030 16507
rect 24860 16473 24894 16507
rect 26709 16473 26743 16507
rect 29745 16473 29779 16507
rect 29929 16473 29963 16507
rect 31217 16473 31251 16507
rect 3233 16405 3267 16439
rect 6009 16405 6043 16439
rect 10241 16405 10275 16439
rect 14473 16405 14507 16439
rect 16681 16405 16715 16439
rect 25973 16405 26007 16439
rect 30113 16405 30147 16439
rect 30297 16405 30331 16439
rect 6745 16201 6779 16235
rect 10977 16201 11011 16235
rect 13553 16201 13587 16235
rect 18705 16201 18739 16235
rect 22661 16201 22695 16235
rect 25973 16201 26007 16235
rect 29009 16201 29043 16235
rect 33701 16201 33735 16235
rect 5733 16133 5767 16167
rect 8953 16133 8987 16167
rect 14105 16133 14139 16167
rect 15200 16133 15234 16167
rect 17785 16133 17819 16167
rect 19993 16133 20027 16167
rect 20729 16133 20763 16167
rect 20821 16133 20855 16167
rect 26341 16133 26375 16167
rect 29285 16133 29319 16167
rect 5549 16065 5583 16099
rect 6561 16065 6595 16099
rect 6745 16065 6779 16099
rect 7389 16065 7423 16099
rect 8861 16065 8895 16099
rect 10425 16065 10459 16099
rect 10977 16065 11011 16099
rect 11161 16065 11195 16099
rect 13369 16065 13403 16099
rect 14289 16065 14323 16099
rect 14473 16065 14507 16099
rect 17417 16065 17451 16099
rect 17601 16065 17635 16099
rect 20453 16065 20487 16099
rect 20546 16065 20580 16099
rect 20959 16065 20993 16099
rect 22017 16065 22051 16099
rect 22110 16065 22144 16099
rect 22293 16065 22327 16099
rect 22385 16065 22419 16099
rect 22523 16065 22557 16099
rect 25145 16065 25179 16099
rect 26157 16065 26191 16099
rect 26433 16065 26467 16099
rect 28181 16065 28215 16099
rect 28457 16065 28491 16099
rect 29193 16065 29227 16099
rect 29377 16065 29411 16099
rect 29561 16065 29595 16099
rect 32588 16065 32622 16099
rect 5365 15997 5399 16031
rect 7665 15997 7699 16031
rect 14933 15997 14967 16031
rect 28273 15997 28307 16031
rect 28365 15997 28399 16031
rect 32321 15997 32355 16031
rect 7941 15929 7975 15963
rect 21097 15929 21131 15963
rect 27997 15929 28031 15963
rect 7757 15861 7791 15895
rect 16313 15861 16347 15895
rect 23857 15861 23891 15895
rect 5273 15657 5307 15691
rect 18061 15657 18095 15691
rect 19901 15657 19935 15691
rect 26525 15657 26559 15691
rect 29101 15657 29135 15691
rect 31677 15657 31711 15691
rect 33885 15657 33919 15691
rect 13645 15589 13679 15623
rect 22569 15521 22603 15555
rect 2697 15453 2731 15487
rect 2881 15453 2915 15487
rect 6101 15453 6135 15487
rect 6285 15453 6319 15487
rect 6745 15453 6779 15487
rect 12541 15453 12575 15487
rect 12633 15453 12667 15487
rect 13369 15453 13403 15487
rect 13645 15453 13679 15487
rect 14289 15453 14323 15487
rect 16221 15453 16255 15487
rect 16405 15453 16439 15487
rect 17969 15453 18003 15487
rect 20821 15453 20855 15487
rect 23397 15453 23431 15487
rect 23673 15453 23707 15487
rect 29193 15453 29227 15487
rect 33425 15453 33459 15487
rect 33701 15453 33735 15487
rect 2973 15385 3007 15419
rect 5457 15385 5491 15419
rect 6193 15385 6227 15419
rect 14565 15385 14599 15419
rect 17785 15385 17819 15419
rect 20177 15385 20211 15419
rect 25237 15385 25271 15419
rect 32965 15385 32999 15419
rect 5089 15317 5123 15351
rect 5257 15317 5291 15351
rect 6837 15317 6871 15351
rect 16405 15317 16439 15351
rect 23213 15317 23247 15351
rect 23581 15317 23615 15351
rect 33517 15317 33551 15351
rect 5448 15113 5482 15147
rect 16037 15113 16071 15147
rect 22937 15113 22971 15147
rect 23305 15113 23339 15147
rect 33609 15113 33643 15147
rect 5825 15045 5859 15079
rect 9689 15045 9723 15079
rect 16865 15045 16899 15079
rect 19993 15045 20027 15079
rect 29929 15045 29963 15079
rect 4169 14977 4203 15011
rect 9045 14977 9079 15011
rect 9229 14977 9263 15011
rect 10517 14977 10551 15011
rect 10701 14977 10735 15011
rect 16129 14977 16163 15011
rect 16313 14977 16347 15011
rect 17049 14977 17083 15011
rect 17417 14977 17451 15011
rect 18245 14977 18279 15011
rect 20453 14977 20487 15011
rect 22201 14977 22235 15011
rect 22385 14977 22419 15011
rect 22477 14977 22511 15011
rect 23121 14977 23155 15011
rect 23397 14977 23431 15011
rect 25062 14977 25096 15011
rect 32321 14977 32355 15011
rect 1685 14909 1719 14943
rect 1961 14909 1995 14943
rect 4077 14909 4111 14943
rect 8953 14909 8987 14943
rect 10425 14909 10459 14943
rect 11161 14909 11195 14943
rect 20729 14909 20763 14943
rect 25329 14909 25363 14943
rect 3433 14841 3467 14875
rect 29745 14841 29779 14875
rect 5273 14773 5307 14807
rect 5457 14773 5491 14807
rect 22017 14773 22051 14807
rect 23949 14773 23983 14807
rect 6193 14569 6227 14603
rect 7205 14569 7239 14603
rect 14381 14569 14415 14603
rect 23765 14569 23799 14603
rect 23949 14569 23983 14603
rect 25973 14569 26007 14603
rect 28733 14569 28767 14603
rect 8493 14501 8527 14535
rect 9229 14501 9263 14535
rect 21005 14501 21039 14535
rect 18521 14433 18555 14467
rect 19625 14433 19659 14467
rect 24593 14433 24627 14467
rect 31401 14433 31435 14467
rect 31861 14433 31895 14467
rect 2697 14365 2731 14399
rect 2881 14365 2915 14399
rect 6101 14365 6135 14399
rect 6377 14365 6411 14399
rect 12817 14365 12851 14399
rect 12909 14365 12943 14399
rect 14289 14365 14323 14399
rect 14473 14365 14507 14399
rect 15577 14365 15611 14399
rect 17785 14365 17819 14399
rect 18245 14365 18279 14399
rect 21649 14365 21683 14399
rect 21741 14365 21775 14399
rect 22017 14365 22051 14399
rect 24849 14365 24883 14399
rect 26433 14365 26467 14399
rect 28273 14365 28307 14399
rect 28549 14365 28583 14399
rect 31125 14365 31159 14399
rect 32137 14365 32171 14399
rect 2973 14297 3007 14331
rect 7021 14297 7055 14331
rect 7941 14297 7975 14331
rect 8217 14297 8251 14331
rect 9505 14297 9539 14331
rect 9689 14297 9723 14331
rect 9781 14297 9815 14331
rect 13093 14297 13127 14331
rect 17325 14297 17359 14331
rect 19892 14297 19926 14331
rect 21833 14297 21867 14331
rect 23581 14297 23615 14331
rect 26700 14297 26734 14331
rect 29745 14297 29779 14331
rect 6561 14229 6595 14263
rect 7221 14229 7255 14263
rect 7389 14229 7423 14263
rect 8033 14229 8067 14263
rect 21465 14229 21499 14263
rect 23765 14229 23799 14263
rect 27813 14229 27847 14263
rect 28365 14229 28399 14263
rect 33241 14229 33275 14263
rect 2605 14025 2639 14059
rect 5917 14025 5951 14059
rect 8309 14025 8343 14059
rect 20729 14025 20763 14059
rect 24685 14025 24719 14059
rect 25053 14025 25087 14059
rect 28917 14025 28951 14059
rect 29101 14025 29135 14059
rect 30113 14025 30147 14059
rect 31401 14025 31435 14059
rect 33701 14025 33735 14059
rect 4445 13957 4479 13991
rect 6561 13957 6595 13991
rect 6745 13957 6779 13991
rect 9597 13957 9631 13991
rect 12081 13957 12115 13991
rect 14657 13957 14691 13991
rect 19441 13957 19475 13991
rect 19625 13957 19659 13991
rect 27629 13957 27663 13991
rect 28733 13957 28767 13991
rect 2697 13889 2731 13923
rect 7021 13889 7055 13923
rect 10149 13889 10183 13923
rect 10241 13889 10275 13923
rect 14105 13889 14139 13923
rect 14289 13889 14323 13923
rect 15209 13889 15243 13923
rect 15577 13889 15611 13923
rect 17141 13889 17175 13923
rect 17325 13889 17359 13923
rect 20545 13889 20579 13923
rect 24593 13889 24627 13923
rect 24869 13889 24903 13923
rect 27399 13889 27433 13923
rect 27537 13889 27571 13923
rect 27721 13889 27755 13923
rect 29653 13889 29687 13923
rect 29745 13889 29779 13923
rect 29929 13889 29963 13923
rect 31309 13889 31343 13923
rect 31585 13889 31619 13923
rect 31769 13889 31803 13923
rect 32597 13889 32631 13923
rect 4169 13821 4203 13855
rect 11805 13821 11839 13855
rect 13553 13821 13587 13855
rect 17601 13821 17635 13855
rect 27261 13821 27295 13855
rect 32321 13821 32355 13855
rect 15761 13753 15795 13787
rect 6745 13685 6779 13719
rect 10149 13685 10183 13719
rect 19625 13685 19659 13719
rect 19809 13685 19843 13719
rect 27905 13685 27939 13719
rect 28917 13685 28951 13719
rect 3433 13481 3467 13515
rect 5457 13481 5491 13515
rect 14381 13481 14415 13515
rect 16313 13481 16347 13515
rect 27353 13481 27387 13515
rect 31677 13481 31711 13515
rect 9137 13345 9171 13379
rect 11805 13345 11839 13379
rect 12081 13345 12115 13379
rect 18613 13345 18647 13379
rect 2329 13277 2363 13311
rect 2513 13277 2547 13311
rect 2973 13277 3007 13311
rect 3065 13277 3099 13311
rect 3249 13277 3283 13311
rect 4629 13277 4663 13311
rect 5273 13277 5307 13311
rect 5457 13277 5491 13311
rect 8309 13277 8343 13311
rect 8401 13277 8435 13311
rect 14289 13277 14323 13311
rect 14841 13277 14875 13311
rect 15669 13277 15703 13311
rect 16589 13277 16623 13311
rect 17969 13277 18003 13311
rect 18337 13277 18371 13311
rect 20637 13277 20671 13311
rect 26065 13277 26099 13311
rect 32965 13277 32999 13311
rect 4261 13209 4295 13243
rect 8585 13209 8619 13243
rect 9413 13209 9447 13243
rect 2421 13141 2455 13175
rect 10885 13141 10919 13175
rect 13553 13141 13587 13175
rect 21925 13141 21959 13175
rect 4445 12937 4479 12971
rect 20453 12937 20487 12971
rect 27905 12937 27939 12971
rect 32321 12937 32355 12971
rect 32689 12937 32723 12971
rect 2421 12869 2455 12903
rect 9505 12869 9539 12903
rect 13001 12869 13035 12903
rect 14749 12869 14783 12903
rect 18429 12869 18463 12903
rect 27629 12869 27663 12903
rect 28733 12869 28767 12903
rect 2145 12801 2179 12835
rect 4353 12801 4387 12835
rect 4537 12801 4571 12835
rect 15393 12801 15427 12835
rect 16037 12801 16071 12835
rect 16957 12801 16991 12835
rect 17141 12801 17175 12835
rect 17693 12801 17727 12835
rect 18245 12801 18279 12835
rect 20637 12801 20671 12835
rect 20729 12801 20763 12835
rect 20913 12801 20947 12835
rect 21005 12801 21039 12835
rect 27261 12801 27295 12835
rect 27409 12801 27443 12835
rect 27537 12801 27571 12835
rect 27726 12801 27760 12835
rect 28549 12801 28583 12835
rect 28825 12801 28859 12835
rect 29745 12801 29779 12835
rect 32505 12801 32539 12835
rect 32781 12801 32815 12835
rect 3893 12733 3927 12767
rect 9781 12733 9815 12767
rect 16129 12733 16163 12767
rect 17233 12733 17267 12767
rect 29561 12733 29595 12767
rect 8033 12597 8067 12631
rect 28365 12597 28399 12631
rect 3157 12393 3191 12427
rect 27905 12325 27939 12359
rect 15301 12257 15335 12291
rect 16681 12257 16715 12291
rect 22569 12257 22603 12291
rect 3157 12189 3191 12223
rect 3341 12189 3375 12223
rect 14565 12189 14599 12223
rect 15209 12189 15243 12223
rect 15945 12189 15979 12223
rect 16589 12189 16623 12223
rect 17601 12189 17635 12223
rect 17969 12189 18003 12223
rect 24777 12189 24811 12223
rect 25053 12189 25087 12223
rect 28084 12189 28118 12223
rect 28456 12189 28490 12223
rect 28549 12189 28583 12223
rect 18245 12121 18279 12155
rect 20821 12121 20855 12155
rect 28181 12121 28215 12155
rect 28273 12121 28307 12155
rect 24593 12053 24627 12087
rect 24961 12053 24995 12087
rect 21097 11849 21131 11883
rect 28733 11849 28767 11883
rect 31309 11849 31343 11883
rect 32689 11849 32723 11883
rect 15761 11781 15795 11815
rect 18521 11781 18555 11815
rect 25697 11781 25731 11815
rect 25881 11781 25915 11815
rect 27620 11781 27654 11815
rect 15945 11713 15979 11747
rect 16957 11713 16991 11747
rect 17141 11713 17175 11747
rect 18061 11713 18095 11747
rect 18245 11713 18279 11747
rect 19717 11713 19751 11747
rect 19984 11713 20018 11747
rect 22017 11713 22051 11747
rect 22273 11713 22307 11747
rect 24124 11713 24158 11747
rect 31217 11713 31251 11747
rect 31493 11713 31527 11747
rect 32505 11713 32539 11747
rect 32781 11713 32815 11747
rect 16221 11645 16255 11679
rect 23857 11645 23891 11679
rect 27353 11645 27387 11679
rect 17233 11577 17267 11611
rect 23397 11509 23431 11543
rect 25237 11509 25271 11543
rect 25881 11509 25915 11543
rect 26065 11509 26099 11543
rect 31677 11509 31711 11543
rect 32321 11509 32355 11543
rect 4169 11305 4203 11339
rect 21557 11305 21591 11339
rect 22845 11305 22879 11339
rect 31493 11305 31527 11339
rect 13645 11237 13679 11271
rect 3249 11101 3283 11135
rect 3433 11101 3467 11135
rect 5549 11101 5583 11135
rect 10333 11101 10367 11135
rect 10600 11101 10634 11135
rect 12725 11101 12759 11135
rect 13093 11101 13127 11135
rect 16865 11101 16899 11135
rect 17049 11101 17083 11135
rect 17601 11101 17635 11135
rect 18061 11101 18095 11135
rect 19993 11101 20027 11135
rect 20086 11101 20120 11135
rect 20269 11101 20303 11135
rect 20361 11101 20395 11135
rect 20499 11101 20533 11135
rect 21097 11101 21131 11135
rect 21373 11101 21407 11135
rect 22201 11101 22235 11135
rect 22294 11101 22328 11135
rect 22707 11101 22741 11135
rect 23581 11101 23615 11135
rect 23857 11101 23891 11135
rect 26065 11101 26099 11135
rect 29929 11101 29963 11135
rect 30205 11101 30239 11135
rect 32873 11101 32907 11135
rect 3985 11033 4019 11067
rect 4185 11033 4219 11067
rect 5816 11033 5850 11067
rect 12633 11033 12667 11067
rect 13461 11033 13495 11067
rect 16773 11033 16807 11067
rect 18337 11033 18371 11067
rect 21189 11033 21223 11067
rect 22477 11033 22511 11067
rect 22569 11033 22603 11067
rect 23673 11033 23707 11067
rect 24041 11033 24075 11067
rect 32606 11033 32640 11067
rect 3249 10965 3283 10999
rect 4353 10965 4387 10999
rect 6929 10965 6963 10999
rect 11713 10965 11747 10999
rect 12357 10965 12391 10999
rect 20637 10965 20671 10999
rect 27353 10965 27387 10999
rect 29745 10965 29779 10999
rect 30113 10965 30147 10999
rect 4195 10761 4229 10795
rect 7849 10761 7883 10795
rect 8769 10761 8803 10795
rect 9873 10761 9907 10795
rect 13645 10761 13679 10795
rect 19717 10761 19751 10795
rect 20453 10761 20487 10795
rect 20821 10761 20855 10795
rect 22385 10761 22419 10795
rect 25973 10761 26007 10795
rect 28733 10761 28767 10795
rect 33701 10761 33735 10795
rect 3985 10693 4019 10727
rect 6745 10693 6779 10727
rect 7021 10693 7055 10727
rect 7481 10693 7515 10727
rect 9137 10693 9171 10727
rect 9505 10693 9539 10727
rect 12541 10693 12575 10727
rect 12909 10693 12943 10727
rect 13277 10693 13311 10727
rect 18245 10693 18279 10727
rect 22753 10693 22787 10727
rect 24860 10693 24894 10727
rect 29377 10693 29411 10727
rect 29561 10693 29595 10727
rect 2513 10625 2547 10659
rect 3157 10625 3191 10659
rect 3341 10625 3375 10659
rect 7113 10625 7147 10659
rect 9045 10625 9079 10659
rect 12817 10625 12851 10659
rect 20637 10625 20671 10659
rect 20913 10625 20947 10659
rect 22569 10625 22603 10659
rect 22661 10625 22695 10659
rect 22937 10625 22971 10659
rect 27620 10625 27654 10659
rect 32577 10625 32611 10659
rect 2421 10557 2455 10591
rect 3249 10557 3283 10591
rect 3433 10557 3467 10591
rect 24593 10557 24627 10591
rect 27353 10557 27387 10591
rect 32321 10557 32355 10591
rect 2973 10421 3007 10455
rect 4169 10421 4203 10455
rect 4353 10421 4387 10455
rect 8033 10421 8067 10455
rect 10057 10421 10091 10455
rect 13829 10421 13863 10455
rect 29561 10421 29595 10455
rect 29745 10421 29779 10455
rect 2697 10217 2731 10251
rect 4169 10217 4203 10251
rect 6745 10217 6779 10251
rect 8585 10217 8619 10251
rect 12633 10217 12667 10251
rect 21281 10217 21315 10251
rect 24961 10217 24995 10251
rect 27353 10217 27387 10251
rect 28273 10217 28307 10251
rect 31677 10217 31711 10251
rect 2881 10081 2915 10115
rect 3249 10081 3283 10115
rect 3341 10081 3375 10115
rect 5365 10081 5399 10115
rect 11253 10081 11287 10115
rect 1777 10013 1811 10047
rect 2053 10013 2087 10047
rect 2973 10013 3007 10047
rect 4445 10013 4479 10047
rect 7205 10013 7239 10047
rect 7472 10013 7506 10047
rect 22569 10013 22603 10047
rect 25099 10013 25133 10047
rect 25329 10013 25363 10047
rect 25512 10013 25546 10047
rect 25605 10013 25639 10047
rect 26065 10013 26099 10047
rect 28413 10013 28447 10047
rect 28641 10013 28675 10047
rect 28824 10013 28858 10047
rect 28917 10013 28951 10047
rect 29929 10013 29963 10047
rect 30113 10013 30147 10047
rect 30297 10013 30331 10047
rect 33425 10013 33459 10047
rect 33701 10013 33735 10047
rect 1869 9945 1903 9979
rect 3985 9945 4019 9979
rect 4169 9945 4203 9979
rect 5632 9945 5666 9979
rect 11520 9945 11554 9979
rect 25237 9945 25271 9979
rect 28549 9945 28583 9979
rect 30021 9945 30055 9979
rect 32965 9945 32999 9979
rect 2237 9877 2271 9911
rect 3065 9877 3099 9911
rect 29745 9877 29779 9911
rect 33517 9877 33551 9911
rect 33885 9877 33919 9911
rect 1961 9673 1995 9707
rect 4169 9673 4203 9707
rect 4813 9673 4847 9707
rect 8493 9673 8527 9707
rect 27721 9673 27755 9707
rect 31401 9673 31435 9707
rect 2329 9605 2363 9639
rect 3249 9605 3283 9639
rect 7380 9605 7414 9639
rect 17233 9605 17267 9639
rect 21005 9605 21039 9639
rect 22385 9605 22419 9639
rect 27353 9605 27387 9639
rect 32321 9605 32355 9639
rect 2145 9537 2179 9571
rect 2421 9537 2455 9571
rect 3341 9537 3375 9571
rect 4077 9537 4111 9571
rect 4721 9537 4755 9571
rect 7113 9537 7147 9571
rect 11969 9537 12003 9571
rect 17049 9537 17083 9571
rect 17325 9537 17359 9571
rect 18245 9537 18279 9571
rect 18429 9537 18463 9571
rect 18521 9537 18555 9571
rect 18613 9537 18647 9571
rect 19441 9537 19475 9571
rect 19625 9537 19659 9571
rect 19717 9537 19751 9571
rect 19855 9537 19889 9571
rect 20637 9537 20671 9571
rect 20730 9537 20764 9571
rect 20913 9537 20947 9571
rect 21143 9537 21177 9571
rect 22201 9537 22235 9571
rect 22477 9537 22511 9571
rect 27169 9537 27203 9571
rect 27445 9537 27479 9571
rect 27537 9537 27571 9571
rect 31309 9537 31343 9571
rect 31585 9537 31619 9571
rect 3433 9469 3467 9503
rect 11713 9469 11747 9503
rect 13093 9401 13127 9435
rect 18797 9401 18831 9435
rect 19993 9401 20027 9435
rect 21281 9401 21315 9435
rect 2881 9333 2915 9367
rect 16865 9333 16899 9367
rect 22017 9333 22051 9367
rect 31769 9333 31803 9367
rect 33609 9333 33643 9367
rect 2973 9129 3007 9163
rect 12173 9129 12207 9163
rect 16405 9129 16439 9163
rect 21281 9129 21315 9163
rect 32321 9129 32355 9163
rect 2789 9061 2823 9095
rect 3985 8993 4019 9027
rect 10793 8993 10827 9027
rect 4169 8925 4203 8959
rect 11060 8925 11094 8959
rect 15025 8925 15059 8959
rect 15292 8925 15326 8959
rect 16865 8925 16899 8959
rect 19901 8925 19935 8959
rect 20168 8925 20202 8959
rect 22661 8925 22695 8959
rect 22845 8925 22879 8959
rect 22937 8925 22971 8959
rect 24593 8925 24627 8959
rect 24869 8925 24903 8959
rect 28733 8925 28767 8959
rect 29009 8925 29043 8959
rect 29929 8925 29963 8959
rect 30205 8925 30239 8959
rect 33701 8925 33735 8959
rect 2927 8857 2961 8891
rect 3341 8857 3375 8891
rect 17132 8857 17166 8891
rect 28825 8857 28859 8891
rect 30113 8857 30147 8891
rect 33456 8857 33490 8891
rect 4353 8789 4387 8823
rect 18245 8789 18279 8823
rect 22477 8789 22511 8823
rect 24685 8789 24719 8823
rect 25053 8789 25087 8823
rect 29193 8789 29227 8823
rect 29745 8789 29779 8823
rect 17693 8585 17727 8619
rect 21005 8585 21039 8619
rect 23673 8585 23707 8619
rect 25881 8585 25915 8619
rect 30021 8585 30055 8619
rect 30849 8585 30883 8619
rect 33701 8585 33735 8619
rect 9597 8517 9631 8551
rect 16068 8517 16102 8551
rect 20637 8517 20671 8551
rect 20729 8517 20763 8551
rect 22753 8517 22787 8551
rect 22937 8517 22971 8551
rect 24808 8517 24842 8551
rect 30481 8517 30515 8551
rect 32566 8517 32600 8551
rect 16313 8449 16347 8483
rect 17509 8449 17543 8483
rect 17785 8449 17819 8483
rect 18245 8449 18279 8483
rect 20453 8449 20487 8483
rect 20821 8449 20855 8483
rect 25513 8449 25547 8483
rect 25697 8449 25731 8483
rect 25973 8449 26007 8483
rect 28641 8449 28675 8483
rect 28908 8449 28942 8483
rect 30665 8449 30699 8483
rect 30941 8449 30975 8483
rect 32321 8449 32355 8483
rect 19993 8381 20027 8415
rect 25053 8381 25087 8415
rect 8309 8313 8343 8347
rect 14933 8313 14967 8347
rect 17325 8313 17359 8347
rect 23121 8313 23155 8347
rect 22937 8245 22971 8279
rect 18613 8041 18647 8075
rect 22937 8041 22971 8075
rect 28273 8041 28307 8075
rect 32413 8041 32447 8075
rect 7113 7837 7147 7871
rect 7297 7837 7331 7871
rect 9873 7837 9907 7871
rect 10057 7837 10091 7871
rect 18889 7837 18923 7871
rect 21649 7837 21683 7871
rect 24593 7837 24627 7871
rect 28549 7837 28583 7871
rect 29745 7837 29779 7871
rect 33701 7837 33735 7871
rect 7389 7769 7423 7803
rect 10241 7769 10275 7803
rect 16221 7769 16255 7803
rect 18429 7769 18463 7803
rect 19441 7769 19475 7803
rect 28089 7769 28123 7803
rect 17509 7701 17543 7735
rect 18613 7701 18647 7735
rect 20729 7701 20763 7735
rect 25881 7701 25915 7735
rect 28273 7701 28307 7735
rect 31033 7701 31067 7735
rect 10701 7497 10735 7531
rect 12173 7497 12207 7531
rect 15577 7497 15611 7531
rect 15761 7497 15795 7531
rect 17693 7497 17727 7531
rect 19533 7497 19567 7531
rect 20821 7497 20855 7531
rect 22385 7497 22419 7531
rect 25973 7497 26007 7531
rect 29101 7497 29135 7531
rect 6837 7429 6871 7463
rect 15945 7429 15979 7463
rect 18245 7429 18279 7463
rect 23397 7429 23431 7463
rect 25053 7429 25087 7463
rect 2513 7361 2547 7395
rect 8953 7361 8987 7395
rect 14749 7361 14783 7395
rect 17509 7361 17543 7395
rect 17785 7361 17819 7395
rect 20637 7361 20671 7395
rect 20913 7361 20947 7395
rect 22201 7361 22235 7395
rect 22477 7361 22511 7395
rect 25789 7361 25823 7395
rect 26065 7361 26099 7395
rect 30389 7361 30423 7395
rect 6561 7293 6595 7327
rect 9229 7293 9263 7327
rect 11897 7293 11931 7327
rect 12081 7293 12115 7327
rect 17325 7293 17359 7327
rect 2605 7157 2639 7191
rect 8309 7157 8343 7191
rect 12541 7157 12575 7191
rect 13461 7157 13495 7191
rect 15761 7157 15795 7191
rect 20453 7157 20487 7191
rect 22017 7157 22051 7191
rect 25605 7157 25639 7191
rect 1685 6953 1719 6987
rect 3169 6953 3203 6987
rect 13093 6953 13127 6987
rect 20821 6953 20855 6987
rect 5457 6817 5491 6851
rect 7941 6817 7975 6851
rect 10149 6817 10183 6851
rect 10701 6817 10735 6851
rect 15577 6817 15611 6851
rect 21281 6817 21315 6851
rect 3433 6749 3467 6783
rect 5724 6749 5758 6783
rect 7665 6749 7699 6783
rect 10241 6749 10275 6783
rect 10563 6749 10597 6783
rect 11713 6749 11747 6783
rect 13553 6749 13587 6783
rect 13737 6749 13771 6783
rect 15844 6749 15878 6783
rect 17417 6749 17451 6783
rect 17601 6749 17635 6783
rect 17877 6749 17911 6783
rect 19441 6749 19475 6783
rect 19708 6749 19742 6783
rect 21548 6749 21582 6783
rect 23765 6749 23799 6783
rect 24041 6749 24075 6783
rect 24593 6749 24627 6783
rect 28926 6749 28960 6783
rect 29193 6749 29227 6783
rect 30113 6749 30147 6783
rect 7757 6681 7791 6715
rect 11958 6681 11992 6715
rect 17785 6681 17819 6715
rect 23949 6681 23983 6715
rect 24860 6681 24894 6715
rect 30358 6681 30392 6715
rect 6837 6613 6871 6647
rect 7297 6613 7331 6647
rect 10977 6613 11011 6647
rect 13645 6613 13679 6647
rect 16957 6613 16991 6647
rect 22661 6613 22695 6647
rect 23581 6613 23615 6647
rect 25973 6613 26007 6647
rect 27813 6613 27847 6647
rect 31493 6613 31527 6647
rect 6929 6409 6963 6443
rect 13001 6409 13035 6443
rect 20913 6409 20947 6443
rect 2789 6341 2823 6375
rect 3709 6341 3743 6375
rect 6837 6341 6871 6375
rect 12909 6341 12943 6375
rect 19800 6341 19834 6375
rect 24694 6341 24728 6375
rect 29570 6341 29604 6375
rect 2973 6273 3007 6307
rect 3157 6273 3191 6307
rect 6653 6205 6687 6239
rect 12725 6205 12759 6239
rect 19533 6205 19567 6239
rect 24961 6205 24995 6239
rect 29837 6205 29871 6239
rect 7297 6137 7331 6171
rect 23581 6137 23615 6171
rect 28457 6137 28491 6171
rect 3801 6069 3835 6103
rect 13369 6069 13403 6103
rect 25973 5865 26007 5899
rect 29193 5865 29227 5899
rect 3985 5729 4019 5763
rect 4353 5729 4387 5763
rect 5733 5729 5767 5763
rect 12909 5729 12943 5763
rect 12633 5661 12667 5695
rect 12725 5661 12759 5695
rect 24593 5661 24627 5695
rect 24860 5661 24894 5695
rect 28733 5661 28767 5695
rect 29009 5661 29043 5695
rect 28825 5593 28859 5627
rect 12909 5525 12943 5559
rect 5641 5321 5675 5355
rect 9505 5321 9539 5355
rect 10425 5321 10459 5355
rect 13093 5321 13127 5355
rect 19533 5321 19567 5355
rect 24685 5321 24719 5355
rect 4353 5253 4387 5287
rect 18245 5253 18279 5287
rect 23397 5253 23431 5287
rect 25789 5253 25823 5287
rect 4077 5185 4111 5219
rect 4261 5185 4295 5219
rect 5733 5185 5767 5219
rect 10333 5185 10367 5219
rect 10517 5185 10551 5219
rect 11969 5185 12003 5219
rect 15209 5185 15243 5219
rect 25973 5185 26007 5219
rect 9229 5117 9263 5151
rect 9413 5117 9447 5151
rect 11713 5117 11747 5151
rect 9873 5049 9907 5083
rect 15117 4981 15151 5015
rect 25605 4981 25639 5015
rect 10885 4777 10919 4811
rect 11989 4777 12023 4811
rect 14565 4709 14599 4743
rect 24961 4709 24995 4743
rect 7205 4641 7239 4675
rect 9137 4641 9171 4675
rect 16221 4641 16255 4675
rect 18705 4641 18739 4675
rect 20453 4641 20487 4675
rect 24593 4641 24627 4675
rect 7472 4573 7506 4607
rect 11897 4573 11931 4607
rect 12265 4573 12299 4607
rect 14289 4573 14323 4607
rect 14565 4573 14599 4607
rect 15945 4573 15979 4607
rect 17417 4573 17451 4607
rect 18429 4573 18463 4607
rect 20177 4573 20211 4607
rect 21649 4573 21683 4607
rect 22293 4573 22327 4607
rect 25881 4573 25915 4607
rect 9413 4505 9447 4539
rect 26148 4505 26182 4539
rect 8585 4437 8619 4471
rect 12449 4437 12483 4471
rect 14381 4437 14415 4471
rect 15577 4437 15611 4471
rect 16037 4437 16071 4471
rect 17509 4437 17543 4471
rect 18061 4437 18095 4471
rect 18521 4437 18555 4471
rect 19809 4437 19843 4471
rect 20269 4437 20303 4471
rect 21557 4437 21591 4471
rect 22201 4437 22235 4471
rect 25053 4437 25087 4471
rect 27261 4437 27295 4471
rect 9689 4233 9723 4267
rect 13369 4233 13403 4267
rect 26157 4233 26191 4267
rect 7297 4165 7331 4199
rect 9597 4165 9631 4199
rect 15200 4165 15234 4199
rect 25452 4165 25486 4199
rect 10425 4097 10459 4131
rect 10517 4097 10551 4131
rect 10793 4097 10827 4131
rect 13461 4097 13495 4131
rect 14933 4097 14967 4131
rect 17049 4097 17083 4131
rect 17693 4097 17727 4131
rect 17960 4097 17994 4131
rect 21198 4097 21232 4131
rect 21465 4097 21499 4131
rect 22017 4097 22051 4131
rect 22284 4097 22318 4131
rect 25697 4097 25731 4131
rect 28282 4097 28316 4131
rect 28549 4097 28583 4131
rect 7021 4029 7055 4063
rect 8769 4029 8803 4063
rect 9873 4029 9907 4063
rect 13645 4029 13679 4063
rect 26617 4029 26651 4063
rect 9229 3961 9263 3995
rect 26249 3961 26283 3995
rect 13001 3893 13035 3927
rect 16313 3893 16347 3927
rect 16957 3893 16991 3927
rect 19073 3893 19107 3927
rect 20085 3893 20119 3927
rect 23397 3893 23431 3927
rect 24317 3893 24351 3927
rect 27169 3893 27203 3927
rect 7941 3689 7975 3723
rect 13737 3689 13771 3723
rect 20913 3689 20947 3723
rect 22109 3689 22143 3723
rect 26801 3689 26835 3723
rect 27813 3689 27847 3723
rect 26433 3621 26467 3655
rect 26893 3621 26927 3655
rect 27905 3621 27939 3655
rect 16681 3553 16715 3587
rect 22753 3553 22787 3587
rect 26985 3553 27019 3587
rect 7941 3485 7975 3519
rect 8125 3485 8159 3519
rect 12357 3485 12391 3519
rect 12624 3485 12658 3519
rect 15669 3485 15703 3519
rect 19533 3485 19567 3519
rect 19800 3485 19834 3519
rect 22477 3485 22511 3519
rect 24593 3485 24627 3519
rect 15402 3417 15436 3451
rect 16948 3417 16982 3451
rect 22569 3417 22603 3451
rect 24860 3417 24894 3451
rect 27353 3417 27387 3451
rect 28273 3417 28307 3451
rect 14289 3349 14323 3383
rect 18061 3349 18095 3383
rect 25973 3349 26007 3383
rect 12541 3145 12575 3179
rect 14381 3145 14415 3179
rect 14749 3145 14783 3179
rect 15301 3145 15335 3179
rect 16957 3145 16991 3179
rect 17325 3145 17359 3179
rect 17417 3145 17451 3179
rect 19717 3145 19751 3179
rect 21097 3145 21131 3179
rect 29101 3145 29135 3179
rect 30389 3077 30423 3111
rect 12633 3009 12667 3043
rect 15209 3009 15243 3043
rect 19809 3009 19843 3043
rect 20913 3009 20947 3043
rect 21189 3009 21223 3043
rect 25145 3009 25179 3043
rect 26065 3009 26099 3043
rect 14197 2941 14231 2975
rect 14289 2941 14323 2975
rect 17601 2941 17635 2975
rect 25513 2941 25547 2975
rect 20729 2873 20763 2907
rect 25605 2873 25639 2907
rect 25697 2873 25731 2907
rect 2053 2397 2087 2431
rect 3065 2397 3099 2431
rect 4445 2397 4479 2431
rect 5641 2397 5675 2431
rect 6561 2397 6595 2431
rect 7757 2397 7791 2431
rect 9137 2397 9171 2431
rect 10333 2397 10367 2431
rect 11713 2397 11747 2431
rect 12909 2397 12943 2431
rect 14289 2397 14323 2431
rect 15485 2397 15519 2431
rect 16865 2397 16899 2431
rect 18061 2397 18095 2431
rect 19441 2397 19475 2431
rect 20637 2397 20671 2431
rect 22017 2397 22051 2431
rect 23213 2397 23247 2431
rect 25053 2397 25087 2431
rect 26249 2397 26283 2431
rect 27629 2397 27663 2431
rect 28365 2397 28399 2431
rect 29745 2397 29779 2431
rect 30941 2397 30975 2431
rect 32321 2397 32355 2431
rect 33517 2397 33551 2431
rect 1777 2329 1811 2363
rect 2789 2329 2823 2363
rect 4169 2329 4203 2363
rect 5365 2329 5399 2363
rect 14565 2329 14599 2363
rect 15761 2329 15795 2363
rect 17141 2329 17175 2363
rect 18337 2329 18371 2363
rect 19717 2329 19751 2363
rect 20913 2329 20947 2363
rect 22293 2329 22327 2363
rect 23489 2329 23523 2363
rect 24777 2329 24811 2363
rect 25973 2329 26007 2363
rect 27353 2329 27387 2363
rect 28641 2329 28675 2363
rect 34345 2261 34379 2295
<< metal1 >>
rect 1104 33754 35027 33776
rect 1104 33702 9390 33754
rect 9442 33702 9454 33754
rect 9506 33702 9518 33754
rect 9570 33702 9582 33754
rect 9634 33702 9646 33754
rect 9698 33702 17831 33754
rect 17883 33702 17895 33754
rect 17947 33702 17959 33754
rect 18011 33702 18023 33754
rect 18075 33702 18087 33754
rect 18139 33702 26272 33754
rect 26324 33702 26336 33754
rect 26388 33702 26400 33754
rect 26452 33702 26464 33754
rect 26516 33702 26528 33754
rect 26580 33702 34713 33754
rect 34765 33702 34777 33754
rect 34829 33702 34841 33754
rect 34893 33702 34905 33754
rect 34957 33702 34969 33754
rect 35021 33702 35027 33754
rect 1104 33680 35027 33702
rect 4890 33572 4896 33584
rect 4851 33544 4896 33572
rect 4890 33532 4896 33544
rect 4948 33532 4954 33584
rect 7834 33572 7840 33584
rect 7795 33544 7840 33572
rect 7834 33532 7840 33544
rect 7892 33532 7898 33584
rect 10594 33532 10600 33584
rect 10652 33572 10658 33584
rect 10781 33575 10839 33581
rect 10781 33572 10793 33575
rect 10652 33544 10793 33572
rect 10652 33532 10658 33544
rect 10781 33541 10793 33544
rect 10827 33541 10839 33575
rect 10781 33535 10839 33541
rect 13814 33532 13820 33584
rect 13872 33572 13878 33584
rect 14461 33575 14519 33581
rect 14461 33572 14473 33575
rect 13872 33544 14473 33572
rect 13872 33532 13878 33544
rect 14461 33541 14473 33544
rect 14507 33541 14519 33575
rect 14461 33535 14519 33541
rect 16574 33532 16580 33584
rect 16632 33572 16638 33584
rect 17037 33575 17095 33581
rect 17037 33572 17049 33575
rect 16632 33544 17049 33572
rect 16632 33532 16638 33544
rect 17037 33541 17049 33544
rect 17083 33541 17095 33575
rect 17037 33535 17095 33541
rect 19426 33532 19432 33584
rect 19484 33572 19490 33584
rect 19705 33575 19763 33581
rect 19705 33572 19717 33575
rect 19484 33544 19717 33572
rect 19484 33532 19490 33544
rect 19705 33541 19717 33544
rect 19751 33541 19763 33575
rect 22646 33572 22652 33584
rect 22607 33544 22652 33572
rect 19705 33535 19763 33541
rect 22646 33532 22652 33544
rect 22704 33532 22710 33584
rect 25590 33572 25596 33584
rect 25551 33544 25596 33572
rect 25590 33532 25596 33544
rect 25648 33532 25654 33584
rect 28258 33532 28264 33584
rect 28316 33572 28322 33584
rect 28537 33575 28595 33581
rect 28537 33572 28549 33575
rect 28316 33544 28549 33572
rect 28316 33532 28322 33544
rect 28537 33541 28549 33544
rect 28583 33541 28595 33575
rect 31478 33572 31484 33584
rect 31439 33544 31484 33572
rect 28537 33535 28595 33541
rect 31478 33532 31484 33544
rect 31536 33532 31542 33584
rect 34238 33572 34244 33584
rect 34199 33544 34244 33572
rect 34238 33532 34244 33544
rect 34296 33532 34302 33584
rect 8018 33368 8024 33380
rect 7979 33340 8024 33368
rect 8018 33328 8024 33340
rect 8076 33328 8082 33380
rect 10965 33371 11023 33377
rect 10965 33337 10977 33371
rect 11011 33368 11023 33371
rect 12250 33368 12256 33380
rect 11011 33340 12256 33368
rect 11011 33337 11023 33340
rect 10965 33331 11023 33337
rect 12250 33328 12256 33340
rect 12308 33328 12314 33380
rect 14274 33368 14280 33380
rect 14235 33340 14280 33368
rect 14274 33328 14280 33340
rect 14332 33328 14338 33380
rect 16850 33368 16856 33380
rect 16811 33340 16856 33368
rect 16850 33328 16856 33340
rect 16908 33328 16914 33380
rect 19518 33368 19524 33380
rect 19479 33340 19524 33368
rect 19518 33328 19524 33340
rect 19576 33328 19582 33380
rect 22462 33368 22468 33380
rect 22423 33340 22468 33368
rect 22462 33328 22468 33340
rect 22520 33328 22526 33380
rect 25406 33368 25412 33380
rect 25367 33340 25412 33368
rect 25406 33328 25412 33340
rect 25464 33328 25470 33380
rect 28350 33368 28356 33380
rect 28311 33340 28356 33368
rect 28350 33328 28356 33340
rect 28408 33328 28414 33380
rect 31294 33368 31300 33380
rect 31255 33340 31300 33368
rect 31294 33328 31300 33340
rect 31352 33328 31358 33380
rect 33410 33328 33416 33380
rect 33468 33368 33474 33380
rect 34057 33371 34115 33377
rect 34057 33368 34069 33371
rect 33468 33340 34069 33368
rect 33468 33328 33474 33340
rect 34057 33337 34069 33340
rect 34103 33337 34115 33371
rect 34057 33331 34115 33337
rect 4982 33300 4988 33312
rect 4943 33272 4988 33300
rect 4982 33260 4988 33272
rect 5040 33260 5046 33312
rect 1104 33210 34868 33232
rect 1104 33158 5170 33210
rect 5222 33158 5234 33210
rect 5286 33158 5298 33210
rect 5350 33158 5362 33210
rect 5414 33158 5426 33210
rect 5478 33158 13611 33210
rect 13663 33158 13675 33210
rect 13727 33158 13739 33210
rect 13791 33158 13803 33210
rect 13855 33158 13867 33210
rect 13919 33158 22052 33210
rect 22104 33158 22116 33210
rect 22168 33158 22180 33210
rect 22232 33158 22244 33210
rect 22296 33158 22308 33210
rect 22360 33158 30493 33210
rect 30545 33158 30557 33210
rect 30609 33158 30621 33210
rect 30673 33158 30685 33210
rect 30737 33158 30749 33210
rect 30801 33158 34868 33210
rect 1104 33136 34868 33158
rect 24578 33028 24584 33040
rect 20732 33000 24584 33028
rect 16850 32960 16856 32972
rect 16500 32932 16856 32960
rect 10229 32895 10287 32901
rect 10229 32861 10241 32895
rect 10275 32892 10287 32895
rect 10502 32892 10508 32904
rect 10275 32864 10508 32892
rect 10275 32861 10287 32864
rect 10229 32855 10287 32861
rect 10502 32852 10508 32864
rect 10560 32852 10566 32904
rect 16500 32901 16528 32932
rect 16850 32920 16856 32932
rect 16908 32920 16914 32972
rect 20622 32960 20628 32972
rect 20583 32932 20628 32960
rect 20622 32920 20628 32932
rect 20680 32920 20686 32972
rect 16301 32895 16359 32901
rect 16301 32861 16313 32895
rect 16347 32861 16359 32895
rect 16301 32855 16359 32861
rect 16485 32895 16543 32901
rect 16485 32861 16497 32895
rect 16531 32861 16543 32895
rect 16485 32855 16543 32861
rect 16577 32895 16635 32901
rect 16577 32861 16589 32895
rect 16623 32892 16635 32895
rect 16623 32864 20484 32892
rect 16623 32861 16635 32864
rect 16577 32855 16635 32861
rect 15841 32827 15899 32833
rect 15841 32793 15853 32827
rect 15887 32824 15899 32827
rect 16206 32824 16212 32836
rect 15887 32796 16212 32824
rect 15887 32793 15899 32796
rect 15841 32787 15899 32793
rect 16206 32784 16212 32796
rect 16264 32784 16270 32836
rect 16316 32824 16344 32855
rect 16758 32824 16764 32836
rect 16316 32796 16764 32824
rect 16758 32784 16764 32796
rect 16816 32784 16822 32836
rect 20456 32824 20484 32864
rect 20530 32852 20536 32904
rect 20588 32892 20594 32904
rect 20732 32892 20760 33000
rect 24578 32988 24584 33000
rect 24636 32988 24642 33040
rect 20806 32920 20812 32972
rect 20864 32960 20870 32972
rect 25406 32960 25412 32972
rect 20864 32932 25412 32960
rect 20864 32920 20870 32932
rect 25406 32920 25412 32932
rect 25464 32920 25470 32972
rect 20588 32864 20760 32892
rect 22465 32895 22523 32901
rect 20588 32852 20594 32864
rect 22465 32861 22477 32895
rect 22511 32892 22523 32895
rect 22922 32892 22928 32904
rect 22511 32864 22928 32892
rect 22511 32861 22523 32864
rect 22465 32855 22523 32861
rect 22922 32852 22928 32864
rect 22980 32852 22986 32904
rect 28350 32824 28356 32836
rect 20456 32796 28356 32824
rect 28350 32784 28356 32796
rect 28408 32784 28414 32836
rect 10134 32756 10140 32768
rect 10095 32728 10140 32756
rect 10134 32716 10140 32728
rect 10192 32716 10198 32768
rect 13262 32716 13268 32768
rect 13320 32756 13326 32768
rect 20806 32756 20812 32768
rect 13320 32728 20812 32756
rect 13320 32716 13326 32728
rect 20806 32716 20812 32728
rect 20864 32716 20870 32768
rect 20901 32759 20959 32765
rect 20901 32725 20913 32759
rect 20947 32756 20959 32759
rect 21266 32756 21272 32768
rect 20947 32728 21272 32756
rect 20947 32725 20959 32728
rect 20901 32719 20959 32725
rect 21266 32716 21272 32728
rect 21324 32716 21330 32768
rect 22002 32716 22008 32768
rect 22060 32756 22066 32768
rect 22373 32759 22431 32765
rect 22373 32756 22385 32759
rect 22060 32728 22385 32756
rect 22060 32716 22066 32728
rect 22373 32725 22385 32728
rect 22419 32725 22431 32759
rect 22373 32719 22431 32725
rect 1104 32666 35027 32688
rect 1104 32614 9390 32666
rect 9442 32614 9454 32666
rect 9506 32614 9518 32666
rect 9570 32614 9582 32666
rect 9634 32614 9646 32666
rect 9698 32614 17831 32666
rect 17883 32614 17895 32666
rect 17947 32614 17959 32666
rect 18011 32614 18023 32666
rect 18075 32614 18087 32666
rect 18139 32614 26272 32666
rect 26324 32614 26336 32666
rect 26388 32614 26400 32666
rect 26452 32614 26464 32666
rect 26516 32614 26528 32666
rect 26580 32614 34713 32666
rect 34765 32614 34777 32666
rect 34829 32614 34841 32666
rect 34893 32614 34905 32666
rect 34957 32614 34969 32666
rect 35021 32614 35027 32666
rect 1104 32592 35027 32614
rect 12250 32552 12256 32564
rect 12211 32524 12256 32552
rect 12250 32512 12256 32524
rect 12308 32512 12314 32564
rect 13449 32555 13507 32561
rect 13449 32521 13461 32555
rect 13495 32552 13507 32555
rect 14274 32552 14280 32564
rect 13495 32524 14280 32552
rect 13495 32521 13507 32524
rect 13449 32515 13507 32521
rect 14274 32512 14280 32524
rect 14332 32512 14338 32564
rect 17313 32555 17371 32561
rect 17313 32521 17325 32555
rect 17359 32552 17371 32555
rect 18049 32555 18107 32561
rect 18049 32552 18061 32555
rect 17359 32524 18061 32552
rect 17359 32521 17371 32524
rect 17313 32515 17371 32521
rect 18049 32521 18061 32524
rect 18095 32521 18107 32555
rect 22462 32552 22468 32564
rect 18049 32515 18107 32521
rect 18156 32524 22468 32552
rect 10686 32484 10692 32496
rect 10428 32456 10692 32484
rect 10428 32425 10456 32456
rect 10686 32444 10692 32456
rect 10744 32444 10750 32496
rect 13262 32484 13268 32496
rect 13223 32456 13268 32484
rect 13262 32444 13268 32456
rect 13320 32444 13326 32496
rect 18156 32484 18184 32524
rect 22462 32512 22468 32524
rect 22520 32512 22526 32564
rect 16546 32456 18184 32484
rect 21177 32487 21235 32493
rect 9861 32419 9919 32425
rect 9861 32385 9873 32419
rect 9907 32416 9919 32419
rect 10413 32419 10471 32425
rect 10413 32416 10425 32419
rect 9907 32388 10425 32416
rect 9907 32385 9919 32388
rect 9861 32379 9919 32385
rect 10413 32385 10425 32388
rect 10459 32385 10471 32419
rect 10413 32379 10471 32385
rect 10502 32376 10508 32428
rect 10560 32416 10566 32428
rect 12069 32419 12127 32425
rect 10560 32388 10605 32416
rect 10560 32376 10566 32388
rect 12069 32385 12081 32419
rect 12115 32416 12127 32419
rect 16546 32416 16574 32456
rect 21177 32453 21189 32487
rect 21223 32484 21235 32487
rect 22097 32487 22155 32493
rect 22097 32484 22109 32487
rect 21223 32456 22109 32484
rect 21223 32453 21235 32456
rect 21177 32447 21235 32453
rect 22097 32453 22109 32456
rect 22143 32453 22155 32487
rect 22097 32447 22155 32453
rect 12115 32388 16574 32416
rect 17221 32419 17279 32425
rect 12115 32385 12127 32388
rect 12069 32379 12127 32385
rect 17221 32385 17233 32419
rect 17267 32416 17279 32419
rect 17862 32416 17868 32428
rect 17267 32388 17868 32416
rect 17267 32385 17279 32388
rect 17221 32379 17279 32385
rect 17862 32376 17868 32388
rect 17920 32416 17926 32428
rect 18049 32419 18107 32425
rect 18049 32416 18061 32419
rect 17920 32388 18061 32416
rect 17920 32376 17926 32388
rect 18049 32385 18061 32388
rect 18095 32385 18107 32419
rect 18049 32379 18107 32385
rect 18230 32376 18236 32428
rect 18288 32416 18294 32428
rect 21085 32419 21143 32425
rect 18288 32388 20760 32416
rect 18288 32376 18294 32388
rect 10689 32351 10747 32357
rect 10689 32317 10701 32351
rect 10735 32317 10747 32351
rect 12342 32348 12348 32360
rect 12255 32320 12348 32348
rect 10689 32311 10747 32317
rect 8570 32240 8576 32292
rect 8628 32280 8634 32292
rect 10704 32280 10732 32311
rect 12342 32308 12348 32320
rect 12400 32348 12406 32360
rect 13541 32351 13599 32357
rect 13541 32348 13553 32351
rect 12400 32320 13553 32348
rect 12400 32308 12406 32320
rect 13541 32317 13553 32320
rect 13587 32317 13599 32351
rect 13541 32311 13599 32317
rect 13446 32280 13452 32292
rect 8628 32252 13452 32280
rect 8628 32240 8634 32252
rect 13446 32240 13452 32252
rect 13504 32240 13510 32292
rect 9861 32215 9919 32221
rect 9861 32181 9873 32215
rect 9907 32212 9919 32215
rect 10042 32212 10048 32224
rect 9907 32184 10048 32212
rect 9907 32181 9919 32184
rect 9861 32175 9919 32181
rect 10042 32172 10048 32184
rect 10100 32172 10106 32224
rect 10594 32172 10600 32224
rect 10652 32212 10658 32224
rect 11793 32215 11851 32221
rect 10652 32184 10697 32212
rect 10652 32172 10658 32184
rect 11793 32181 11805 32215
rect 11839 32212 11851 32215
rect 11974 32212 11980 32224
rect 11839 32184 11980 32212
rect 11839 32181 11851 32184
rect 11793 32175 11851 32181
rect 11974 32172 11980 32184
rect 12032 32172 12038 32224
rect 12989 32215 13047 32221
rect 12989 32181 13001 32215
rect 13035 32212 13047 32215
rect 13170 32212 13176 32224
rect 13035 32184 13176 32212
rect 13035 32181 13047 32184
rect 12989 32175 13047 32181
rect 13170 32172 13176 32184
rect 13228 32172 13234 32224
rect 13556 32212 13584 32311
rect 13998 32308 14004 32360
rect 14056 32348 14062 32360
rect 17402 32348 17408 32360
rect 14056 32320 17264 32348
rect 17363 32320 17408 32348
rect 14056 32308 14062 32320
rect 13630 32240 13636 32292
rect 13688 32280 13694 32292
rect 16853 32283 16911 32289
rect 16853 32280 16865 32283
rect 13688 32252 16865 32280
rect 13688 32240 13694 32252
rect 16853 32249 16865 32252
rect 16899 32249 16911 32283
rect 17236 32280 17264 32320
rect 17402 32308 17408 32320
rect 17460 32308 17466 32360
rect 19518 32280 19524 32292
rect 17236 32252 19524 32280
rect 16853 32243 16911 32249
rect 19518 32240 19524 32252
rect 19576 32240 19582 32292
rect 20732 32289 20760 32388
rect 21085 32385 21097 32419
rect 21131 32416 21143 32419
rect 22002 32416 22008 32428
rect 21131 32388 22008 32416
rect 21131 32385 21143 32388
rect 21085 32379 21143 32385
rect 22002 32376 22008 32388
rect 22060 32376 22066 32428
rect 22189 32419 22247 32425
rect 22189 32385 22201 32419
rect 22235 32416 22247 32419
rect 22554 32416 22560 32428
rect 22235 32388 22560 32416
rect 22235 32385 22247 32388
rect 22189 32379 22247 32385
rect 22554 32376 22560 32388
rect 22612 32376 22618 32428
rect 23109 32419 23167 32425
rect 23109 32385 23121 32419
rect 23155 32385 23167 32419
rect 23290 32416 23296 32428
rect 23251 32388 23296 32416
rect 23109 32379 23167 32385
rect 21266 32348 21272 32360
rect 21227 32320 21272 32348
rect 21266 32308 21272 32320
rect 21324 32308 21330 32360
rect 23124 32348 23152 32379
rect 23290 32376 23296 32388
rect 23348 32376 23354 32428
rect 24489 32419 24547 32425
rect 24489 32385 24501 32419
rect 24535 32385 24547 32419
rect 24489 32379 24547 32385
rect 23382 32348 23388 32360
rect 23124 32320 23388 32348
rect 23382 32308 23388 32320
rect 23440 32308 23446 32360
rect 24504 32348 24532 32379
rect 24578 32376 24584 32428
rect 24636 32416 24642 32428
rect 24673 32419 24731 32425
rect 24673 32416 24685 32419
rect 24636 32388 24685 32416
rect 24636 32376 24642 32388
rect 24673 32385 24685 32388
rect 24719 32385 24731 32419
rect 27706 32416 27712 32428
rect 27667 32388 27712 32416
rect 24673 32379 24731 32385
rect 27706 32376 27712 32388
rect 27764 32376 27770 32428
rect 28626 32416 28632 32428
rect 28587 32388 28632 32416
rect 28626 32376 28632 32388
rect 28684 32376 28690 32428
rect 30469 32419 30527 32425
rect 30469 32385 30481 32419
rect 30515 32416 30527 32419
rect 31294 32416 31300 32428
rect 30515 32388 31300 32416
rect 30515 32385 30527 32388
rect 30469 32379 30527 32385
rect 31294 32376 31300 32388
rect 31352 32376 31358 32428
rect 33410 32416 33416 32428
rect 33371 32388 33416 32416
rect 33410 32376 33416 32388
rect 33468 32376 33474 32428
rect 24762 32348 24768 32360
rect 24504 32320 24768 32348
rect 24762 32308 24768 32320
rect 24820 32308 24826 32360
rect 20717 32283 20775 32289
rect 20717 32249 20729 32283
rect 20763 32249 20775 32283
rect 20717 32243 20775 32249
rect 21174 32240 21180 32292
rect 21232 32280 21238 32292
rect 23017 32283 23075 32289
rect 23017 32280 23029 32283
rect 21232 32252 23029 32280
rect 21232 32240 21238 32252
rect 23017 32249 23029 32252
rect 23063 32249 23075 32283
rect 27157 32283 27215 32289
rect 27157 32280 27169 32283
rect 23017 32243 23075 32249
rect 23124 32252 27169 32280
rect 16758 32212 16764 32224
rect 13556 32184 16764 32212
rect 16758 32172 16764 32184
rect 16816 32172 16822 32224
rect 18506 32172 18512 32224
rect 18564 32212 18570 32224
rect 22738 32212 22744 32224
rect 18564 32184 22744 32212
rect 18564 32172 18570 32184
rect 22738 32172 22744 32184
rect 22796 32172 22802 32224
rect 22922 32172 22928 32224
rect 22980 32212 22986 32224
rect 23124 32212 23152 32252
rect 27157 32249 27169 32252
rect 27203 32249 27215 32283
rect 27157 32243 27215 32249
rect 22980 32184 23152 32212
rect 24581 32215 24639 32221
rect 22980 32172 22986 32184
rect 24581 32181 24593 32215
rect 24627 32212 24639 32215
rect 25038 32212 25044 32224
rect 24627 32184 25044 32212
rect 24627 32181 24639 32184
rect 24581 32175 24639 32181
rect 25038 32172 25044 32184
rect 25096 32172 25102 32224
rect 30190 32172 30196 32224
rect 30248 32212 30254 32224
rect 30285 32215 30343 32221
rect 30285 32212 30297 32215
rect 30248 32184 30297 32212
rect 30248 32172 30254 32184
rect 30285 32181 30297 32184
rect 30331 32181 30343 32215
rect 33226 32212 33232 32224
rect 33187 32184 33232 32212
rect 30285 32175 30343 32181
rect 33226 32172 33232 32184
rect 33284 32172 33290 32224
rect 1104 32122 34868 32144
rect 1104 32070 5170 32122
rect 5222 32070 5234 32122
rect 5286 32070 5298 32122
rect 5350 32070 5362 32122
rect 5414 32070 5426 32122
rect 5478 32070 13611 32122
rect 13663 32070 13675 32122
rect 13727 32070 13739 32122
rect 13791 32070 13803 32122
rect 13855 32070 13867 32122
rect 13919 32070 22052 32122
rect 22104 32070 22116 32122
rect 22168 32070 22180 32122
rect 22232 32070 22244 32122
rect 22296 32070 22308 32122
rect 22360 32070 30493 32122
rect 30545 32070 30557 32122
rect 30609 32070 30621 32122
rect 30673 32070 30685 32122
rect 30737 32070 30749 32122
rect 30801 32070 34868 32122
rect 1104 32048 34868 32070
rect 8496 31980 9812 32008
rect 8496 31881 8524 31980
rect 8570 31900 8576 31952
rect 8628 31900 8634 31952
rect 8754 31900 8760 31952
rect 8812 31940 8818 31952
rect 9309 31943 9367 31949
rect 9309 31940 9321 31943
rect 8812 31912 9321 31940
rect 8812 31900 8818 31912
rect 9309 31909 9321 31912
rect 9355 31909 9367 31943
rect 9309 31903 9367 31909
rect 8481 31875 8539 31881
rect 8481 31841 8493 31875
rect 8527 31841 8539 31875
rect 8481 31835 8539 31841
rect 8588 31813 8616 31900
rect 9784 31881 9812 31980
rect 10502 31968 10508 32020
rect 10560 32008 10566 32020
rect 15749 32011 15807 32017
rect 10560 31980 12664 32008
rect 10560 31968 10566 31980
rect 11149 31943 11207 31949
rect 11149 31909 11161 31943
rect 11195 31940 11207 31943
rect 11698 31940 11704 31952
rect 11195 31912 11704 31940
rect 11195 31909 11207 31912
rect 11149 31903 11207 31909
rect 11698 31900 11704 31912
rect 11756 31900 11762 31952
rect 12360 31912 12572 31940
rect 9769 31875 9827 31881
rect 9769 31841 9781 31875
rect 9815 31841 9827 31875
rect 9769 31835 9827 31841
rect 9858 31832 9864 31884
rect 9916 31872 9922 31884
rect 11609 31875 11667 31881
rect 9916 31844 9961 31872
rect 9916 31832 9922 31844
rect 11609 31841 11621 31875
rect 11655 31872 11667 31875
rect 12360 31872 12388 31912
rect 11655 31844 12388 31872
rect 11655 31841 11667 31844
rect 11609 31835 11667 31841
rect 8389 31807 8447 31813
rect 8389 31773 8401 31807
rect 8435 31804 8447 31807
rect 8573 31807 8631 31813
rect 8435 31776 8524 31804
rect 8435 31773 8447 31776
rect 8389 31767 8447 31773
rect 8496 31736 8524 31776
rect 8573 31773 8585 31807
rect 8619 31773 8631 31807
rect 9677 31807 9735 31813
rect 9677 31804 9689 31807
rect 8573 31767 8631 31773
rect 8772 31776 9689 31804
rect 8772 31736 8800 31776
rect 9677 31773 9689 31776
rect 9723 31804 9735 31807
rect 10134 31804 10140 31816
rect 9723 31776 10140 31804
rect 9723 31773 9735 31776
rect 9677 31767 9735 31773
rect 10134 31764 10140 31776
rect 10192 31764 10198 31816
rect 11701 31807 11759 31813
rect 11701 31773 11713 31807
rect 11747 31804 11759 31807
rect 12342 31804 12348 31816
rect 11747 31776 12348 31804
rect 11747 31773 11759 31776
rect 11701 31767 11759 31773
rect 12342 31764 12348 31776
rect 12400 31764 12406 31816
rect 12544 31804 12572 31912
rect 12636 31872 12664 31980
rect 15749 31977 15761 32011
rect 15795 32008 15807 32011
rect 16114 32008 16120 32020
rect 15795 31980 16120 32008
rect 15795 31977 15807 31980
rect 15749 31971 15807 31977
rect 16114 31968 16120 31980
rect 16172 31968 16178 32020
rect 18049 32011 18107 32017
rect 18049 31977 18061 32011
rect 18095 32008 18107 32011
rect 18230 32008 18236 32020
rect 18095 31980 18236 32008
rect 18095 31977 18107 31980
rect 18049 31971 18107 31977
rect 18230 31968 18236 31980
rect 18288 31968 18294 32020
rect 20622 31968 20628 32020
rect 20680 32008 20686 32020
rect 21269 32011 21327 32017
rect 21269 32008 21281 32011
rect 20680 31980 21281 32008
rect 20680 31968 20686 31980
rect 21269 31977 21281 31980
rect 21315 31977 21327 32011
rect 21269 31971 21327 31977
rect 23290 31968 23296 32020
rect 23348 32008 23354 32020
rect 23753 32011 23811 32017
rect 23753 32008 23765 32011
rect 23348 31980 23765 32008
rect 23348 31968 23354 31980
rect 23753 31977 23765 31980
rect 23799 31977 23811 32011
rect 23753 31971 23811 31977
rect 13998 31940 14004 31952
rect 12820 31912 14004 31940
rect 12713 31875 12771 31881
rect 12713 31872 12725 31875
rect 12636 31844 12725 31872
rect 12713 31841 12725 31844
rect 12759 31841 12771 31875
rect 12713 31835 12771 31841
rect 12820 31804 12848 31912
rect 13998 31900 14004 31912
rect 14056 31900 14062 31952
rect 15933 31943 15991 31949
rect 15933 31909 15945 31943
rect 15979 31940 15991 31943
rect 16666 31940 16672 31952
rect 15979 31912 16672 31940
rect 15979 31909 15991 31912
rect 15933 31903 15991 31909
rect 16666 31900 16672 31912
rect 16724 31900 16730 31952
rect 18325 31943 18383 31949
rect 18325 31940 18337 31943
rect 16868 31912 18337 31940
rect 13541 31875 13599 31881
rect 13541 31841 13553 31875
rect 13587 31872 13599 31875
rect 14369 31875 14427 31881
rect 14369 31872 14381 31875
rect 13587 31844 14381 31872
rect 13587 31841 13599 31844
rect 13541 31835 13599 31841
rect 14369 31841 14381 31844
rect 14415 31841 14427 31875
rect 14369 31835 14427 31841
rect 12544 31776 12848 31804
rect 13449 31807 13507 31813
rect 13449 31773 13461 31807
rect 13495 31804 13507 31807
rect 13998 31804 14004 31816
rect 13495 31776 14004 31804
rect 13495 31773 13507 31776
rect 13449 31767 13507 31773
rect 13998 31764 14004 31776
rect 14056 31764 14062 31816
rect 14274 31804 14280 31816
rect 14235 31776 14280 31804
rect 14274 31764 14280 31776
rect 14332 31764 14338 31816
rect 14461 31807 14519 31813
rect 14461 31773 14473 31807
rect 14507 31804 14519 31807
rect 14642 31804 14648 31816
rect 14507 31776 14648 31804
rect 14507 31773 14519 31776
rect 14461 31767 14519 31773
rect 14642 31764 14648 31776
rect 14700 31804 14706 31816
rect 16868 31813 16896 31912
rect 18325 31909 18337 31912
rect 18371 31909 18383 31943
rect 18325 31903 18383 31909
rect 20530 31900 20536 31952
rect 20588 31940 20594 31952
rect 22554 31940 22560 31952
rect 20588 31912 22140 31940
rect 22467 31912 22560 31940
rect 20588 31900 20594 31912
rect 17126 31872 17132 31884
rect 17087 31844 17132 31872
rect 17126 31832 17132 31844
rect 17184 31832 17190 31884
rect 22112 31881 22140 31912
rect 22554 31900 22560 31912
rect 22612 31940 22618 31952
rect 24581 31943 24639 31949
rect 24581 31940 24593 31943
rect 22612 31912 24593 31940
rect 22612 31900 22618 31912
rect 24581 31909 24593 31912
rect 24627 31909 24639 31943
rect 24581 31903 24639 31909
rect 19429 31875 19487 31881
rect 19429 31872 19441 31875
rect 18340 31844 19441 31872
rect 16393 31807 16451 31813
rect 16393 31804 16405 31807
rect 14700 31776 16405 31804
rect 14700 31764 14706 31776
rect 16393 31773 16405 31776
rect 16439 31773 16451 31807
rect 16393 31767 16451 31773
rect 16853 31807 16911 31813
rect 16853 31773 16865 31807
rect 16899 31773 16911 31807
rect 17310 31804 17316 31816
rect 17271 31776 17316 31804
rect 16853 31767 16911 31773
rect 17310 31764 17316 31776
rect 17368 31764 17374 31816
rect 17862 31764 17868 31816
rect 17920 31804 17926 31816
rect 18340 31813 18368 31844
rect 19429 31841 19441 31844
rect 19475 31841 19487 31875
rect 22097 31875 22155 31881
rect 19429 31835 19487 31841
rect 20272 31844 21220 31872
rect 18325 31807 18383 31813
rect 18325 31804 18337 31807
rect 17920 31776 18337 31804
rect 17920 31764 17926 31776
rect 18325 31773 18337 31776
rect 18371 31773 18383 31807
rect 18506 31804 18512 31816
rect 18467 31776 18512 31804
rect 18325 31767 18383 31773
rect 18506 31764 18512 31776
rect 18564 31764 18570 31816
rect 20272 31813 20300 31844
rect 21192 31816 21220 31844
rect 22097 31841 22109 31875
rect 22143 31841 22155 31875
rect 22572 31872 22600 31900
rect 22649 31875 22707 31881
rect 22649 31872 22661 31875
rect 22572 31844 22661 31872
rect 22097 31835 22155 31841
rect 22649 31841 22661 31844
rect 22695 31841 22707 31875
rect 22649 31835 22707 31841
rect 22738 31832 22744 31884
rect 22796 31872 22802 31884
rect 23109 31875 23167 31881
rect 23109 31872 23121 31875
rect 22796 31844 23121 31872
rect 22796 31832 22802 31844
rect 23109 31841 23121 31844
rect 23155 31841 23167 31875
rect 25038 31872 25044 31884
rect 24999 31844 25044 31872
rect 23109 31835 23167 31841
rect 25038 31832 25044 31844
rect 25096 31832 25102 31884
rect 25130 31832 25136 31884
rect 25188 31872 25194 31884
rect 25188 31844 25233 31872
rect 25188 31832 25194 31844
rect 20257 31807 20315 31813
rect 20257 31773 20269 31807
rect 20303 31773 20315 31807
rect 20257 31767 20315 31773
rect 20441 31807 20499 31813
rect 20441 31773 20453 31807
rect 20487 31804 20499 31807
rect 20806 31804 20812 31816
rect 20487 31776 20812 31804
rect 20487 31773 20499 31776
rect 20441 31767 20499 31773
rect 20806 31764 20812 31776
rect 20864 31764 20870 31816
rect 20993 31807 21051 31813
rect 20993 31773 21005 31807
rect 21039 31804 21051 31807
rect 21082 31804 21088 31816
rect 21039 31776 21088 31804
rect 21039 31773 21051 31776
rect 20993 31767 21051 31773
rect 21082 31764 21088 31776
rect 21140 31764 21146 31816
rect 21174 31764 21180 31816
rect 21232 31764 21238 31816
rect 22922 31804 22928 31816
rect 22883 31776 22928 31804
rect 22922 31764 22928 31776
rect 22980 31764 22986 31816
rect 23750 31804 23756 31816
rect 23711 31776 23756 31804
rect 23750 31764 23756 31776
rect 23808 31764 23814 31816
rect 23937 31807 23995 31813
rect 23937 31773 23949 31807
rect 23983 31773 23995 31807
rect 26602 31804 26608 31816
rect 26563 31776 26608 31804
rect 23937 31767 23995 31773
rect 8496 31708 8800 31736
rect 10042 31696 10048 31748
rect 10100 31736 10106 31748
rect 15562 31736 15568 31748
rect 10100 31708 15568 31736
rect 10100 31696 10106 31708
rect 15562 31696 15568 31708
rect 15620 31696 15626 31748
rect 16114 31696 16120 31748
rect 16172 31736 16178 31748
rect 17221 31739 17279 31745
rect 17221 31736 17233 31739
rect 16172 31708 17233 31736
rect 16172 31696 16178 31708
rect 17221 31705 17233 31708
rect 17267 31705 17279 31739
rect 17221 31699 17279 31705
rect 8018 31628 8024 31680
rect 8076 31668 8082 31680
rect 11609 31671 11667 31677
rect 11609 31668 11621 31671
rect 8076 31640 11621 31668
rect 8076 31628 8082 31640
rect 11609 31637 11621 31640
rect 11655 31637 11667 31671
rect 11609 31631 11667 31637
rect 15746 31628 15752 31680
rect 15804 31677 15810 31680
rect 15804 31671 15823 31677
rect 15811 31637 15823 31671
rect 15804 31631 15823 31637
rect 21085 31671 21143 31677
rect 21085 31637 21097 31671
rect 21131 31668 21143 31671
rect 21192 31668 21220 31764
rect 21266 31696 21272 31748
rect 21324 31736 21330 31748
rect 21324 31708 21369 31736
rect 21324 31696 21330 31708
rect 22646 31696 22652 31748
rect 22704 31736 22710 31748
rect 22940 31736 22968 31764
rect 22704 31708 22968 31736
rect 22704 31696 22710 31708
rect 23382 31696 23388 31748
rect 23440 31736 23446 31748
rect 23952 31736 23980 31767
rect 26602 31764 26608 31776
rect 26660 31764 26666 31816
rect 27338 31804 27344 31816
rect 27299 31776 27344 31804
rect 27338 31764 27344 31776
rect 27396 31764 27402 31816
rect 27706 31736 27712 31748
rect 23440 31708 23980 31736
rect 27554 31708 27712 31736
rect 23440 31696 23446 31708
rect 27706 31696 27712 31708
rect 27764 31696 27770 31748
rect 23566 31668 23572 31680
rect 21131 31640 21220 31668
rect 23527 31640 23572 31668
rect 21131 31637 21143 31640
rect 21085 31631 21143 31637
rect 15804 31628 15810 31631
rect 23566 31628 23572 31640
rect 23624 31628 23630 31680
rect 24578 31628 24584 31680
rect 24636 31668 24642 31680
rect 24762 31668 24768 31680
rect 24636 31640 24768 31668
rect 24636 31628 24642 31640
rect 24762 31628 24768 31640
rect 24820 31668 24826 31680
rect 24949 31671 25007 31677
rect 24949 31668 24961 31671
rect 24820 31640 24961 31668
rect 24820 31628 24826 31640
rect 24949 31637 24961 31640
rect 24995 31637 25007 31671
rect 24949 31631 25007 31637
rect 1104 31578 35027 31600
rect 1104 31526 9390 31578
rect 9442 31526 9454 31578
rect 9506 31526 9518 31578
rect 9570 31526 9582 31578
rect 9634 31526 9646 31578
rect 9698 31526 17831 31578
rect 17883 31526 17895 31578
rect 17947 31526 17959 31578
rect 18011 31526 18023 31578
rect 18075 31526 18087 31578
rect 18139 31526 26272 31578
rect 26324 31526 26336 31578
rect 26388 31526 26400 31578
rect 26452 31526 26464 31578
rect 26516 31526 26528 31578
rect 26580 31526 34713 31578
rect 34765 31526 34777 31578
rect 34829 31526 34841 31578
rect 34893 31526 34905 31578
rect 34957 31526 34969 31578
rect 35021 31526 35027 31578
rect 1104 31504 35027 31526
rect 9493 31467 9551 31473
rect 9493 31433 9505 31467
rect 9539 31464 9551 31467
rect 9858 31464 9864 31476
rect 9539 31436 9864 31464
rect 9539 31433 9551 31436
rect 9493 31427 9551 31433
rect 9858 31424 9864 31436
rect 9916 31424 9922 31476
rect 13541 31467 13599 31473
rect 13541 31433 13553 31467
rect 13587 31464 13599 31467
rect 14274 31464 14280 31476
rect 13587 31436 14280 31464
rect 13587 31433 13599 31436
rect 13541 31427 13599 31433
rect 14274 31424 14280 31436
rect 14332 31424 14338 31476
rect 16114 31464 16120 31476
rect 16075 31436 16120 31464
rect 16114 31424 16120 31436
rect 16172 31464 16178 31476
rect 17037 31467 17095 31473
rect 17037 31464 17049 31467
rect 16172 31436 17049 31464
rect 16172 31424 16178 31436
rect 17037 31433 17049 31436
rect 17083 31433 17095 31467
rect 17037 31427 17095 31433
rect 17310 31424 17316 31476
rect 17368 31464 17374 31476
rect 17589 31467 17647 31473
rect 17589 31464 17601 31467
rect 17368 31436 17601 31464
rect 17368 31424 17374 31436
rect 17589 31433 17601 31436
rect 17635 31433 17647 31467
rect 17589 31427 17647 31433
rect 20806 31424 20812 31476
rect 20864 31473 20870 31476
rect 20864 31467 20892 31473
rect 20880 31433 20892 31467
rect 20864 31427 20892 31433
rect 24765 31467 24823 31473
rect 24765 31433 24777 31467
rect 24811 31464 24823 31467
rect 25130 31464 25136 31476
rect 24811 31436 25136 31464
rect 24811 31433 24823 31436
rect 24765 31427 24823 31433
rect 20864 31424 20870 31427
rect 25130 31424 25136 31436
rect 25188 31424 25194 31476
rect 25869 31467 25927 31473
rect 25869 31433 25881 31467
rect 25915 31464 25927 31467
rect 26602 31464 26608 31476
rect 25915 31436 26608 31464
rect 25915 31433 25927 31436
rect 25869 31427 25927 31433
rect 26602 31424 26608 31436
rect 26660 31424 26666 31476
rect 28626 31424 28632 31476
rect 28684 31464 28690 31476
rect 28813 31467 28871 31473
rect 28813 31464 28825 31467
rect 28684 31436 28825 31464
rect 28684 31424 28690 31436
rect 28813 31433 28825 31436
rect 28859 31433 28871 31467
rect 28813 31427 28871 31433
rect 10042 31356 10048 31408
rect 10100 31356 10106 31408
rect 10594 31356 10600 31408
rect 10652 31396 10658 31408
rect 10689 31399 10747 31405
rect 10689 31396 10701 31399
rect 10652 31368 10701 31396
rect 10652 31356 10658 31368
rect 10689 31365 10701 31368
rect 10735 31365 10747 31399
rect 10689 31359 10747 31365
rect 13188 31368 15516 31396
rect 9125 31331 9183 31337
rect 9125 31297 9137 31331
rect 9171 31328 9183 31331
rect 9858 31328 9864 31340
rect 9171 31300 9864 31328
rect 9171 31297 9183 31300
rect 9125 31291 9183 31297
rect 9858 31288 9864 31300
rect 9916 31328 9922 31340
rect 10060 31328 10088 31356
rect 10226 31328 10232 31340
rect 9916 31300 10088 31328
rect 10187 31300 10232 31328
rect 9916 31288 9922 31300
rect 10226 31288 10232 31300
rect 10284 31288 10290 31340
rect 10321 31331 10379 31337
rect 10321 31297 10333 31331
rect 10367 31297 10379 31331
rect 10321 31291 10379 31297
rect 9217 31263 9275 31269
rect 9217 31229 9229 31263
rect 9263 31260 9275 31263
rect 9398 31260 9404 31272
rect 9263 31232 9404 31260
rect 9263 31229 9275 31232
rect 9217 31223 9275 31229
rect 9398 31220 9404 31232
rect 9456 31220 9462 31272
rect 10042 31220 10048 31272
rect 10100 31260 10106 31272
rect 10336 31260 10364 31291
rect 13078 31288 13084 31340
rect 13136 31328 13142 31340
rect 13188 31337 13216 31368
rect 15488 31340 15516 31368
rect 15562 31356 15568 31408
rect 15620 31396 15626 31408
rect 16853 31399 16911 31405
rect 16853 31396 16865 31399
rect 15620 31368 16865 31396
rect 15620 31356 15626 31368
rect 16853 31365 16865 31368
rect 16899 31396 16911 31399
rect 20438 31396 20444 31408
rect 16899 31368 20444 31396
rect 16899 31365 16911 31368
rect 16853 31359 16911 31365
rect 20438 31356 20444 31368
rect 20496 31356 20502 31408
rect 22189 31399 22247 31405
rect 22189 31396 22201 31399
rect 20640 31368 22201 31396
rect 13173 31331 13231 31337
rect 13173 31328 13185 31331
rect 13136 31300 13185 31328
rect 13136 31288 13142 31300
rect 13173 31297 13185 31300
rect 13219 31297 13231 31331
rect 14090 31328 14096 31340
rect 14051 31300 14096 31328
rect 13173 31291 13231 31297
rect 14090 31288 14096 31300
rect 14148 31288 14154 31340
rect 14826 31328 14832 31340
rect 14787 31300 14832 31328
rect 14826 31288 14832 31300
rect 14884 31288 14890 31340
rect 14921 31331 14979 31337
rect 14921 31297 14933 31331
rect 14967 31297 14979 31331
rect 14921 31291 14979 31297
rect 10100 31232 10364 31260
rect 10100 31220 10106 31232
rect 10410 31220 10416 31272
rect 10468 31260 10474 31272
rect 13262 31260 13268 31272
rect 10468 31232 10513 31260
rect 13223 31232 13268 31260
rect 10468 31220 10474 31232
rect 13262 31220 13268 31232
rect 13320 31220 13326 31272
rect 13924 31232 14596 31260
rect 10962 31192 10968 31204
rect 10923 31164 10968 31192
rect 10962 31152 10968 31164
rect 11020 31152 11026 31204
rect 13924 31192 13952 31232
rect 11072 31164 13952 31192
rect 10686 31084 10692 31136
rect 10744 31124 10750 31136
rect 11072 31124 11100 31164
rect 14274 31124 14280 31136
rect 10744 31096 11100 31124
rect 14235 31096 14280 31124
rect 10744 31084 10750 31096
rect 14274 31084 14280 31096
rect 14332 31084 14338 31136
rect 14568 31124 14596 31232
rect 14642 31220 14648 31272
rect 14700 31260 14706 31272
rect 14936 31260 14964 31291
rect 15470 31288 15476 31340
rect 15528 31328 15534 31340
rect 16117 31331 16175 31337
rect 16117 31328 16129 31331
rect 15528 31300 16129 31328
rect 15528 31288 15534 31300
rect 16117 31297 16129 31300
rect 16163 31297 16175 31331
rect 16298 31328 16304 31340
rect 16259 31300 16304 31328
rect 16117 31291 16175 31297
rect 16298 31288 16304 31300
rect 16356 31288 16362 31340
rect 17126 31328 17132 31340
rect 17039 31300 17132 31328
rect 17126 31288 17132 31300
rect 17184 31288 17190 31340
rect 17589 31331 17647 31337
rect 17589 31297 17601 31331
rect 17635 31297 17647 31331
rect 17589 31291 17647 31297
rect 14700 31232 14964 31260
rect 14700 31220 14706 31232
rect 15746 31220 15752 31272
rect 15804 31260 15810 31272
rect 17144 31260 17172 31288
rect 15804 31232 17172 31260
rect 15804 31220 15810 31232
rect 17604 31192 17632 31291
rect 17678 31288 17684 31340
rect 17736 31328 17742 31340
rect 17773 31331 17831 31337
rect 17773 31328 17785 31331
rect 17736 31300 17785 31328
rect 17736 31288 17742 31300
rect 17773 31297 17785 31300
rect 17819 31297 17831 31331
rect 17773 31291 17831 31297
rect 20162 31288 20168 31340
rect 20220 31328 20226 31340
rect 20640 31337 20668 31368
rect 22189 31365 22201 31368
rect 22235 31365 22247 31399
rect 22189 31359 22247 31365
rect 24596 31368 25636 31396
rect 20625 31331 20683 31337
rect 20625 31328 20637 31331
rect 20220 31300 20637 31328
rect 20220 31288 20226 31300
rect 20625 31297 20637 31300
rect 20671 31297 20683 31331
rect 20625 31291 20683 31297
rect 20990 31288 20996 31340
rect 21048 31328 21054 31340
rect 21085 31331 21143 31337
rect 21085 31328 21097 31331
rect 21048 31300 21097 31328
rect 21048 31288 21054 31300
rect 21085 31297 21097 31300
rect 21131 31297 21143 31331
rect 22646 31328 22652 31340
rect 22607 31300 22652 31328
rect 21085 31291 21143 31297
rect 22646 31288 22652 31300
rect 22704 31288 22710 31340
rect 22738 31288 22744 31340
rect 22796 31328 22802 31340
rect 23014 31328 23020 31340
rect 22796 31300 22841 31328
rect 22975 31300 23020 31328
rect 22796 31288 22802 31300
rect 23014 31288 23020 31300
rect 23072 31288 23078 31340
rect 23293 31331 23351 31337
rect 23293 31297 23305 31331
rect 23339 31297 23351 31331
rect 23566 31328 23572 31340
rect 23527 31300 23572 31328
rect 23293 31291 23351 31297
rect 20530 31260 20536 31272
rect 20491 31232 20536 31260
rect 20530 31220 20536 31232
rect 20588 31220 20594 31272
rect 20898 31192 20904 31204
rect 16776 31164 20904 31192
rect 16776 31124 16804 31164
rect 20898 31152 20904 31164
rect 20956 31152 20962 31204
rect 21266 31152 21272 31204
rect 21324 31192 21330 31204
rect 21376 31192 21404 31246
rect 21450 31220 21456 31272
rect 21508 31260 21514 31272
rect 23308 31260 23336 31291
rect 23566 31288 23572 31300
rect 23624 31288 23630 31340
rect 24213 31331 24271 31337
rect 24213 31297 24225 31331
rect 24259 31328 24271 31331
rect 24486 31328 24492 31340
rect 24259 31300 24492 31328
rect 24259 31297 24271 31300
rect 24213 31291 24271 31297
rect 24486 31288 24492 31300
rect 24544 31288 24550 31340
rect 24596 31337 24624 31368
rect 24581 31331 24639 31337
rect 24581 31297 24593 31331
rect 24627 31297 24639 31331
rect 24581 31291 24639 31297
rect 25038 31288 25044 31340
rect 25096 31328 25102 31340
rect 25225 31331 25283 31337
rect 25225 31328 25237 31331
rect 25096 31300 25237 31328
rect 25096 31288 25102 31300
rect 25225 31297 25237 31300
rect 25271 31297 25283 31331
rect 25225 31291 25283 31297
rect 25314 31288 25320 31340
rect 25372 31328 25378 31340
rect 25409 31331 25467 31337
rect 25409 31328 25421 31331
rect 25372 31300 25421 31328
rect 25372 31288 25378 31300
rect 25409 31297 25421 31300
rect 25455 31297 25467 31331
rect 25409 31291 25467 31297
rect 25608 31269 25636 31368
rect 25685 31331 25743 31337
rect 25685 31297 25697 31331
rect 25731 31328 25743 31331
rect 26050 31328 26056 31340
rect 25731 31300 26056 31328
rect 25731 31297 25743 31300
rect 25685 31291 25743 31297
rect 26050 31288 26056 31300
rect 26108 31288 26114 31340
rect 27338 31328 27344 31340
rect 27299 31300 27344 31328
rect 27338 31288 27344 31300
rect 27396 31288 27402 31340
rect 27522 31288 27528 31340
rect 27580 31328 27586 31340
rect 27617 31331 27675 31337
rect 27617 31328 27629 31331
rect 27580 31300 27629 31328
rect 27580 31288 27586 31300
rect 27617 31297 27629 31300
rect 27663 31297 27675 31331
rect 27617 31291 27675 31297
rect 27706 31288 27712 31340
rect 27764 31328 27770 31340
rect 28353 31331 28411 31337
rect 28353 31328 28365 31331
rect 27764 31300 28365 31328
rect 27764 31288 27770 31300
rect 28353 31297 28365 31300
rect 28399 31297 28411 31331
rect 28353 31291 28411 31297
rect 28534 31288 28540 31340
rect 28592 31328 28598 31340
rect 28629 31331 28687 31337
rect 28629 31328 28641 31331
rect 28592 31300 28641 31328
rect 28592 31288 28598 31300
rect 28629 31297 28641 31300
rect 28675 31297 28687 31331
rect 28629 31291 28687 31297
rect 21508 31232 23336 31260
rect 25593 31263 25651 31269
rect 21508 31220 21514 31232
rect 25593 31229 25605 31263
rect 25639 31260 25651 31263
rect 25774 31260 25780 31272
rect 25639 31232 25780 31260
rect 25639 31229 25651 31232
rect 25593 31223 25651 31229
rect 25774 31220 25780 31232
rect 25832 31260 25838 31272
rect 27157 31263 27215 31269
rect 27157 31260 27169 31263
rect 25832 31232 27169 31260
rect 25832 31220 25838 31232
rect 27157 31229 27169 31232
rect 27203 31229 27215 31263
rect 27157 31223 27215 31229
rect 21726 31192 21732 31204
rect 21324 31164 21732 31192
rect 21324 31152 21330 31164
rect 21726 31152 21732 31164
rect 21784 31152 21790 31204
rect 22738 31152 22744 31204
rect 22796 31192 22802 31204
rect 23566 31192 23572 31204
rect 22796 31164 23572 31192
rect 22796 31152 22802 31164
rect 23566 31152 23572 31164
rect 23624 31152 23630 31204
rect 25501 31195 25559 31201
rect 25501 31161 25513 31195
rect 25547 31161 25559 31195
rect 28442 31192 28448 31204
rect 28403 31164 28448 31192
rect 25501 31155 25559 31161
rect 14568 31096 16804 31124
rect 16853 31127 16911 31133
rect 16853 31093 16865 31127
rect 16899 31124 16911 31127
rect 17034 31124 17040 31136
rect 16899 31096 17040 31124
rect 16899 31093 16911 31096
rect 16853 31087 16911 31093
rect 17034 31084 17040 31096
rect 17092 31084 17098 31136
rect 24581 31127 24639 31133
rect 24581 31093 24593 31127
rect 24627 31124 24639 31127
rect 25516 31124 25544 31155
rect 28442 31152 28448 31164
rect 28500 31152 28506 31204
rect 25590 31124 25596 31136
rect 24627 31096 25596 31124
rect 24627 31093 24639 31096
rect 24581 31087 24639 31093
rect 25590 31084 25596 31096
rect 25648 31084 25654 31136
rect 1104 31034 34868 31056
rect 1104 30982 5170 31034
rect 5222 30982 5234 31034
rect 5286 30982 5298 31034
rect 5350 30982 5362 31034
rect 5414 30982 5426 31034
rect 5478 30982 13611 31034
rect 13663 30982 13675 31034
rect 13727 30982 13739 31034
rect 13791 30982 13803 31034
rect 13855 30982 13867 31034
rect 13919 30982 22052 31034
rect 22104 30982 22116 31034
rect 22168 30982 22180 31034
rect 22232 30982 22244 31034
rect 22296 30982 22308 31034
rect 22360 30982 30493 31034
rect 30545 30982 30557 31034
rect 30609 30982 30621 31034
rect 30673 30982 30685 31034
rect 30737 30982 30749 31034
rect 30801 30982 34868 31034
rect 1104 30960 34868 30982
rect 9398 30920 9404 30932
rect 9359 30892 9404 30920
rect 9398 30880 9404 30892
rect 9456 30880 9462 30932
rect 10042 30920 10048 30932
rect 10003 30892 10048 30920
rect 10042 30880 10048 30892
rect 10100 30880 10106 30932
rect 10226 30880 10232 30932
rect 10284 30920 10290 30932
rect 10689 30923 10747 30929
rect 10689 30920 10701 30923
rect 10284 30892 10701 30920
rect 10284 30880 10290 30892
rect 10689 30889 10701 30892
rect 10735 30889 10747 30923
rect 10689 30883 10747 30889
rect 13262 30880 13268 30932
rect 13320 30920 13326 30932
rect 13541 30923 13599 30929
rect 13541 30920 13553 30923
rect 13320 30892 13553 30920
rect 13320 30880 13326 30892
rect 13541 30889 13553 30892
rect 13587 30889 13599 30923
rect 13541 30883 13599 30889
rect 17037 30923 17095 30929
rect 17037 30889 17049 30923
rect 17083 30920 17095 30923
rect 17402 30920 17408 30932
rect 17083 30892 17408 30920
rect 17083 30889 17095 30892
rect 17037 30883 17095 30889
rect 17402 30880 17408 30892
rect 17460 30880 17466 30932
rect 20990 30920 20996 30932
rect 20951 30892 20996 30920
rect 20990 30880 20996 30892
rect 21048 30880 21054 30932
rect 22833 30923 22891 30929
rect 22833 30889 22845 30923
rect 22879 30920 22891 30923
rect 23014 30920 23020 30932
rect 22879 30892 23020 30920
rect 22879 30889 22891 30892
rect 22833 30883 22891 30889
rect 23014 30880 23020 30892
rect 23072 30880 23078 30932
rect 10060 30784 10088 30880
rect 14826 30812 14832 30864
rect 14884 30852 14890 30864
rect 24946 30852 24952 30864
rect 14884 30824 16160 30852
rect 24907 30824 24952 30852
rect 14884 30812 14890 30824
rect 9324 30756 10088 30784
rect 9324 30725 9352 30756
rect 10502 30744 10508 30796
rect 10560 30784 10566 30796
rect 13449 30787 13507 30793
rect 10560 30756 10824 30784
rect 10560 30744 10566 30756
rect 9309 30719 9367 30725
rect 9309 30685 9321 30719
rect 9355 30685 9367 30719
rect 9309 30679 9367 30685
rect 9493 30719 9551 30725
rect 9493 30685 9505 30719
rect 9539 30685 9551 30719
rect 9950 30716 9956 30728
rect 9911 30688 9956 30716
rect 9493 30679 9551 30685
rect 9508 30648 9536 30679
rect 9950 30676 9956 30688
rect 10008 30676 10014 30728
rect 10137 30719 10195 30725
rect 10137 30685 10149 30719
rect 10183 30716 10195 30719
rect 10597 30719 10655 30725
rect 10183 30688 10548 30716
rect 10183 30685 10195 30688
rect 10137 30679 10195 30685
rect 10520 30660 10548 30688
rect 10597 30685 10609 30719
rect 10643 30716 10655 30719
rect 10686 30716 10692 30728
rect 10643 30688 10692 30716
rect 10643 30685 10655 30688
rect 10597 30679 10655 30685
rect 10686 30676 10692 30688
rect 10744 30676 10750 30728
rect 10796 30725 10824 30756
rect 13449 30753 13461 30787
rect 13495 30784 13507 30787
rect 14844 30784 14872 30812
rect 15746 30784 15752 30796
rect 13495 30756 14872 30784
rect 15707 30756 15752 30784
rect 13495 30753 13507 30756
rect 13449 30747 13507 30753
rect 15746 30744 15752 30756
rect 15804 30744 15810 30796
rect 10781 30719 10839 30725
rect 10781 30685 10793 30719
rect 10827 30685 10839 30719
rect 10781 30679 10839 30685
rect 13633 30719 13691 30725
rect 13633 30685 13645 30719
rect 13679 30685 13691 30719
rect 13633 30679 13691 30685
rect 13725 30719 13783 30725
rect 13725 30685 13737 30719
rect 13771 30716 13783 30719
rect 14090 30716 14096 30728
rect 13771 30688 14096 30716
rect 13771 30685 13783 30688
rect 13725 30679 13783 30685
rect 10410 30648 10416 30660
rect 9508 30620 10416 30648
rect 10410 30608 10416 30620
rect 10468 30608 10474 30660
rect 10502 30608 10508 30660
rect 10560 30608 10566 30660
rect 13648 30648 13676 30679
rect 14090 30676 14096 30688
rect 14148 30716 14154 30728
rect 14550 30716 14556 30728
rect 14148 30688 14556 30716
rect 14148 30676 14154 30688
rect 14550 30676 14556 30688
rect 14608 30676 14614 30728
rect 14918 30716 14924 30728
rect 14879 30688 14924 30716
rect 14918 30676 14924 30688
rect 14976 30676 14982 30728
rect 15470 30716 15476 30728
rect 15431 30688 15476 30716
rect 15470 30676 15476 30688
rect 15528 30676 15534 30728
rect 16132 30725 16160 30824
rect 24946 30812 24952 30824
rect 25004 30852 25010 30864
rect 25004 30824 27660 30852
rect 25004 30812 25010 30824
rect 20625 30787 20683 30793
rect 20625 30753 20637 30787
rect 20671 30784 20683 30787
rect 23201 30787 23259 30793
rect 20671 30756 22094 30784
rect 20671 30753 20683 30756
rect 20625 30747 20683 30753
rect 15933 30719 15991 30725
rect 15933 30685 15945 30719
rect 15979 30685 15991 30719
rect 15933 30679 15991 30685
rect 16117 30719 16175 30725
rect 16117 30685 16129 30719
rect 16163 30685 16175 30719
rect 16117 30679 16175 30685
rect 14936 30648 14964 30676
rect 13648 30620 14964 30648
rect 15948 30648 15976 30679
rect 16666 30676 16672 30728
rect 16724 30716 16730 30728
rect 16853 30719 16911 30725
rect 16853 30716 16865 30719
rect 16724 30688 16865 30716
rect 16724 30676 16730 30688
rect 16853 30685 16865 30688
rect 16899 30685 16911 30719
rect 17034 30716 17040 30728
rect 16995 30688 17040 30716
rect 16853 30679 16911 30685
rect 17034 30676 17040 30688
rect 17092 30676 17098 30728
rect 20809 30719 20867 30725
rect 20809 30685 20821 30719
rect 20855 30716 20867 30719
rect 21450 30716 21456 30728
rect 20855 30688 21456 30716
rect 20855 30685 20867 30688
rect 20809 30679 20867 30685
rect 21450 30676 21456 30688
rect 21508 30676 21514 30728
rect 22066 30716 22094 30756
rect 23201 30753 23213 30787
rect 23247 30784 23259 30787
rect 23382 30784 23388 30796
rect 23247 30756 23388 30784
rect 23247 30753 23259 30756
rect 23201 30747 23259 30753
rect 23382 30744 23388 30756
rect 23440 30784 23446 30796
rect 27433 30787 27491 30793
rect 27433 30784 27445 30787
rect 23440 30756 27445 30784
rect 23440 30744 23446 30756
rect 27433 30753 27445 30756
rect 27479 30753 27491 30787
rect 27433 30747 27491 30753
rect 23017 30719 23075 30725
rect 23017 30716 23029 30719
rect 22066 30688 23029 30716
rect 23017 30685 23029 30688
rect 23063 30685 23075 30719
rect 23290 30716 23296 30728
rect 23251 30688 23296 30716
rect 23017 30679 23075 30685
rect 16298 30648 16304 30660
rect 15948 30620 16304 30648
rect 13998 30540 14004 30592
rect 14056 30580 14062 30592
rect 15948 30580 15976 30620
rect 16298 30608 16304 30620
rect 16356 30648 16362 30660
rect 18782 30648 18788 30660
rect 16356 30620 18788 30648
rect 16356 30608 16362 30620
rect 18782 30608 18788 30620
rect 18840 30608 18846 30660
rect 23032 30648 23060 30679
rect 23290 30676 23296 30688
rect 23348 30676 23354 30728
rect 25133 30719 25191 30725
rect 25133 30685 25145 30719
rect 25179 30716 25191 30719
rect 25314 30716 25320 30728
rect 25179 30688 25320 30716
rect 25179 30685 25191 30688
rect 25133 30679 25191 30685
rect 25314 30676 25320 30688
rect 25372 30676 25378 30728
rect 25590 30716 25596 30728
rect 25551 30688 25596 30716
rect 25590 30676 25596 30688
rect 25648 30676 25654 30728
rect 25774 30716 25780 30728
rect 25735 30688 25780 30716
rect 25774 30676 25780 30688
rect 25832 30676 25838 30728
rect 26050 30676 26056 30728
rect 26108 30716 26114 30728
rect 27632 30725 27660 30824
rect 26145 30719 26203 30725
rect 26145 30716 26157 30719
rect 26108 30688 26157 30716
rect 26108 30676 26114 30688
rect 26145 30685 26157 30688
rect 26191 30685 26203 30719
rect 26145 30679 26203 30685
rect 27617 30719 27675 30725
rect 27617 30685 27629 30719
rect 27663 30716 27675 30719
rect 27706 30716 27712 30728
rect 27663 30688 27712 30716
rect 27663 30685 27675 30688
rect 27617 30679 27675 30685
rect 27706 30676 27712 30688
rect 27764 30676 27770 30728
rect 28074 30716 28080 30728
rect 28035 30688 28080 30716
rect 28074 30676 28080 30688
rect 28132 30676 28138 30728
rect 28445 30719 28503 30725
rect 28445 30685 28457 30719
rect 28491 30685 28503 30719
rect 28626 30716 28632 30728
rect 28587 30688 28632 30716
rect 28445 30679 28503 30685
rect 23750 30648 23756 30660
rect 23032 30620 23756 30648
rect 23750 30608 23756 30620
rect 23808 30648 23814 30660
rect 25038 30648 25044 30660
rect 23808 30620 25044 30648
rect 23808 30608 23814 30620
rect 25038 30608 25044 30620
rect 25096 30608 25102 30660
rect 28460 30648 28488 30679
rect 28626 30676 28632 30688
rect 28684 30676 28690 30728
rect 28534 30648 28540 30660
rect 28460 30620 28540 30648
rect 28534 30608 28540 30620
rect 28592 30608 28598 30660
rect 14056 30552 15976 30580
rect 14056 30540 14062 30552
rect 1104 30490 35027 30512
rect 1104 30438 9390 30490
rect 9442 30438 9454 30490
rect 9506 30438 9518 30490
rect 9570 30438 9582 30490
rect 9634 30438 9646 30490
rect 9698 30438 17831 30490
rect 17883 30438 17895 30490
rect 17947 30438 17959 30490
rect 18011 30438 18023 30490
rect 18075 30438 18087 30490
rect 18139 30438 26272 30490
rect 26324 30438 26336 30490
rect 26388 30438 26400 30490
rect 26452 30438 26464 30490
rect 26516 30438 26528 30490
rect 26580 30438 34713 30490
rect 34765 30438 34777 30490
rect 34829 30438 34841 30490
rect 34893 30438 34905 30490
rect 34957 30438 34969 30490
rect 35021 30438 35027 30490
rect 1104 30416 35027 30438
rect 25038 30336 25044 30388
rect 25096 30376 25102 30388
rect 25096 30348 26280 30376
rect 25096 30336 25102 30348
rect 18788 30320 18840 30326
rect 21542 30308 21548 30320
rect 18788 30262 18840 30268
rect 19628 30280 21548 30308
rect 14274 30240 14280 30252
rect 14235 30212 14280 30240
rect 14274 30200 14280 30212
rect 14332 30200 14338 30252
rect 14918 30240 14924 30252
rect 14879 30212 14924 30240
rect 14918 30200 14924 30212
rect 14976 30200 14982 30252
rect 19153 30243 19211 30249
rect 19153 30209 19165 30243
rect 19199 30240 19211 30243
rect 19628 30240 19656 30280
rect 21542 30268 21548 30280
rect 21600 30268 21606 30320
rect 19199 30212 19656 30240
rect 19705 30243 19763 30249
rect 19199 30209 19211 30212
rect 19153 30203 19211 30209
rect 19705 30209 19717 30243
rect 19751 30240 19763 30243
rect 20254 30240 20260 30252
rect 19751 30212 20260 30240
rect 19751 30209 19763 30212
rect 19705 30203 19763 30209
rect 20254 30200 20260 30212
rect 20312 30200 20318 30252
rect 20993 30243 21051 30249
rect 20993 30209 21005 30243
rect 21039 30240 21051 30243
rect 21266 30240 21272 30252
rect 21039 30212 21272 30240
rect 21039 30209 21051 30212
rect 20993 30203 21051 30209
rect 21266 30200 21272 30212
rect 21324 30200 21330 30252
rect 24670 30240 24676 30252
rect 24631 30212 24676 30240
rect 24670 30200 24676 30212
rect 24728 30200 24734 30252
rect 25225 30243 25283 30249
rect 25225 30209 25237 30243
rect 25271 30209 25283 30243
rect 25225 30203 25283 30209
rect 25240 30172 25268 30203
rect 25314 30200 25320 30252
rect 25372 30240 25378 30252
rect 25372 30212 25417 30240
rect 25372 30200 25378 30212
rect 25590 30200 25596 30252
rect 25648 30240 25654 30252
rect 25685 30243 25743 30249
rect 25685 30240 25697 30243
rect 25648 30212 25697 30240
rect 25648 30200 25654 30212
rect 25685 30209 25697 30212
rect 25731 30209 25743 30243
rect 25685 30203 25743 30209
rect 25406 30172 25412 30184
rect 25240 30144 25412 30172
rect 25406 30132 25412 30144
rect 25464 30132 25470 30184
rect 25700 30172 25728 30203
rect 25774 30200 25780 30252
rect 25832 30240 25838 30252
rect 25869 30243 25927 30249
rect 25869 30240 25881 30243
rect 25832 30212 25881 30240
rect 25832 30200 25838 30212
rect 25869 30209 25881 30212
rect 25915 30209 25927 30243
rect 26050 30240 26056 30252
rect 26011 30212 26056 30240
rect 25869 30203 25927 30209
rect 26050 30200 26056 30212
rect 26108 30200 26114 30252
rect 26252 30240 26280 30348
rect 27154 30336 27160 30388
rect 27212 30376 27218 30388
rect 27338 30376 27344 30388
rect 27212 30348 27344 30376
rect 27212 30336 27218 30348
rect 27338 30336 27344 30348
rect 27396 30376 27402 30388
rect 27433 30379 27491 30385
rect 27433 30376 27445 30379
rect 27396 30348 27445 30376
rect 27396 30336 27402 30348
rect 27433 30345 27445 30348
rect 27479 30345 27491 30379
rect 27433 30339 27491 30345
rect 28353 30379 28411 30385
rect 28353 30345 28365 30379
rect 28399 30376 28411 30379
rect 28442 30376 28448 30388
rect 28399 30348 28448 30376
rect 28399 30345 28411 30348
rect 28353 30339 28411 30345
rect 28442 30336 28448 30348
rect 28500 30336 28506 30388
rect 28074 30268 28080 30320
rect 28132 30308 28138 30320
rect 29549 30311 29607 30317
rect 29549 30308 29561 30311
rect 28132 30280 29561 30308
rect 28132 30268 28138 30280
rect 27371 30243 27429 30249
rect 27371 30240 27383 30243
rect 26252 30212 27383 30240
rect 27371 30209 27383 30212
rect 27417 30240 27429 30243
rect 27522 30240 27528 30252
rect 27417 30212 27528 30240
rect 27417 30209 27429 30212
rect 27371 30203 27429 30209
rect 27522 30200 27528 30212
rect 27580 30200 27586 30252
rect 28552 30249 28580 30280
rect 29549 30277 29561 30280
rect 29595 30277 29607 30311
rect 30745 30311 30803 30317
rect 30745 30308 30757 30311
rect 29549 30271 29607 30277
rect 29656 30280 30757 30308
rect 28537 30243 28595 30249
rect 28537 30209 28549 30243
rect 28583 30209 28595 30243
rect 28537 30203 28595 30209
rect 28813 30243 28871 30249
rect 28813 30209 28825 30243
rect 28859 30209 28871 30243
rect 28813 30203 28871 30209
rect 27890 30172 27896 30184
rect 25700 30144 27292 30172
rect 27803 30144 27896 30172
rect 27264 30113 27292 30144
rect 27890 30132 27896 30144
rect 27948 30172 27954 30184
rect 28828 30172 28856 30203
rect 28902 30200 28908 30252
rect 28960 30240 28966 30252
rect 28997 30243 29055 30249
rect 28997 30240 29009 30243
rect 28960 30212 29009 30240
rect 28960 30200 28966 30212
rect 28997 30209 29009 30212
rect 29043 30209 29055 30243
rect 28997 30203 29055 30209
rect 29086 30172 29092 30184
rect 27948 30144 28580 30172
rect 28828 30144 29092 30172
rect 27948 30132 27954 30144
rect 28552 30116 28580 30144
rect 29086 30132 29092 30144
rect 29144 30132 29150 30184
rect 27249 30107 27307 30113
rect 27249 30073 27261 30107
rect 27295 30073 27307 30107
rect 27249 30067 27307 30073
rect 27801 30107 27859 30113
rect 27801 30073 27813 30107
rect 27847 30104 27859 30107
rect 28442 30104 28448 30116
rect 27847 30076 28448 30104
rect 27847 30073 27859 30076
rect 27801 30067 27859 30073
rect 28442 30064 28448 30076
rect 28500 30064 28506 30116
rect 28534 30064 28540 30116
rect 28592 30104 28598 30116
rect 29656 30104 29684 30280
rect 30745 30277 30757 30280
rect 30791 30277 30803 30311
rect 30745 30271 30803 30277
rect 29733 30243 29791 30249
rect 29733 30209 29745 30243
rect 29779 30240 29791 30243
rect 29779 30212 29868 30240
rect 29779 30209 29791 30212
rect 29733 30203 29791 30209
rect 28592 30076 29684 30104
rect 29840 30172 29868 30212
rect 29914 30200 29920 30252
rect 29972 30240 29978 30252
rect 30377 30243 30435 30249
rect 30377 30240 30389 30243
rect 29972 30212 30389 30240
rect 29972 30200 29978 30212
rect 30377 30209 30389 30212
rect 30423 30209 30435 30243
rect 30377 30203 30435 30209
rect 30561 30243 30619 30249
rect 30561 30209 30573 30243
rect 30607 30209 30619 30243
rect 30561 30203 30619 30209
rect 30576 30172 30604 30203
rect 29840 30144 30604 30172
rect 28592 30064 28598 30076
rect 12894 29996 12900 30048
rect 12952 30036 12958 30048
rect 13449 30039 13507 30045
rect 13449 30036 13461 30039
rect 12952 30008 13461 30036
rect 12952 29996 12958 30008
rect 13449 30005 13461 30008
rect 13495 30005 13507 30039
rect 13449 29999 13507 30005
rect 20714 29996 20720 30048
rect 20772 30036 20778 30048
rect 20901 30039 20959 30045
rect 20901 30036 20913 30039
rect 20772 30008 20913 30036
rect 20772 29996 20778 30008
rect 20901 30005 20913 30008
rect 20947 30005 20959 30039
rect 20901 29999 20959 30005
rect 27522 29996 27528 30048
rect 27580 30036 27586 30048
rect 29840 30036 29868 30144
rect 27580 30008 29868 30036
rect 27580 29996 27586 30008
rect 1104 29946 34868 29968
rect 1104 29894 5170 29946
rect 5222 29894 5234 29946
rect 5286 29894 5298 29946
rect 5350 29894 5362 29946
rect 5414 29894 5426 29946
rect 5478 29894 13611 29946
rect 13663 29894 13675 29946
rect 13727 29894 13739 29946
rect 13791 29894 13803 29946
rect 13855 29894 13867 29946
rect 13919 29894 22052 29946
rect 22104 29894 22116 29946
rect 22168 29894 22180 29946
rect 22232 29894 22244 29946
rect 22296 29894 22308 29946
rect 22360 29894 30493 29946
rect 30545 29894 30557 29946
rect 30609 29894 30621 29946
rect 30673 29894 30685 29946
rect 30737 29894 30749 29946
rect 30801 29894 34868 29946
rect 1104 29872 34868 29894
rect 10502 29832 10508 29844
rect 9600 29804 10508 29832
rect 9600 29637 9628 29804
rect 10502 29792 10508 29804
rect 10560 29792 10566 29844
rect 14826 29832 14832 29844
rect 14787 29804 14832 29832
rect 14826 29792 14832 29804
rect 14884 29792 14890 29844
rect 25133 29835 25191 29841
rect 25133 29801 25145 29835
rect 25179 29832 25191 29835
rect 26050 29832 26056 29844
rect 25179 29804 26056 29832
rect 25179 29801 25191 29804
rect 25133 29795 25191 29801
rect 26050 29792 26056 29804
rect 26108 29792 26114 29844
rect 27430 29792 27436 29844
rect 27488 29832 27494 29844
rect 29914 29832 29920 29844
rect 27488 29804 29920 29832
rect 27488 29792 27494 29804
rect 29914 29792 29920 29804
rect 29972 29792 29978 29844
rect 19628 29736 22094 29764
rect 9950 29696 9956 29708
rect 9784 29668 9956 29696
rect 9784 29637 9812 29668
rect 9950 29656 9956 29668
rect 10008 29696 10014 29708
rect 12618 29696 12624 29708
rect 10008 29668 12624 29696
rect 10008 29656 10014 29668
rect 9585 29631 9643 29637
rect 9585 29597 9597 29631
rect 9631 29597 9643 29631
rect 9585 29591 9643 29597
rect 9769 29631 9827 29637
rect 9769 29597 9781 29631
rect 9815 29597 9827 29631
rect 9769 29591 9827 29597
rect 9861 29631 9919 29637
rect 9861 29597 9873 29631
rect 9907 29597 9919 29631
rect 10244 29630 10272 29668
rect 12618 29656 12624 29668
rect 12676 29696 12682 29708
rect 13078 29696 13084 29708
rect 12676 29668 13084 29696
rect 12676 29656 12682 29668
rect 13078 29656 13084 29668
rect 13136 29656 13142 29708
rect 10321 29631 10379 29637
rect 10321 29630 10333 29631
rect 10244 29602 10333 29630
rect 9861 29591 9919 29597
rect 10321 29597 10333 29602
rect 10367 29597 10379 29631
rect 10321 29591 10379 29597
rect 10413 29631 10471 29637
rect 10413 29597 10425 29631
rect 10459 29628 10471 29631
rect 10502 29628 10508 29640
rect 10459 29600 10508 29628
rect 10459 29597 10471 29600
rect 10413 29591 10471 29597
rect 9876 29560 9904 29591
rect 10502 29588 10508 29600
rect 10560 29628 10566 29640
rect 12894 29628 12900 29640
rect 10560 29600 12900 29628
rect 10560 29588 10566 29600
rect 12894 29588 12900 29600
rect 12952 29588 12958 29640
rect 12989 29631 13047 29637
rect 12989 29597 13001 29631
rect 13035 29597 13047 29631
rect 12989 29591 13047 29597
rect 13173 29631 13231 29637
rect 13173 29597 13185 29631
rect 13219 29628 13231 29631
rect 14921 29631 14979 29637
rect 14921 29628 14933 29631
rect 13219 29600 14933 29628
rect 13219 29597 13231 29600
rect 13173 29591 13231 29597
rect 14921 29597 14933 29600
rect 14967 29628 14979 29631
rect 15010 29628 15016 29640
rect 14967 29600 15016 29628
rect 14967 29597 14979 29600
rect 14921 29591 14979 29597
rect 10597 29563 10655 29569
rect 10597 29560 10609 29563
rect 9876 29532 10609 29560
rect 10597 29529 10609 29532
rect 10643 29560 10655 29563
rect 10962 29560 10968 29572
rect 10643 29532 10968 29560
rect 10643 29529 10655 29532
rect 10597 29523 10655 29529
rect 10962 29520 10968 29532
rect 11020 29520 11026 29572
rect 13004 29560 13032 29591
rect 15010 29588 15016 29600
rect 15068 29588 15074 29640
rect 19242 29588 19248 29640
rect 19300 29628 19306 29640
rect 19628 29637 19656 29736
rect 20441 29699 20499 29705
rect 20441 29665 20453 29699
rect 20487 29696 20499 29699
rect 20530 29696 20536 29708
rect 20487 29668 20536 29696
rect 20487 29665 20499 29668
rect 20441 29659 20499 29665
rect 20530 29656 20536 29668
rect 20588 29656 20594 29708
rect 21542 29696 21548 29708
rect 21503 29668 21548 29696
rect 21542 29656 21548 29668
rect 21600 29656 21606 29708
rect 22066 29696 22094 29736
rect 23290 29724 23296 29776
rect 23348 29764 23354 29776
rect 27341 29767 27399 29773
rect 27341 29764 27353 29767
rect 23348 29736 27353 29764
rect 23348 29724 23354 29736
rect 27341 29733 27353 29736
rect 27387 29733 27399 29767
rect 27890 29764 27896 29776
rect 27341 29727 27399 29733
rect 27540 29736 27896 29764
rect 27430 29696 27436 29708
rect 22066 29668 27436 29696
rect 27430 29656 27436 29668
rect 27488 29656 27494 29708
rect 19613 29631 19671 29637
rect 19613 29628 19625 29631
rect 19300 29600 19625 29628
rect 19300 29588 19306 29600
rect 19613 29597 19625 29600
rect 19659 29597 19671 29631
rect 20162 29628 20168 29640
rect 20123 29600 20168 29628
rect 19613 29591 19671 29597
rect 20162 29588 20168 29600
rect 20220 29588 20226 29640
rect 20806 29588 20812 29640
rect 20864 29628 20870 29640
rect 20993 29631 21051 29637
rect 20993 29628 21005 29631
rect 20864 29600 21005 29628
rect 20864 29588 20870 29600
rect 20993 29597 21005 29600
rect 21039 29597 21051 29631
rect 20993 29591 21051 29597
rect 21266 29588 21272 29640
rect 21324 29628 21330 29640
rect 21361 29631 21419 29637
rect 21361 29628 21373 29631
rect 21324 29600 21373 29628
rect 21324 29588 21330 29600
rect 21361 29597 21373 29600
rect 21407 29628 21419 29631
rect 21634 29628 21640 29640
rect 21407 29600 21640 29628
rect 21407 29597 21419 29600
rect 21361 29591 21419 29597
rect 21634 29588 21640 29600
rect 21692 29588 21698 29640
rect 24762 29628 24768 29640
rect 24723 29600 24768 29628
rect 24762 29588 24768 29600
rect 24820 29588 24826 29640
rect 27540 29637 27568 29736
rect 27890 29724 27896 29736
rect 27948 29724 27954 29776
rect 27621 29699 27679 29705
rect 27621 29665 27633 29699
rect 27667 29696 27679 29699
rect 28074 29696 28080 29708
rect 27667 29668 28080 29696
rect 27667 29665 27679 29668
rect 27621 29659 27679 29665
rect 28074 29656 28080 29668
rect 28132 29656 28138 29708
rect 28626 29696 28632 29708
rect 28184 29668 28632 29696
rect 24949 29631 25007 29637
rect 24949 29597 24961 29631
rect 24995 29597 25007 29631
rect 24949 29591 25007 29597
rect 27525 29631 27583 29637
rect 27525 29597 27537 29631
rect 27571 29597 27583 29631
rect 27706 29628 27712 29640
rect 27667 29600 27712 29628
rect 27525 29591 27583 29597
rect 14274 29560 14280 29572
rect 13004 29532 14280 29560
rect 14274 29520 14280 29532
rect 14332 29520 14338 29572
rect 15102 29560 15108 29572
rect 15063 29532 15108 29560
rect 15102 29520 15108 29532
rect 15160 29520 15166 29572
rect 24578 29520 24584 29572
rect 24636 29560 24642 29572
rect 24964 29560 24992 29591
rect 27706 29588 27712 29600
rect 27764 29588 27770 29640
rect 27801 29631 27859 29637
rect 27801 29597 27813 29631
rect 27847 29628 27859 29631
rect 28184 29628 28212 29668
rect 28626 29656 28632 29668
rect 28684 29656 28690 29708
rect 27847 29600 28212 29628
rect 27847 29597 27859 29600
rect 27801 29591 27859 29597
rect 28258 29588 28264 29640
rect 28316 29628 28322 29640
rect 28353 29631 28411 29637
rect 28353 29628 28365 29631
rect 28316 29600 28365 29628
rect 28316 29588 28322 29600
rect 28353 29597 28365 29600
rect 28399 29597 28411 29631
rect 28353 29591 28411 29597
rect 28537 29631 28595 29637
rect 28537 29597 28549 29631
rect 28583 29597 28595 29631
rect 28537 29591 28595 29597
rect 24636 29532 24992 29560
rect 24636 29520 24642 29532
rect 25406 29520 25412 29572
rect 25464 29560 25470 29572
rect 26050 29560 26056 29572
rect 25464 29532 26056 29560
rect 25464 29520 25470 29532
rect 26050 29520 26056 29532
rect 26108 29560 26114 29572
rect 28552 29560 28580 29591
rect 28810 29588 28816 29640
rect 28868 29628 28874 29640
rect 28905 29631 28963 29637
rect 28905 29628 28917 29631
rect 28868 29600 28917 29628
rect 28868 29588 28874 29600
rect 28905 29597 28917 29600
rect 28951 29597 28963 29631
rect 28905 29591 28963 29597
rect 26108 29532 28580 29560
rect 26108 29520 26114 29532
rect 9306 29452 9312 29504
rect 9364 29492 9370 29504
rect 9401 29495 9459 29501
rect 9401 29492 9413 29495
rect 9364 29464 9413 29492
rect 9364 29452 9370 29464
rect 9401 29461 9413 29464
rect 9447 29461 9459 29495
rect 10318 29492 10324 29504
rect 10279 29464 10324 29492
rect 9401 29455 9459 29461
rect 10318 29452 10324 29464
rect 10376 29452 10382 29504
rect 12802 29492 12808 29504
rect 12763 29464 12808 29492
rect 12802 29452 12808 29464
rect 12860 29452 12866 29504
rect 19426 29452 19432 29504
rect 19484 29492 19490 29504
rect 19521 29495 19579 29501
rect 19521 29492 19533 29495
rect 19484 29464 19533 29492
rect 19484 29452 19490 29464
rect 19521 29461 19533 29464
rect 19567 29461 19579 29495
rect 19521 29455 19579 29461
rect 21361 29495 21419 29501
rect 21361 29461 21373 29495
rect 21407 29492 21419 29495
rect 21450 29492 21456 29504
rect 21407 29464 21456 29492
rect 21407 29461 21419 29464
rect 21361 29455 21419 29461
rect 21450 29452 21456 29464
rect 21508 29452 21514 29504
rect 28813 29495 28871 29501
rect 28813 29461 28825 29495
rect 28859 29492 28871 29495
rect 29086 29492 29092 29504
rect 28859 29464 29092 29492
rect 28859 29461 28871 29464
rect 28813 29455 28871 29461
rect 29086 29452 29092 29464
rect 29144 29452 29150 29504
rect 1104 29402 35027 29424
rect 1104 29350 9390 29402
rect 9442 29350 9454 29402
rect 9506 29350 9518 29402
rect 9570 29350 9582 29402
rect 9634 29350 9646 29402
rect 9698 29350 17831 29402
rect 17883 29350 17895 29402
rect 17947 29350 17959 29402
rect 18011 29350 18023 29402
rect 18075 29350 18087 29402
rect 18139 29350 26272 29402
rect 26324 29350 26336 29402
rect 26388 29350 26400 29402
rect 26452 29350 26464 29402
rect 26516 29350 26528 29402
rect 26580 29350 34713 29402
rect 34765 29350 34777 29402
rect 34829 29350 34841 29402
rect 34893 29350 34905 29402
rect 34957 29350 34969 29402
rect 35021 29350 35027 29402
rect 1104 29328 35027 29350
rect 8128 29260 9536 29288
rect 8128 29161 8156 29260
rect 8297 29223 8355 29229
rect 8297 29189 8309 29223
rect 8343 29220 8355 29223
rect 8343 29192 9352 29220
rect 8343 29189 8355 29192
rect 8297 29183 8355 29189
rect 9324 29164 9352 29192
rect 8113 29155 8171 29161
rect 8113 29121 8125 29155
rect 8159 29121 8171 29155
rect 8113 29115 8171 29121
rect 8389 29155 8447 29161
rect 8389 29121 8401 29155
rect 8435 29152 8447 29155
rect 9033 29155 9091 29161
rect 9033 29152 9045 29155
rect 8435 29124 9045 29152
rect 8435 29121 8447 29124
rect 8389 29115 8447 29121
rect 9033 29121 9045 29124
rect 9079 29121 9091 29155
rect 9306 29152 9312 29164
rect 9267 29124 9312 29152
rect 9033 29115 9091 29121
rect 9048 29084 9076 29115
rect 9306 29112 9312 29124
rect 9364 29112 9370 29164
rect 9508 29161 9536 29260
rect 12894 29248 12900 29300
rect 12952 29248 12958 29300
rect 14550 29288 14556 29300
rect 14511 29260 14556 29288
rect 14550 29248 14556 29260
rect 14608 29248 14614 29300
rect 14918 29248 14924 29300
rect 14976 29288 14982 29300
rect 20254 29288 20260 29300
rect 14976 29260 17816 29288
rect 20215 29260 20260 29288
rect 14976 29248 14982 29260
rect 12912 29220 12940 29248
rect 12544 29192 12940 29220
rect 9493 29155 9551 29161
rect 9493 29121 9505 29155
rect 9539 29152 9551 29155
rect 11054 29152 11060 29164
rect 9539 29124 11060 29152
rect 9539 29121 9551 29124
rect 9493 29115 9551 29121
rect 11054 29112 11060 29124
rect 11112 29112 11118 29164
rect 11790 29152 11796 29164
rect 11751 29124 11796 29152
rect 11790 29112 11796 29124
rect 11848 29112 11854 29164
rect 12544 29161 12572 29192
rect 15102 29180 15108 29232
rect 15160 29220 15166 29232
rect 17788 29229 17816 29260
rect 20254 29248 20260 29260
rect 20312 29248 20318 29300
rect 21726 29248 21732 29300
rect 21784 29288 21790 29300
rect 22097 29291 22155 29297
rect 22097 29288 22109 29291
rect 21784 29260 22109 29288
rect 21784 29248 21790 29260
rect 22097 29257 22109 29260
rect 22143 29257 22155 29291
rect 25314 29288 25320 29300
rect 22097 29251 22155 29257
rect 25240 29260 25320 29288
rect 15381 29223 15439 29229
rect 15381 29220 15393 29223
rect 15160 29192 15393 29220
rect 15160 29180 15166 29192
rect 15381 29189 15393 29192
rect 15427 29189 15439 29223
rect 15381 29183 15439 29189
rect 17773 29223 17831 29229
rect 17773 29189 17785 29223
rect 17819 29189 17831 29223
rect 19334 29220 19340 29232
rect 17773 29183 17831 29189
rect 19260 29192 19340 29220
rect 12529 29155 12587 29161
rect 12529 29121 12541 29155
rect 12575 29121 12587 29155
rect 12529 29115 12587 29121
rect 12618 29112 12624 29164
rect 12676 29152 12682 29164
rect 12676 29124 12721 29152
rect 12676 29112 12682 29124
rect 12802 29112 12808 29164
rect 12860 29152 12866 29164
rect 12897 29155 12955 29161
rect 12897 29152 12909 29155
rect 12860 29124 12909 29152
rect 12860 29112 12866 29124
rect 12897 29121 12909 29124
rect 12943 29121 12955 29155
rect 12897 29115 12955 29121
rect 13173 29155 13231 29161
rect 13173 29121 13185 29155
rect 13219 29152 13231 29155
rect 13354 29152 13360 29164
rect 13219 29124 13360 29152
rect 13219 29121 13231 29124
rect 13173 29115 13231 29121
rect 13354 29112 13360 29124
rect 13412 29112 13418 29164
rect 14737 29155 14795 29161
rect 14737 29121 14749 29155
rect 14783 29152 14795 29155
rect 15120 29152 15148 29180
rect 15562 29152 15568 29164
rect 14783 29124 15148 29152
rect 15523 29124 15568 29152
rect 14783 29121 14795 29124
rect 14737 29115 14795 29121
rect 15562 29112 15568 29124
rect 15620 29112 15626 29164
rect 15746 29152 15752 29164
rect 15707 29124 15752 29152
rect 15746 29112 15752 29124
rect 15804 29112 15810 29164
rect 19260 29161 19288 29192
rect 19334 29180 19340 29192
rect 19392 29180 19398 29232
rect 20456 29192 21496 29220
rect 20456 29164 20484 29192
rect 19245 29155 19303 29161
rect 19245 29121 19257 29155
rect 19291 29121 19303 29155
rect 19426 29152 19432 29164
rect 19387 29124 19432 29152
rect 19245 29115 19303 29121
rect 19426 29112 19432 29124
rect 19484 29112 19490 29164
rect 20438 29152 20444 29164
rect 20399 29124 20444 29152
rect 20438 29112 20444 29124
rect 20496 29112 20502 29164
rect 20533 29155 20591 29161
rect 20533 29121 20545 29155
rect 20579 29121 20591 29155
rect 20714 29152 20720 29164
rect 20675 29124 20720 29152
rect 20533 29115 20591 29121
rect 10318 29084 10324 29096
rect 9048 29056 10324 29084
rect 10318 29044 10324 29056
rect 10376 29044 10382 29096
rect 14921 29087 14979 29093
rect 14921 29053 14933 29087
rect 14967 29084 14979 29087
rect 15010 29084 15016 29096
rect 14967 29056 15016 29084
rect 14967 29053 14979 29056
rect 14921 29047 14979 29053
rect 15010 29044 15016 29056
rect 15068 29044 15074 29096
rect 20162 29044 20168 29096
rect 20220 29084 20226 29096
rect 20548 29084 20576 29115
rect 20714 29112 20720 29124
rect 20772 29112 20778 29164
rect 20806 29112 20812 29164
rect 20864 29152 20870 29164
rect 21468 29161 21496 29192
rect 21634 29180 21640 29232
rect 21692 29220 21698 29232
rect 21692 29192 22600 29220
rect 21692 29180 21698 29192
rect 21269 29155 21327 29161
rect 21269 29152 21281 29155
rect 20864 29124 20909 29152
rect 21008 29124 21281 29152
rect 20864 29112 20870 29124
rect 21008 29084 21036 29124
rect 21269 29121 21281 29124
rect 21315 29121 21327 29155
rect 21269 29115 21327 29121
rect 21453 29155 21511 29161
rect 21453 29121 21465 29155
rect 21499 29121 21511 29155
rect 22278 29152 22284 29164
rect 22239 29124 22284 29152
rect 21453 29115 21511 29121
rect 22278 29112 22284 29124
rect 22336 29112 22342 29164
rect 22572 29161 22600 29192
rect 23474 29180 23480 29232
rect 23532 29220 23538 29232
rect 23661 29223 23719 29229
rect 23661 29220 23673 29223
rect 23532 29192 23673 29220
rect 23532 29180 23538 29192
rect 23661 29189 23673 29192
rect 23707 29220 23719 29223
rect 24670 29220 24676 29232
rect 23707 29192 24676 29220
rect 23707 29189 23719 29192
rect 23661 29183 23719 29189
rect 24670 29180 24676 29192
rect 24728 29180 24734 29232
rect 25240 29229 25268 29260
rect 25314 29248 25320 29260
rect 25372 29248 25378 29300
rect 27522 29288 27528 29300
rect 27483 29260 27528 29288
rect 27522 29248 27528 29260
rect 27580 29248 27586 29300
rect 27614 29248 27620 29300
rect 27672 29288 27678 29300
rect 28258 29288 28264 29300
rect 28316 29297 28322 29300
rect 28316 29291 28335 29297
rect 27672 29260 28264 29288
rect 27672 29248 27678 29260
rect 28258 29248 28264 29260
rect 28323 29257 28335 29291
rect 28316 29251 28335 29257
rect 28445 29291 28503 29297
rect 28445 29257 28457 29291
rect 28491 29288 28503 29291
rect 28902 29288 28908 29300
rect 28491 29260 28908 29288
rect 28491 29257 28503 29260
rect 28445 29251 28503 29257
rect 28316 29248 28322 29251
rect 28902 29248 28908 29260
rect 28960 29248 28966 29300
rect 25225 29223 25283 29229
rect 25225 29189 25237 29223
rect 25271 29189 25283 29223
rect 27982 29220 27988 29232
rect 25225 29183 25283 29189
rect 27448 29192 27988 29220
rect 27448 29164 27476 29192
rect 27982 29180 27988 29192
rect 28040 29180 28046 29232
rect 28074 29180 28080 29232
rect 28132 29220 28138 29232
rect 28132 29192 28177 29220
rect 28132 29180 28138 29192
rect 22557 29155 22615 29161
rect 22557 29121 22569 29155
rect 22603 29121 22615 29155
rect 22738 29152 22744 29164
rect 22699 29124 22744 29152
rect 22557 29115 22615 29121
rect 22738 29112 22744 29124
rect 22796 29112 22802 29164
rect 23566 29112 23572 29164
rect 23624 29152 23630 29164
rect 25317 29155 25375 29161
rect 25317 29152 25329 29155
rect 23624 29124 25329 29152
rect 23624 29112 23630 29124
rect 25317 29121 25329 29124
rect 25363 29121 25375 29155
rect 25317 29115 25375 29121
rect 25593 29155 25651 29161
rect 25593 29121 25605 29155
rect 25639 29152 25651 29155
rect 25774 29152 25780 29164
rect 25639 29124 25780 29152
rect 25639 29121 25651 29124
rect 25593 29115 25651 29121
rect 25774 29112 25780 29124
rect 25832 29112 25838 29164
rect 27430 29152 27436 29164
rect 27391 29124 27436 29152
rect 27430 29112 27436 29124
rect 27488 29112 27494 29164
rect 27617 29155 27675 29161
rect 27617 29121 27629 29155
rect 27663 29152 27675 29155
rect 28902 29152 28908 29164
rect 27663 29124 28120 29152
rect 28863 29124 28908 29152
rect 27663 29121 27675 29124
rect 27617 29115 27675 29121
rect 20220 29056 21036 29084
rect 20220 29044 20226 29056
rect 21634 29044 21640 29096
rect 21692 29084 21698 29096
rect 22373 29087 22431 29093
rect 22373 29084 22385 29087
rect 21692 29056 22385 29084
rect 21692 29044 21698 29056
rect 22373 29053 22385 29056
rect 22419 29053 22431 29087
rect 22373 29047 22431 29053
rect 21361 29019 21419 29025
rect 21361 28985 21373 29019
rect 21407 29016 21419 29019
rect 21450 29016 21456 29028
rect 21407 28988 21456 29016
rect 21407 28985 21419 28988
rect 21361 28979 21419 28985
rect 21450 28976 21456 28988
rect 21508 28976 21514 29028
rect 22465 29019 22523 29025
rect 22465 28985 22477 29019
rect 22511 29016 22523 29019
rect 23201 29019 23259 29025
rect 23201 29016 23213 29019
rect 22511 28988 23213 29016
rect 22511 28985 22523 28988
rect 22465 28979 22523 28985
rect 23201 28985 23213 28988
rect 23247 28985 23259 29019
rect 23201 28979 23259 28985
rect 23290 28976 23296 29028
rect 23348 29016 23354 29028
rect 23385 29019 23443 29025
rect 23385 29016 23397 29019
rect 23348 28988 23397 29016
rect 23348 28976 23354 28988
rect 23385 28985 23397 28988
rect 23431 29016 23443 29019
rect 27632 29016 27660 29115
rect 23431 28988 27660 29016
rect 27890 28994 27896 29028
rect 23431 28985 23443 28988
rect 23385 28979 23443 28985
rect 27724 28976 27896 28994
rect 27948 28976 27954 29028
rect 28092 29016 28120 29124
rect 28902 29112 28908 29124
rect 28960 29112 28966 29164
rect 29086 29152 29092 29164
rect 29047 29124 29092 29152
rect 29086 29112 29092 29124
rect 29144 29112 29150 29164
rect 28626 29044 28632 29096
rect 28684 29084 28690 29096
rect 29181 29087 29239 29093
rect 29181 29084 29193 29087
rect 28684 29056 29193 29084
rect 28684 29044 28690 29056
rect 29181 29053 29193 29056
rect 29227 29053 29239 29087
rect 29181 29047 29239 29053
rect 30282 29016 30288 29028
rect 28092 28988 30288 29016
rect 30282 28976 30288 28988
rect 30340 28976 30346 29028
rect 27724 28966 27936 28976
rect 7742 28908 7748 28960
rect 7800 28948 7806 28960
rect 7929 28951 7987 28957
rect 7929 28948 7941 28951
rect 7800 28920 7941 28948
rect 7800 28908 7806 28920
rect 7929 28917 7941 28920
rect 7975 28917 7987 28951
rect 7929 28911 7987 28917
rect 9306 28908 9312 28960
rect 9364 28948 9370 28960
rect 9401 28951 9459 28957
rect 9401 28948 9413 28951
rect 9364 28920 9413 28948
rect 9364 28908 9370 28920
rect 9401 28917 9413 28920
rect 9447 28917 9459 28951
rect 9401 28911 9459 28917
rect 10410 28908 10416 28960
rect 10468 28948 10474 28960
rect 11793 28951 11851 28957
rect 11793 28948 11805 28951
rect 10468 28920 11805 28948
rect 10468 28908 10474 28920
rect 11793 28917 11805 28920
rect 11839 28917 11851 28951
rect 11793 28911 11851 28917
rect 27522 28908 27528 28960
rect 27580 28948 27586 28960
rect 27724 28948 27752 28966
rect 27580 28920 27752 28948
rect 28261 28951 28319 28957
rect 27580 28908 27586 28920
rect 28261 28917 28273 28951
rect 28307 28948 28319 28951
rect 28810 28948 28816 28960
rect 28307 28920 28816 28948
rect 28307 28917 28319 28920
rect 28261 28911 28319 28917
rect 28810 28908 28816 28920
rect 28868 28908 28874 28960
rect 1104 28858 34868 28880
rect 1104 28806 5170 28858
rect 5222 28806 5234 28858
rect 5286 28806 5298 28858
rect 5350 28806 5362 28858
rect 5414 28806 5426 28858
rect 5478 28806 13611 28858
rect 13663 28806 13675 28858
rect 13727 28806 13739 28858
rect 13791 28806 13803 28858
rect 13855 28806 13867 28858
rect 13919 28806 22052 28858
rect 22104 28806 22116 28858
rect 22168 28806 22180 28858
rect 22232 28806 22244 28858
rect 22296 28806 22308 28858
rect 22360 28806 30493 28858
rect 30545 28806 30557 28858
rect 30609 28806 30621 28858
rect 30673 28806 30685 28858
rect 30737 28806 30749 28858
rect 30801 28806 34868 28858
rect 1104 28784 34868 28806
rect 13354 28704 13360 28756
rect 13412 28744 13418 28756
rect 21082 28744 21088 28756
rect 13412 28716 15240 28744
rect 21043 28716 21088 28744
rect 13412 28704 13418 28716
rect 10965 28679 11023 28685
rect 10965 28645 10977 28679
rect 11011 28676 11023 28679
rect 11054 28676 11060 28688
rect 11011 28648 11060 28676
rect 11011 28645 11023 28648
rect 10965 28639 11023 28645
rect 11054 28636 11060 28648
rect 11112 28636 11118 28688
rect 15212 28685 15240 28716
rect 21082 28704 21088 28716
rect 21140 28704 21146 28756
rect 28810 28704 28816 28756
rect 28868 28744 28874 28756
rect 28905 28747 28963 28753
rect 28905 28744 28917 28747
rect 28868 28716 28917 28744
rect 28868 28704 28874 28716
rect 28905 28713 28917 28716
rect 28951 28713 28963 28747
rect 28905 28707 28963 28713
rect 15197 28679 15255 28685
rect 15197 28645 15209 28679
rect 15243 28645 15255 28679
rect 20806 28676 20812 28688
rect 15197 28639 15255 28645
rect 20640 28648 20812 28676
rect 11609 28611 11667 28617
rect 11609 28577 11621 28611
rect 11655 28608 11667 28611
rect 11790 28608 11796 28620
rect 11655 28580 11796 28608
rect 11655 28577 11667 28580
rect 11609 28571 11667 28577
rect 11790 28568 11796 28580
rect 11848 28608 11854 28620
rect 12526 28608 12532 28620
rect 11848 28580 12532 28608
rect 11848 28568 11854 28580
rect 12526 28568 12532 28580
rect 12584 28608 12590 28620
rect 13173 28611 13231 28617
rect 13173 28608 13185 28611
rect 12584 28580 13185 28608
rect 12584 28568 12590 28580
rect 13173 28577 13185 28580
rect 13219 28577 13231 28611
rect 13354 28608 13360 28620
rect 13315 28580 13360 28608
rect 13173 28571 13231 28577
rect 13354 28568 13360 28580
rect 13412 28568 13418 28620
rect 15010 28568 15016 28620
rect 15068 28608 15074 28620
rect 15930 28608 15936 28620
rect 15068 28580 15936 28608
rect 15068 28568 15074 28580
rect 15930 28568 15936 28580
rect 15988 28608 15994 28620
rect 20073 28611 20131 28617
rect 15988 28580 19748 28608
rect 15988 28568 15994 28580
rect 19720 28552 19748 28580
rect 20073 28577 20085 28611
rect 20119 28608 20131 28611
rect 20640 28608 20668 28648
rect 20806 28636 20812 28648
rect 20864 28676 20870 28688
rect 21634 28676 21640 28688
rect 20864 28648 21640 28676
rect 20864 28636 20870 28648
rect 21634 28636 21640 28648
rect 21692 28636 21698 28688
rect 21266 28608 21272 28620
rect 20119 28580 20668 28608
rect 20119 28577 20131 28580
rect 20073 28571 20131 28577
rect 7742 28500 7748 28552
rect 7800 28540 7806 28552
rect 9030 28540 9036 28552
rect 7800 28512 9036 28540
rect 7800 28500 7806 28512
rect 9030 28500 9036 28512
rect 9088 28540 9094 28552
rect 9125 28543 9183 28549
rect 9125 28540 9137 28543
rect 9088 28512 9137 28540
rect 9088 28500 9094 28512
rect 9125 28509 9137 28512
rect 9171 28509 9183 28543
rect 9306 28540 9312 28552
rect 9267 28512 9312 28540
rect 9125 28503 9183 28509
rect 9306 28500 9312 28512
rect 9364 28500 9370 28552
rect 10962 28500 10968 28552
rect 11020 28540 11026 28552
rect 11241 28543 11299 28549
rect 11241 28540 11253 28543
rect 11020 28512 11253 28540
rect 11020 28500 11026 28512
rect 11241 28509 11253 28512
rect 11287 28509 11299 28543
rect 11241 28503 11299 28509
rect 12069 28543 12127 28549
rect 12069 28509 12081 28543
rect 12115 28509 12127 28543
rect 12069 28503 12127 28509
rect 12345 28543 12403 28549
rect 12345 28509 12357 28543
rect 12391 28540 12403 28543
rect 12802 28540 12808 28552
rect 12391 28512 12808 28540
rect 12391 28509 12403 28512
rect 12345 28503 12403 28509
rect 12084 28472 12112 28503
rect 12802 28500 12808 28512
rect 12860 28500 12866 28552
rect 12986 28500 12992 28552
rect 13044 28540 13050 28552
rect 13081 28543 13139 28549
rect 13081 28540 13093 28543
rect 13044 28512 13093 28540
rect 13044 28500 13050 28512
rect 13081 28509 13093 28512
rect 13127 28509 13139 28543
rect 13081 28503 13139 28509
rect 13262 28500 13268 28552
rect 13320 28540 13326 28552
rect 14550 28540 14556 28552
rect 13320 28512 13365 28540
rect 14511 28512 14556 28540
rect 13320 28500 13326 28512
rect 14550 28500 14556 28512
rect 14608 28500 14614 28552
rect 14921 28543 14979 28549
rect 14921 28509 14933 28543
rect 14967 28540 14979 28543
rect 15102 28540 15108 28552
rect 14967 28512 15108 28540
rect 14967 28509 14979 28512
rect 14921 28503 14979 28509
rect 15102 28500 15108 28512
rect 15160 28500 15166 28552
rect 15378 28540 15384 28552
rect 15339 28512 15384 28540
rect 15378 28500 15384 28512
rect 15436 28500 15442 28552
rect 15470 28500 15476 28552
rect 15528 28540 15534 28552
rect 16301 28543 16359 28549
rect 16301 28540 16313 28543
rect 15528 28512 16313 28540
rect 15528 28500 15534 28512
rect 16301 28509 16313 28512
rect 16347 28509 16359 28543
rect 19702 28540 19708 28552
rect 19663 28512 19708 28540
rect 16301 28503 16359 28509
rect 19702 28500 19708 28512
rect 19760 28500 19766 28552
rect 19886 28540 19892 28552
rect 19847 28512 19892 28540
rect 19886 28500 19892 28512
rect 19944 28500 19950 28552
rect 20640 28549 20668 28580
rect 20824 28580 21272 28608
rect 20824 28549 20852 28580
rect 21266 28568 21272 28580
rect 21324 28568 21330 28620
rect 26237 28611 26295 28617
rect 26237 28577 26249 28611
rect 26283 28608 26295 28611
rect 27154 28608 27160 28620
rect 26283 28580 27160 28608
rect 26283 28577 26295 28580
rect 26237 28571 26295 28577
rect 27154 28568 27160 28580
rect 27212 28568 27218 28620
rect 27614 28568 27620 28620
rect 27672 28568 27678 28620
rect 20533 28543 20591 28549
rect 20533 28509 20545 28543
rect 20579 28509 20591 28543
rect 20533 28503 20591 28509
rect 20625 28543 20683 28549
rect 20625 28509 20637 28543
rect 20671 28509 20683 28543
rect 20809 28543 20867 28549
rect 20809 28540 20821 28543
rect 20625 28503 20683 28509
rect 20732 28512 20821 28540
rect 13354 28472 13360 28484
rect 12084 28444 13360 28472
rect 13354 28432 13360 28444
rect 13412 28432 13418 28484
rect 15746 28432 15752 28484
rect 15804 28472 15810 28484
rect 16669 28475 16727 28481
rect 16669 28472 16681 28475
rect 15804 28444 16681 28472
rect 15804 28432 15810 28444
rect 16669 28441 16681 28444
rect 16715 28472 16727 28475
rect 19242 28472 19248 28484
rect 16715 28444 19248 28472
rect 16715 28441 16727 28444
rect 16669 28435 16727 28441
rect 19242 28432 19248 28444
rect 19300 28432 19306 28484
rect 20548 28416 20576 28503
rect 20732 28484 20760 28512
rect 20809 28509 20821 28512
rect 20855 28509 20867 28543
rect 20809 28503 20867 28509
rect 20901 28543 20959 28549
rect 20901 28509 20913 28543
rect 20947 28540 20959 28543
rect 22830 28540 22836 28552
rect 20947 28512 21588 28540
rect 22743 28512 22836 28540
rect 20947 28509 20959 28512
rect 20901 28503 20959 28509
rect 21560 28484 21588 28512
rect 22830 28500 22836 28512
rect 22888 28540 22894 28552
rect 23290 28540 23296 28552
rect 22888 28512 23296 28540
rect 22888 28500 22894 28512
rect 23290 28500 23296 28512
rect 23348 28500 23354 28552
rect 23385 28543 23443 28549
rect 23385 28509 23397 28543
rect 23431 28540 23443 28543
rect 23474 28540 23480 28552
rect 23431 28512 23480 28540
rect 23431 28509 23443 28512
rect 23385 28503 23443 28509
rect 23474 28500 23480 28512
rect 23532 28500 23538 28552
rect 27890 28540 27896 28552
rect 27738 28512 27896 28540
rect 27890 28500 27896 28512
rect 27948 28500 27954 28552
rect 28994 28540 29000 28552
rect 28955 28512 29000 28540
rect 28994 28500 29000 28512
rect 29052 28500 29058 28552
rect 20714 28432 20720 28484
rect 20772 28432 20778 28484
rect 21542 28432 21548 28484
rect 21600 28472 21606 28484
rect 21600 28444 22494 28472
rect 21600 28432 21606 28444
rect 9214 28404 9220 28416
rect 9175 28376 9220 28404
rect 9214 28364 9220 28376
rect 9272 28364 9278 28416
rect 12894 28404 12900 28416
rect 12855 28376 12900 28404
rect 12894 28364 12900 28376
rect 12952 28364 12958 28416
rect 20530 28404 20536 28416
rect 20443 28376 20536 28404
rect 20530 28364 20536 28376
rect 20588 28404 20594 28416
rect 22738 28404 22744 28416
rect 20588 28376 22744 28404
rect 20588 28364 20594 28376
rect 22738 28364 22744 28376
rect 22796 28364 22802 28416
rect 27246 28404 27252 28416
rect 27207 28376 27252 28404
rect 27246 28364 27252 28376
rect 27304 28364 27310 28416
rect 1104 28314 35027 28336
rect 1104 28262 9390 28314
rect 9442 28262 9454 28314
rect 9506 28262 9518 28314
rect 9570 28262 9582 28314
rect 9634 28262 9646 28314
rect 9698 28262 17831 28314
rect 17883 28262 17895 28314
rect 17947 28262 17959 28314
rect 18011 28262 18023 28314
rect 18075 28262 18087 28314
rect 18139 28262 26272 28314
rect 26324 28262 26336 28314
rect 26388 28262 26400 28314
rect 26452 28262 26464 28314
rect 26516 28262 26528 28314
rect 26580 28262 34713 28314
rect 34765 28262 34777 28314
rect 34829 28262 34841 28314
rect 34893 28262 34905 28314
rect 34957 28262 34969 28314
rect 35021 28262 35027 28314
rect 1104 28240 35027 28262
rect 9858 28200 9864 28212
rect 8864 28172 9864 28200
rect 7742 28064 7748 28076
rect 7703 28036 7748 28064
rect 7742 28024 7748 28036
rect 7800 28024 7806 28076
rect 7837 28067 7895 28073
rect 7837 28033 7849 28067
rect 7883 28064 7895 28067
rect 8021 28067 8079 28073
rect 7883 28036 7972 28064
rect 7883 28033 7895 28036
rect 7837 28027 7895 28033
rect 7944 27928 7972 28036
rect 8021 28033 8033 28067
rect 8067 28033 8079 28067
rect 8754 28064 8760 28076
rect 8715 28036 8760 28064
rect 8021 28027 8079 28033
rect 8036 27996 8064 28027
rect 8754 28024 8760 28036
rect 8812 28024 8818 28076
rect 8864 28073 8892 28172
rect 9858 28160 9864 28172
rect 9916 28160 9922 28212
rect 12986 28200 12992 28212
rect 12406 28172 12992 28200
rect 10962 28092 10968 28144
rect 11020 28132 11026 28144
rect 12406 28132 12434 28172
rect 12986 28160 12992 28172
rect 13044 28160 13050 28212
rect 13354 28160 13360 28212
rect 13412 28160 13418 28212
rect 15378 28200 15384 28212
rect 15339 28172 15384 28200
rect 15378 28160 15384 28172
rect 15436 28160 15442 28212
rect 22370 28200 22376 28212
rect 22331 28172 22376 28200
rect 22370 28160 22376 28172
rect 22428 28160 22434 28212
rect 13372 28132 13400 28160
rect 15010 28132 15016 28144
rect 11020 28104 12434 28132
rect 12912 28104 13400 28132
rect 14016 28104 15016 28132
rect 11020 28092 11026 28104
rect 8849 28067 8907 28073
rect 8849 28033 8861 28067
rect 8895 28033 8907 28067
rect 9030 28064 9036 28076
rect 8991 28036 9036 28064
rect 8849 28027 8907 28033
rect 8864 27996 8892 28027
rect 9030 28024 9036 28036
rect 9088 28024 9094 28076
rect 12176 28073 12204 28104
rect 12161 28067 12219 28073
rect 12161 28033 12173 28067
rect 12207 28033 12219 28067
rect 12526 28064 12532 28076
rect 12487 28036 12532 28064
rect 12161 28027 12219 28033
rect 12526 28024 12532 28036
rect 12584 28024 12590 28076
rect 12912 28073 12940 28104
rect 14016 28076 14044 28104
rect 15010 28092 15016 28104
rect 15068 28092 15074 28144
rect 15562 28092 15568 28144
rect 15620 28132 15626 28144
rect 15933 28135 15991 28141
rect 15933 28132 15945 28135
rect 15620 28104 15945 28132
rect 15620 28092 15626 28104
rect 15933 28101 15945 28104
rect 15979 28132 15991 28135
rect 16022 28132 16028 28144
rect 15979 28104 16028 28132
rect 15979 28101 15991 28104
rect 15933 28095 15991 28101
rect 16022 28092 16028 28104
rect 16080 28092 16086 28144
rect 19337 28135 19395 28141
rect 19337 28101 19349 28135
rect 19383 28132 19395 28135
rect 19886 28132 19892 28144
rect 19383 28104 19892 28132
rect 19383 28101 19395 28104
rect 19337 28095 19395 28101
rect 19886 28092 19892 28104
rect 19944 28132 19950 28144
rect 20625 28135 20683 28141
rect 19944 28104 20300 28132
rect 19944 28092 19950 28104
rect 12897 28067 12955 28073
rect 12897 28033 12909 28067
rect 12943 28033 12955 28067
rect 12897 28027 12955 28033
rect 13262 28024 13268 28076
rect 13320 28064 13326 28076
rect 13357 28067 13415 28073
rect 13357 28064 13369 28067
rect 13320 28036 13369 28064
rect 13320 28024 13326 28036
rect 13357 28033 13369 28036
rect 13403 28064 13415 28067
rect 13817 28067 13875 28073
rect 13817 28064 13829 28067
rect 13403 28036 13829 28064
rect 13403 28033 13415 28036
rect 13357 28027 13415 28033
rect 13817 28033 13829 28036
rect 13863 28033 13875 28067
rect 13817 28027 13875 28033
rect 13998 28024 14004 28076
rect 14056 28064 14062 28076
rect 14185 28067 14243 28073
rect 14056 28036 14149 28064
rect 14056 28024 14062 28036
rect 14185 28033 14197 28067
rect 14231 28064 14243 28067
rect 14274 28064 14280 28076
rect 14231 28036 14280 28064
rect 14231 28033 14243 28036
rect 14185 28027 14243 28033
rect 14274 28024 14280 28036
rect 14332 28024 14338 28076
rect 15381 28067 15439 28073
rect 15381 28033 15393 28067
rect 15427 28064 15439 28067
rect 15470 28064 15476 28076
rect 15427 28036 15476 28064
rect 15427 28033 15439 28036
rect 15381 28027 15439 28033
rect 15470 28024 15476 28036
rect 15528 28024 15534 28076
rect 19242 28064 19248 28076
rect 19203 28036 19248 28064
rect 19242 28024 19248 28036
rect 19300 28024 19306 28076
rect 20272 28073 20300 28104
rect 20625 28101 20637 28135
rect 20671 28132 20683 28135
rect 20714 28132 20720 28144
rect 20671 28104 20720 28132
rect 20671 28101 20683 28104
rect 20625 28095 20683 28101
rect 20714 28092 20720 28104
rect 20772 28092 20778 28144
rect 22830 28132 22836 28144
rect 22791 28104 22836 28132
rect 22830 28092 22836 28104
rect 22888 28092 22894 28144
rect 19429 28067 19487 28073
rect 19429 28033 19441 28067
rect 19475 28033 19487 28067
rect 19429 28027 19487 28033
rect 20257 28067 20315 28073
rect 20257 28033 20269 28067
rect 20303 28033 20315 28067
rect 20257 28027 20315 28033
rect 20533 28067 20591 28073
rect 20533 28033 20545 28067
rect 20579 28064 20591 28067
rect 24670 28064 24676 28076
rect 20579 28036 24676 28064
rect 20579 28033 20591 28036
rect 20533 28027 20591 28033
rect 8036 27968 8892 27996
rect 8941 27999 8999 28005
rect 8941 27965 8953 27999
rect 8987 27996 8999 27999
rect 9306 27996 9312 28008
rect 8987 27968 9312 27996
rect 8987 27965 8999 27968
rect 8941 27959 8999 27965
rect 8956 27928 8984 27959
rect 9306 27956 9312 27968
rect 9364 27956 9370 28008
rect 12434 27956 12440 28008
rect 12492 27996 12498 28008
rect 12492 27968 12537 27996
rect 12492 27956 12498 27968
rect 14550 27956 14556 28008
rect 14608 27996 14614 28008
rect 15289 27999 15347 28005
rect 15289 27996 15301 27999
rect 14608 27968 15301 27996
rect 14608 27956 14614 27968
rect 15289 27965 15301 27968
rect 15335 27965 15347 27999
rect 15289 27959 15347 27965
rect 19334 27956 19340 28008
rect 19392 27996 19398 28008
rect 19444 27996 19472 28027
rect 24670 28024 24676 28036
rect 24728 28024 24734 28076
rect 25038 28064 25044 28076
rect 24999 28036 25044 28064
rect 25038 28024 25044 28036
rect 25096 28024 25102 28076
rect 25222 28024 25228 28076
rect 25280 28064 25286 28076
rect 25685 28067 25743 28073
rect 25685 28064 25697 28067
rect 25280 28036 25697 28064
rect 25280 28024 25286 28036
rect 25685 28033 25697 28036
rect 25731 28033 25743 28067
rect 25685 28027 25743 28033
rect 27062 28024 27068 28076
rect 27120 28064 27126 28076
rect 27249 28067 27307 28073
rect 27249 28064 27261 28067
rect 27120 28036 27261 28064
rect 27120 28024 27126 28036
rect 27249 28033 27261 28036
rect 27295 28033 27307 28067
rect 27249 28027 27307 28033
rect 27525 28067 27583 28073
rect 27525 28033 27537 28067
rect 27571 28064 27583 28067
rect 27706 28064 27712 28076
rect 27571 28036 27712 28064
rect 27571 28033 27583 28036
rect 27525 28027 27583 28033
rect 27706 28024 27712 28036
rect 27764 28024 27770 28076
rect 29270 28024 29276 28076
rect 29328 28064 29334 28076
rect 30101 28067 30159 28073
rect 30101 28064 30113 28067
rect 29328 28036 30113 28064
rect 29328 28024 29334 28036
rect 30101 28033 30113 28036
rect 30147 28033 30159 28067
rect 30282 28064 30288 28076
rect 30243 28036 30288 28064
rect 30101 28027 30159 28033
rect 30282 28024 30288 28036
rect 30340 28024 30346 28076
rect 30377 28067 30435 28073
rect 30377 28033 30389 28067
rect 30423 28064 30435 28067
rect 32306 28064 32312 28076
rect 30423 28036 32312 28064
rect 30423 28033 30435 28036
rect 30377 28027 30435 28033
rect 32306 28024 32312 28036
rect 32364 28024 32370 28076
rect 19392 27968 19472 27996
rect 19392 27956 19398 27968
rect 25130 27956 25136 28008
rect 25188 27956 25194 28008
rect 25774 27996 25780 28008
rect 25735 27968 25780 27996
rect 25774 27956 25780 27968
rect 25832 27956 25838 28008
rect 26234 27956 26240 28008
rect 26292 27996 26298 28008
rect 27157 27999 27215 28005
rect 27157 27996 27169 27999
rect 26292 27968 27169 27996
rect 26292 27956 26298 27968
rect 27157 27965 27169 27968
rect 27203 27965 27215 27999
rect 27157 27959 27215 27965
rect 7944 27900 8984 27928
rect 12986 27888 12992 27940
rect 13044 27928 13050 27940
rect 15378 27928 15384 27940
rect 13044 27900 15384 27928
rect 13044 27888 13050 27900
rect 15378 27888 15384 27900
rect 15436 27888 15442 27940
rect 22557 27931 22615 27937
rect 22557 27897 22569 27931
rect 22603 27928 22615 27931
rect 23474 27928 23480 27940
rect 22603 27900 23480 27928
rect 22603 27897 22615 27900
rect 22557 27891 22615 27897
rect 23474 27888 23480 27900
rect 23532 27888 23538 27940
rect 24857 27931 24915 27937
rect 24857 27897 24869 27931
rect 24903 27928 24915 27931
rect 25866 27928 25872 27940
rect 24903 27900 25872 27928
rect 24903 27897 24915 27900
rect 24857 27891 24915 27897
rect 25866 27888 25872 27900
rect 25924 27888 25930 27940
rect 8205 27863 8263 27869
rect 8205 27829 8217 27863
rect 8251 27860 8263 27863
rect 9122 27860 9128 27872
rect 8251 27832 9128 27860
rect 8251 27829 8263 27832
rect 8205 27823 8263 27829
rect 9122 27820 9128 27832
rect 9180 27820 9186 27872
rect 9217 27863 9275 27869
rect 9217 27829 9229 27863
rect 9263 27860 9275 27863
rect 9306 27860 9312 27872
rect 9263 27832 9312 27860
rect 9263 27829 9275 27832
rect 9217 27823 9275 27829
rect 9306 27820 9312 27832
rect 9364 27860 9370 27872
rect 9582 27860 9588 27872
rect 9364 27832 9588 27860
rect 9364 27820 9370 27832
rect 9582 27820 9588 27832
rect 9640 27820 9646 27872
rect 19702 27820 19708 27872
rect 19760 27860 19766 27872
rect 26602 27860 26608 27872
rect 19760 27832 26608 27860
rect 19760 27820 19766 27832
rect 26602 27820 26608 27832
rect 26660 27820 26666 27872
rect 29917 27863 29975 27869
rect 29917 27829 29929 27863
rect 29963 27860 29975 27863
rect 30006 27860 30012 27872
rect 29963 27832 30012 27860
rect 29963 27829 29975 27832
rect 29917 27823 29975 27829
rect 30006 27820 30012 27832
rect 30064 27820 30070 27872
rect 1104 27770 34868 27792
rect 1104 27718 5170 27770
rect 5222 27718 5234 27770
rect 5286 27718 5298 27770
rect 5350 27718 5362 27770
rect 5414 27718 5426 27770
rect 5478 27718 13611 27770
rect 13663 27718 13675 27770
rect 13727 27718 13739 27770
rect 13791 27718 13803 27770
rect 13855 27718 13867 27770
rect 13919 27718 22052 27770
rect 22104 27718 22116 27770
rect 22168 27718 22180 27770
rect 22232 27718 22244 27770
rect 22296 27718 22308 27770
rect 22360 27718 30493 27770
rect 30545 27718 30557 27770
rect 30609 27718 30621 27770
rect 30673 27718 30685 27770
rect 30737 27718 30749 27770
rect 30801 27718 34868 27770
rect 1104 27696 34868 27718
rect 16022 27548 16028 27600
rect 16080 27588 16086 27600
rect 16853 27591 16911 27597
rect 16853 27588 16865 27591
rect 16080 27560 16865 27588
rect 16080 27548 16086 27560
rect 16853 27557 16865 27560
rect 16899 27557 16911 27591
rect 16853 27551 16911 27557
rect 24578 27548 24584 27600
rect 24636 27588 24642 27600
rect 25225 27591 25283 27597
rect 25225 27588 25237 27591
rect 24636 27560 25237 27588
rect 24636 27548 24642 27560
rect 25225 27557 25237 27560
rect 25271 27557 25283 27591
rect 27890 27588 27896 27600
rect 27851 27560 27896 27588
rect 25225 27551 25283 27557
rect 27890 27548 27896 27560
rect 27948 27548 27954 27600
rect 12526 27480 12532 27532
rect 12584 27520 12590 27532
rect 12805 27523 12863 27529
rect 12805 27520 12817 27523
rect 12584 27492 12817 27520
rect 12584 27480 12590 27492
rect 12805 27489 12817 27492
rect 12851 27489 12863 27523
rect 12805 27483 12863 27489
rect 13078 27480 13084 27532
rect 13136 27520 13142 27532
rect 14369 27523 14427 27529
rect 14369 27520 14381 27523
rect 13136 27492 14381 27520
rect 13136 27480 13142 27492
rect 14369 27489 14381 27492
rect 14415 27489 14427 27523
rect 22373 27523 22431 27529
rect 22373 27520 22385 27523
rect 14369 27483 14427 27489
rect 22020 27492 22385 27520
rect 9122 27412 9128 27464
rect 9180 27452 9186 27464
rect 9309 27455 9367 27461
rect 9309 27452 9321 27455
rect 9180 27424 9321 27452
rect 9180 27412 9186 27424
rect 9309 27421 9321 27424
rect 9355 27421 9367 27455
rect 9309 27415 9367 27421
rect 9493 27455 9551 27461
rect 9493 27421 9505 27455
rect 9539 27421 9551 27455
rect 9493 27415 9551 27421
rect 9508 27384 9536 27415
rect 9582 27412 9588 27464
rect 9640 27452 9646 27464
rect 9677 27455 9735 27461
rect 9677 27452 9689 27455
rect 9640 27424 9689 27452
rect 9640 27412 9646 27424
rect 9677 27421 9689 27424
rect 9723 27421 9735 27455
rect 9677 27415 9735 27421
rect 13173 27455 13231 27461
rect 13173 27421 13185 27455
rect 13219 27421 13231 27455
rect 13173 27415 13231 27421
rect 13357 27455 13415 27461
rect 13357 27421 13369 27455
rect 13403 27452 13415 27455
rect 13814 27452 13820 27464
rect 13403 27424 13820 27452
rect 13403 27421 13415 27424
rect 13357 27415 13415 27421
rect 9766 27384 9772 27396
rect 9508 27356 9772 27384
rect 9766 27344 9772 27356
rect 9824 27344 9830 27396
rect 10137 27387 10195 27393
rect 10137 27353 10149 27387
rect 10183 27384 10195 27387
rect 12342 27384 12348 27396
rect 10183 27356 12348 27384
rect 10183 27353 10195 27356
rect 10137 27347 10195 27353
rect 8202 27276 8208 27328
rect 8260 27316 8266 27328
rect 10152 27316 10180 27347
rect 12342 27344 12348 27356
rect 12400 27344 12406 27396
rect 13188 27384 13216 27415
rect 13814 27412 13820 27424
rect 13872 27412 13878 27464
rect 14921 27455 14979 27461
rect 14921 27421 14933 27455
rect 14967 27421 14979 27455
rect 14921 27415 14979 27421
rect 13998 27384 14004 27396
rect 13188 27356 14004 27384
rect 13998 27344 14004 27356
rect 14056 27344 14062 27396
rect 8260 27288 10180 27316
rect 14936 27316 14964 27415
rect 15838 27412 15844 27464
rect 15896 27452 15902 27464
rect 15933 27455 15991 27461
rect 15933 27452 15945 27455
rect 15896 27424 15945 27452
rect 15896 27412 15902 27424
rect 15933 27421 15945 27424
rect 15979 27421 15991 27455
rect 15933 27415 15991 27421
rect 16022 27412 16028 27464
rect 16080 27452 16086 27464
rect 16209 27455 16267 27461
rect 16080 27424 16125 27452
rect 16080 27412 16086 27424
rect 16209 27421 16221 27455
rect 16255 27452 16267 27455
rect 18230 27452 18236 27464
rect 16255 27424 18138 27452
rect 18191 27424 18236 27452
rect 16255 27421 16267 27424
rect 16209 27415 16267 27421
rect 16393 27387 16451 27393
rect 16393 27353 16405 27387
rect 16439 27384 16451 27387
rect 17966 27387 18024 27393
rect 17966 27384 17978 27387
rect 16439 27356 17978 27384
rect 16439 27353 16451 27356
rect 16393 27347 16451 27353
rect 17966 27353 17978 27356
rect 18012 27353 18024 27387
rect 18110 27384 18138 27424
rect 18230 27412 18236 27424
rect 18288 27412 18294 27464
rect 19242 27384 19248 27396
rect 18110 27356 19248 27384
rect 17966 27347 18024 27353
rect 19242 27344 19248 27356
rect 19300 27344 19306 27396
rect 20990 27344 20996 27396
rect 21048 27384 21054 27396
rect 22020 27384 22048 27492
rect 22373 27489 22385 27492
rect 22419 27489 22431 27523
rect 22373 27483 22431 27489
rect 25866 27480 25872 27532
rect 25924 27520 25930 27532
rect 28445 27523 28503 27529
rect 28445 27520 28457 27523
rect 25924 27492 26740 27520
rect 25924 27480 25930 27492
rect 22097 27455 22155 27461
rect 22097 27421 22109 27455
rect 22143 27452 22155 27455
rect 23566 27452 23572 27464
rect 22143 27424 23572 27452
rect 22143 27421 22155 27424
rect 22097 27415 22155 27421
rect 23566 27412 23572 27424
rect 23624 27412 23630 27464
rect 25409 27455 25467 27461
rect 25409 27421 25421 27455
rect 25455 27452 25467 27455
rect 25682 27452 25688 27464
rect 25455 27424 25544 27452
rect 25643 27424 25688 27452
rect 25455 27421 25467 27424
rect 25409 27415 25467 27421
rect 25038 27384 25044 27396
rect 21048 27356 25044 27384
rect 21048 27344 21054 27356
rect 25038 27344 25044 27356
rect 25096 27344 25102 27396
rect 19794 27316 19800 27328
rect 14936 27288 19800 27316
rect 8260 27276 8266 27288
rect 19794 27276 19800 27288
rect 19852 27276 19858 27328
rect 25516 27316 25544 27424
rect 25682 27412 25688 27424
rect 25740 27412 25746 27464
rect 26053 27455 26111 27461
rect 26053 27421 26065 27455
rect 26099 27421 26111 27455
rect 26053 27415 26111 27421
rect 25590 27344 25596 27396
rect 25648 27384 25654 27396
rect 26068 27384 26096 27415
rect 26142 27412 26148 27464
rect 26200 27452 26206 27464
rect 26712 27461 26740 27492
rect 27724 27492 28457 27520
rect 27724 27464 27752 27492
rect 28445 27489 28457 27492
rect 28491 27489 28503 27523
rect 28445 27483 28503 27489
rect 26329 27455 26387 27461
rect 26329 27452 26341 27455
rect 26200 27424 26341 27452
rect 26200 27412 26206 27424
rect 26329 27421 26341 27424
rect 26375 27421 26387 27455
rect 26329 27415 26387 27421
rect 26697 27455 26755 27461
rect 26697 27421 26709 27455
rect 26743 27421 26755 27455
rect 26697 27415 26755 27421
rect 27433 27455 27491 27461
rect 27433 27421 27445 27455
rect 27479 27421 27491 27455
rect 27706 27452 27712 27464
rect 27667 27424 27712 27452
rect 27433 27415 27491 27421
rect 26234 27384 26240 27396
rect 25648 27356 26240 27384
rect 25648 27344 25654 27356
rect 26234 27344 26240 27356
rect 26292 27344 26298 27396
rect 26344 27384 26372 27415
rect 27448 27384 27476 27415
rect 27706 27412 27712 27424
rect 27764 27412 27770 27464
rect 27982 27412 27988 27464
rect 28040 27452 28046 27464
rect 28353 27455 28411 27461
rect 28353 27452 28365 27455
rect 28040 27424 28365 27452
rect 28040 27412 28046 27424
rect 28353 27421 28365 27424
rect 28399 27421 28411 27455
rect 28353 27415 28411 27421
rect 28537 27455 28595 27461
rect 28537 27421 28549 27455
rect 28583 27452 28595 27455
rect 28994 27452 29000 27464
rect 28583 27424 29000 27452
rect 28583 27421 28595 27424
rect 28537 27415 28595 27421
rect 28994 27412 29000 27424
rect 29052 27452 29058 27464
rect 29730 27452 29736 27464
rect 29052 27424 29132 27452
rect 29691 27424 29736 27452
rect 29052 27412 29058 27424
rect 26344 27356 27476 27384
rect 25774 27316 25780 27328
rect 25516 27288 25780 27316
rect 25774 27276 25780 27288
rect 25832 27316 25838 27328
rect 26694 27316 26700 27328
rect 25832 27288 26700 27316
rect 25832 27276 25838 27288
rect 26694 27276 26700 27288
rect 26752 27276 26758 27328
rect 27062 27276 27068 27328
rect 27120 27316 27126 27328
rect 27525 27319 27583 27325
rect 27525 27316 27537 27319
rect 27120 27288 27537 27316
rect 27120 27276 27126 27288
rect 27525 27285 27537 27288
rect 27571 27285 27583 27319
rect 29104 27316 29132 27424
rect 29730 27412 29736 27424
rect 29788 27412 29794 27464
rect 29178 27344 29184 27396
rect 29236 27384 29242 27396
rect 29978 27387 30036 27393
rect 29978 27384 29990 27387
rect 29236 27356 29990 27384
rect 29236 27344 29242 27356
rect 29978 27353 29990 27356
rect 30024 27353 30036 27387
rect 29978 27347 30036 27353
rect 31113 27319 31171 27325
rect 31113 27316 31125 27319
rect 29104 27288 31125 27316
rect 27525 27279 27583 27285
rect 31113 27285 31125 27288
rect 31159 27285 31171 27319
rect 31113 27279 31171 27285
rect 1104 27226 35027 27248
rect 1104 27174 9390 27226
rect 9442 27174 9454 27226
rect 9506 27174 9518 27226
rect 9570 27174 9582 27226
rect 9634 27174 9646 27226
rect 9698 27174 17831 27226
rect 17883 27174 17895 27226
rect 17947 27174 17959 27226
rect 18011 27174 18023 27226
rect 18075 27174 18087 27226
rect 18139 27174 26272 27226
rect 26324 27174 26336 27226
rect 26388 27174 26400 27226
rect 26452 27174 26464 27226
rect 26516 27174 26528 27226
rect 26580 27174 34713 27226
rect 34765 27174 34777 27226
rect 34829 27174 34841 27226
rect 34893 27174 34905 27226
rect 34957 27174 34969 27226
rect 35021 27174 35027 27226
rect 1104 27152 35027 27174
rect 8297 27115 8355 27121
rect 8297 27081 8309 27115
rect 8343 27112 8355 27115
rect 12069 27115 12127 27121
rect 8343 27084 9444 27112
rect 8343 27081 8355 27084
rect 8297 27075 8355 27081
rect 8754 27004 8760 27056
rect 8812 27044 8818 27056
rect 8812 27016 9352 27044
rect 8812 27004 8818 27016
rect 8202 26976 8208 26988
rect 8163 26948 8208 26976
rect 8202 26936 8208 26948
rect 8260 26936 8266 26988
rect 8481 26979 8539 26985
rect 8481 26945 8493 26979
rect 8527 26976 8539 26979
rect 9214 26976 9220 26988
rect 8527 26948 9220 26976
rect 8527 26945 8539 26948
rect 8481 26939 8539 26945
rect 9214 26936 9220 26948
rect 9272 26936 9278 26988
rect 9324 26985 9352 27016
rect 9309 26979 9367 26985
rect 9309 26945 9321 26979
rect 9355 26945 9367 26979
rect 9309 26939 9367 26945
rect 9033 26911 9091 26917
rect 9033 26877 9045 26911
rect 9079 26877 9091 26911
rect 9033 26871 9091 26877
rect 9125 26911 9183 26917
rect 9125 26877 9137 26911
rect 9171 26908 9183 26911
rect 9416 26908 9444 27084
rect 12069 27081 12081 27115
rect 12115 27112 12127 27115
rect 12894 27112 12900 27124
rect 12115 27084 12900 27112
rect 12115 27081 12127 27084
rect 12069 27075 12127 27081
rect 12894 27072 12900 27084
rect 12952 27072 12958 27124
rect 18230 27072 18236 27124
rect 18288 27112 18294 27124
rect 19521 27115 19579 27121
rect 19521 27112 19533 27115
rect 18288 27084 19533 27112
rect 18288 27072 18294 27084
rect 19521 27081 19533 27084
rect 19567 27081 19579 27115
rect 19521 27075 19579 27081
rect 20809 27115 20867 27121
rect 20809 27081 20821 27115
rect 20855 27112 20867 27115
rect 20990 27112 20996 27124
rect 20855 27084 20996 27112
rect 20855 27081 20867 27084
rect 20809 27075 20867 27081
rect 20990 27072 20996 27084
rect 21048 27072 21054 27124
rect 30282 27072 30288 27124
rect 30340 27112 30346 27124
rect 31113 27115 31171 27121
rect 31113 27112 31125 27115
rect 30340 27084 31125 27112
rect 30340 27072 30346 27084
rect 31113 27081 31125 27084
rect 31159 27081 31171 27115
rect 31113 27075 31171 27081
rect 13078 27044 13084 27056
rect 11900 27016 13084 27044
rect 11900 26985 11928 27016
rect 13078 27004 13084 27016
rect 13136 27004 13142 27056
rect 13814 27004 13820 27056
rect 13872 27044 13878 27056
rect 14274 27044 14280 27056
rect 13872 27016 14280 27044
rect 13872 27004 13878 27016
rect 14274 27004 14280 27016
rect 14332 27044 14338 27056
rect 15473 27047 15531 27053
rect 15473 27044 15485 27047
rect 14332 27016 15485 27044
rect 14332 27004 14338 27016
rect 15473 27013 15485 27016
rect 15519 27013 15531 27047
rect 15473 27007 15531 27013
rect 19794 27004 19800 27056
rect 19852 27044 19858 27056
rect 26142 27044 26148 27056
rect 19852 27016 22140 27044
rect 19852 27004 19858 27016
rect 11885 26979 11943 26985
rect 11885 26945 11897 26979
rect 11931 26945 11943 26979
rect 11885 26939 11943 26945
rect 12161 26979 12219 26985
rect 12161 26945 12173 26979
rect 12207 26976 12219 26979
rect 12434 26976 12440 26988
rect 12207 26948 12440 26976
rect 12207 26945 12219 26948
rect 12161 26939 12219 26945
rect 12434 26936 12440 26948
rect 12492 26936 12498 26988
rect 13096 26976 13124 27004
rect 13633 26979 13691 26985
rect 13633 26976 13645 26979
rect 13096 26948 13645 26976
rect 13633 26945 13645 26948
rect 13679 26945 13691 26979
rect 15654 26976 15660 26988
rect 15615 26948 15660 26976
rect 13633 26939 13691 26945
rect 15654 26936 15660 26948
rect 15712 26936 15718 26988
rect 15746 26936 15752 26988
rect 15804 26976 15810 26988
rect 18233 26979 18291 26985
rect 15804 26948 15849 26976
rect 15804 26936 15810 26948
rect 18233 26945 18245 26979
rect 18279 26976 18291 26979
rect 18322 26976 18328 26988
rect 18279 26948 18328 26976
rect 18279 26945 18291 26948
rect 18233 26939 18291 26945
rect 18322 26936 18328 26948
rect 18380 26936 18386 26988
rect 20717 26979 20775 26985
rect 20717 26945 20729 26979
rect 20763 26945 20775 26979
rect 20990 26976 20996 26988
rect 20951 26948 20996 26976
rect 20717 26939 20775 26945
rect 10686 26908 10692 26920
rect 9171 26880 10692 26908
rect 9171 26877 9183 26880
rect 9125 26871 9183 26877
rect 8481 26843 8539 26849
rect 8481 26809 8493 26843
rect 8527 26840 8539 26843
rect 9048 26840 9076 26871
rect 10686 26868 10692 26880
rect 10744 26868 10750 26920
rect 12618 26868 12624 26920
rect 12676 26908 12682 26920
rect 13725 26911 13783 26917
rect 13725 26908 13737 26911
rect 12676 26880 13737 26908
rect 12676 26868 12682 26880
rect 13725 26877 13737 26880
rect 13771 26908 13783 26911
rect 20530 26908 20536 26920
rect 13771 26880 20536 26908
rect 13771 26877 13783 26880
rect 13725 26871 13783 26877
rect 20530 26868 20536 26880
rect 20588 26868 20594 26920
rect 8527 26812 9076 26840
rect 20732 26840 20760 26939
rect 20990 26936 20996 26948
rect 21048 26936 21054 26988
rect 22112 26985 22140 27016
rect 25700 27016 26148 27044
rect 22097 26979 22155 26985
rect 22097 26945 22109 26979
rect 22143 26945 22155 26979
rect 22097 26939 22155 26945
rect 24762 26936 24768 26988
rect 24820 26976 24826 26988
rect 24949 26979 25007 26985
rect 24949 26976 24961 26979
rect 24820 26948 24961 26976
rect 24820 26936 24826 26948
rect 24949 26945 24961 26948
rect 24995 26945 25007 26979
rect 25130 26976 25136 26988
rect 25091 26948 25136 26976
rect 24949 26939 25007 26945
rect 25130 26936 25136 26948
rect 25188 26936 25194 26988
rect 25590 26976 25596 26988
rect 25551 26948 25596 26976
rect 25590 26936 25596 26948
rect 25648 26936 25654 26988
rect 25700 26985 25728 27016
rect 26142 27004 26148 27016
rect 26200 27044 26206 27056
rect 27525 27047 27583 27053
rect 27525 27044 27537 27047
rect 26200 27016 27537 27044
rect 26200 27004 26206 27016
rect 27525 27013 27537 27016
rect 27571 27013 27583 27047
rect 27525 27007 27583 27013
rect 25685 26979 25743 26985
rect 25685 26945 25697 26979
rect 25731 26945 25743 26979
rect 25866 26976 25872 26988
rect 25827 26948 25872 26976
rect 25685 26939 25743 26945
rect 25866 26936 25872 26948
rect 25924 26936 25930 26988
rect 27246 26976 27252 26988
rect 27207 26948 27252 26976
rect 27246 26936 27252 26948
rect 27304 26936 27310 26988
rect 27338 26936 27344 26988
rect 27396 26976 27402 26988
rect 30006 26976 30012 26988
rect 27396 26948 27441 26976
rect 29967 26948 30012 26976
rect 27396 26936 27402 26948
rect 30006 26936 30012 26948
rect 30064 26936 30070 26988
rect 22646 26908 22652 26920
rect 22607 26880 22652 26908
rect 22646 26868 22652 26880
rect 22704 26868 22710 26920
rect 26142 26868 26148 26920
rect 26200 26908 26206 26920
rect 26421 26911 26479 26917
rect 26421 26908 26433 26911
rect 26200 26880 26433 26908
rect 26200 26868 26206 26880
rect 26421 26877 26433 26880
rect 26467 26908 26479 26911
rect 27614 26908 27620 26920
rect 26467 26880 27620 26908
rect 26467 26877 26479 26880
rect 26421 26871 26479 26877
rect 27614 26868 27620 26880
rect 27672 26868 27678 26920
rect 29730 26908 29736 26920
rect 29643 26880 29736 26908
rect 29730 26868 29736 26880
rect 29788 26908 29794 26920
rect 29914 26908 29920 26920
rect 29788 26880 29920 26908
rect 29788 26868 29794 26880
rect 29914 26868 29920 26880
rect 29972 26868 29978 26920
rect 21542 26840 21548 26852
rect 20732 26812 21548 26840
rect 8527 26809 8539 26812
rect 8481 26803 8539 26809
rect 21542 26800 21548 26812
rect 21600 26800 21606 26852
rect 9214 26732 9220 26784
rect 9272 26772 9278 26784
rect 9493 26775 9551 26781
rect 9493 26772 9505 26775
rect 9272 26744 9505 26772
rect 9272 26732 9278 26744
rect 9493 26741 9505 26744
rect 9539 26741 9551 26775
rect 9493 26735 9551 26741
rect 11146 26732 11152 26784
rect 11204 26772 11210 26784
rect 11701 26775 11759 26781
rect 11701 26772 11713 26775
rect 11204 26744 11713 26772
rect 11204 26732 11210 26744
rect 11701 26741 11713 26744
rect 11747 26741 11759 26775
rect 11701 26735 11759 26741
rect 21177 26775 21235 26781
rect 21177 26741 21189 26775
rect 21223 26772 21235 26775
rect 22370 26772 22376 26784
rect 21223 26744 22376 26772
rect 21223 26741 21235 26744
rect 21177 26735 21235 26741
rect 22370 26732 22376 26744
rect 22428 26732 22434 26784
rect 24578 26732 24584 26784
rect 24636 26772 24642 26784
rect 27154 26772 27160 26784
rect 24636 26744 27160 26772
rect 24636 26732 24642 26744
rect 27154 26732 27160 26744
rect 27212 26732 27218 26784
rect 1104 26682 34868 26704
rect 1104 26630 5170 26682
rect 5222 26630 5234 26682
rect 5286 26630 5298 26682
rect 5350 26630 5362 26682
rect 5414 26630 5426 26682
rect 5478 26630 13611 26682
rect 13663 26630 13675 26682
rect 13727 26630 13739 26682
rect 13791 26630 13803 26682
rect 13855 26630 13867 26682
rect 13919 26630 22052 26682
rect 22104 26630 22116 26682
rect 22168 26630 22180 26682
rect 22232 26630 22244 26682
rect 22296 26630 22308 26682
rect 22360 26630 30493 26682
rect 30545 26630 30557 26682
rect 30609 26630 30621 26682
rect 30673 26630 30685 26682
rect 30737 26630 30749 26682
rect 30801 26630 34868 26682
rect 1104 26608 34868 26630
rect 12345 26571 12403 26577
rect 12345 26537 12357 26571
rect 12391 26568 12403 26571
rect 12434 26568 12440 26580
rect 12391 26540 12440 26568
rect 12391 26537 12403 26540
rect 12345 26531 12403 26537
rect 12434 26528 12440 26540
rect 12492 26528 12498 26580
rect 12894 26528 12900 26580
rect 12952 26568 12958 26580
rect 13354 26568 13360 26580
rect 12952 26540 13360 26568
rect 12952 26528 12958 26540
rect 13354 26528 13360 26540
rect 13412 26568 13418 26580
rect 13449 26571 13507 26577
rect 13449 26568 13461 26571
rect 13412 26540 13461 26568
rect 13412 26528 13418 26540
rect 13449 26537 13461 26540
rect 13495 26537 13507 26571
rect 13449 26531 13507 26537
rect 25130 26528 25136 26580
rect 25188 26568 25194 26580
rect 25225 26571 25283 26577
rect 25225 26568 25237 26571
rect 25188 26540 25237 26568
rect 25188 26528 25194 26540
rect 25225 26537 25237 26540
rect 25271 26537 25283 26571
rect 25958 26568 25964 26580
rect 25225 26531 25283 26537
rect 25608 26540 25964 26568
rect 9306 26460 9312 26512
rect 9364 26500 9370 26512
rect 25608 26509 25636 26540
rect 25958 26528 25964 26540
rect 26016 26528 26022 26580
rect 26602 26528 26608 26580
rect 26660 26568 26666 26580
rect 26786 26568 26792 26580
rect 26660 26540 26792 26568
rect 26660 26528 26666 26540
rect 26786 26528 26792 26540
rect 26844 26528 26850 26580
rect 27062 26568 27068 26580
rect 27023 26540 27068 26568
rect 27062 26528 27068 26540
rect 27120 26528 27126 26580
rect 29178 26568 29184 26580
rect 29139 26540 29184 26568
rect 29178 26528 29184 26540
rect 29236 26528 29242 26580
rect 9401 26503 9459 26509
rect 9401 26500 9413 26503
rect 9364 26472 9413 26500
rect 9364 26460 9370 26472
rect 9401 26469 9413 26472
rect 9447 26469 9459 26503
rect 13265 26503 13323 26509
rect 13265 26500 13277 26503
rect 9401 26463 9459 26469
rect 11716 26472 13277 26500
rect 11146 26432 11152 26444
rect 11107 26404 11152 26432
rect 11146 26392 11152 26404
rect 11204 26392 11210 26444
rect 11716 26441 11744 26472
rect 13265 26469 13277 26472
rect 13311 26469 13323 26503
rect 13265 26463 13323 26469
rect 25593 26503 25651 26509
rect 25593 26469 25605 26503
rect 25639 26469 25651 26503
rect 25593 26463 25651 26469
rect 27522 26460 27528 26512
rect 27580 26460 27586 26512
rect 28626 26460 28632 26512
rect 28684 26500 28690 26512
rect 31297 26503 31355 26509
rect 31297 26500 31309 26503
rect 28684 26472 31309 26500
rect 28684 26460 28690 26472
rect 31297 26469 31309 26472
rect 31343 26469 31355 26503
rect 31297 26463 31355 26469
rect 11701 26435 11759 26441
rect 11701 26401 11713 26435
rect 11747 26401 11759 26435
rect 12713 26435 12771 26441
rect 12713 26432 12725 26435
rect 11701 26395 11759 26401
rect 12406 26404 12725 26432
rect 11333 26367 11391 26373
rect 11333 26333 11345 26367
rect 11379 26364 11391 26367
rect 12406 26364 12434 26404
rect 12713 26401 12725 26404
rect 12759 26432 12771 26435
rect 12802 26432 12808 26444
rect 12759 26404 12808 26432
rect 12759 26401 12771 26404
rect 12713 26395 12771 26401
rect 12802 26392 12808 26404
rect 12860 26392 12866 26444
rect 17957 26435 18015 26441
rect 17957 26401 17969 26435
rect 18003 26432 18015 26435
rect 18230 26432 18236 26444
rect 18003 26404 18236 26432
rect 18003 26401 18015 26404
rect 17957 26395 18015 26401
rect 18230 26392 18236 26404
rect 18288 26392 18294 26444
rect 20990 26432 20996 26444
rect 18616 26404 20996 26432
rect 12618 26364 12624 26376
rect 11379 26336 12434 26364
rect 12579 26336 12624 26364
rect 11379 26333 11391 26336
rect 11333 26327 11391 26333
rect 12618 26324 12624 26336
rect 12676 26324 12682 26376
rect 13078 26324 13084 26376
rect 13136 26364 13142 26376
rect 15657 26367 15715 26373
rect 13136 26336 13676 26364
rect 13136 26324 13142 26336
rect 9125 26299 9183 26305
rect 9125 26265 9137 26299
rect 9171 26296 9183 26299
rect 9766 26296 9772 26308
rect 9171 26268 9772 26296
rect 9171 26265 9183 26268
rect 9125 26259 9183 26265
rect 9766 26256 9772 26268
rect 9824 26296 9830 26308
rect 11609 26299 11667 26305
rect 11609 26296 11621 26299
rect 9824 26268 11621 26296
rect 9824 26256 9830 26268
rect 11609 26265 11621 26268
rect 11655 26265 11667 26299
rect 11609 26259 11667 26265
rect 12526 26256 12532 26308
rect 12584 26296 12590 26308
rect 13446 26305 13452 26308
rect 13417 26299 13452 26305
rect 13417 26296 13429 26299
rect 12584 26268 13429 26296
rect 12584 26256 12590 26268
rect 13417 26265 13429 26268
rect 13504 26296 13510 26308
rect 13648 26305 13676 26336
rect 15657 26333 15669 26367
rect 15703 26364 15715 26367
rect 15838 26364 15844 26376
rect 15703 26336 15844 26364
rect 15703 26333 15715 26336
rect 15657 26327 15715 26333
rect 15838 26324 15844 26336
rect 15896 26324 15902 26376
rect 15933 26367 15991 26373
rect 15933 26333 15945 26367
rect 15979 26364 15991 26367
rect 17218 26364 17224 26376
rect 15979 26336 17224 26364
rect 15979 26333 15991 26336
rect 15933 26327 15991 26333
rect 17218 26324 17224 26336
rect 17276 26324 17282 26376
rect 18616 26373 18644 26404
rect 20990 26392 20996 26404
rect 21048 26432 21054 26444
rect 21634 26432 21640 26444
rect 21048 26404 21640 26432
rect 21048 26392 21054 26404
rect 21634 26392 21640 26404
rect 21692 26392 21698 26444
rect 22738 26392 22744 26444
rect 22796 26432 22802 26444
rect 27540 26432 27568 26460
rect 22796 26404 25728 26432
rect 22796 26392 22802 26404
rect 18601 26367 18659 26373
rect 18601 26333 18613 26367
rect 18647 26333 18659 26367
rect 18601 26327 18659 26333
rect 18877 26367 18935 26373
rect 18877 26333 18889 26367
rect 18923 26364 18935 26367
rect 21542 26364 21548 26376
rect 18923 26336 21548 26364
rect 18923 26333 18935 26336
rect 18877 26327 18935 26333
rect 21542 26324 21548 26336
rect 21600 26324 21606 26376
rect 25038 26324 25044 26376
rect 25096 26364 25102 26376
rect 25314 26364 25320 26376
rect 25096 26336 25320 26364
rect 25096 26324 25102 26336
rect 25314 26324 25320 26336
rect 25372 26364 25378 26376
rect 25409 26367 25467 26373
rect 25409 26364 25421 26367
rect 25372 26336 25421 26364
rect 25372 26324 25378 26336
rect 25409 26333 25421 26336
rect 25455 26333 25467 26367
rect 25409 26327 25467 26333
rect 25498 26324 25504 26376
rect 25556 26364 25562 26376
rect 25700 26373 25728 26404
rect 26804 26404 27568 26432
rect 25684 26367 25742 26373
rect 25556 26336 25601 26364
rect 25556 26324 25562 26336
rect 25684 26333 25696 26367
rect 25730 26333 25742 26367
rect 25866 26364 25872 26376
rect 25827 26336 25872 26364
rect 25684 26327 25742 26333
rect 25866 26324 25872 26336
rect 25924 26324 25930 26376
rect 26510 26364 26516 26376
rect 26471 26336 26516 26364
rect 26510 26324 26516 26336
rect 26568 26324 26574 26376
rect 26804 26373 26832 26404
rect 26605 26367 26663 26373
rect 26605 26333 26617 26367
rect 26651 26333 26663 26367
rect 26605 26327 26663 26333
rect 26789 26367 26847 26373
rect 26789 26333 26801 26367
rect 26835 26333 26847 26367
rect 26789 26327 26847 26333
rect 13633 26299 13691 26305
rect 13504 26268 13565 26296
rect 13417 26259 13452 26265
rect 13446 26256 13452 26259
rect 13504 26256 13510 26268
rect 13633 26265 13645 26299
rect 13679 26265 13691 26299
rect 13633 26259 13691 26265
rect 16117 26299 16175 26305
rect 16117 26265 16129 26299
rect 16163 26296 16175 26299
rect 17690 26299 17748 26305
rect 17690 26296 17702 26299
rect 16163 26268 17702 26296
rect 16163 26265 16175 26268
rect 16117 26259 16175 26265
rect 17690 26265 17702 26268
rect 17736 26265 17748 26299
rect 18414 26296 18420 26308
rect 18375 26268 18420 26296
rect 17690 26259 17748 26265
rect 18414 26256 18420 26268
rect 18472 26256 18478 26308
rect 18785 26299 18843 26305
rect 18785 26265 18797 26299
rect 18831 26296 18843 26299
rect 19334 26296 19340 26308
rect 18831 26268 19340 26296
rect 18831 26265 18843 26268
rect 18785 26259 18843 26265
rect 19334 26256 19340 26268
rect 19392 26256 19398 26308
rect 22554 26296 22560 26308
rect 22515 26268 22560 26296
rect 22554 26256 22560 26268
rect 22612 26256 22618 26308
rect 22646 26256 22652 26308
rect 22704 26296 22710 26308
rect 25130 26296 25136 26308
rect 22704 26268 25136 26296
rect 22704 26256 22710 26268
rect 25130 26256 25136 26268
rect 25188 26256 25194 26308
rect 26620 26296 26648 26327
rect 26878 26324 26884 26376
rect 26936 26364 26942 26376
rect 26936 26336 26981 26364
rect 26936 26324 26942 26336
rect 27154 26324 27160 26376
rect 27212 26364 27218 26376
rect 27525 26367 27583 26373
rect 27525 26364 27537 26367
rect 27212 26336 27537 26364
rect 27212 26324 27218 26336
rect 27525 26333 27537 26336
rect 27571 26333 27583 26367
rect 28718 26364 28724 26376
rect 28679 26336 28724 26364
rect 27525 26327 27583 26333
rect 28718 26324 28724 26336
rect 28776 26324 28782 26376
rect 28813 26367 28871 26373
rect 28813 26333 28825 26367
rect 28859 26364 28871 26367
rect 28902 26364 28908 26376
rect 28859 26336 28908 26364
rect 28859 26333 28871 26336
rect 28813 26327 28871 26333
rect 28902 26324 28908 26336
rect 28960 26324 28966 26376
rect 28997 26367 29055 26373
rect 28997 26333 29009 26367
rect 29043 26333 29055 26367
rect 28997 26327 29055 26333
rect 27614 26296 27620 26308
rect 26620 26268 27620 26296
rect 27614 26256 27620 26268
rect 27672 26256 27678 26308
rect 27801 26299 27859 26305
rect 27801 26296 27813 26299
rect 27724 26268 27813 26296
rect 9306 26188 9312 26240
rect 9364 26228 9370 26240
rect 9585 26231 9643 26237
rect 9585 26228 9597 26231
rect 9364 26200 9597 26228
rect 9364 26188 9370 26200
rect 9585 26197 9597 26200
rect 9631 26197 9643 26231
rect 9585 26191 9643 26197
rect 15654 26188 15660 26240
rect 15712 26228 15718 26240
rect 15749 26231 15807 26237
rect 15749 26228 15761 26231
rect 15712 26200 15761 26228
rect 15712 26188 15718 26200
rect 15749 26197 15761 26200
rect 15795 26228 15807 26231
rect 16577 26231 16635 26237
rect 16577 26228 16589 26231
rect 15795 26200 16589 26228
rect 15795 26197 15807 26200
rect 15749 26191 15807 26197
rect 16577 26197 16589 26200
rect 16623 26197 16635 26231
rect 16577 26191 16635 26197
rect 21085 26231 21143 26237
rect 21085 26197 21097 26231
rect 21131 26228 21143 26231
rect 21174 26228 21180 26240
rect 21131 26200 21180 26228
rect 21131 26197 21143 26200
rect 21085 26191 21143 26197
rect 21174 26188 21180 26200
rect 21232 26188 21238 26240
rect 26786 26188 26792 26240
rect 26844 26228 26850 26240
rect 27724 26228 27752 26268
rect 27801 26265 27813 26268
rect 27847 26265 27859 26299
rect 27801 26259 27859 26265
rect 29012 26240 29040 26327
rect 29086 26256 29092 26308
rect 29144 26296 29150 26308
rect 30009 26299 30067 26305
rect 30009 26296 30021 26299
rect 29144 26268 30021 26296
rect 29144 26256 29150 26268
rect 30009 26265 30021 26268
rect 30055 26265 30067 26299
rect 30009 26259 30067 26265
rect 26844 26200 27752 26228
rect 26844 26188 26850 26200
rect 28994 26188 29000 26240
rect 29052 26188 29058 26240
rect 1104 26138 35027 26160
rect 1104 26086 9390 26138
rect 9442 26086 9454 26138
rect 9506 26086 9518 26138
rect 9570 26086 9582 26138
rect 9634 26086 9646 26138
rect 9698 26086 17831 26138
rect 17883 26086 17895 26138
rect 17947 26086 17959 26138
rect 18011 26086 18023 26138
rect 18075 26086 18087 26138
rect 18139 26086 26272 26138
rect 26324 26086 26336 26138
rect 26388 26086 26400 26138
rect 26452 26086 26464 26138
rect 26516 26086 26528 26138
rect 26580 26086 34713 26138
rect 34765 26086 34777 26138
rect 34829 26086 34841 26138
rect 34893 26086 34905 26138
rect 34957 26086 34969 26138
rect 35021 26086 35027 26138
rect 1104 26064 35027 26086
rect 9766 25984 9772 26036
rect 9824 26024 9830 26036
rect 10590 26027 10648 26033
rect 10590 26024 10602 26027
rect 9824 25996 10602 26024
rect 9824 25984 9830 25996
rect 10590 25993 10602 25996
rect 10636 25993 10648 26027
rect 10590 25987 10648 25993
rect 12253 26027 12311 26033
rect 12253 25993 12265 26027
rect 12299 26024 12311 26027
rect 12526 26024 12532 26036
rect 12299 25996 12532 26024
rect 12299 25993 12311 25996
rect 12253 25987 12311 25993
rect 12526 25984 12532 25996
rect 12584 25984 12590 26036
rect 14734 26024 14740 26036
rect 13188 25996 14740 26024
rect 9306 25916 9312 25968
rect 9364 25956 9370 25968
rect 10505 25959 10563 25965
rect 10505 25956 10517 25959
rect 9364 25928 10517 25956
rect 9364 25916 9370 25928
rect 9508 25897 9536 25928
rect 10505 25925 10517 25928
rect 10551 25925 10563 25959
rect 10505 25919 10563 25925
rect 12434 25916 12440 25968
rect 12492 25956 12498 25968
rect 13081 25959 13139 25965
rect 13081 25956 13093 25959
rect 12492 25928 13093 25956
rect 12492 25916 12498 25928
rect 13081 25925 13093 25928
rect 13127 25925 13139 25959
rect 13081 25919 13139 25925
rect 9493 25891 9551 25897
rect 9493 25857 9505 25891
rect 9539 25857 9551 25891
rect 9766 25888 9772 25900
rect 9727 25860 9772 25888
rect 9493 25851 9551 25857
rect 9766 25848 9772 25860
rect 9824 25848 9830 25900
rect 10410 25888 10416 25900
rect 10371 25860 10416 25888
rect 10410 25848 10416 25860
rect 10468 25848 10474 25900
rect 10689 25891 10747 25897
rect 10689 25857 10701 25891
rect 10735 25888 10747 25891
rect 12250 25888 12256 25900
rect 10735 25860 12256 25888
rect 10735 25857 10747 25860
rect 10689 25851 10747 25857
rect 12250 25848 12256 25860
rect 12308 25848 12314 25900
rect 12342 25848 12348 25900
rect 12400 25888 12406 25900
rect 13188 25888 13216 25996
rect 14734 25984 14740 25996
rect 14792 25984 14798 26036
rect 21361 26027 21419 26033
rect 21361 25993 21373 26027
rect 21407 26024 21419 26027
rect 22646 26024 22652 26036
rect 21407 25996 22652 26024
rect 21407 25993 21419 25996
rect 21361 25987 21419 25993
rect 22646 25984 22652 25996
rect 22704 25984 22710 26036
rect 23566 26024 23572 26036
rect 23527 25996 23572 26024
rect 23566 25984 23572 25996
rect 23624 25984 23630 26036
rect 25593 26027 25651 26033
rect 25593 25993 25605 26027
rect 25639 26024 25651 26027
rect 25682 26024 25688 26036
rect 25639 25996 25688 26024
rect 25639 25993 25651 25996
rect 25593 25987 25651 25993
rect 25682 25984 25688 25996
rect 25740 25984 25746 26036
rect 27157 26027 27215 26033
rect 27157 25993 27169 26027
rect 27203 26024 27215 26027
rect 27246 26024 27252 26036
rect 27203 25996 27252 26024
rect 27203 25993 27215 25996
rect 27157 25987 27215 25993
rect 27246 25984 27252 25996
rect 27304 25984 27310 26036
rect 29914 26024 29920 26036
rect 29875 25996 29920 26024
rect 29914 25984 29920 25996
rect 29972 25984 29978 26036
rect 13354 25956 13360 25968
rect 13315 25928 13360 25956
rect 13354 25916 13360 25928
rect 13412 25916 13418 25968
rect 19242 25916 19248 25968
rect 19300 25956 19306 25968
rect 20990 25956 20996 25968
rect 19300 25928 20996 25956
rect 19300 25916 19306 25928
rect 20990 25916 20996 25928
rect 21048 25956 21054 25968
rect 24581 25959 24639 25965
rect 21048 25928 21220 25956
rect 21048 25916 21054 25928
rect 13265 25891 13323 25897
rect 13265 25888 13277 25891
rect 12400 25860 13277 25888
rect 12400 25848 12406 25860
rect 13265 25857 13277 25860
rect 13311 25857 13323 25891
rect 13265 25851 13323 25857
rect 9214 25780 9220 25832
rect 9272 25820 9278 25832
rect 9585 25823 9643 25829
rect 9585 25820 9597 25823
rect 9272 25792 9597 25820
rect 9272 25780 9278 25792
rect 9585 25789 9597 25792
rect 9631 25789 9643 25823
rect 9585 25783 9643 25789
rect 12069 25823 12127 25829
rect 12069 25789 12081 25823
rect 12115 25820 12127 25823
rect 13372 25820 13400 25916
rect 13446 25848 13452 25900
rect 13504 25897 13510 25900
rect 13504 25888 13512 25897
rect 16942 25888 16948 25900
rect 13504 25860 13549 25888
rect 16903 25860 16948 25888
rect 13504 25851 13512 25860
rect 13504 25848 13510 25851
rect 16942 25848 16948 25860
rect 17000 25848 17006 25900
rect 19610 25888 19616 25900
rect 19571 25860 19616 25888
rect 19610 25848 19616 25860
rect 19668 25848 19674 25900
rect 21192 25897 21220 25928
rect 24581 25925 24593 25959
rect 24627 25956 24639 25959
rect 25133 25959 25191 25965
rect 25133 25956 25145 25959
rect 24627 25928 25145 25956
rect 24627 25925 24639 25928
rect 24581 25919 24639 25925
rect 25133 25925 25145 25928
rect 25179 25956 25191 25959
rect 25498 25956 25504 25968
rect 25179 25928 25504 25956
rect 25179 25925 25191 25928
rect 25133 25919 25191 25925
rect 25498 25916 25504 25928
rect 25556 25916 25562 25968
rect 28626 25956 28632 25968
rect 28587 25928 28632 25956
rect 28626 25916 28632 25928
rect 28684 25916 28690 25968
rect 21177 25891 21235 25897
rect 21177 25857 21189 25891
rect 21223 25857 21235 25891
rect 21177 25851 21235 25857
rect 21453 25891 21511 25897
rect 21453 25857 21465 25891
rect 21499 25888 21511 25891
rect 21542 25888 21548 25900
rect 21499 25860 21548 25888
rect 21499 25857 21511 25860
rect 21453 25851 21511 25857
rect 21542 25848 21548 25860
rect 21600 25848 21606 25900
rect 22281 25891 22339 25897
rect 22281 25857 22293 25891
rect 22327 25888 22339 25891
rect 22370 25888 22376 25900
rect 22327 25860 22376 25888
rect 22327 25857 22339 25860
rect 22281 25851 22339 25857
rect 22370 25848 22376 25860
rect 22428 25848 22434 25900
rect 24489 25891 24547 25897
rect 24489 25857 24501 25891
rect 24535 25857 24547 25891
rect 24670 25888 24676 25900
rect 24631 25860 24676 25888
rect 24489 25851 24547 25857
rect 22005 25823 22063 25829
rect 22005 25820 22017 25823
rect 12115 25792 13400 25820
rect 21192 25792 22017 25820
rect 12115 25789 12127 25792
rect 12069 25783 12127 25789
rect 9600 25752 9628 25783
rect 21192 25764 21220 25792
rect 22005 25789 22017 25792
rect 22051 25789 22063 25823
rect 22005 25783 22063 25789
rect 23658 25780 23664 25832
rect 23716 25820 23722 25832
rect 24504 25820 24532 25851
rect 24670 25848 24676 25860
rect 24728 25848 24734 25900
rect 25866 25848 25872 25900
rect 25924 25888 25930 25900
rect 26510 25888 26516 25900
rect 25924 25860 26516 25888
rect 25924 25848 25930 25860
rect 26510 25848 26516 25860
rect 26568 25848 26574 25900
rect 27614 25888 27620 25900
rect 27575 25860 27620 25888
rect 27614 25848 27620 25860
rect 27672 25848 27678 25900
rect 32306 25888 32312 25900
rect 32267 25860 32312 25888
rect 32306 25848 32312 25860
rect 32364 25848 32370 25900
rect 32398 25848 32404 25900
rect 32456 25888 32462 25900
rect 32585 25891 32643 25897
rect 32456 25860 32501 25888
rect 32456 25848 32462 25860
rect 32585 25857 32597 25891
rect 32631 25857 32643 25891
rect 32585 25851 32643 25857
rect 26050 25820 26056 25832
rect 23716 25792 26056 25820
rect 23716 25780 23722 25792
rect 26050 25780 26056 25792
rect 26108 25780 26114 25832
rect 26605 25823 26663 25829
rect 26605 25789 26617 25823
rect 26651 25820 26663 25823
rect 26694 25820 26700 25832
rect 26651 25792 26700 25820
rect 26651 25789 26663 25792
rect 26605 25783 26663 25789
rect 26694 25780 26700 25792
rect 26752 25780 26758 25832
rect 27062 25780 27068 25832
rect 27120 25820 27126 25832
rect 27341 25823 27399 25829
rect 27341 25820 27353 25823
rect 27120 25792 27353 25820
rect 27120 25780 27126 25792
rect 27341 25789 27353 25792
rect 27387 25789 27399 25823
rect 27341 25783 27399 25789
rect 27433 25823 27491 25829
rect 27433 25789 27445 25823
rect 27479 25789 27491 25823
rect 27433 25783 27491 25789
rect 10410 25752 10416 25764
rect 9600 25724 10416 25752
rect 10410 25712 10416 25724
rect 10468 25712 10474 25764
rect 14458 25752 14464 25764
rect 12406 25724 14464 25752
rect 9953 25687 10011 25693
rect 9953 25653 9965 25687
rect 9999 25684 10011 25687
rect 12406 25684 12434 25724
rect 14458 25712 14464 25724
rect 14516 25712 14522 25764
rect 21174 25712 21180 25764
rect 21232 25712 21238 25764
rect 24854 25712 24860 25764
rect 24912 25752 24918 25764
rect 25409 25755 25467 25761
rect 25409 25752 25421 25755
rect 24912 25724 25421 25752
rect 24912 25712 24918 25724
rect 25409 25721 25421 25724
rect 25455 25752 25467 25755
rect 26878 25752 26884 25764
rect 25455 25724 26884 25752
rect 25455 25721 25467 25724
rect 25409 25715 25467 25721
rect 26878 25712 26884 25724
rect 26936 25752 26942 25764
rect 27448 25752 27476 25783
rect 27522 25780 27528 25832
rect 27580 25820 27586 25832
rect 27580 25792 27625 25820
rect 27580 25780 27586 25792
rect 32490 25780 32496 25832
rect 32548 25820 32554 25832
rect 32600 25820 32628 25851
rect 32548 25792 32628 25820
rect 32548 25780 32554 25792
rect 26936 25724 27476 25752
rect 26936 25712 26942 25724
rect 9999 25656 12434 25684
rect 12621 25687 12679 25693
rect 9999 25653 10011 25656
rect 9953 25647 10011 25653
rect 12621 25653 12633 25687
rect 12667 25684 12679 25687
rect 12710 25684 12716 25696
rect 12667 25656 12716 25684
rect 12667 25653 12679 25656
rect 12621 25647 12679 25653
rect 12710 25644 12716 25656
rect 12768 25644 12774 25696
rect 13078 25684 13084 25696
rect 13039 25656 13084 25684
rect 13078 25644 13084 25656
rect 13136 25644 13142 25696
rect 17218 25684 17224 25696
rect 17179 25656 17224 25684
rect 17218 25644 17224 25656
rect 17276 25644 17282 25696
rect 18322 25684 18328 25696
rect 18283 25656 18328 25684
rect 18322 25644 18328 25656
rect 18380 25644 18386 25696
rect 20898 25644 20904 25696
rect 20956 25684 20962 25696
rect 20993 25687 21051 25693
rect 20993 25684 21005 25687
rect 20956 25656 21005 25684
rect 20956 25644 20962 25656
rect 20993 25653 21005 25656
rect 21039 25653 21051 25687
rect 32766 25684 32772 25696
rect 32727 25656 32772 25684
rect 20993 25647 21051 25653
rect 32766 25644 32772 25656
rect 32824 25644 32830 25696
rect 1104 25594 34868 25616
rect 1104 25542 5170 25594
rect 5222 25542 5234 25594
rect 5286 25542 5298 25594
rect 5350 25542 5362 25594
rect 5414 25542 5426 25594
rect 5478 25542 13611 25594
rect 13663 25542 13675 25594
rect 13727 25542 13739 25594
rect 13791 25542 13803 25594
rect 13855 25542 13867 25594
rect 13919 25542 22052 25594
rect 22104 25542 22116 25594
rect 22168 25542 22180 25594
rect 22232 25542 22244 25594
rect 22296 25542 22308 25594
rect 22360 25542 30493 25594
rect 30545 25542 30557 25594
rect 30609 25542 30621 25594
rect 30673 25542 30685 25594
rect 30737 25542 30749 25594
rect 30801 25542 34868 25594
rect 1104 25520 34868 25542
rect 15381 25483 15439 25489
rect 15381 25449 15393 25483
rect 15427 25480 15439 25483
rect 15654 25480 15660 25492
rect 15427 25452 15660 25480
rect 15427 25449 15439 25452
rect 15381 25443 15439 25449
rect 15654 25440 15660 25452
rect 15712 25440 15718 25492
rect 19794 25480 19800 25492
rect 19755 25452 19800 25480
rect 19794 25440 19800 25452
rect 19852 25440 19858 25492
rect 25958 25440 25964 25492
rect 26016 25480 26022 25492
rect 26053 25483 26111 25489
rect 26053 25480 26065 25483
rect 26016 25452 26065 25480
rect 26016 25440 26022 25452
rect 26053 25449 26065 25452
rect 26099 25449 26111 25483
rect 26053 25443 26111 25449
rect 26237 25483 26295 25489
rect 26237 25449 26249 25483
rect 26283 25480 26295 25483
rect 26786 25480 26792 25492
rect 26283 25452 26792 25480
rect 26283 25449 26295 25452
rect 26237 25443 26295 25449
rect 26786 25440 26792 25452
rect 26844 25440 26850 25492
rect 27614 25440 27620 25492
rect 27672 25480 27678 25492
rect 28261 25483 28319 25489
rect 28261 25480 28273 25483
rect 27672 25452 28273 25480
rect 27672 25440 27678 25452
rect 28261 25449 28273 25452
rect 28307 25449 28319 25483
rect 31481 25483 31539 25489
rect 31481 25480 31493 25483
rect 28261 25443 28319 25449
rect 29012 25452 31493 25480
rect 3326 25304 3332 25356
rect 3384 25344 3390 25356
rect 3973 25347 4031 25353
rect 3973 25344 3985 25347
rect 3384 25316 3985 25344
rect 3384 25304 3390 25316
rect 3973 25313 3985 25316
rect 4019 25313 4031 25347
rect 13078 25344 13084 25356
rect 3973 25307 4031 25313
rect 12544 25316 13084 25344
rect 4154 25276 4160 25288
rect 4115 25248 4160 25276
rect 4154 25236 4160 25248
rect 4212 25236 4218 25288
rect 4249 25279 4307 25285
rect 4249 25245 4261 25279
rect 4295 25245 4307 25279
rect 4249 25239 4307 25245
rect 6733 25279 6791 25285
rect 6733 25245 6745 25279
rect 6779 25276 6791 25279
rect 6822 25276 6828 25288
rect 6779 25248 6828 25276
rect 6779 25245 6791 25248
rect 6733 25239 6791 25245
rect 4264 25208 4292 25239
rect 6822 25236 6828 25248
rect 6880 25236 6886 25288
rect 6917 25279 6975 25285
rect 6917 25245 6929 25279
rect 6963 25276 6975 25279
rect 7466 25276 7472 25288
rect 6963 25248 7472 25276
rect 6963 25245 6975 25248
rect 6917 25239 6975 25245
rect 7466 25236 7472 25248
rect 7524 25236 7530 25288
rect 12250 25276 12256 25288
rect 12211 25248 12256 25276
rect 12250 25236 12256 25248
rect 12308 25236 12314 25288
rect 12544 25285 12572 25316
rect 13078 25304 13084 25316
rect 13136 25304 13142 25356
rect 15672 25344 15700 25440
rect 16298 25412 16304 25424
rect 16259 25384 16304 25412
rect 16298 25372 16304 25384
rect 16356 25372 16362 25424
rect 21174 25344 21180 25356
rect 15672 25316 16344 25344
rect 21135 25316 21180 25344
rect 12529 25279 12587 25285
rect 12529 25245 12541 25279
rect 12575 25245 12587 25279
rect 12710 25276 12716 25288
rect 12671 25248 12716 25276
rect 12529 25239 12587 25245
rect 12710 25236 12716 25248
rect 12768 25236 12774 25288
rect 15286 25236 15292 25288
rect 15344 25236 15350 25288
rect 15378 25236 15384 25288
rect 15436 25276 15442 25288
rect 16316 25285 16344 25316
rect 21174 25304 21180 25316
rect 21232 25304 21238 25356
rect 24670 25304 24676 25356
rect 24728 25344 24734 25356
rect 24765 25347 24823 25353
rect 24765 25344 24777 25347
rect 24728 25316 24777 25344
rect 24728 25304 24734 25316
rect 24765 25313 24777 25316
rect 24811 25313 24823 25347
rect 26602 25344 26608 25356
rect 26515 25316 26608 25344
rect 24765 25307 24823 25313
rect 16025 25279 16083 25285
rect 16025 25276 16037 25279
rect 15436 25248 16037 25276
rect 15436 25236 15442 25248
rect 16025 25245 16037 25248
rect 16071 25245 16083 25279
rect 16025 25239 16083 25245
rect 16301 25279 16359 25285
rect 16301 25245 16313 25279
rect 16347 25245 16359 25279
rect 16301 25239 16359 25245
rect 20898 25236 20904 25288
rect 20956 25285 20962 25288
rect 20956 25276 20968 25285
rect 20956 25248 21001 25276
rect 20956 25239 20968 25248
rect 20956 25236 20962 25239
rect 23474 25236 23480 25288
rect 23532 25276 23538 25288
rect 24578 25276 24584 25288
rect 23532 25248 24584 25276
rect 23532 25236 23538 25248
rect 24578 25236 24584 25248
rect 24636 25236 24642 25288
rect 24780 25276 24808 25307
rect 26602 25304 26608 25316
rect 26660 25344 26666 25356
rect 26660 25316 28396 25344
rect 26660 25304 26666 25316
rect 27246 25276 27252 25288
rect 27304 25285 27310 25288
rect 28368 25285 28396 25316
rect 27304 25279 27337 25285
rect 24780 25248 27252 25276
rect 27246 25236 27252 25248
rect 27325 25245 27337 25279
rect 27304 25239 27337 25245
rect 27426 25279 27484 25285
rect 27426 25245 27438 25279
rect 27472 25245 27484 25279
rect 27426 25239 27484 25245
rect 28353 25279 28411 25285
rect 28353 25245 28365 25279
rect 28399 25276 28411 25279
rect 28902 25276 28908 25288
rect 28399 25248 28908 25276
rect 28399 25245 28411 25248
rect 28353 25239 28411 25245
rect 27304 25236 27310 25239
rect 10226 25208 10232 25220
rect 4264 25180 10232 25208
rect 10226 25168 10232 25180
rect 10284 25168 10290 25220
rect 12268 25208 12296 25236
rect 15304 25208 15332 25236
rect 12268 25180 15332 25208
rect 15470 25168 15476 25220
rect 15528 25208 15534 25220
rect 15565 25211 15623 25217
rect 15565 25208 15577 25211
rect 15528 25180 15577 25208
rect 15528 25168 15534 25180
rect 15565 25177 15577 25180
rect 15611 25177 15623 25211
rect 15565 25171 15623 25177
rect 3970 25140 3976 25152
rect 3931 25112 3976 25140
rect 3970 25100 3976 25112
rect 4028 25100 4034 25152
rect 5074 25100 5080 25152
rect 5132 25140 5138 25152
rect 6733 25143 6791 25149
rect 6733 25140 6745 25143
rect 5132 25112 6745 25140
rect 5132 25100 5138 25112
rect 6733 25109 6745 25112
rect 6779 25109 6791 25143
rect 6733 25103 6791 25109
rect 12069 25143 12127 25149
rect 12069 25109 12081 25143
rect 12115 25140 12127 25143
rect 13446 25140 13452 25152
rect 12115 25112 13452 25140
rect 12115 25109 12127 25112
rect 12069 25103 12127 25109
rect 13446 25100 13452 25112
rect 13504 25100 13510 25152
rect 15194 25140 15200 25152
rect 15155 25112 15200 25140
rect 15194 25100 15200 25112
rect 15252 25100 15258 25152
rect 15378 25149 15384 25152
rect 15365 25143 15384 25149
rect 15365 25109 15377 25143
rect 15365 25103 15384 25109
rect 15378 25100 15384 25103
rect 15436 25100 15442 25152
rect 15580 25140 15608 25171
rect 21082 25168 21088 25220
rect 21140 25208 21146 25220
rect 21637 25211 21695 25217
rect 21637 25208 21649 25211
rect 21140 25180 21649 25208
rect 21140 25168 21146 25180
rect 21637 25177 21649 25180
rect 21683 25177 21695 25211
rect 21637 25171 21695 25177
rect 26050 25168 26056 25220
rect 26108 25208 26114 25220
rect 26237 25211 26295 25217
rect 26237 25208 26249 25211
rect 26108 25180 26249 25208
rect 26108 25168 26114 25180
rect 26237 25177 26249 25180
rect 26283 25177 26295 25211
rect 26237 25171 26295 25177
rect 26510 25168 26516 25220
rect 26568 25208 26574 25220
rect 27448 25208 27476 25239
rect 28902 25236 28908 25248
rect 28960 25236 28966 25288
rect 29012 25208 29040 25452
rect 31481 25449 31493 25452
rect 31527 25480 31539 25483
rect 32398 25480 32404 25492
rect 31527 25452 32404 25480
rect 31527 25449 31539 25452
rect 31481 25443 31539 25449
rect 32398 25440 32404 25452
rect 32456 25440 32462 25492
rect 30098 25276 30104 25288
rect 30059 25248 30104 25276
rect 30098 25236 30104 25248
rect 30156 25236 30162 25288
rect 30368 25279 30426 25285
rect 30368 25245 30380 25279
rect 30414 25276 30426 25279
rect 32766 25276 32772 25288
rect 30414 25248 32772 25276
rect 30414 25245 30426 25248
rect 30368 25239 30426 25245
rect 32766 25236 32772 25248
rect 32824 25236 32830 25288
rect 26568 25180 29040 25208
rect 26568 25168 26574 25180
rect 16117 25143 16175 25149
rect 16117 25140 16129 25143
rect 15580 25112 16129 25140
rect 16117 25109 16129 25112
rect 16163 25140 16175 25143
rect 16390 25140 16396 25152
rect 16163 25112 16396 25140
rect 16163 25109 16175 25112
rect 16117 25103 16175 25109
rect 16390 25100 16396 25112
rect 16448 25100 16454 25152
rect 22554 25100 22560 25152
rect 22612 25140 22618 25152
rect 22925 25143 22983 25149
rect 22925 25140 22937 25143
rect 22612 25112 22937 25140
rect 22612 25100 22618 25112
rect 22925 25109 22937 25112
rect 22971 25109 22983 25143
rect 27062 25140 27068 25152
rect 27023 25112 27068 25140
rect 22925 25103 22983 25109
rect 27062 25100 27068 25112
rect 27120 25100 27126 25152
rect 1104 25050 35027 25072
rect 1104 24998 9390 25050
rect 9442 24998 9454 25050
rect 9506 24998 9518 25050
rect 9570 24998 9582 25050
rect 9634 24998 9646 25050
rect 9698 24998 17831 25050
rect 17883 24998 17895 25050
rect 17947 24998 17959 25050
rect 18011 24998 18023 25050
rect 18075 24998 18087 25050
rect 18139 24998 26272 25050
rect 26324 24998 26336 25050
rect 26388 24998 26400 25050
rect 26452 24998 26464 25050
rect 26516 24998 26528 25050
rect 26580 24998 34713 25050
rect 34765 24998 34777 25050
rect 34829 24998 34841 25050
rect 34893 24998 34905 25050
rect 34957 24998 34969 25050
rect 35021 24998 35027 25050
rect 1104 24976 35027 24998
rect 17218 24896 17224 24948
rect 17276 24936 17282 24948
rect 23382 24936 23388 24948
rect 17276 24908 23388 24936
rect 17276 24896 17282 24908
rect 23382 24896 23388 24908
rect 23440 24896 23446 24948
rect 4706 24828 4712 24880
rect 4764 24868 4770 24880
rect 5261 24871 5319 24877
rect 5261 24868 5273 24871
rect 4764 24840 5273 24868
rect 4764 24828 4770 24840
rect 5261 24837 5273 24840
rect 5307 24837 5319 24871
rect 21453 24871 21511 24877
rect 5261 24831 5319 24837
rect 15212 24840 15976 24868
rect 15212 24812 15240 24840
rect 3326 24760 3332 24812
rect 3384 24800 3390 24812
rect 3384 24772 4646 24800
rect 3384 24760 3390 24772
rect 6822 24760 6828 24812
rect 6880 24800 6886 24812
rect 6917 24803 6975 24809
rect 6917 24800 6929 24803
rect 6880 24772 6929 24800
rect 6880 24760 6886 24772
rect 6917 24769 6929 24772
rect 6963 24769 6975 24803
rect 6917 24763 6975 24769
rect 7466 24760 7472 24812
rect 7524 24760 7530 24812
rect 12802 24760 12808 24812
rect 12860 24800 12866 24812
rect 14829 24803 14887 24809
rect 14829 24800 14841 24803
rect 12860 24772 14841 24800
rect 12860 24760 12866 24772
rect 14829 24769 14841 24772
rect 14875 24769 14887 24803
rect 14829 24763 14887 24769
rect 15105 24803 15163 24809
rect 15105 24769 15117 24803
rect 15151 24769 15163 24803
rect 15105 24763 15163 24769
rect 3694 24732 3700 24744
rect 3655 24704 3700 24732
rect 3694 24692 3700 24704
rect 3752 24692 3758 24744
rect 3973 24735 4031 24741
rect 3973 24701 3985 24735
rect 4019 24732 4031 24735
rect 4062 24732 4068 24744
rect 4019 24704 4068 24732
rect 4019 24701 4031 24704
rect 3973 24695 4031 24701
rect 4062 24692 4068 24704
rect 4120 24692 4126 24744
rect 4522 24692 4528 24744
rect 4580 24732 4586 24744
rect 4709 24735 4767 24741
rect 4709 24732 4721 24735
rect 4580 24704 4721 24732
rect 4580 24692 4586 24704
rect 4709 24701 4721 24704
rect 4755 24701 4767 24735
rect 4709 24695 4767 24701
rect 7929 24735 7987 24741
rect 7929 24701 7941 24735
rect 7975 24732 7987 24735
rect 8478 24732 8484 24744
rect 7975 24704 8484 24732
rect 7975 24701 7987 24704
rect 7929 24695 7987 24701
rect 8478 24692 8484 24704
rect 8536 24692 8542 24744
rect 15120 24732 15148 24763
rect 15194 24760 15200 24812
rect 15252 24800 15258 24812
rect 15252 24772 15297 24800
rect 15252 24760 15258 24772
rect 15378 24760 15384 24812
rect 15436 24800 15442 24812
rect 15948 24809 15976 24840
rect 21453 24837 21465 24871
rect 21499 24868 21511 24871
rect 23658 24868 23664 24880
rect 21499 24840 22140 24868
rect 23619 24840 23664 24868
rect 21499 24837 21511 24840
rect 21453 24831 21511 24837
rect 15933 24803 15991 24809
rect 15436 24772 15481 24800
rect 15436 24760 15442 24772
rect 15933 24769 15945 24803
rect 15979 24769 15991 24803
rect 15933 24763 15991 24769
rect 16117 24803 16175 24809
rect 16117 24769 16129 24803
rect 16163 24800 16175 24803
rect 16298 24800 16304 24812
rect 16163 24772 16304 24800
rect 16163 24769 16175 24772
rect 16117 24763 16175 24769
rect 15289 24735 15347 24741
rect 15120 24704 15240 24732
rect 15212 24664 15240 24704
rect 15289 24701 15301 24735
rect 15335 24732 15347 24735
rect 16132 24732 16160 24763
rect 16298 24760 16304 24772
rect 16356 24760 16362 24812
rect 18141 24803 18199 24809
rect 18141 24769 18153 24803
rect 18187 24800 18199 24803
rect 18414 24800 18420 24812
rect 18187 24772 18420 24800
rect 18187 24769 18199 24772
rect 18141 24763 18199 24769
rect 18414 24760 18420 24772
rect 18472 24760 18478 24812
rect 20438 24760 20444 24812
rect 20496 24800 20502 24812
rect 20993 24803 21051 24809
rect 20993 24800 21005 24803
rect 20496 24772 21005 24800
rect 20496 24760 20502 24772
rect 20993 24769 21005 24772
rect 21039 24769 21051 24803
rect 20993 24763 21051 24769
rect 21085 24803 21143 24809
rect 21085 24769 21097 24803
rect 21131 24769 21143 24803
rect 21085 24763 21143 24769
rect 15335 24704 16160 24732
rect 15335 24701 15347 24704
rect 15289 24695 15347 24701
rect 17310 24692 17316 24744
rect 17368 24732 17374 24744
rect 17865 24735 17923 24741
rect 17865 24732 17877 24735
rect 17368 24704 17877 24732
rect 17368 24692 17374 24704
rect 17865 24701 17877 24704
rect 17911 24701 17923 24735
rect 19334 24732 19340 24744
rect 19295 24704 19340 24732
rect 17865 24695 17923 24701
rect 19334 24692 19340 24704
rect 19392 24692 19398 24744
rect 20622 24692 20628 24744
rect 20680 24732 20686 24744
rect 21100 24732 21128 24763
rect 21174 24760 21180 24812
rect 21232 24800 21238 24812
rect 21269 24803 21327 24809
rect 21269 24800 21281 24803
rect 21232 24772 21281 24800
rect 21232 24760 21238 24772
rect 21269 24769 21281 24772
rect 21315 24769 21327 24803
rect 21269 24763 21327 24769
rect 22005 24735 22063 24741
rect 22005 24732 22017 24735
rect 20680 24704 21128 24732
rect 21284 24704 22017 24732
rect 20680 24692 20686 24704
rect 15562 24664 15568 24676
rect 15212 24636 15568 24664
rect 15562 24624 15568 24636
rect 15620 24624 15626 24676
rect 20640 24664 20668 24692
rect 21284 24676 21312 24704
rect 22005 24701 22017 24704
rect 22051 24701 22063 24735
rect 22112 24732 22140 24840
rect 23658 24828 23664 24840
rect 23716 24828 23722 24880
rect 24854 24828 24860 24880
rect 24912 24868 24918 24880
rect 25041 24871 25099 24877
rect 25041 24868 25053 24871
rect 24912 24840 25053 24868
rect 24912 24828 24918 24840
rect 25041 24837 25053 24840
rect 25087 24837 25099 24871
rect 27062 24868 27068 24880
rect 25041 24831 25099 24837
rect 26160 24840 27068 24868
rect 25130 24760 25136 24812
rect 25188 24800 25194 24812
rect 25314 24800 25320 24812
rect 25188 24772 25233 24800
rect 25275 24772 25320 24800
rect 25188 24760 25194 24772
rect 25314 24760 25320 24772
rect 25372 24760 25378 24812
rect 26160 24809 26188 24840
rect 27062 24828 27068 24840
rect 27120 24828 27126 24880
rect 27154 24828 27160 24880
rect 27212 24868 27218 24880
rect 28629 24871 28687 24877
rect 28629 24868 28641 24871
rect 27212 24840 28641 24868
rect 27212 24828 27218 24840
rect 28629 24837 28641 24840
rect 28675 24837 28687 24871
rect 28810 24868 28816 24880
rect 28771 24840 28816 24868
rect 28629 24831 28687 24837
rect 28810 24828 28816 24840
rect 28868 24828 28874 24880
rect 26145 24803 26203 24809
rect 26145 24769 26157 24803
rect 26191 24769 26203 24803
rect 29086 24800 29092 24812
rect 29047 24772 29092 24800
rect 26145 24763 26203 24769
rect 29086 24760 29092 24772
rect 29144 24760 29150 24812
rect 30374 24809 30380 24812
rect 30368 24763 30380 24809
rect 30432 24800 30438 24812
rect 30432 24772 30468 24800
rect 30374 24760 30380 24763
rect 30432 24760 30438 24772
rect 22281 24735 22339 24741
rect 22281 24732 22293 24735
rect 22112 24704 22293 24732
rect 22005 24695 22063 24701
rect 22281 24701 22293 24704
rect 22327 24701 22339 24735
rect 22281 24695 22339 24701
rect 26421 24735 26479 24741
rect 26421 24701 26433 24735
rect 26467 24732 26479 24735
rect 27982 24732 27988 24744
rect 26467 24704 27988 24732
rect 26467 24701 26479 24704
rect 26421 24695 26479 24701
rect 27982 24692 27988 24704
rect 28040 24692 28046 24744
rect 30098 24732 30104 24744
rect 30059 24704 30104 24732
rect 30098 24692 30104 24704
rect 30156 24692 30162 24744
rect 18800 24636 20668 24664
rect 2593 24599 2651 24605
rect 2593 24565 2605 24599
rect 2639 24596 2651 24599
rect 3234 24596 3240 24608
rect 2639 24568 3240 24596
rect 2639 24565 2651 24568
rect 2593 24559 2651 24565
rect 3234 24556 3240 24568
rect 3292 24556 3298 24608
rect 15194 24556 15200 24608
rect 15252 24596 15258 24608
rect 16117 24599 16175 24605
rect 16117 24596 16129 24599
rect 15252 24568 16129 24596
rect 15252 24556 15258 24568
rect 16117 24565 16129 24568
rect 16163 24565 16175 24599
rect 16117 24559 16175 24565
rect 16390 24556 16396 24608
rect 16448 24596 16454 24608
rect 18800 24596 18828 24636
rect 21266 24624 21272 24676
rect 21324 24624 21330 24676
rect 23308 24636 23520 24664
rect 16448 24568 18828 24596
rect 16448 24556 16454 24568
rect 20530 24556 20536 24608
rect 20588 24596 20594 24608
rect 23308 24596 23336 24636
rect 20588 24568 23336 24596
rect 23492 24596 23520 24636
rect 25424 24636 28856 24664
rect 25424 24596 25452 24636
rect 25958 24596 25964 24608
rect 23492 24568 25452 24596
rect 25919 24568 25964 24596
rect 20588 24556 20594 24568
rect 25958 24556 25964 24568
rect 26016 24556 26022 24608
rect 26329 24599 26387 24605
rect 26329 24565 26341 24599
rect 26375 24596 26387 24599
rect 26602 24596 26608 24608
rect 26375 24568 26608 24596
rect 26375 24565 26387 24568
rect 26329 24559 26387 24565
rect 26602 24556 26608 24568
rect 26660 24556 26666 24608
rect 28828 24605 28856 24636
rect 28813 24599 28871 24605
rect 28813 24565 28825 24599
rect 28859 24565 28871 24599
rect 28813 24559 28871 24565
rect 28902 24556 28908 24608
rect 28960 24596 28966 24608
rect 31478 24596 31484 24608
rect 28960 24568 31484 24596
rect 28960 24556 28966 24568
rect 31478 24556 31484 24568
rect 31536 24556 31542 24608
rect 1104 24506 34868 24528
rect 1104 24454 5170 24506
rect 5222 24454 5234 24506
rect 5286 24454 5298 24506
rect 5350 24454 5362 24506
rect 5414 24454 5426 24506
rect 5478 24454 13611 24506
rect 13663 24454 13675 24506
rect 13727 24454 13739 24506
rect 13791 24454 13803 24506
rect 13855 24454 13867 24506
rect 13919 24454 22052 24506
rect 22104 24454 22116 24506
rect 22168 24454 22180 24506
rect 22232 24454 22244 24506
rect 22296 24454 22308 24506
rect 22360 24454 30493 24506
rect 30545 24454 30557 24506
rect 30609 24454 30621 24506
rect 30673 24454 30685 24506
rect 30737 24454 30749 24506
rect 30801 24454 34868 24506
rect 1104 24432 34868 24454
rect 3326 24392 3332 24404
rect 3287 24364 3332 24392
rect 3326 24352 3332 24364
rect 3384 24352 3390 24404
rect 3694 24352 3700 24404
rect 3752 24392 3758 24404
rect 4617 24395 4675 24401
rect 4617 24392 4629 24395
rect 3752 24364 4629 24392
rect 3752 24352 3758 24364
rect 4617 24361 4629 24364
rect 4663 24361 4675 24395
rect 6822 24392 6828 24404
rect 6783 24364 6828 24392
rect 4617 24355 4675 24361
rect 6822 24352 6828 24364
rect 6880 24352 6886 24404
rect 14642 24352 14648 24404
rect 14700 24392 14706 24404
rect 20530 24392 20536 24404
rect 14700 24364 20536 24392
rect 14700 24352 14706 24364
rect 20530 24352 20536 24364
rect 20588 24352 20594 24404
rect 20640 24364 23704 24392
rect 2593 24327 2651 24333
rect 2593 24293 2605 24327
rect 2639 24324 2651 24327
rect 9214 24324 9220 24336
rect 2639 24296 4108 24324
rect 2639 24293 2651 24296
rect 2593 24287 2651 24293
rect 3970 24256 3976 24268
rect 3931 24228 3976 24256
rect 3970 24216 3976 24228
rect 4028 24216 4034 24268
rect 4080 24265 4108 24296
rect 4264 24296 9220 24324
rect 4065 24259 4123 24265
rect 4065 24225 4077 24259
rect 4111 24225 4123 24259
rect 4065 24219 4123 24225
rect 2317 24191 2375 24197
rect 2317 24157 2329 24191
rect 2363 24188 2375 24191
rect 3234 24188 3240 24200
rect 2363 24160 3096 24188
rect 3195 24160 3240 24188
rect 2363 24157 2375 24160
rect 2317 24151 2375 24157
rect 2590 24120 2596 24132
rect 2551 24092 2596 24120
rect 2590 24080 2596 24092
rect 2648 24080 2654 24132
rect 3068 24120 3096 24160
rect 3234 24148 3240 24160
rect 3292 24148 3298 24200
rect 3421 24191 3479 24197
rect 3421 24157 3433 24191
rect 3467 24188 3479 24191
rect 3786 24188 3792 24200
rect 3467 24160 3792 24188
rect 3467 24157 3479 24160
rect 3421 24151 3479 24157
rect 3786 24148 3792 24160
rect 3844 24188 3850 24200
rect 4264 24188 4292 24296
rect 9214 24284 9220 24296
rect 9272 24284 9278 24336
rect 15746 24284 15752 24336
rect 15804 24284 15810 24336
rect 15838 24284 15844 24336
rect 15896 24324 15902 24336
rect 17954 24324 17960 24336
rect 15896 24296 17960 24324
rect 15896 24284 15902 24296
rect 17954 24284 17960 24296
rect 18012 24324 18018 24336
rect 20438 24324 20444 24336
rect 18012 24296 20444 24324
rect 18012 24284 18018 24296
rect 20438 24284 20444 24296
rect 20496 24324 20502 24336
rect 20640 24324 20668 24364
rect 21174 24324 21180 24336
rect 20496 24296 20668 24324
rect 20824 24296 21180 24324
rect 20496 24284 20502 24296
rect 5077 24259 5135 24265
rect 5077 24256 5089 24259
rect 4356 24228 5089 24256
rect 4356 24197 4384 24228
rect 5077 24225 5089 24228
rect 5123 24225 5135 24259
rect 5077 24219 5135 24225
rect 5166 24216 5172 24268
rect 5224 24256 5230 24268
rect 5445 24259 5503 24265
rect 5445 24256 5457 24259
rect 5224 24228 5457 24256
rect 5224 24216 5230 24228
rect 5445 24225 5457 24228
rect 5491 24225 5503 24259
rect 5445 24219 5503 24225
rect 13446 24216 13452 24268
rect 13504 24256 13510 24268
rect 15764 24256 15792 24284
rect 18046 24256 18052 24268
rect 13504 24228 14780 24256
rect 15764 24228 17080 24256
rect 13504 24216 13510 24228
rect 3844 24160 4292 24188
rect 4341 24191 4399 24197
rect 3844 24148 3850 24160
rect 4341 24157 4353 24191
rect 4387 24157 4399 24191
rect 4341 24151 4399 24157
rect 4430 24148 4436 24200
rect 4488 24188 4494 24200
rect 4488 24160 4533 24188
rect 4488 24148 4494 24160
rect 4706 24148 4712 24200
rect 4764 24188 4770 24200
rect 5261 24191 5319 24197
rect 5261 24188 5273 24191
rect 4764 24160 5273 24188
rect 4764 24148 4770 24160
rect 5261 24157 5273 24160
rect 5307 24157 5319 24191
rect 5261 24151 5319 24157
rect 5353 24191 5411 24197
rect 5353 24157 5365 24191
rect 5399 24157 5411 24191
rect 5353 24151 5411 24157
rect 5537 24191 5595 24197
rect 5537 24157 5549 24191
rect 5583 24188 5595 24191
rect 7190 24188 7196 24200
rect 5583 24160 7196 24188
rect 5583 24157 5595 24160
rect 5537 24151 5595 24157
rect 4154 24120 4160 24132
rect 3068 24092 4160 24120
rect 4154 24080 4160 24092
rect 4212 24080 4218 24132
rect 4246 24080 4252 24132
rect 4304 24120 4310 24132
rect 5368 24120 5396 24151
rect 7190 24148 7196 24160
rect 7248 24148 7254 24200
rect 7561 24191 7619 24197
rect 7561 24157 7573 24191
rect 7607 24157 7619 24191
rect 7561 24151 7619 24157
rect 8481 24191 8539 24197
rect 8481 24157 8493 24191
rect 8527 24188 8539 24191
rect 9306 24188 9312 24200
rect 8527 24160 9312 24188
rect 8527 24157 8539 24160
rect 8481 24151 8539 24157
rect 7282 24120 7288 24132
rect 4304 24092 7288 24120
rect 4304 24080 4310 24092
rect 7282 24080 7288 24092
rect 7340 24080 7346 24132
rect 7576 24064 7604 24151
rect 9306 24148 9312 24160
rect 9364 24148 9370 24200
rect 11974 24188 11980 24200
rect 11935 24160 11980 24188
rect 11974 24148 11980 24160
rect 12032 24148 12038 24200
rect 12161 24191 12219 24197
rect 12161 24157 12173 24191
rect 12207 24188 12219 24191
rect 13078 24188 13084 24200
rect 12207 24160 13084 24188
rect 12207 24157 12219 24160
rect 12161 24151 12219 24157
rect 13078 24148 13084 24160
rect 13136 24148 13142 24200
rect 14461 24191 14519 24197
rect 14461 24157 14473 24191
rect 14507 24157 14519 24191
rect 14461 24151 14519 24157
rect 8294 24080 8300 24132
rect 8352 24120 8358 24132
rect 12250 24120 12256 24132
rect 8352 24092 12256 24120
rect 8352 24080 8358 24092
rect 12250 24080 12256 24092
rect 12308 24080 12314 24132
rect 14476 24120 14504 24151
rect 14550 24148 14556 24200
rect 14608 24188 14614 24200
rect 14752 24197 14780 24228
rect 14737 24191 14795 24197
rect 14608 24160 14653 24188
rect 14608 24148 14614 24160
rect 14737 24157 14749 24191
rect 14783 24157 14795 24191
rect 14737 24151 14795 24157
rect 14826 24148 14832 24200
rect 14884 24188 14890 24200
rect 15749 24191 15807 24197
rect 14884 24160 14929 24188
rect 14884 24148 14890 24160
rect 15749 24157 15761 24191
rect 15795 24157 15807 24191
rect 15930 24188 15936 24200
rect 15891 24160 15936 24188
rect 15749 24151 15807 24157
rect 15654 24120 15660 24132
rect 14476 24092 15660 24120
rect 15654 24080 15660 24092
rect 15712 24080 15718 24132
rect 2409 24055 2467 24061
rect 2409 24021 2421 24055
rect 2455 24052 2467 24055
rect 4890 24052 4896 24064
rect 2455 24024 4896 24052
rect 2455 24021 2467 24024
rect 2409 24015 2467 24021
rect 4890 24012 4896 24024
rect 4948 24052 4954 24064
rect 7558 24052 7564 24064
rect 4948 24024 7564 24052
rect 4948 24012 4954 24024
rect 7558 24012 7564 24024
rect 7616 24012 7622 24064
rect 12161 24055 12219 24061
rect 12161 24021 12173 24055
rect 12207 24052 12219 24055
rect 12618 24052 12624 24064
rect 12207 24024 12624 24052
rect 12207 24021 12219 24024
rect 12161 24015 12219 24021
rect 12618 24012 12624 24024
rect 12676 24012 12682 24064
rect 12894 24012 12900 24064
rect 12952 24052 12958 24064
rect 14277 24055 14335 24061
rect 14277 24052 14289 24055
rect 12952 24024 14289 24052
rect 12952 24012 12958 24024
rect 14277 24021 14289 24024
rect 14323 24021 14335 24055
rect 15562 24052 15568 24064
rect 15523 24024 15568 24052
rect 14277 24015 14335 24021
rect 15562 24012 15568 24024
rect 15620 24012 15626 24064
rect 15761 24052 15789 24151
rect 15930 24148 15936 24160
rect 15988 24148 15994 24200
rect 17052 24197 17080 24228
rect 17880 24228 18052 24256
rect 17880 24197 17908 24228
rect 18046 24216 18052 24228
rect 18104 24216 18110 24268
rect 18230 24216 18236 24268
rect 18288 24256 18294 24268
rect 20824 24256 20852 24296
rect 21174 24284 21180 24296
rect 21232 24284 21238 24336
rect 22741 24327 22799 24333
rect 22741 24293 22753 24327
rect 22787 24324 22799 24327
rect 23474 24324 23480 24336
rect 22787 24296 23480 24324
rect 22787 24293 22799 24296
rect 22741 24287 22799 24293
rect 23474 24284 23480 24296
rect 23532 24284 23538 24336
rect 18288 24228 20852 24256
rect 20901 24259 20959 24265
rect 18288 24216 18294 24228
rect 20901 24225 20913 24259
rect 20947 24256 20959 24259
rect 21082 24256 21088 24268
rect 20947 24228 21088 24256
rect 20947 24225 20959 24228
rect 20901 24219 20959 24225
rect 21082 24216 21088 24228
rect 21140 24216 21146 24268
rect 17037 24191 17095 24197
rect 17037 24157 17049 24191
rect 17083 24157 17095 24191
rect 17037 24151 17095 24157
rect 17221 24191 17279 24197
rect 17221 24157 17233 24191
rect 17267 24157 17279 24191
rect 17221 24151 17279 24157
rect 17865 24191 17923 24197
rect 17865 24157 17877 24191
rect 17911 24157 17923 24191
rect 17865 24151 17923 24157
rect 17236 24120 17264 24151
rect 17954 24148 17960 24200
rect 18012 24188 18018 24200
rect 20364 24197 20576 24198
rect 18141 24191 18199 24197
rect 18141 24188 18153 24191
rect 18012 24160 18153 24188
rect 18012 24148 18018 24160
rect 18141 24157 18153 24160
rect 18187 24157 18199 24191
rect 18141 24151 18199 24157
rect 20364 24191 20591 24197
rect 20364 24170 20545 24191
rect 18049 24123 18107 24129
rect 18049 24120 18061 24123
rect 17236 24092 18061 24120
rect 18049 24089 18061 24092
rect 18095 24120 18107 24123
rect 18690 24120 18696 24132
rect 18095 24092 18696 24120
rect 18095 24089 18107 24092
rect 18049 24083 18107 24089
rect 18690 24080 18696 24092
rect 18748 24080 18754 24132
rect 17129 24055 17187 24061
rect 17129 24052 17141 24055
rect 15761 24024 17141 24052
rect 17129 24021 17141 24024
rect 17175 24052 17187 24055
rect 17402 24052 17408 24064
rect 17175 24024 17408 24052
rect 17175 24021 17187 24024
rect 17129 24015 17187 24021
rect 17402 24012 17408 24024
rect 17460 24012 17466 24064
rect 17586 24012 17592 24064
rect 17644 24052 17650 24064
rect 17681 24055 17739 24061
rect 17681 24052 17693 24055
rect 17644 24024 17693 24052
rect 17644 24012 17650 24024
rect 17681 24021 17693 24024
rect 17727 24021 17739 24055
rect 20364 24052 20392 24170
rect 20533 24157 20545 24170
rect 20579 24157 20591 24191
rect 20533 24151 20591 24157
rect 20714 24148 20720 24200
rect 20772 24188 20778 24200
rect 20772 24160 20817 24188
rect 20772 24148 20778 24160
rect 21192 24120 21220 24284
rect 21266 24148 21272 24200
rect 21324 24188 21330 24200
rect 21361 24191 21419 24197
rect 21361 24188 21373 24191
rect 21324 24160 21373 24188
rect 21324 24148 21330 24160
rect 21361 24157 21373 24160
rect 21407 24157 21419 24191
rect 23382 24188 23388 24200
rect 23295 24160 23388 24188
rect 21361 24151 21419 24157
rect 23382 24148 23388 24160
rect 23440 24148 23446 24200
rect 23676 24197 23704 24364
rect 30374 24352 30380 24404
rect 30432 24392 30438 24404
rect 30469 24395 30527 24401
rect 30469 24392 30481 24395
rect 30432 24364 30481 24392
rect 30432 24352 30438 24364
rect 30469 24361 30481 24364
rect 30515 24361 30527 24395
rect 30469 24355 30527 24361
rect 27522 24256 27528 24268
rect 25240 24228 27528 24256
rect 23661 24191 23719 24197
rect 23661 24157 23673 24191
rect 23707 24157 23719 24191
rect 23661 24151 23719 24157
rect 23750 24148 23756 24200
rect 23808 24188 23814 24200
rect 25240 24197 25268 24228
rect 27522 24216 27528 24228
rect 27580 24216 27586 24268
rect 28718 24216 28724 24268
rect 28776 24256 28782 24268
rect 32306 24256 32312 24268
rect 28776 24228 32312 24256
rect 28776 24216 28782 24228
rect 25225 24191 25283 24197
rect 25225 24188 25237 24191
rect 23808 24160 25237 24188
rect 23808 24148 23814 24160
rect 25225 24157 25237 24160
rect 25271 24157 25283 24191
rect 25225 24151 25283 24157
rect 25409 24191 25467 24197
rect 25409 24157 25421 24191
rect 25455 24188 25467 24191
rect 26694 24188 26700 24200
rect 25455 24160 26700 24188
rect 25455 24157 25467 24160
rect 25409 24151 25467 24157
rect 26694 24148 26700 24160
rect 26752 24148 26758 24200
rect 30653 24191 30711 24197
rect 30653 24157 30665 24191
rect 30699 24188 30711 24191
rect 30834 24188 30840 24200
rect 30699 24160 30840 24188
rect 30699 24157 30711 24160
rect 30653 24151 30711 24157
rect 30834 24148 30840 24160
rect 30892 24148 30898 24200
rect 30939 24191 30997 24197
rect 30939 24157 30951 24191
rect 30985 24188 30997 24191
rect 31036 24188 31064 24228
rect 32306 24216 32312 24228
rect 32364 24216 32370 24268
rect 30985 24160 31064 24188
rect 30985 24157 30997 24160
rect 30939 24151 30997 24157
rect 21628 24123 21686 24129
rect 21192 24092 21312 24120
rect 21174 24052 21180 24064
rect 20364 24024 21180 24052
rect 17681 24015 17739 24021
rect 21174 24012 21180 24024
rect 21232 24012 21238 24064
rect 21284 24052 21312 24092
rect 21628 24089 21640 24123
rect 21674 24120 21686 24123
rect 23201 24123 23259 24129
rect 23201 24120 23213 24123
rect 21674 24092 23213 24120
rect 21674 24089 21686 24092
rect 21628 24083 21686 24089
rect 23201 24089 23213 24092
rect 23247 24089 23259 24123
rect 23400 24120 23428 24148
rect 24486 24120 24492 24132
rect 23400 24092 24492 24120
rect 23201 24083 23259 24089
rect 24486 24080 24492 24092
rect 24544 24120 24550 24132
rect 28994 24120 29000 24132
rect 24544 24092 29000 24120
rect 24544 24080 24550 24092
rect 28994 24080 29000 24092
rect 29052 24080 29058 24132
rect 21726 24052 21732 24064
rect 21284 24024 21732 24052
rect 21726 24012 21732 24024
rect 21784 24052 21790 24064
rect 23474 24052 23480 24064
rect 21784 24024 23480 24052
rect 21784 24012 21790 24024
rect 23474 24012 23480 24024
rect 23532 24012 23538 24064
rect 23569 24055 23627 24061
rect 23569 24021 23581 24055
rect 23615 24052 23627 24055
rect 24670 24052 24676 24064
rect 23615 24024 24676 24052
rect 23615 24021 23627 24024
rect 23569 24015 23627 24021
rect 24670 24012 24676 24024
rect 24728 24012 24734 24064
rect 25222 24052 25228 24064
rect 25183 24024 25228 24052
rect 25222 24012 25228 24024
rect 25280 24012 25286 24064
rect 30837 24055 30895 24061
rect 30837 24021 30849 24055
rect 30883 24052 30895 24055
rect 31478 24052 31484 24064
rect 30883 24024 31484 24052
rect 30883 24021 30895 24024
rect 30837 24015 30895 24021
rect 31478 24012 31484 24024
rect 31536 24012 31542 24064
rect 1104 23962 35027 23984
rect 1104 23910 9390 23962
rect 9442 23910 9454 23962
rect 9506 23910 9518 23962
rect 9570 23910 9582 23962
rect 9634 23910 9646 23962
rect 9698 23910 17831 23962
rect 17883 23910 17895 23962
rect 17947 23910 17959 23962
rect 18011 23910 18023 23962
rect 18075 23910 18087 23962
rect 18139 23910 26272 23962
rect 26324 23910 26336 23962
rect 26388 23910 26400 23962
rect 26452 23910 26464 23962
rect 26516 23910 26528 23962
rect 26580 23910 34713 23962
rect 34765 23910 34777 23962
rect 34829 23910 34841 23962
rect 34893 23910 34905 23962
rect 34957 23910 34969 23962
rect 35021 23910 35027 23962
rect 1104 23888 35027 23910
rect 2590 23808 2596 23860
rect 2648 23848 2654 23860
rect 5077 23851 5135 23857
rect 5077 23848 5089 23851
rect 2648 23820 5089 23848
rect 2648 23808 2654 23820
rect 5077 23817 5089 23820
rect 5123 23817 5135 23851
rect 8294 23848 8300 23860
rect 5077 23811 5135 23817
rect 5276 23820 8300 23848
rect 4338 23780 4344 23792
rect 3344 23752 4344 23780
rect 3344 23721 3372 23752
rect 4338 23740 4344 23752
rect 4396 23740 4402 23792
rect 4522 23740 4528 23792
rect 4580 23780 4586 23792
rect 4617 23783 4675 23789
rect 4617 23780 4629 23783
rect 4580 23752 4629 23780
rect 4580 23740 4586 23752
rect 4617 23749 4629 23752
rect 4663 23749 4675 23783
rect 4617 23743 4675 23749
rect 3329 23715 3387 23721
rect 3329 23681 3341 23715
rect 3375 23681 3387 23715
rect 3329 23675 3387 23681
rect 3418 23672 3424 23724
rect 3476 23712 3482 23724
rect 5276 23721 5304 23820
rect 8294 23808 8300 23820
rect 8352 23808 8358 23860
rect 8389 23851 8447 23857
rect 8389 23817 8401 23851
rect 8435 23848 8447 23851
rect 8570 23848 8576 23860
rect 8435 23820 8576 23848
rect 8435 23817 8447 23820
rect 8389 23811 8447 23817
rect 8570 23808 8576 23820
rect 8628 23848 8634 23860
rect 9398 23848 9404 23860
rect 8628 23820 9404 23848
rect 8628 23808 8634 23820
rect 9398 23808 9404 23820
rect 9456 23808 9462 23860
rect 15105 23851 15163 23857
rect 15105 23817 15117 23851
rect 15151 23848 15163 23851
rect 15378 23848 15384 23860
rect 15151 23820 15384 23848
rect 15151 23817 15163 23820
rect 15105 23811 15163 23817
rect 15378 23808 15384 23820
rect 15436 23848 15442 23860
rect 15933 23851 15991 23857
rect 15933 23848 15945 23851
rect 15436 23820 15945 23848
rect 15436 23808 15442 23820
rect 15933 23817 15945 23820
rect 15979 23817 15991 23851
rect 15933 23811 15991 23817
rect 20622 23808 20628 23860
rect 20680 23848 20686 23860
rect 20680 23820 22094 23848
rect 20680 23808 20686 23820
rect 5460 23752 6914 23780
rect 4065 23715 4123 23721
rect 4065 23712 4077 23715
rect 3476 23684 4077 23712
rect 3476 23672 3482 23684
rect 4065 23681 4077 23684
rect 4111 23712 4123 23715
rect 5261 23715 5319 23721
rect 5261 23712 5273 23715
rect 4111 23684 5273 23712
rect 4111 23681 4123 23684
rect 4065 23675 4123 23681
rect 5261 23681 5273 23684
rect 5307 23681 5319 23715
rect 5460 23712 5488 23752
rect 5261 23675 5319 23681
rect 5368 23684 5488 23712
rect 5537 23715 5595 23721
rect 5368 23653 5396 23684
rect 5537 23681 5549 23715
rect 5583 23712 5595 23715
rect 6730 23712 6736 23724
rect 5583 23684 6736 23712
rect 5583 23681 5595 23684
rect 5537 23675 5595 23681
rect 6730 23672 6736 23684
rect 6788 23672 6794 23724
rect 6886 23712 6914 23752
rect 8478 23740 8484 23792
rect 8536 23780 8542 23792
rect 14642 23780 14648 23792
rect 8536 23752 9904 23780
rect 8536 23740 8542 23752
rect 8938 23712 8944 23724
rect 6886 23684 8944 23712
rect 8938 23672 8944 23684
rect 8996 23672 9002 23724
rect 9214 23712 9220 23724
rect 9175 23684 9220 23712
rect 9214 23672 9220 23684
rect 9272 23672 9278 23724
rect 9876 23721 9904 23752
rect 13004 23752 14648 23780
rect 9861 23715 9919 23721
rect 9861 23681 9873 23715
rect 9907 23681 9919 23715
rect 9861 23675 9919 23681
rect 10045 23715 10103 23721
rect 10045 23681 10057 23715
rect 10091 23681 10103 23715
rect 12894 23712 12900 23724
rect 12855 23684 12900 23712
rect 10045 23675 10103 23681
rect 5353 23647 5411 23653
rect 5353 23613 5365 23647
rect 5399 23613 5411 23647
rect 5353 23607 5411 23613
rect 5445 23647 5503 23653
rect 5445 23613 5457 23647
rect 5491 23644 5503 23647
rect 6638 23644 6644 23656
rect 5491 23616 6644 23644
rect 5491 23613 5503 23616
rect 5445 23607 5503 23613
rect 3234 23536 3240 23588
rect 3292 23576 3298 23588
rect 5368 23576 5396 23607
rect 6638 23604 6644 23616
rect 6696 23604 6702 23656
rect 6825 23647 6883 23653
rect 6825 23613 6837 23647
rect 6871 23613 6883 23647
rect 7098 23644 7104 23656
rect 7059 23616 7104 23644
rect 6825 23607 6883 23613
rect 3292 23548 5396 23576
rect 3292 23536 3298 23548
rect 4062 23468 4068 23520
rect 4120 23508 4126 23520
rect 6840 23508 6868 23607
rect 7098 23604 7104 23616
rect 7156 23604 7162 23656
rect 7466 23604 7472 23656
rect 7524 23644 7530 23656
rect 9033 23647 9091 23653
rect 9033 23644 9045 23647
rect 7524 23616 9045 23644
rect 7524 23604 7530 23616
rect 9033 23613 9045 23616
rect 9079 23613 9091 23647
rect 9398 23644 9404 23656
rect 9359 23616 9404 23644
rect 9033 23607 9091 23613
rect 9398 23604 9404 23616
rect 9456 23604 9462 23656
rect 9953 23579 10011 23585
rect 9953 23576 9965 23579
rect 7760 23548 9965 23576
rect 4120 23480 6868 23508
rect 4120 23468 4126 23480
rect 7282 23468 7288 23520
rect 7340 23508 7346 23520
rect 7760 23508 7788 23548
rect 9953 23545 9965 23548
rect 9999 23545 10011 23579
rect 9953 23539 10011 23545
rect 7340 23480 7788 23508
rect 7340 23468 7346 23480
rect 8294 23468 8300 23520
rect 8352 23508 8358 23520
rect 10060 23508 10088 23675
rect 12894 23672 12900 23684
rect 12952 23672 12958 23724
rect 12250 23644 12256 23656
rect 12211 23616 12256 23644
rect 12250 23604 12256 23616
rect 12308 23604 12314 23656
rect 13004 23653 13032 23752
rect 14642 23740 14648 23752
rect 14700 23740 14706 23792
rect 14921 23783 14979 23789
rect 14921 23749 14933 23783
rect 14967 23780 14979 23783
rect 15194 23780 15200 23792
rect 14967 23752 15200 23780
rect 14967 23749 14979 23752
rect 14921 23743 14979 23749
rect 15194 23740 15200 23752
rect 15252 23740 15258 23792
rect 19981 23783 20039 23789
rect 19981 23749 19993 23783
rect 20027 23780 20039 23783
rect 20898 23780 20904 23792
rect 20027 23752 20904 23780
rect 20027 23749 20039 23752
rect 19981 23743 20039 23749
rect 20898 23740 20904 23752
rect 20956 23780 20962 23792
rect 21910 23780 21916 23792
rect 20956 23752 21916 23780
rect 20956 23740 20962 23752
rect 21910 23740 21916 23752
rect 21968 23740 21974 23792
rect 22066 23780 22094 23820
rect 23474 23808 23480 23860
rect 23532 23848 23538 23860
rect 29270 23848 29276 23860
rect 23532 23820 29276 23848
rect 23532 23808 23538 23820
rect 29270 23808 29276 23820
rect 29328 23808 29334 23860
rect 30098 23848 30104 23860
rect 30059 23820 30104 23848
rect 30098 23808 30104 23820
rect 30156 23808 30162 23860
rect 22281 23783 22339 23789
rect 22281 23780 22293 23783
rect 22066 23752 22293 23780
rect 22281 23749 22293 23752
rect 22327 23780 22339 23783
rect 23750 23780 23756 23792
rect 22327 23752 23756 23780
rect 22327 23749 22339 23752
rect 22281 23743 22339 23749
rect 23750 23740 23756 23752
rect 23808 23740 23814 23792
rect 28626 23780 28632 23792
rect 28587 23752 28632 23780
rect 28626 23740 28632 23752
rect 28684 23740 28690 23792
rect 13078 23672 13084 23724
rect 13136 23712 13142 23724
rect 13265 23715 13323 23721
rect 13265 23712 13277 23715
rect 13136 23684 13277 23712
rect 13136 23672 13142 23684
rect 13265 23681 13277 23684
rect 13311 23681 13323 23715
rect 13265 23675 13323 23681
rect 14369 23715 14427 23721
rect 14369 23681 14381 23715
rect 14415 23712 14427 23715
rect 15562 23712 15568 23724
rect 14415 23684 15568 23712
rect 14415 23681 14427 23684
rect 14369 23675 14427 23681
rect 15562 23672 15568 23684
rect 15620 23672 15626 23724
rect 15930 23672 15936 23724
rect 15988 23712 15994 23724
rect 16117 23715 16175 23721
rect 16117 23712 16129 23715
rect 15988 23684 16129 23712
rect 15988 23672 15994 23684
rect 16117 23681 16129 23684
rect 16163 23681 16175 23715
rect 16117 23675 16175 23681
rect 16301 23715 16359 23721
rect 16301 23681 16313 23715
rect 16347 23712 16359 23715
rect 17402 23712 17408 23724
rect 16347 23684 17408 23712
rect 16347 23681 16359 23684
rect 16301 23675 16359 23681
rect 17402 23672 17408 23684
rect 17460 23672 17466 23724
rect 20530 23712 20536 23724
rect 20491 23684 20536 23712
rect 20530 23672 20536 23684
rect 20588 23672 20594 23724
rect 20714 23672 20720 23724
rect 20772 23712 20778 23724
rect 22649 23715 22707 23721
rect 20772 23684 22600 23712
rect 20772 23672 20778 23684
rect 12989 23647 13047 23653
rect 12989 23613 13001 23647
rect 13035 23613 13047 23647
rect 13170 23644 13176 23656
rect 13131 23616 13176 23644
rect 12989 23607 13047 23613
rect 13170 23604 13176 23616
rect 13228 23604 13234 23656
rect 14734 23604 14740 23656
rect 14792 23644 14798 23656
rect 14829 23647 14887 23653
rect 14829 23644 14841 23647
rect 14792 23616 14841 23644
rect 14792 23604 14798 23616
rect 14829 23613 14841 23616
rect 14875 23613 14887 23647
rect 14829 23607 14887 23613
rect 15197 23647 15255 23653
rect 15197 23613 15209 23647
rect 15243 23613 15255 23647
rect 15197 23607 15255 23613
rect 14277 23579 14335 23585
rect 14277 23545 14289 23579
rect 14323 23576 14335 23579
rect 15212 23576 15240 23607
rect 15286 23604 15292 23656
rect 15344 23644 15350 23656
rect 18414 23644 18420 23656
rect 15344 23616 18420 23644
rect 15344 23604 15350 23616
rect 18414 23604 18420 23616
rect 18472 23604 18478 23656
rect 20806 23644 20812 23656
rect 20767 23616 20812 23644
rect 20806 23604 20812 23616
rect 20864 23604 20870 23656
rect 22572 23644 22600 23684
rect 22649 23681 22661 23715
rect 22695 23712 22707 23715
rect 23658 23712 23664 23724
rect 22695 23684 23664 23712
rect 22695 23681 22707 23684
rect 22649 23675 22707 23681
rect 23658 23672 23664 23684
rect 23716 23672 23722 23724
rect 27154 23644 27160 23656
rect 22572 23616 27160 23644
rect 27154 23604 27160 23616
rect 27212 23604 27218 23656
rect 14323 23548 15240 23576
rect 14323 23545 14335 23548
rect 14277 23539 14335 23545
rect 8352 23480 10088 23508
rect 15212 23508 15240 23548
rect 15473 23579 15531 23585
rect 15473 23545 15485 23579
rect 15519 23576 15531 23579
rect 16574 23576 16580 23588
rect 15519 23548 16580 23576
rect 15519 23545 15531 23548
rect 15473 23539 15531 23545
rect 16574 23536 16580 23548
rect 16632 23536 16638 23588
rect 18693 23579 18751 23585
rect 18693 23545 18705 23579
rect 18739 23576 18751 23579
rect 19702 23576 19708 23588
rect 18739 23548 19708 23576
rect 18739 23545 18751 23548
rect 18693 23539 18751 23545
rect 19702 23536 19708 23548
rect 19760 23536 19766 23588
rect 20070 23536 20076 23588
rect 20128 23576 20134 23588
rect 28810 23576 28816 23588
rect 20128 23548 28816 23576
rect 20128 23536 20134 23548
rect 28810 23536 28816 23548
rect 28868 23536 28874 23588
rect 15286 23508 15292 23520
rect 15212 23480 15292 23508
rect 8352 23468 8358 23480
rect 15286 23468 15292 23480
rect 15344 23468 15350 23520
rect 24946 23468 24952 23520
rect 25004 23508 25010 23520
rect 25958 23508 25964 23520
rect 25004 23480 25964 23508
rect 25004 23468 25010 23480
rect 25958 23468 25964 23480
rect 26016 23468 26022 23520
rect 1104 23418 34868 23440
rect 1104 23366 5170 23418
rect 5222 23366 5234 23418
rect 5286 23366 5298 23418
rect 5350 23366 5362 23418
rect 5414 23366 5426 23418
rect 5478 23366 13611 23418
rect 13663 23366 13675 23418
rect 13727 23366 13739 23418
rect 13791 23366 13803 23418
rect 13855 23366 13867 23418
rect 13919 23366 22052 23418
rect 22104 23366 22116 23418
rect 22168 23366 22180 23418
rect 22232 23366 22244 23418
rect 22296 23366 22308 23418
rect 22360 23366 30493 23418
rect 30545 23366 30557 23418
rect 30609 23366 30621 23418
rect 30673 23366 30685 23418
rect 30737 23366 30749 23418
rect 30801 23366 34868 23418
rect 1104 23344 34868 23366
rect 3329 23307 3387 23313
rect 3329 23273 3341 23307
rect 3375 23304 3387 23307
rect 4154 23304 4160 23316
rect 3375 23276 4160 23304
rect 3375 23273 3387 23276
rect 3329 23267 3387 23273
rect 4154 23264 4160 23276
rect 4212 23264 4218 23316
rect 6917 23307 6975 23313
rect 6917 23273 6929 23307
rect 6963 23304 6975 23307
rect 7098 23304 7104 23316
rect 6963 23276 7104 23304
rect 6963 23273 6975 23276
rect 6917 23267 6975 23273
rect 7098 23264 7104 23276
rect 7156 23264 7162 23316
rect 7558 23264 7564 23316
rect 7616 23304 7622 23316
rect 7616 23276 9260 23304
rect 7616 23264 7622 23276
rect 4430 23196 4436 23248
rect 4488 23236 4494 23248
rect 4617 23239 4675 23245
rect 4617 23236 4629 23239
rect 4488 23208 4629 23236
rect 4488 23196 4494 23208
rect 4617 23205 4629 23208
rect 4663 23205 4675 23239
rect 4617 23199 4675 23205
rect 6638 23196 6644 23248
rect 6696 23236 6702 23248
rect 8570 23236 8576 23248
rect 6696 23208 6914 23236
rect 6696 23196 6702 23208
rect 4157 23171 4215 23177
rect 4157 23137 4169 23171
rect 4203 23168 4215 23171
rect 4246 23168 4252 23180
rect 4203 23140 4252 23168
rect 4203 23137 4215 23140
rect 4157 23131 4215 23137
rect 4246 23128 4252 23140
rect 4304 23128 4310 23180
rect 4706 23168 4712 23180
rect 4667 23140 4712 23168
rect 4706 23128 4712 23140
rect 4764 23128 4770 23180
rect 6886 23168 6914 23208
rect 8312 23208 8576 23236
rect 8312 23177 8340 23208
rect 8570 23196 8576 23208
rect 8628 23196 8634 23248
rect 9125 23239 9183 23245
rect 9125 23205 9137 23239
rect 9171 23205 9183 23239
rect 9125 23199 9183 23205
rect 8205 23171 8263 23177
rect 8205 23168 8217 23171
rect 6886 23140 8217 23168
rect 8205 23137 8217 23140
rect 8251 23137 8263 23171
rect 8205 23131 8263 23137
rect 8297 23171 8355 23177
rect 8297 23137 8309 23171
rect 8343 23137 8355 23171
rect 8297 23131 8355 23137
rect 8389 23171 8447 23177
rect 8389 23137 8401 23171
rect 8435 23168 8447 23171
rect 8846 23168 8852 23180
rect 8435 23140 8852 23168
rect 8435 23137 8447 23140
rect 8389 23131 8447 23137
rect 8846 23128 8852 23140
rect 8904 23128 8910 23180
rect 3418 23100 3424 23112
rect 3379 23072 3424 23100
rect 3418 23060 3424 23072
rect 3476 23060 3482 23112
rect 4341 23103 4399 23109
rect 4341 23069 4353 23103
rect 4387 23100 4399 23103
rect 5074 23100 5080 23112
rect 4387 23072 5080 23100
rect 4387 23069 4399 23072
rect 4341 23063 4399 23069
rect 5074 23060 5080 23072
rect 5132 23060 5138 23112
rect 7098 23100 7104 23112
rect 7059 23072 7104 23100
rect 7098 23060 7104 23072
rect 7156 23060 7162 23112
rect 7282 23100 7288 23112
rect 7243 23072 7288 23100
rect 7282 23060 7288 23072
rect 7340 23060 7346 23112
rect 7558 23100 7564 23112
rect 7519 23072 7564 23100
rect 7558 23060 7564 23072
rect 7616 23060 7622 23112
rect 8110 23100 8116 23112
rect 8071 23072 8116 23100
rect 8110 23060 8116 23072
rect 8168 23060 8174 23112
rect 9140 23100 9168 23199
rect 8496 23072 9168 23100
rect 7006 22992 7012 23044
rect 7064 23032 7070 23044
rect 7193 23035 7251 23041
rect 7193 23032 7205 23035
rect 7064 23004 7205 23032
rect 7064 22992 7070 23004
rect 7193 23001 7205 23004
rect 7239 23001 7251 23035
rect 7193 22995 7251 23001
rect 7423 23035 7481 23041
rect 7423 23001 7435 23035
rect 7469 23032 7481 23035
rect 8496 23032 8524 23072
rect 7469 23004 8524 23032
rect 9125 23035 9183 23041
rect 7469 23001 7481 23004
rect 7423 22995 7481 23001
rect 9125 23001 9137 23035
rect 9171 23001 9183 23035
rect 9125 22995 9183 23001
rect 7208 22964 7236 22995
rect 8110 22964 8116 22976
rect 7208 22936 8116 22964
rect 8110 22924 8116 22936
rect 8168 22924 8174 22976
rect 8573 22967 8631 22973
rect 8573 22933 8585 22967
rect 8619 22964 8631 22967
rect 9140 22964 9168 22995
rect 8619 22936 9168 22964
rect 9232 22964 9260 23276
rect 9398 23264 9404 23316
rect 9456 23304 9462 23316
rect 9858 23304 9864 23316
rect 9456 23276 9864 23304
rect 9456 23264 9462 23276
rect 9858 23264 9864 23276
rect 9916 23304 9922 23316
rect 13998 23304 14004 23316
rect 9916 23276 14004 23304
rect 9916 23264 9922 23276
rect 13998 23264 14004 23276
rect 14056 23264 14062 23316
rect 18690 23304 18696 23316
rect 18651 23276 18696 23304
rect 18690 23264 18696 23276
rect 18748 23264 18754 23316
rect 21910 23304 21916 23316
rect 21871 23276 21916 23304
rect 21910 23264 21916 23276
rect 21968 23264 21974 23316
rect 15657 23239 15715 23245
rect 15657 23205 15669 23239
rect 15703 23236 15715 23239
rect 16209 23239 16267 23245
rect 16209 23236 16221 23239
rect 15703 23208 16221 23236
rect 15703 23205 15715 23208
rect 15657 23199 15715 23205
rect 16209 23205 16221 23208
rect 16255 23205 16267 23239
rect 16209 23199 16267 23205
rect 19610 23196 19616 23248
rect 19668 23236 19674 23248
rect 19705 23239 19763 23245
rect 19705 23236 19717 23239
rect 19668 23208 19717 23236
rect 19668 23196 19674 23208
rect 19705 23205 19717 23208
rect 19751 23205 19763 23239
rect 19705 23199 19763 23205
rect 24670 23196 24676 23248
rect 24728 23236 24734 23248
rect 24728 23208 25544 23236
rect 24728 23196 24734 23208
rect 15286 23168 15292 23180
rect 15247 23140 15292 23168
rect 15286 23128 15292 23140
rect 15344 23128 15350 23180
rect 15378 23128 15384 23180
rect 15436 23168 15442 23180
rect 16574 23168 16580 23180
rect 15436 23140 15481 23168
rect 16535 23140 16580 23168
rect 15436 23128 15442 23140
rect 16574 23128 16580 23140
rect 16632 23128 16638 23180
rect 17310 23168 17316 23180
rect 17271 23140 17316 23168
rect 17310 23128 17316 23140
rect 17368 23128 17374 23180
rect 25222 23168 25228 23180
rect 25183 23140 25228 23168
rect 25222 23128 25228 23140
rect 25280 23128 25286 23180
rect 25516 23168 25544 23208
rect 25516 23140 25912 23168
rect 9306 23060 9312 23112
rect 9364 23100 9370 23112
rect 9401 23103 9459 23109
rect 9401 23100 9413 23103
rect 9364 23072 9413 23100
rect 9364 23060 9370 23072
rect 9401 23069 9413 23072
rect 9447 23069 9459 23103
rect 9401 23063 9459 23069
rect 12066 23060 12072 23112
rect 12124 23100 12130 23112
rect 12124 23072 12169 23100
rect 12124 23060 12130 23072
rect 14734 23060 14740 23112
rect 14792 23060 14798 23112
rect 15194 23100 15200 23112
rect 15155 23072 15200 23100
rect 15194 23060 15200 23072
rect 15252 23060 15258 23112
rect 17586 23109 17592 23112
rect 15473 23103 15531 23109
rect 15473 23069 15485 23103
rect 15519 23069 15531 23103
rect 17580 23100 17592 23109
rect 17547 23072 17592 23100
rect 15473 23063 15531 23069
rect 17580 23063 17592 23072
rect 9766 22992 9772 23044
rect 9824 23032 9830 23044
rect 11793 23035 11851 23041
rect 9824 23004 10626 23032
rect 9824 22992 9830 23004
rect 11793 23001 11805 23035
rect 11839 23032 11851 23035
rect 11882 23032 11888 23044
rect 11839 23004 11888 23032
rect 11839 23001 11851 23004
rect 11793 22995 11851 23001
rect 11882 22992 11888 23004
rect 11940 22992 11946 23044
rect 12434 22992 12440 23044
rect 12492 23032 12498 23044
rect 12529 23035 12587 23041
rect 12529 23032 12541 23035
rect 12492 23004 12541 23032
rect 12492 22992 12498 23004
rect 12529 23001 12541 23004
rect 12575 23001 12587 23035
rect 12529 22995 12587 23001
rect 13265 23035 13323 23041
rect 13265 23001 13277 23035
rect 13311 23001 13323 23035
rect 14752 23032 14780 23060
rect 15488 23032 15516 23063
rect 17586 23060 17592 23063
rect 17644 23060 17650 23112
rect 19426 23100 19432 23112
rect 19387 23072 19432 23100
rect 19426 23060 19432 23072
rect 19484 23060 19490 23112
rect 19702 23100 19708 23112
rect 19663 23072 19708 23100
rect 19702 23060 19708 23072
rect 19760 23060 19766 23112
rect 20625 23103 20683 23109
rect 20625 23069 20637 23103
rect 20671 23100 20683 23103
rect 20806 23100 20812 23112
rect 20671 23072 20812 23100
rect 20671 23069 20683 23072
rect 20625 23063 20683 23069
rect 20806 23060 20812 23072
rect 20864 23060 20870 23112
rect 20990 23060 20996 23112
rect 21048 23100 21054 23112
rect 25884 23109 25912 23140
rect 27706 23128 27712 23180
rect 27764 23168 27770 23180
rect 28721 23171 28779 23177
rect 28721 23168 28733 23171
rect 27764 23140 28733 23168
rect 27764 23128 27770 23140
rect 28721 23137 28733 23140
rect 28767 23168 28779 23171
rect 31021 23171 31079 23177
rect 31021 23168 31033 23171
rect 28767 23140 31033 23168
rect 28767 23137 28779 23140
rect 28721 23131 28779 23137
rect 31021 23137 31033 23140
rect 31067 23137 31079 23171
rect 32674 23168 32680 23180
rect 32635 23140 32680 23168
rect 31021 23131 31079 23137
rect 32674 23128 32680 23140
rect 32732 23128 32738 23180
rect 33134 23168 33140 23180
rect 33047 23140 33140 23168
rect 33134 23128 33140 23140
rect 33192 23168 33198 23180
rect 33192 23140 33824 23168
rect 33192 23128 33198 23140
rect 24765 23103 24823 23109
rect 24765 23100 24777 23103
rect 21048 23072 24777 23100
rect 21048 23060 21054 23072
rect 24765 23069 24777 23072
rect 24811 23069 24823 23103
rect 24765 23063 24823 23069
rect 24857 23103 24915 23109
rect 24857 23069 24869 23103
rect 24903 23100 24915 23103
rect 25777 23103 25835 23109
rect 25777 23100 25789 23103
rect 24903 23072 25789 23100
rect 24903 23069 24915 23072
rect 24857 23063 24915 23069
rect 25777 23069 25789 23072
rect 25823 23069 25835 23103
rect 25777 23063 25835 23069
rect 25869 23103 25927 23109
rect 25869 23069 25881 23103
rect 25915 23069 25927 23103
rect 27522 23100 27528 23112
rect 27483 23072 27528 23100
rect 25869 23063 25927 23069
rect 27522 23060 27528 23072
rect 27580 23060 27586 23112
rect 27982 23100 27988 23112
rect 27943 23072 27988 23100
rect 27982 23060 27988 23072
rect 28040 23060 28046 23112
rect 28258 23100 28264 23112
rect 28219 23072 28264 23100
rect 28258 23060 28264 23072
rect 28316 23060 28322 23112
rect 28905 23103 28963 23109
rect 28905 23069 28917 23103
rect 28951 23069 28963 23103
rect 31754 23100 31760 23112
rect 31715 23072 31760 23100
rect 28905 23063 28963 23069
rect 17494 23032 17500 23044
rect 14752 23004 17500 23032
rect 13265 22995 13323 23001
rect 9309 22967 9367 22973
rect 9309 22964 9321 22967
rect 9232 22936 9321 22964
rect 8619 22933 8631 22936
rect 8573 22927 8631 22933
rect 9309 22933 9321 22936
rect 9355 22964 9367 22967
rect 10134 22964 10140 22976
rect 9355 22936 10140 22964
rect 9355 22933 9367 22936
rect 9309 22927 9367 22933
rect 10134 22924 10140 22936
rect 10192 22924 10198 22976
rect 10318 22964 10324 22976
rect 10279 22936 10324 22964
rect 10318 22924 10324 22936
rect 10376 22924 10382 22976
rect 10410 22924 10416 22976
rect 10468 22964 10474 22976
rect 12802 22964 12808 22976
rect 10468 22936 12808 22964
rect 10468 22924 10474 22936
rect 12802 22924 12808 22936
rect 12860 22964 12866 22976
rect 13280 22964 13308 22995
rect 17494 22992 17500 23004
rect 17552 22992 17558 23044
rect 24581 23035 24639 23041
rect 24581 23001 24593 23035
rect 24627 23032 24639 23035
rect 25314 23032 25320 23044
rect 24627 23004 25320 23032
rect 24627 23001 24639 23004
rect 24581 22995 24639 23001
rect 25314 22992 25320 23004
rect 25372 22992 25378 23044
rect 27614 22992 27620 23044
rect 27672 23032 27678 23044
rect 27801 23035 27859 23041
rect 27801 23032 27813 23035
rect 27672 23004 27813 23032
rect 27672 22992 27678 23004
rect 27801 23001 27813 23004
rect 27847 23032 27859 23035
rect 28920 23032 28948 23063
rect 31754 23060 31760 23072
rect 31812 23060 31818 23112
rect 32030 23100 32036 23112
rect 31991 23072 32036 23100
rect 32030 23060 32036 23072
rect 32088 23060 32094 23112
rect 32398 23060 32404 23112
rect 32456 23100 32462 23112
rect 32769 23103 32827 23109
rect 32769 23100 32781 23103
rect 32456 23072 32781 23100
rect 32456 23060 32462 23072
rect 32769 23069 32781 23072
rect 32815 23069 32827 23103
rect 32769 23063 32827 23069
rect 33318 23060 33324 23112
rect 33376 23100 33382 23112
rect 33796 23109 33824 23140
rect 33597 23103 33655 23109
rect 33597 23100 33609 23103
rect 33376 23072 33609 23100
rect 33376 23060 33382 23072
rect 33597 23069 33609 23072
rect 33643 23069 33655 23103
rect 33597 23063 33655 23069
rect 33781 23103 33839 23109
rect 33781 23069 33793 23103
rect 33827 23069 33839 23103
rect 33781 23063 33839 23069
rect 27847 23004 28948 23032
rect 29089 23035 29147 23041
rect 27847 23001 27859 23004
rect 27801 22995 27859 23001
rect 29089 23001 29101 23035
rect 29135 23032 29147 23035
rect 31294 23032 31300 23044
rect 29135 23004 31300 23032
rect 29135 23001 29147 23004
rect 29089 22995 29147 23001
rect 31294 22992 31300 23004
rect 31352 22992 31358 23044
rect 12860 22936 13308 22964
rect 12860 22924 12866 22936
rect 14734 22924 14740 22976
rect 14792 22964 14798 22976
rect 16117 22967 16175 22973
rect 16117 22964 16129 22967
rect 14792 22936 16129 22964
rect 14792 22924 14798 22936
rect 16117 22933 16129 22936
rect 16163 22933 16175 22967
rect 16117 22927 16175 22933
rect 18506 22924 18512 22976
rect 18564 22964 18570 22976
rect 20622 22964 20628 22976
rect 18564 22936 20628 22964
rect 18564 22924 18570 22936
rect 20622 22924 20628 22936
rect 20680 22924 20686 22976
rect 24854 22924 24860 22976
rect 24912 22964 24918 22976
rect 24949 22967 25007 22973
rect 24949 22964 24961 22967
rect 24912 22936 24961 22964
rect 24912 22924 24918 22936
rect 24949 22933 24961 22936
rect 24995 22933 25007 22967
rect 25130 22964 25136 22976
rect 25091 22936 25136 22964
rect 24949 22927 25007 22933
rect 25130 22924 25136 22936
rect 25188 22924 25194 22976
rect 31110 22924 31116 22976
rect 31168 22964 31174 22976
rect 33226 22964 33232 22976
rect 31168 22936 33232 22964
rect 31168 22924 31174 22936
rect 33226 22924 33232 22936
rect 33284 22924 33290 22976
rect 33502 22924 33508 22976
rect 33560 22964 33566 22976
rect 33689 22967 33747 22973
rect 33689 22964 33701 22967
rect 33560 22936 33701 22964
rect 33560 22924 33566 22936
rect 33689 22933 33701 22936
rect 33735 22933 33747 22967
rect 33689 22927 33747 22933
rect 1104 22874 35027 22896
rect 1104 22822 9390 22874
rect 9442 22822 9454 22874
rect 9506 22822 9518 22874
rect 9570 22822 9582 22874
rect 9634 22822 9646 22874
rect 9698 22822 17831 22874
rect 17883 22822 17895 22874
rect 17947 22822 17959 22874
rect 18011 22822 18023 22874
rect 18075 22822 18087 22874
rect 18139 22822 26272 22874
rect 26324 22822 26336 22874
rect 26388 22822 26400 22874
rect 26452 22822 26464 22874
rect 26516 22822 26528 22874
rect 26580 22822 34713 22874
rect 34765 22822 34777 22874
rect 34829 22822 34841 22874
rect 34893 22822 34905 22874
rect 34957 22822 34969 22874
rect 35021 22822 35027 22874
rect 1104 22800 35027 22822
rect 3773 22763 3831 22769
rect 3773 22729 3785 22763
rect 3819 22760 3831 22763
rect 4522 22760 4528 22772
rect 3819 22732 4528 22760
rect 3819 22729 3831 22732
rect 3773 22723 3831 22729
rect 4522 22720 4528 22732
rect 4580 22720 4586 22772
rect 7193 22763 7251 22769
rect 7193 22729 7205 22763
rect 7239 22760 7251 22763
rect 7558 22760 7564 22772
rect 7239 22732 7564 22760
rect 7239 22729 7251 22732
rect 7193 22723 7251 22729
rect 7558 22720 7564 22732
rect 7616 22720 7622 22772
rect 12434 22760 12440 22772
rect 9324 22732 12440 22760
rect 3234 22652 3240 22704
rect 3292 22692 3298 22704
rect 3973 22695 4031 22701
rect 3973 22692 3985 22695
rect 3292 22664 3985 22692
rect 3292 22652 3298 22664
rect 3973 22661 3985 22664
rect 4019 22661 4031 22695
rect 3973 22655 4031 22661
rect 7098 22652 7104 22704
rect 7156 22692 7162 22704
rect 8113 22695 8171 22701
rect 8113 22692 8125 22695
rect 7156 22664 8125 22692
rect 7156 22652 7162 22664
rect 8113 22661 8125 22664
rect 8159 22661 8171 22695
rect 8294 22692 8300 22704
rect 8255 22664 8300 22692
rect 8113 22655 8171 22661
rect 8294 22652 8300 22664
rect 8352 22652 8358 22704
rect 8478 22692 8484 22704
rect 8439 22664 8484 22692
rect 8478 22652 8484 22664
rect 8536 22652 8542 22704
rect 4890 22624 4896 22636
rect 4851 22596 4896 22624
rect 4890 22584 4896 22596
rect 4948 22584 4954 22636
rect 7377 22627 7435 22633
rect 7377 22593 7389 22627
rect 7423 22624 7435 22627
rect 7466 22624 7472 22636
rect 7423 22596 7472 22624
rect 7423 22593 7435 22596
rect 7377 22587 7435 22593
rect 7466 22584 7472 22596
rect 7524 22584 7530 22636
rect 7561 22627 7619 22633
rect 7561 22593 7573 22627
rect 7607 22593 7619 22627
rect 7561 22587 7619 22593
rect 7653 22627 7711 22633
rect 7653 22593 7665 22627
rect 7699 22624 7711 22627
rect 8846 22624 8852 22636
rect 7699 22596 8852 22624
rect 7699 22593 7711 22596
rect 7653 22587 7711 22593
rect 7576 22556 7604 22587
rect 8846 22584 8852 22596
rect 8904 22584 8910 22636
rect 4632 22528 7604 22556
rect 4632 22432 4660 22528
rect 4982 22448 4988 22500
rect 5040 22488 5046 22500
rect 9324 22488 9352 22732
rect 12434 22720 12440 22732
rect 12492 22720 12498 22772
rect 31110 22760 31116 22772
rect 14568 22732 31116 22760
rect 9677 22695 9735 22701
rect 9677 22661 9689 22695
rect 9723 22692 9735 22695
rect 9766 22692 9772 22704
rect 9723 22664 9772 22692
rect 9723 22661 9735 22664
rect 9677 22655 9735 22661
rect 9766 22652 9772 22664
rect 9824 22652 9830 22704
rect 12529 22695 12587 22701
rect 12529 22692 12541 22695
rect 9876 22664 12541 22692
rect 9401 22627 9459 22633
rect 9401 22593 9413 22627
rect 9447 22593 9459 22627
rect 9401 22587 9459 22593
rect 9493 22627 9551 22633
rect 9493 22593 9505 22627
rect 9539 22593 9551 22627
rect 9493 22587 9551 22593
rect 5040 22460 9352 22488
rect 9416 22488 9444 22587
rect 9508 22556 9536 22587
rect 9582 22584 9588 22636
rect 9640 22624 9646 22636
rect 9876 22624 9904 22664
rect 12529 22661 12541 22664
rect 12575 22661 12587 22695
rect 14461 22695 14519 22701
rect 14461 22692 14473 22695
rect 12529 22655 12587 22661
rect 13188 22664 14473 22692
rect 9640 22596 9904 22624
rect 10321 22627 10379 22633
rect 9640 22584 9646 22596
rect 10321 22593 10333 22627
rect 10367 22624 10379 22627
rect 10410 22624 10416 22636
rect 10367 22596 10416 22624
rect 10367 22593 10379 22596
rect 10321 22587 10379 22593
rect 10410 22584 10416 22596
rect 10468 22584 10474 22636
rect 11698 22624 11704 22636
rect 11659 22596 11704 22624
rect 11698 22584 11704 22596
rect 11756 22584 11762 22636
rect 11885 22627 11943 22633
rect 11885 22593 11897 22627
rect 11931 22593 11943 22627
rect 11885 22587 11943 22593
rect 10965 22559 11023 22565
rect 10965 22556 10977 22559
rect 9508 22528 10977 22556
rect 10965 22525 10977 22528
rect 11011 22556 11023 22559
rect 11790 22556 11796 22568
rect 11011 22528 11796 22556
rect 11011 22525 11023 22528
rect 10965 22519 11023 22525
rect 11790 22516 11796 22528
rect 11848 22516 11854 22568
rect 11900 22556 11928 22587
rect 12618 22584 12624 22636
rect 12676 22624 12682 22636
rect 13188 22633 13216 22664
rect 14461 22661 14473 22664
rect 14507 22661 14519 22695
rect 14461 22655 14519 22661
rect 12897 22627 12955 22633
rect 12897 22624 12909 22627
rect 12676 22596 12909 22624
rect 12676 22584 12682 22596
rect 12897 22593 12909 22596
rect 12943 22593 12955 22627
rect 12897 22587 12955 22593
rect 13173 22627 13231 22633
rect 13173 22593 13185 22627
rect 13219 22593 13231 22627
rect 13173 22587 13231 22593
rect 13262 22584 13268 22636
rect 13320 22624 13326 22636
rect 13357 22627 13415 22633
rect 13357 22624 13369 22627
rect 13320 22596 13369 22624
rect 13320 22584 13326 22596
rect 13357 22593 13369 22596
rect 13403 22593 13415 22627
rect 13357 22587 13415 22593
rect 13633 22627 13691 22633
rect 13633 22593 13645 22627
rect 13679 22593 13691 22627
rect 13633 22587 13691 22593
rect 13909 22627 13967 22633
rect 13909 22593 13921 22627
rect 13955 22624 13967 22627
rect 14568 22624 14596 22732
rect 31110 22720 31116 22732
rect 31168 22720 31174 22772
rect 32030 22720 32036 22772
rect 32088 22760 32094 22772
rect 32401 22763 32459 22769
rect 32401 22760 32413 22763
rect 32088 22732 32413 22760
rect 32088 22720 32094 22732
rect 32401 22729 32413 22732
rect 32447 22729 32459 22763
rect 32401 22723 32459 22729
rect 15470 22652 15476 22704
rect 15528 22692 15534 22704
rect 15565 22695 15623 22701
rect 15565 22692 15577 22695
rect 15528 22664 15577 22692
rect 15528 22652 15534 22664
rect 15565 22661 15577 22664
rect 15611 22661 15623 22695
rect 18506 22692 18512 22704
rect 15565 22655 15623 22661
rect 18340 22664 18512 22692
rect 14734 22624 14740 22636
rect 13955 22596 14596 22624
rect 14695 22596 14740 22624
rect 13955 22593 13967 22596
rect 13909 22587 13967 22593
rect 12710 22556 12716 22568
rect 11900 22528 12716 22556
rect 12710 22516 12716 22528
rect 12768 22556 12774 22568
rect 13078 22556 13084 22568
rect 12768 22528 13084 22556
rect 12768 22516 12774 22528
rect 13078 22516 13084 22528
rect 13136 22556 13142 22568
rect 13648 22556 13676 22587
rect 14734 22584 14740 22596
rect 14792 22584 14798 22636
rect 15381 22627 15439 22633
rect 15381 22593 15393 22627
rect 15427 22593 15439 22627
rect 15654 22624 15660 22636
rect 15615 22596 15660 22624
rect 15381 22587 15439 22593
rect 13136 22528 13676 22556
rect 13136 22516 13142 22528
rect 14090 22516 14096 22568
rect 14148 22556 14154 22568
rect 14461 22559 14519 22565
rect 14461 22556 14473 22559
rect 14148 22528 14473 22556
rect 14148 22516 14154 22528
rect 14461 22525 14473 22528
rect 14507 22556 14519 22559
rect 14642 22556 14648 22568
rect 14507 22528 14648 22556
rect 14507 22525 14519 22528
rect 14461 22519 14519 22525
rect 14642 22516 14648 22528
rect 14700 22516 14706 22568
rect 15396 22556 15424 22587
rect 15654 22584 15660 22596
rect 15712 22624 15718 22636
rect 16390 22624 16396 22636
rect 15712 22596 16396 22624
rect 15712 22584 15718 22596
rect 16390 22584 16396 22596
rect 16448 22584 16454 22636
rect 17402 22624 17408 22636
rect 17363 22596 17408 22624
rect 17402 22584 17408 22596
rect 17460 22584 17466 22636
rect 17494 22584 17500 22636
rect 17552 22624 17558 22636
rect 18340 22633 18368 22664
rect 18506 22652 18512 22664
rect 18564 22652 18570 22704
rect 18690 22692 18696 22704
rect 18651 22664 18696 22692
rect 18690 22652 18696 22664
rect 18748 22652 18754 22704
rect 23661 22695 23719 22701
rect 23661 22661 23673 22695
rect 23707 22692 23719 22695
rect 25130 22692 25136 22704
rect 23707 22664 25136 22692
rect 23707 22661 23719 22664
rect 23661 22655 23719 22661
rect 25130 22652 25136 22664
rect 25188 22692 25194 22704
rect 25225 22695 25283 22701
rect 25225 22692 25237 22695
rect 25188 22664 25237 22692
rect 25188 22652 25194 22664
rect 25225 22661 25237 22664
rect 25271 22661 25283 22695
rect 32048 22692 32076 22720
rect 25225 22655 25283 22661
rect 31036 22664 32076 22692
rect 33045 22695 33103 22701
rect 17589 22627 17647 22633
rect 17589 22624 17601 22627
rect 17552 22596 17601 22624
rect 17552 22584 17558 22596
rect 17589 22593 17601 22596
rect 17635 22624 17647 22627
rect 18325 22627 18383 22633
rect 17635 22596 18276 22624
rect 17635 22593 17647 22596
rect 17589 22587 17647 22593
rect 17972 22556 18092 22567
rect 18248 22565 18276 22596
rect 18325 22593 18337 22627
rect 18371 22593 18383 22627
rect 20070 22624 20076 22636
rect 20031 22596 20076 22624
rect 18325 22587 18383 22593
rect 20070 22584 20076 22596
rect 20128 22584 20134 22636
rect 20165 22627 20223 22633
rect 20165 22593 20177 22627
rect 20211 22593 20223 22627
rect 20165 22587 20223 22593
rect 20349 22627 20407 22633
rect 20349 22593 20361 22627
rect 20395 22593 20407 22627
rect 20349 22587 20407 22593
rect 20441 22627 20499 22633
rect 20441 22593 20453 22627
rect 20487 22624 20499 22627
rect 20622 22624 20628 22636
rect 20487 22596 20628 22624
rect 20487 22593 20499 22596
rect 20441 22587 20499 22593
rect 18233 22559 18291 22565
rect 15396 22539 18138 22556
rect 15396 22528 18000 22539
rect 18064 22528 18138 22539
rect 11974 22488 11980 22500
rect 9416 22460 11980 22488
rect 5040 22448 5046 22460
rect 11974 22448 11980 22460
rect 12032 22448 12038 22500
rect 17497 22491 17555 22497
rect 17497 22457 17509 22491
rect 17543 22488 17555 22491
rect 17954 22488 17960 22500
rect 17543 22460 17960 22488
rect 17543 22457 17555 22460
rect 17497 22451 17555 22457
rect 17954 22448 17960 22460
rect 18012 22448 18018 22500
rect 18110 22488 18138 22528
rect 18233 22525 18245 22559
rect 18279 22556 18291 22559
rect 20180 22556 20208 22587
rect 18279 22528 20208 22556
rect 18279 22525 18291 22528
rect 18233 22519 18291 22525
rect 20364 22488 20392 22587
rect 20622 22584 20628 22596
rect 20680 22584 20686 22636
rect 21174 22584 21180 22636
rect 21232 22624 21238 22636
rect 21818 22624 21824 22636
rect 21232 22596 21824 22624
rect 21232 22584 21238 22596
rect 21818 22584 21824 22596
rect 21876 22624 21882 22636
rect 22005 22627 22063 22633
rect 22005 22624 22017 22627
rect 21876 22596 22017 22624
rect 21876 22584 21882 22596
rect 22005 22593 22017 22596
rect 22051 22593 22063 22627
rect 22186 22624 22192 22636
rect 22147 22596 22192 22624
rect 22005 22587 22063 22593
rect 22020 22556 22048 22587
rect 22186 22584 22192 22596
rect 22244 22584 22250 22636
rect 23569 22627 23627 22633
rect 23569 22593 23581 22627
rect 23615 22593 23627 22627
rect 23569 22587 23627 22593
rect 24857 22627 24915 22633
rect 24857 22593 24869 22627
rect 24903 22624 24915 22627
rect 27154 22624 27160 22636
rect 24903 22596 27160 22624
rect 24903 22593 24915 22596
rect 24857 22587 24915 22593
rect 23584 22556 23612 22587
rect 27154 22584 27160 22596
rect 27212 22584 27218 22636
rect 27982 22624 27988 22636
rect 27943 22596 27988 22624
rect 27982 22584 27988 22596
rect 28040 22584 28046 22636
rect 28258 22584 28264 22636
rect 28316 22624 28322 22636
rect 31036 22633 31064 22664
rect 33045 22661 33057 22695
rect 33091 22692 33103 22695
rect 33134 22692 33140 22704
rect 33091 22664 33140 22692
rect 33091 22661 33103 22664
rect 33045 22655 33103 22661
rect 33134 22652 33140 22664
rect 33192 22652 33198 22704
rect 33502 22692 33508 22704
rect 33463 22664 33508 22692
rect 33502 22652 33508 22664
rect 33560 22652 33566 22704
rect 28813 22627 28871 22633
rect 28813 22624 28825 22627
rect 28316 22596 28825 22624
rect 28316 22584 28322 22596
rect 28813 22593 28825 22596
rect 28859 22624 28871 22627
rect 31021 22627 31079 22633
rect 28859 22596 30972 22624
rect 28859 22593 28871 22596
rect 28813 22587 28871 22593
rect 22020 22528 23612 22556
rect 23842 22516 23848 22568
rect 23900 22556 23906 22568
rect 24765 22559 24823 22565
rect 24765 22556 24777 22559
rect 23900 22528 24777 22556
rect 23900 22516 23906 22528
rect 24765 22525 24777 22528
rect 24811 22525 24823 22559
rect 24765 22519 24823 22525
rect 25133 22559 25191 22565
rect 25133 22525 25145 22559
rect 25179 22556 25191 22559
rect 26142 22556 26148 22568
rect 25179 22528 26148 22556
rect 25179 22525 25191 22528
rect 25133 22519 25191 22525
rect 26142 22516 26148 22528
rect 26200 22516 26206 22568
rect 22005 22491 22063 22497
rect 22005 22488 22017 22491
rect 18110 22460 20024 22488
rect 20364 22460 22017 22488
rect 3602 22420 3608 22432
rect 3563 22392 3608 22420
rect 3602 22380 3608 22392
rect 3660 22380 3666 22432
rect 3786 22420 3792 22432
rect 3747 22392 3792 22420
rect 3786 22380 3792 22392
rect 3844 22380 3850 22432
rect 4338 22380 4344 22432
rect 4396 22420 4402 22432
rect 4525 22423 4583 22429
rect 4525 22420 4537 22423
rect 4396 22392 4537 22420
rect 4396 22380 4402 22392
rect 4525 22389 4537 22392
rect 4571 22420 4583 22423
rect 4614 22420 4620 22432
rect 4571 22392 4620 22420
rect 4571 22389 4583 22392
rect 4525 22383 4583 22389
rect 4614 22380 4620 22392
rect 4672 22380 4678 22432
rect 11793 22423 11851 22429
rect 11793 22389 11805 22423
rect 11839 22420 11851 22423
rect 13170 22420 13176 22432
rect 11839 22392 13176 22420
rect 11839 22389 11851 22392
rect 11793 22383 11851 22389
rect 13170 22380 13176 22392
rect 13228 22380 13234 22432
rect 14645 22423 14703 22429
rect 14645 22389 14657 22423
rect 14691 22420 14703 22423
rect 15197 22423 15255 22429
rect 15197 22420 15209 22423
rect 14691 22392 15209 22420
rect 14691 22389 14703 22392
rect 14645 22383 14703 22389
rect 15197 22389 15209 22392
rect 15243 22389 15255 22423
rect 18046 22420 18052 22432
rect 18007 22392 18052 22420
rect 15197 22383 15255 22389
rect 18046 22380 18052 22392
rect 18104 22380 18110 22432
rect 19886 22420 19892 22432
rect 19847 22392 19892 22420
rect 19886 22380 19892 22392
rect 19944 22380 19950 22432
rect 19996 22420 20024 22460
rect 22005 22457 22017 22460
rect 22051 22457 22063 22491
rect 22005 22451 22063 22457
rect 23014 22420 23020 22432
rect 19996 22392 23020 22420
rect 23014 22380 23020 22392
rect 23072 22380 23078 22432
rect 24578 22420 24584 22432
rect 24539 22392 24584 22420
rect 24578 22380 24584 22392
rect 24636 22380 24642 22432
rect 26970 22380 26976 22432
rect 27028 22420 27034 22432
rect 27341 22423 27399 22429
rect 27341 22420 27353 22423
rect 27028 22392 27353 22420
rect 27028 22380 27034 22392
rect 27341 22389 27353 22392
rect 27387 22389 27399 22423
rect 27341 22383 27399 22389
rect 30374 22380 30380 22432
rect 30432 22420 30438 22432
rect 30837 22423 30895 22429
rect 30837 22420 30849 22423
rect 30432 22392 30849 22420
rect 30432 22380 30438 22392
rect 30837 22389 30849 22392
rect 30883 22389 30895 22423
rect 30944 22420 30972 22596
rect 31021 22593 31033 22627
rect 31067 22593 31079 22627
rect 31021 22587 31079 22593
rect 31205 22627 31263 22633
rect 31205 22593 31217 22627
rect 31251 22624 31263 22627
rect 31386 22624 31392 22636
rect 31251 22596 31392 22624
rect 31251 22593 31263 22596
rect 31205 22587 31263 22593
rect 31386 22584 31392 22596
rect 31444 22584 31450 22636
rect 32674 22624 32680 22636
rect 32635 22596 32680 22624
rect 32674 22584 32680 22596
rect 32732 22584 32738 22636
rect 33686 22624 33692 22636
rect 33647 22596 33692 22624
rect 33686 22584 33692 22596
rect 33744 22584 33750 22636
rect 31113 22559 31171 22565
rect 31113 22525 31125 22559
rect 31159 22525 31171 22559
rect 31294 22556 31300 22568
rect 31255 22528 31300 22556
rect 31113 22519 31171 22525
rect 31128 22488 31156 22519
rect 31294 22516 31300 22528
rect 31352 22516 31358 22568
rect 32398 22516 32404 22568
rect 32456 22556 32462 22568
rect 32539 22559 32597 22565
rect 32539 22556 32551 22559
rect 32456 22528 32551 22556
rect 32456 22516 32462 22528
rect 32539 22525 32551 22528
rect 32585 22525 32597 22559
rect 32539 22519 32597 22525
rect 32953 22559 33011 22565
rect 32953 22525 32965 22559
rect 32999 22556 33011 22559
rect 33318 22556 33324 22568
rect 32999 22528 33324 22556
rect 32999 22525 33011 22528
rect 32953 22519 33011 22525
rect 33318 22516 33324 22528
rect 33376 22516 33382 22568
rect 31478 22488 31484 22500
rect 31128 22460 31484 22488
rect 31478 22448 31484 22460
rect 31536 22448 31542 22500
rect 31726 22460 33824 22488
rect 31726 22420 31754 22460
rect 33796 22429 33824 22460
rect 30944 22392 31754 22420
rect 33781 22423 33839 22429
rect 30837 22383 30895 22389
rect 33781 22389 33793 22423
rect 33827 22389 33839 22423
rect 33781 22383 33839 22389
rect 1104 22330 34868 22352
rect 1104 22278 5170 22330
rect 5222 22278 5234 22330
rect 5286 22278 5298 22330
rect 5350 22278 5362 22330
rect 5414 22278 5426 22330
rect 5478 22278 13611 22330
rect 13663 22278 13675 22330
rect 13727 22278 13739 22330
rect 13791 22278 13803 22330
rect 13855 22278 13867 22330
rect 13919 22278 22052 22330
rect 22104 22278 22116 22330
rect 22168 22278 22180 22330
rect 22232 22278 22244 22330
rect 22296 22278 22308 22330
rect 22360 22278 30493 22330
rect 30545 22278 30557 22330
rect 30609 22278 30621 22330
rect 30673 22278 30685 22330
rect 30737 22278 30749 22330
rect 30801 22278 34868 22330
rect 1104 22256 34868 22278
rect 11698 22176 11704 22228
rect 11756 22216 11762 22228
rect 11805 22219 11863 22225
rect 11805 22216 11817 22219
rect 11756 22188 11817 22216
rect 11756 22176 11762 22188
rect 11805 22185 11817 22188
rect 11851 22185 11863 22219
rect 11805 22179 11863 22185
rect 16390 22176 16396 22228
rect 16448 22216 16454 22228
rect 20070 22216 20076 22228
rect 16448 22188 20076 22216
rect 16448 22176 16454 22188
rect 20070 22176 20076 22188
rect 20128 22176 20134 22228
rect 20898 22176 20904 22228
rect 20956 22176 20962 22228
rect 23014 22216 23020 22228
rect 22975 22188 23020 22216
rect 23014 22176 23020 22188
rect 23072 22176 23078 22228
rect 23201 22219 23259 22225
rect 23201 22185 23213 22219
rect 23247 22185 23259 22219
rect 23201 22179 23259 22185
rect 33505 22219 33563 22225
rect 33505 22185 33517 22219
rect 33551 22216 33563 22219
rect 33686 22216 33692 22228
rect 33551 22188 33692 22216
rect 33551 22185 33563 22188
rect 33505 22179 33563 22185
rect 6638 22108 6644 22160
rect 6696 22148 6702 22160
rect 10318 22148 10324 22160
rect 6696 22120 10324 22148
rect 6696 22108 6702 22120
rect 10318 22108 10324 22120
rect 10376 22108 10382 22160
rect 12710 22108 12716 22160
rect 12768 22148 12774 22160
rect 12901 22151 12959 22157
rect 12901 22148 12913 22151
rect 12768 22120 12913 22148
rect 12768 22108 12774 22120
rect 12901 22117 12913 22120
rect 12947 22117 12959 22151
rect 12901 22111 12959 22117
rect 12989 22151 13047 22157
rect 12989 22117 13001 22151
rect 13035 22148 13047 22151
rect 13078 22148 13084 22160
rect 13035 22120 13084 22148
rect 13035 22117 13047 22120
rect 12989 22111 13047 22117
rect 13078 22108 13084 22120
rect 13136 22148 13142 22160
rect 13262 22148 13268 22160
rect 13136 22120 13268 22148
rect 13136 22108 13142 22120
rect 13262 22108 13268 22120
rect 13320 22108 13326 22160
rect 20916 22148 20944 22176
rect 20824 22120 20944 22148
rect 10778 22040 10784 22092
rect 10836 22080 10842 22092
rect 10836 22052 12434 22080
rect 10836 22040 10842 22052
rect 7098 21972 7104 22024
rect 7156 22012 7162 22024
rect 7193 22015 7251 22021
rect 7193 22012 7205 22015
rect 7156 21984 7205 22012
rect 7156 21972 7162 21984
rect 7193 21981 7205 21984
rect 7239 22012 7251 22015
rect 7466 22012 7472 22024
rect 7239 21984 7472 22012
rect 7239 21981 7251 21984
rect 7193 21975 7251 21981
rect 7466 21972 7472 21984
rect 7524 21972 7530 22024
rect 9306 22012 9312 22024
rect 9267 21984 9312 22012
rect 9306 21972 9312 21984
rect 9364 21972 9370 22024
rect 12066 21972 12072 22024
rect 12124 22012 12130 22024
rect 12124 21984 12169 22012
rect 12124 21972 12130 21984
rect 11698 21944 11704 21956
rect 11362 21916 11704 21944
rect 11698 21904 11704 21916
rect 11756 21904 11762 21956
rect 7190 21876 7196 21888
rect 7151 21848 7196 21876
rect 7190 21836 7196 21848
rect 7248 21836 7254 21888
rect 8846 21836 8852 21888
rect 8904 21876 8910 21888
rect 9030 21876 9036 21888
rect 8904 21848 9036 21876
rect 8904 21836 8910 21848
rect 9030 21836 9036 21848
rect 9088 21876 9094 21888
rect 9217 21879 9275 21885
rect 9217 21876 9229 21879
rect 9088 21848 9229 21876
rect 9088 21836 9094 21848
rect 9217 21845 9229 21848
rect 9263 21845 9275 21879
rect 9217 21839 9275 21845
rect 10226 21836 10232 21888
rect 10284 21876 10290 21888
rect 10321 21879 10379 21885
rect 10321 21876 10333 21879
rect 10284 21848 10333 21876
rect 10284 21836 10290 21848
rect 10321 21845 10333 21848
rect 10367 21876 10379 21879
rect 11054 21876 11060 21888
rect 10367 21848 11060 21876
rect 10367 21845 10379 21848
rect 10321 21839 10379 21845
rect 11054 21836 11060 21848
rect 11112 21836 11118 21888
rect 12406 21876 12434 22052
rect 18046 22040 18052 22092
rect 18104 22089 18110 22092
rect 18104 22083 18153 22089
rect 18104 22049 18107 22083
rect 18141 22049 18153 22083
rect 20438 22080 20444 22092
rect 18104 22043 18153 22049
rect 18248 22052 20444 22080
rect 18104 22040 18110 22043
rect 12805 22015 12863 22021
rect 12805 21981 12817 22015
rect 12851 21981 12863 22015
rect 12805 21975 12863 21981
rect 13081 22015 13139 22021
rect 13081 21981 13093 22015
rect 13127 22012 13139 22015
rect 13170 22012 13176 22024
rect 13127 21984 13176 22012
rect 13127 21981 13139 21984
rect 13081 21975 13139 21981
rect 12820 21944 12848 21975
rect 13170 21972 13176 21984
rect 13228 21972 13234 22024
rect 17954 22012 17960 22024
rect 17915 21984 17960 22012
rect 17954 21972 17960 21984
rect 18012 21972 18018 22024
rect 18248 22012 18276 22052
rect 20438 22040 20444 22052
rect 20496 22040 20502 22092
rect 18156 21984 18276 22012
rect 18325 22015 18383 22021
rect 18156 21944 18184 21984
rect 18325 21981 18337 22015
rect 18371 22012 18383 22015
rect 18414 22012 18420 22024
rect 18371 21984 18420 22012
rect 18371 21981 18383 21984
rect 18325 21975 18383 21981
rect 18414 21972 18420 21984
rect 18472 21972 18478 22024
rect 18782 21972 18788 22024
rect 18840 22012 18846 22024
rect 20824 22021 20852 22120
rect 22646 22108 22652 22160
rect 22704 22148 22710 22160
rect 23216 22148 23244 22179
rect 33686 22176 33692 22188
rect 33744 22176 33750 22228
rect 30374 22148 30380 22160
rect 22704 22120 23244 22148
rect 30024 22120 30380 22148
rect 22704 22108 22710 22120
rect 24854 22080 24860 22092
rect 24815 22052 24860 22080
rect 24854 22040 24860 22052
rect 24912 22040 24918 22092
rect 24946 22040 24952 22092
rect 25004 22080 25010 22092
rect 26970 22080 26976 22092
rect 25004 22052 25049 22080
rect 26931 22052 26976 22080
rect 25004 22040 25010 22052
rect 26970 22040 26976 22052
rect 27028 22040 27034 22092
rect 27246 22040 27252 22092
rect 27304 22080 27310 22092
rect 29914 22080 29920 22092
rect 27304 22052 29920 22080
rect 27304 22040 27310 22052
rect 29914 22040 29920 22052
rect 29972 22040 29978 22092
rect 30024 22089 30052 22120
rect 30374 22108 30380 22120
rect 30432 22108 30438 22160
rect 30009 22083 30067 22089
rect 30009 22049 30021 22083
rect 30055 22080 30067 22083
rect 33134 22080 33140 22092
rect 30055 22052 30089 22080
rect 33095 22052 33140 22080
rect 30055 22049 30067 22052
rect 30009 22043 30067 22049
rect 33134 22040 33140 22052
rect 33192 22040 33198 22092
rect 19613 22015 19671 22021
rect 19613 22012 19625 22015
rect 18840 21984 19625 22012
rect 18840 21972 18846 21984
rect 19613 21981 19625 21984
rect 19659 21981 19671 22015
rect 19613 21975 19671 21981
rect 19889 22015 19947 22021
rect 19889 21981 19901 22015
rect 19935 22006 19947 22015
rect 20809 22015 20867 22021
rect 19996 22006 20760 22012
rect 19935 21984 20760 22006
rect 19935 21981 20024 21984
rect 19889 21978 20024 21981
rect 19889 21975 19947 21978
rect 12820 21916 18184 21944
rect 18230 21904 18236 21956
rect 18288 21944 18294 21956
rect 19628 21944 19656 21975
rect 20732 21944 20760 21984
rect 20809 21981 20821 22015
rect 20855 21981 20867 22015
rect 20809 21975 20867 21981
rect 22830 21972 22836 22024
rect 22888 22012 22894 22024
rect 23201 22015 23259 22021
rect 23201 22012 23213 22015
rect 22888 21984 23213 22012
rect 22888 21972 22894 21984
rect 23201 21981 23213 21984
rect 23247 21981 23259 22015
rect 23201 21975 23259 21981
rect 23385 22015 23443 22021
rect 23385 21981 23397 22015
rect 23431 22012 23443 22015
rect 24578 22012 24584 22024
rect 23431 21984 24584 22012
rect 23431 21981 23443 21984
rect 23385 21975 23443 21981
rect 24578 21972 24584 21984
rect 24636 21972 24642 22024
rect 24762 22012 24768 22024
rect 24723 21984 24768 22012
rect 24762 21972 24768 21984
rect 24820 21972 24826 22024
rect 25041 22015 25099 22021
rect 25041 21981 25053 22015
rect 25087 22012 25099 22015
rect 25130 22012 25136 22024
rect 25087 21984 25136 22012
rect 25087 21981 25099 21984
rect 25041 21975 25099 21981
rect 25130 21972 25136 21984
rect 25188 21972 25194 22024
rect 26053 22015 26111 22021
rect 26053 21981 26065 22015
rect 26099 21981 26111 22015
rect 26053 21975 26111 21981
rect 26237 22015 26295 22021
rect 26237 21981 26249 22015
rect 26283 22012 26295 22015
rect 26988 22012 27016 22040
rect 26283 21984 27016 22012
rect 26283 21981 26295 21984
rect 26237 21975 26295 21981
rect 21082 21944 21088 21956
rect 18288 21916 18333 21944
rect 19628 21916 20668 21944
rect 20732 21916 21088 21944
rect 18288 21904 18294 21916
rect 12621 21879 12679 21885
rect 12621 21876 12633 21879
rect 12406 21848 12633 21876
rect 12621 21845 12633 21848
rect 12667 21845 12679 21879
rect 12621 21839 12679 21845
rect 18966 21836 18972 21888
rect 19024 21876 19030 21888
rect 19429 21879 19487 21885
rect 19429 21876 19441 21879
rect 19024 21848 19441 21876
rect 19024 21836 19030 21848
rect 19429 21845 19441 21848
rect 19475 21845 19487 21879
rect 19794 21876 19800 21888
rect 19755 21848 19800 21876
rect 19429 21839 19487 21845
rect 19794 21836 19800 21848
rect 19852 21836 19858 21888
rect 20640 21876 20668 21916
rect 21082 21904 21088 21916
rect 21140 21944 21146 21956
rect 21542 21944 21548 21956
rect 21140 21916 21548 21944
rect 21140 21904 21146 21916
rect 21542 21904 21548 21916
rect 21600 21904 21606 21956
rect 26068 21944 26096 21975
rect 27062 21972 27068 22024
rect 27120 22012 27126 22024
rect 27801 22015 27859 22021
rect 27120 21984 27165 22012
rect 27120 21972 27126 21984
rect 27801 21981 27813 22015
rect 27847 22012 27859 22015
rect 28629 22015 28687 22021
rect 28629 22012 28641 22015
rect 27847 21984 28641 22012
rect 27847 21981 27859 21984
rect 27801 21975 27859 21981
rect 28629 21981 28641 21984
rect 28675 21981 28687 22015
rect 28629 21975 28687 21981
rect 30101 22015 30159 22021
rect 30101 21981 30113 22015
rect 30147 21981 30159 22015
rect 31018 22012 31024 22024
rect 30979 21984 31024 22012
rect 30101 21975 30159 21981
rect 27080 21944 27108 21972
rect 26068 21916 27108 21944
rect 27522 21904 27528 21956
rect 27580 21944 27586 21956
rect 28261 21947 28319 21953
rect 28261 21944 28273 21947
rect 27580 21916 28273 21944
rect 27580 21904 27586 21916
rect 28261 21913 28273 21916
rect 28307 21913 28319 21947
rect 28442 21944 28448 21956
rect 28403 21916 28448 21944
rect 28261 21907 28319 21913
rect 28442 21904 28448 21916
rect 28500 21904 28506 21956
rect 30116 21944 30144 21975
rect 31018 21972 31024 21984
rect 31076 22012 31082 22024
rect 31386 22012 31392 22024
rect 31076 21984 31248 22012
rect 31347 21984 31392 22012
rect 31076 21972 31082 21984
rect 30374 21944 30380 21956
rect 30116 21916 30380 21944
rect 30374 21904 30380 21916
rect 30432 21944 30438 21956
rect 31113 21947 31171 21953
rect 31113 21944 31125 21947
rect 30432 21916 31125 21944
rect 30432 21904 30438 21916
rect 31113 21913 31125 21916
rect 31159 21913 31171 21947
rect 31220 21944 31248 21984
rect 31386 21972 31392 21984
rect 31444 21972 31450 22024
rect 31570 22012 31576 22024
rect 31531 21984 31576 22012
rect 31570 21972 31576 21984
rect 31628 22012 31634 22024
rect 32033 22015 32091 22021
rect 32033 22012 32045 22015
rect 31628 21984 32045 22012
rect 31628 21972 31634 21984
rect 32033 21981 32045 21984
rect 32079 21981 32091 22015
rect 32398 22012 32404 22024
rect 32359 21984 32404 22012
rect 32033 21975 32091 21981
rect 32398 21972 32404 21984
rect 32456 21972 32462 22024
rect 32582 22012 32588 22024
rect 32543 21984 32588 22012
rect 32582 21972 32588 21984
rect 32640 21972 32646 22024
rect 33318 22012 33324 22024
rect 33279 21984 33324 22012
rect 33318 21972 33324 21984
rect 33376 21972 33382 22024
rect 32125 21947 32183 21953
rect 32125 21944 32137 21947
rect 31220 21916 32137 21944
rect 31113 21907 31171 21913
rect 32125 21913 32137 21916
rect 32171 21913 32183 21947
rect 32125 21907 32183 21913
rect 21174 21876 21180 21888
rect 20640 21848 21180 21876
rect 21174 21836 21180 21848
rect 21232 21836 21238 21888
rect 22278 21876 22284 21888
rect 22239 21848 22284 21876
rect 22278 21836 22284 21848
rect 22336 21836 22342 21888
rect 25038 21836 25044 21888
rect 25096 21876 25102 21888
rect 25225 21879 25283 21885
rect 25225 21876 25237 21879
rect 25096 21848 25237 21876
rect 25096 21836 25102 21848
rect 25225 21845 25237 21848
rect 25271 21845 25283 21879
rect 25225 21839 25283 21845
rect 26145 21879 26203 21885
rect 26145 21845 26157 21879
rect 26191 21876 26203 21879
rect 26878 21876 26884 21888
rect 26191 21848 26884 21876
rect 26191 21845 26203 21848
rect 26145 21839 26203 21845
rect 26878 21836 26884 21848
rect 26936 21836 26942 21888
rect 26970 21836 26976 21888
rect 27028 21876 27034 21888
rect 27709 21879 27767 21885
rect 27709 21876 27721 21879
rect 27028 21848 27721 21876
rect 27028 21836 27034 21848
rect 27709 21845 27721 21848
rect 27755 21845 27767 21879
rect 29730 21876 29736 21888
rect 29691 21848 29736 21876
rect 27709 21839 27767 21845
rect 29730 21836 29736 21848
rect 29788 21836 29794 21888
rect 1104 21786 35027 21808
rect 1104 21734 9390 21786
rect 9442 21734 9454 21786
rect 9506 21734 9518 21786
rect 9570 21734 9582 21786
rect 9634 21734 9646 21786
rect 9698 21734 17831 21786
rect 17883 21734 17895 21786
rect 17947 21734 17959 21786
rect 18011 21734 18023 21786
rect 18075 21734 18087 21786
rect 18139 21734 26272 21786
rect 26324 21734 26336 21786
rect 26388 21734 26400 21786
rect 26452 21734 26464 21786
rect 26516 21734 26528 21786
rect 26580 21734 34713 21786
rect 34765 21734 34777 21786
rect 34829 21734 34841 21786
rect 34893 21734 34905 21786
rect 34957 21734 34969 21786
rect 35021 21734 35027 21786
rect 1104 21712 35027 21734
rect 18414 21632 18420 21684
rect 18472 21672 18478 21684
rect 19426 21672 19432 21684
rect 18472 21644 19432 21672
rect 18472 21632 18478 21644
rect 19426 21632 19432 21644
rect 19484 21632 19490 21684
rect 20530 21672 20536 21684
rect 19720 21644 20536 21672
rect 11698 21604 11704 21616
rect 11659 21576 11704 21604
rect 11698 21564 11704 21576
rect 11756 21564 11762 21616
rect 2869 21539 2927 21545
rect 2869 21505 2881 21539
rect 2915 21536 2927 21539
rect 3602 21536 3608 21548
rect 2915 21508 3608 21536
rect 2915 21505 2927 21508
rect 2869 21499 2927 21505
rect 3602 21496 3608 21508
rect 3660 21536 3666 21548
rect 3789 21539 3847 21545
rect 3789 21536 3801 21539
rect 3660 21508 3801 21536
rect 3660 21496 3666 21508
rect 3789 21505 3801 21508
rect 3835 21505 3847 21539
rect 3789 21499 3847 21505
rect 4065 21539 4123 21545
rect 4065 21505 4077 21539
rect 4111 21536 4123 21539
rect 7466 21536 7472 21548
rect 4111 21508 7472 21536
rect 4111 21505 4123 21508
rect 4065 21499 4123 21505
rect 7466 21496 7472 21508
rect 7524 21496 7530 21548
rect 11790 21536 11796 21548
rect 11751 21508 11796 21536
rect 11790 21496 11796 21508
rect 11848 21496 11854 21548
rect 11974 21536 11980 21548
rect 11935 21508 11980 21536
rect 11974 21496 11980 21508
rect 12032 21496 12038 21548
rect 13998 21496 14004 21548
rect 14056 21536 14062 21548
rect 14461 21539 14519 21545
rect 14461 21536 14473 21539
rect 14056 21508 14473 21536
rect 14056 21496 14062 21508
rect 14461 21505 14473 21508
rect 14507 21505 14519 21539
rect 15286 21536 15292 21548
rect 15247 21508 15292 21536
rect 14461 21499 14519 21505
rect 15286 21496 15292 21508
rect 15344 21496 15350 21548
rect 15473 21539 15531 21545
rect 15473 21505 15485 21539
rect 15519 21536 15531 21539
rect 15746 21536 15752 21548
rect 15519 21508 15752 21536
rect 15519 21505 15531 21508
rect 15473 21499 15531 21505
rect 15746 21496 15752 21508
rect 15804 21536 15810 21548
rect 17678 21536 17684 21548
rect 15804 21508 17684 21536
rect 15804 21496 15810 21508
rect 17678 21496 17684 21508
rect 17736 21496 17742 21548
rect 19613 21539 19671 21545
rect 19613 21505 19625 21539
rect 19659 21536 19671 21539
rect 19720 21536 19748 21644
rect 20530 21632 20536 21644
rect 20588 21632 20594 21684
rect 26970 21672 26976 21684
rect 22066 21644 26976 21672
rect 22066 21604 22094 21644
rect 26970 21632 26976 21644
rect 27028 21632 27034 21684
rect 27154 21672 27160 21684
rect 27115 21644 27160 21672
rect 27154 21632 27160 21644
rect 27212 21632 27218 21684
rect 27522 21632 27528 21684
rect 27580 21632 27586 21684
rect 30374 21672 30380 21684
rect 30335 21644 30380 21672
rect 30374 21632 30380 21644
rect 30432 21632 30438 21684
rect 31665 21675 31723 21681
rect 31665 21641 31677 21675
rect 31711 21672 31723 21675
rect 31754 21672 31760 21684
rect 31711 21644 31760 21672
rect 31711 21641 31723 21644
rect 31665 21635 31723 21641
rect 31754 21632 31760 21644
rect 31812 21632 31818 21684
rect 20548 21576 22094 21604
rect 19886 21536 19892 21548
rect 19659 21508 19748 21536
rect 19847 21508 19892 21536
rect 19659 21505 19671 21508
rect 19613 21499 19671 21505
rect 19886 21496 19892 21508
rect 19944 21496 19950 21548
rect 20548 21545 20576 21576
rect 26878 21564 26884 21616
rect 26936 21604 26942 21616
rect 27540 21604 27568 21632
rect 28442 21604 28448 21616
rect 26936 21576 27568 21604
rect 28184 21576 28448 21604
rect 26936 21564 26942 21576
rect 20533 21539 20591 21545
rect 20533 21505 20545 21539
rect 20579 21505 20591 21539
rect 20533 21499 20591 21505
rect 20625 21539 20683 21545
rect 20625 21505 20637 21539
rect 20671 21505 20683 21539
rect 20625 21499 20683 21505
rect 22005 21539 22063 21545
rect 22005 21505 22017 21539
rect 22051 21505 22063 21539
rect 22278 21536 22284 21548
rect 22239 21508 22284 21536
rect 22005 21499 22063 21505
rect 3145 21471 3203 21477
rect 3145 21437 3157 21471
rect 3191 21468 3203 21471
rect 3694 21468 3700 21480
rect 3191 21440 3700 21468
rect 3191 21437 3203 21440
rect 3145 21431 3203 21437
rect 3694 21428 3700 21440
rect 3752 21428 3758 21480
rect 3881 21471 3939 21477
rect 3881 21437 3893 21471
rect 3927 21468 3939 21471
rect 4430 21468 4436 21480
rect 3927 21440 4436 21468
rect 3927 21437 3939 21440
rect 3881 21431 3939 21437
rect 2961 21403 3019 21409
rect 2961 21369 2973 21403
rect 3007 21400 3019 21403
rect 3896 21400 3924 21431
rect 4430 21428 4436 21440
rect 4488 21428 4494 21480
rect 18230 21428 18236 21480
rect 18288 21468 18294 21480
rect 20640 21468 20668 21499
rect 18288 21440 20668 21468
rect 18288 21428 18294 21440
rect 3007 21372 3924 21400
rect 3973 21403 4031 21409
rect 3007 21369 3019 21372
rect 2961 21363 3019 21369
rect 3973 21369 3985 21403
rect 4019 21400 4031 21403
rect 4062 21400 4068 21412
rect 4019 21372 4068 21400
rect 4019 21369 4031 21372
rect 3973 21363 4031 21369
rect 3050 21292 3056 21344
rect 3108 21332 3114 21344
rect 3602 21332 3608 21344
rect 3108 21304 3153 21332
rect 3563 21304 3608 21332
rect 3108 21292 3114 21304
rect 3602 21292 3608 21304
rect 3660 21292 3666 21344
rect 3694 21292 3700 21344
rect 3752 21332 3758 21344
rect 3988 21332 4016 21363
rect 4062 21360 4068 21372
rect 4120 21360 4126 21412
rect 19242 21360 19248 21412
rect 19300 21400 19306 21412
rect 22020 21400 22048 21499
rect 22278 21496 22284 21508
rect 22336 21496 22342 21548
rect 27525 21539 27583 21545
rect 27525 21505 27537 21539
rect 27571 21536 27583 21539
rect 27706 21536 27712 21548
rect 27571 21508 27712 21536
rect 27571 21505 27583 21508
rect 27525 21499 27583 21505
rect 27706 21496 27712 21508
rect 27764 21496 27770 21548
rect 28184 21545 28212 21576
rect 28442 21564 28448 21576
rect 28500 21564 28506 21616
rect 30466 21604 30472 21616
rect 30300 21576 30472 21604
rect 28169 21539 28227 21545
rect 28169 21505 28181 21539
rect 28215 21505 28227 21539
rect 28169 21499 28227 21505
rect 28353 21539 28411 21545
rect 28353 21505 28365 21539
rect 28399 21536 28411 21539
rect 29730 21536 29736 21548
rect 28399 21508 29736 21536
rect 28399 21505 28411 21508
rect 28353 21499 28411 21505
rect 22370 21468 22376 21480
rect 22331 21440 22376 21468
rect 22370 21428 22376 21440
rect 22428 21428 22434 21480
rect 23198 21468 23204 21480
rect 23159 21440 23204 21468
rect 23198 21428 23204 21440
rect 23256 21428 23262 21480
rect 23477 21471 23535 21477
rect 23477 21437 23489 21471
rect 23523 21468 23535 21471
rect 23566 21468 23572 21480
rect 23523 21440 23572 21468
rect 23523 21437 23535 21440
rect 23477 21431 23535 21437
rect 23566 21428 23572 21440
rect 23624 21428 23630 21480
rect 23934 21428 23940 21480
rect 23992 21468 23998 21480
rect 24581 21471 24639 21477
rect 24581 21468 24593 21471
rect 23992 21440 24593 21468
rect 23992 21428 23998 21440
rect 24581 21437 24593 21440
rect 24627 21468 24639 21471
rect 27338 21468 27344 21480
rect 24627 21440 27344 21468
rect 24627 21437 24639 21440
rect 24581 21431 24639 21437
rect 27338 21428 27344 21440
rect 27396 21428 27402 21480
rect 27433 21471 27491 21477
rect 27433 21437 27445 21471
rect 27479 21468 27491 21471
rect 27614 21468 27620 21480
rect 27479 21440 27620 21468
rect 27479 21437 27491 21440
rect 27433 21431 27491 21437
rect 27614 21428 27620 21440
rect 27672 21428 27678 21480
rect 28184 21400 28212 21499
rect 29730 21496 29736 21508
rect 29788 21496 29794 21548
rect 30300 21545 30328 21576
rect 30466 21564 30472 21576
rect 30524 21564 30530 21616
rect 30561 21607 30619 21613
rect 30561 21573 30573 21607
rect 30607 21604 30619 21607
rect 31018 21604 31024 21616
rect 30607 21576 31024 21604
rect 30607 21573 30619 21576
rect 30561 21567 30619 21573
rect 31018 21564 31024 21576
rect 31076 21564 31082 21616
rect 31386 21564 31392 21616
rect 31444 21604 31450 21616
rect 31444 21576 31708 21604
rect 31444 21564 31450 21576
rect 30285 21539 30343 21545
rect 30285 21505 30297 21539
rect 30331 21505 30343 21539
rect 31478 21536 31484 21548
rect 31439 21508 31484 21536
rect 30285 21499 30343 21505
rect 31478 21496 31484 21508
rect 31536 21496 31542 21548
rect 31680 21545 31708 21576
rect 31665 21539 31723 21545
rect 31665 21505 31677 21539
rect 31711 21536 31723 21539
rect 32582 21536 32588 21548
rect 31711 21508 32588 21536
rect 31711 21505 31723 21508
rect 31665 21499 31723 21505
rect 32582 21496 32588 21508
rect 32640 21496 32646 21548
rect 19300 21372 22094 21400
rect 19300 21360 19306 21372
rect 3752 21304 4016 21332
rect 14553 21335 14611 21341
rect 3752 21292 3758 21304
rect 14553 21301 14565 21335
rect 14599 21332 14611 21335
rect 15378 21332 15384 21344
rect 14599 21304 15384 21332
rect 14599 21301 14611 21304
rect 14553 21295 14611 21301
rect 15378 21292 15384 21304
rect 15436 21292 15442 21344
rect 15473 21335 15531 21341
rect 15473 21301 15485 21335
rect 15519 21332 15531 21335
rect 15838 21332 15844 21344
rect 15519 21304 15844 21332
rect 15519 21301 15531 21304
rect 15473 21295 15531 21301
rect 15838 21292 15844 21304
rect 15896 21292 15902 21344
rect 15930 21292 15936 21344
rect 15988 21332 15994 21344
rect 19429 21335 19487 21341
rect 19429 21332 19441 21335
rect 15988 21304 19441 21332
rect 15988 21292 15994 21304
rect 19429 21301 19441 21304
rect 19475 21301 19487 21335
rect 22066 21332 22094 21372
rect 24504 21372 28212 21400
rect 23842 21332 23848 21344
rect 22066 21304 23848 21332
rect 19429 21295 19487 21301
rect 23842 21292 23848 21304
rect 23900 21332 23906 21344
rect 24504 21332 24532 21372
rect 23900 21304 24532 21332
rect 23900 21292 23906 21304
rect 27890 21292 27896 21344
rect 27948 21332 27954 21344
rect 28353 21335 28411 21341
rect 28353 21332 28365 21335
rect 27948 21304 28365 21332
rect 27948 21292 27954 21304
rect 28353 21301 28365 21304
rect 28399 21301 28411 21335
rect 28353 21295 28411 21301
rect 28442 21292 28448 21344
rect 28500 21332 28506 21344
rect 30561 21335 30619 21341
rect 30561 21332 30573 21335
rect 28500 21304 30573 21332
rect 28500 21292 28506 21304
rect 30561 21301 30573 21304
rect 30607 21301 30619 21335
rect 30561 21295 30619 21301
rect 1104 21242 34868 21264
rect 1104 21190 5170 21242
rect 5222 21190 5234 21242
rect 5286 21190 5298 21242
rect 5350 21190 5362 21242
rect 5414 21190 5426 21242
rect 5478 21190 13611 21242
rect 13663 21190 13675 21242
rect 13727 21190 13739 21242
rect 13791 21190 13803 21242
rect 13855 21190 13867 21242
rect 13919 21190 22052 21242
rect 22104 21190 22116 21242
rect 22168 21190 22180 21242
rect 22232 21190 22244 21242
rect 22296 21190 22308 21242
rect 22360 21190 30493 21242
rect 30545 21190 30557 21242
rect 30609 21190 30621 21242
rect 30673 21190 30685 21242
rect 30737 21190 30749 21242
rect 30801 21190 34868 21242
rect 1104 21168 34868 21190
rect 13078 21088 13084 21140
rect 13136 21128 13142 21140
rect 13449 21131 13507 21137
rect 13449 21128 13461 21131
rect 13136 21100 13461 21128
rect 13136 21088 13142 21100
rect 13449 21097 13461 21100
rect 13495 21097 13507 21131
rect 13449 21091 13507 21097
rect 14645 21131 14703 21137
rect 14645 21097 14657 21131
rect 14691 21097 14703 21131
rect 14645 21091 14703 21097
rect 16117 21131 16175 21137
rect 16117 21097 16129 21131
rect 16163 21128 16175 21131
rect 17310 21128 17316 21140
rect 16163 21100 17316 21128
rect 16163 21097 16175 21100
rect 16117 21091 16175 21097
rect 14660 21060 14688 21091
rect 17310 21088 17316 21100
rect 17368 21088 17374 21140
rect 18782 21128 18788 21140
rect 18743 21100 18788 21128
rect 18782 21088 18788 21100
rect 18840 21088 18846 21140
rect 21266 21128 21272 21140
rect 21227 21100 21272 21128
rect 21266 21088 21272 21100
rect 21324 21088 21330 21140
rect 23566 21128 23572 21140
rect 23527 21100 23572 21128
rect 23566 21088 23572 21100
rect 23624 21088 23630 21140
rect 23750 21088 23756 21140
rect 23808 21128 23814 21140
rect 30926 21128 30932 21140
rect 23808 21100 30932 21128
rect 23808 21088 23814 21100
rect 30926 21088 30932 21100
rect 30984 21088 30990 21140
rect 31478 21128 31484 21140
rect 31439 21100 31484 21128
rect 31478 21088 31484 21100
rect 31536 21088 31542 21140
rect 32398 21128 32404 21140
rect 32359 21100 32404 21128
rect 32398 21088 32404 21100
rect 32456 21088 32462 21140
rect 25866 21060 25872 21072
rect 14660 21032 25872 21060
rect 25866 21020 25872 21032
rect 25924 21020 25930 21072
rect 25958 21020 25964 21072
rect 26016 21060 26022 21072
rect 32490 21060 32496 21072
rect 26016 21032 32496 21060
rect 26016 21020 26022 21032
rect 32490 21020 32496 21032
rect 32548 21020 32554 21072
rect 7377 20995 7435 21001
rect 7377 20961 7389 20995
rect 7423 20992 7435 20995
rect 7466 20992 7472 21004
rect 7423 20964 7472 20992
rect 7423 20961 7435 20964
rect 7377 20955 7435 20961
rect 7466 20952 7472 20964
rect 7524 20952 7530 21004
rect 14660 20964 18644 20992
rect 3234 20924 3240 20936
rect 3195 20896 3240 20924
rect 3234 20884 3240 20896
rect 3292 20884 3298 20936
rect 3421 20927 3479 20933
rect 3421 20893 3433 20927
rect 3467 20924 3479 20927
rect 4430 20924 4436 20936
rect 3467 20896 4436 20924
rect 3467 20893 3479 20896
rect 3421 20887 3479 20893
rect 4430 20884 4436 20896
rect 4488 20884 4494 20936
rect 7282 20884 7288 20936
rect 7340 20924 7346 20936
rect 7561 20927 7619 20933
rect 7561 20924 7573 20927
rect 7340 20896 7573 20924
rect 7340 20884 7346 20896
rect 7561 20893 7573 20896
rect 7607 20893 7619 20927
rect 7561 20887 7619 20893
rect 7650 20884 7656 20936
rect 7708 20924 7714 20936
rect 7708 20896 7753 20924
rect 7708 20884 7714 20896
rect 10134 20884 10140 20936
rect 10192 20924 10198 20936
rect 10410 20924 10416 20936
rect 10192 20896 10416 20924
rect 10192 20884 10198 20896
rect 10410 20884 10416 20896
rect 10468 20884 10474 20936
rect 10689 20927 10747 20933
rect 10689 20893 10701 20927
rect 10735 20924 10747 20927
rect 10778 20924 10784 20936
rect 10735 20896 10784 20924
rect 10735 20893 10747 20896
rect 10689 20887 10747 20893
rect 10778 20884 10784 20896
rect 10836 20884 10842 20936
rect 13446 20884 13452 20936
rect 13504 20924 13510 20936
rect 13541 20927 13599 20933
rect 13541 20924 13553 20927
rect 13504 20896 13553 20924
rect 13504 20884 13510 20896
rect 13541 20893 13553 20896
rect 13587 20893 13599 20927
rect 14458 20924 14464 20936
rect 14419 20896 14464 20924
rect 13541 20887 13599 20893
rect 14458 20884 14464 20896
rect 14516 20884 14522 20936
rect 14660 20933 14688 20964
rect 14645 20927 14703 20933
rect 14645 20893 14657 20927
rect 14691 20893 14703 20927
rect 14645 20887 14703 20893
rect 17405 20927 17463 20933
rect 17405 20893 17417 20927
rect 17451 20924 17463 20927
rect 18322 20924 18328 20936
rect 17451 20896 18328 20924
rect 17451 20893 17463 20896
rect 17405 20887 17463 20893
rect 18322 20884 18328 20896
rect 18380 20884 18386 20936
rect 10597 20859 10655 20865
rect 10597 20825 10609 20859
rect 10643 20856 10655 20859
rect 11882 20856 11888 20868
rect 10643 20828 11888 20856
rect 10643 20825 10655 20828
rect 10597 20819 10655 20825
rect 11882 20816 11888 20828
rect 11940 20856 11946 20868
rect 15930 20856 15936 20868
rect 11940 20828 15936 20856
rect 11940 20816 11946 20828
rect 15930 20816 15936 20828
rect 15988 20816 15994 20868
rect 18509 20859 18567 20865
rect 18509 20825 18521 20859
rect 18555 20825 18567 20859
rect 18616 20856 18644 20964
rect 20070 20952 20076 21004
rect 20128 20992 20134 21004
rect 20165 20995 20223 21001
rect 20165 20992 20177 20995
rect 20128 20964 20177 20992
rect 20128 20952 20134 20964
rect 20165 20961 20177 20964
rect 20211 20961 20223 20995
rect 20165 20955 20223 20961
rect 20257 20995 20315 21001
rect 20257 20961 20269 20995
rect 20303 20992 20315 20995
rect 21450 20992 21456 21004
rect 20303 20964 21456 20992
rect 20303 20961 20315 20964
rect 20257 20955 20315 20961
rect 21450 20952 21456 20964
rect 21508 20952 21514 21004
rect 28442 20992 28448 21004
rect 22066 20964 28448 20992
rect 19242 20884 19248 20936
rect 19300 20924 19306 20936
rect 19797 20927 19855 20933
rect 19797 20924 19809 20927
rect 19300 20896 19809 20924
rect 19300 20884 19306 20896
rect 19797 20893 19809 20896
rect 19843 20893 19855 20927
rect 19797 20887 19855 20893
rect 19889 20927 19947 20933
rect 19889 20893 19901 20927
rect 19935 20924 19947 20927
rect 22066 20924 22094 20964
rect 28442 20952 28448 20964
rect 28500 20952 28506 21004
rect 33045 20995 33103 21001
rect 33045 20992 33057 20995
rect 31680 20964 33057 20992
rect 22554 20924 22560 20936
rect 19935 20896 22094 20924
rect 22515 20896 22560 20924
rect 19935 20893 19947 20896
rect 19889 20887 19947 20893
rect 22554 20884 22560 20896
rect 22612 20884 22618 20936
rect 23750 20924 23756 20936
rect 23308 20896 23756 20924
rect 18616 20828 19656 20856
rect 18509 20819 18567 20825
rect 3142 20748 3148 20800
rect 3200 20788 3206 20800
rect 3329 20791 3387 20797
rect 3329 20788 3341 20791
rect 3200 20760 3341 20788
rect 3200 20748 3206 20760
rect 3329 20757 3341 20760
rect 3375 20757 3387 20791
rect 7374 20788 7380 20800
rect 7335 20760 7380 20788
rect 3329 20751 3387 20757
rect 7374 20748 7380 20760
rect 7432 20748 7438 20800
rect 10226 20788 10232 20800
rect 10187 20760 10232 20788
rect 10226 20748 10232 20760
rect 10284 20748 10290 20800
rect 14274 20788 14280 20800
rect 14235 20760 14280 20788
rect 14274 20748 14280 20760
rect 14332 20748 14338 20800
rect 15838 20748 15844 20800
rect 15896 20788 15902 20800
rect 18524 20788 18552 20819
rect 19628 20797 19656 20828
rect 21174 20816 21180 20868
rect 21232 20856 21238 20868
rect 23308 20856 23336 20896
rect 23750 20884 23756 20896
rect 23808 20884 23814 20936
rect 23934 20924 23940 20936
rect 23895 20896 23940 20924
rect 23934 20884 23940 20896
rect 23992 20884 23998 20936
rect 24029 20927 24087 20933
rect 24029 20893 24041 20927
rect 24075 20893 24087 20927
rect 24029 20887 24087 20893
rect 21232 20828 23336 20856
rect 21232 20816 21238 20828
rect 15896 20760 18552 20788
rect 19613 20791 19671 20797
rect 15896 20748 15902 20760
rect 19613 20757 19625 20791
rect 19659 20757 19671 20791
rect 19613 20751 19671 20757
rect 23382 20748 23388 20800
rect 23440 20788 23446 20800
rect 23934 20788 23940 20800
rect 23440 20760 23940 20788
rect 23440 20748 23446 20760
rect 23934 20748 23940 20760
rect 23992 20748 23998 20800
rect 24044 20788 24072 20887
rect 24670 20884 24676 20936
rect 24728 20924 24734 20936
rect 24765 20927 24823 20933
rect 24765 20924 24777 20927
rect 24728 20896 24777 20924
rect 24728 20884 24734 20896
rect 24765 20893 24777 20896
rect 24811 20893 24823 20927
rect 25041 20927 25099 20933
rect 25041 20924 25053 20927
rect 24765 20887 24823 20893
rect 24872 20896 25053 20924
rect 24118 20816 24124 20868
rect 24176 20856 24182 20868
rect 24581 20859 24639 20865
rect 24581 20856 24593 20859
rect 24176 20828 24593 20856
rect 24176 20816 24182 20828
rect 24581 20825 24593 20828
rect 24627 20825 24639 20859
rect 24872 20856 24900 20896
rect 25041 20893 25053 20896
rect 25087 20924 25099 20927
rect 25498 20924 25504 20936
rect 25087 20896 25504 20924
rect 25087 20893 25099 20896
rect 25041 20887 25099 20893
rect 25498 20884 25504 20896
rect 25556 20924 25562 20936
rect 28718 20924 28724 20936
rect 25556 20896 28724 20924
rect 25556 20884 25562 20896
rect 28718 20884 28724 20896
rect 28776 20884 28782 20936
rect 31680 20933 31708 20964
rect 33045 20961 33057 20964
rect 33091 20961 33103 20995
rect 33045 20955 33103 20961
rect 31572 20927 31630 20933
rect 31572 20893 31584 20927
rect 31618 20893 31630 20927
rect 31572 20887 31630 20893
rect 31665 20927 31723 20933
rect 31665 20893 31677 20927
rect 31711 20893 31723 20927
rect 32214 20924 32220 20936
rect 32175 20896 32220 20924
rect 31665 20887 31723 20893
rect 24581 20819 24639 20825
rect 24688 20828 24900 20856
rect 24688 20788 24716 20828
rect 27338 20816 27344 20868
rect 27396 20856 27402 20868
rect 29086 20856 29092 20868
rect 27396 20828 29092 20856
rect 27396 20816 27402 20828
rect 29086 20816 29092 20828
rect 29144 20816 29150 20868
rect 31588 20856 31616 20887
rect 32214 20884 32220 20896
rect 32272 20884 32278 20936
rect 32306 20884 32312 20936
rect 32364 20924 32370 20936
rect 32401 20927 32459 20933
rect 32401 20924 32413 20927
rect 32364 20896 32413 20924
rect 32364 20884 32370 20896
rect 32401 20893 32413 20896
rect 32447 20893 32459 20927
rect 32950 20924 32956 20936
rect 32911 20896 32956 20924
rect 32401 20887 32459 20893
rect 32950 20884 32956 20896
rect 33008 20884 33014 20936
rect 33137 20927 33195 20933
rect 33137 20924 33149 20927
rect 33060 20896 33149 20924
rect 33060 20868 33088 20896
rect 33137 20893 33149 20896
rect 33183 20893 33195 20927
rect 33137 20887 33195 20893
rect 32766 20856 32772 20868
rect 31588 20828 32772 20856
rect 32766 20816 32772 20828
rect 32824 20816 32830 20868
rect 33042 20816 33048 20868
rect 33100 20816 33106 20868
rect 24946 20788 24952 20800
rect 24044 20760 24716 20788
rect 24907 20760 24952 20788
rect 24946 20748 24952 20760
rect 25004 20748 25010 20800
rect 29104 20788 29132 20816
rect 32214 20788 32220 20800
rect 29104 20760 32220 20788
rect 32214 20748 32220 20760
rect 32272 20788 32278 20800
rect 32398 20788 32404 20800
rect 32272 20760 32404 20788
rect 32272 20748 32278 20760
rect 32398 20748 32404 20760
rect 32456 20748 32462 20800
rect 1104 20698 35027 20720
rect 1104 20646 9390 20698
rect 9442 20646 9454 20698
rect 9506 20646 9518 20698
rect 9570 20646 9582 20698
rect 9634 20646 9646 20698
rect 9698 20646 17831 20698
rect 17883 20646 17895 20698
rect 17947 20646 17959 20698
rect 18011 20646 18023 20698
rect 18075 20646 18087 20698
rect 18139 20646 26272 20698
rect 26324 20646 26336 20698
rect 26388 20646 26400 20698
rect 26452 20646 26464 20698
rect 26516 20646 26528 20698
rect 26580 20646 34713 20698
rect 34765 20646 34777 20698
rect 34829 20646 34841 20698
rect 34893 20646 34905 20698
rect 34957 20646 34969 20698
rect 35021 20646 35027 20698
rect 1104 20624 35027 20646
rect 7837 20587 7895 20593
rect 7837 20553 7849 20587
rect 7883 20584 7895 20587
rect 8294 20584 8300 20596
rect 7883 20556 8300 20584
rect 7883 20553 7895 20556
rect 7837 20547 7895 20553
rect 8294 20544 8300 20556
rect 8352 20544 8358 20596
rect 8389 20587 8447 20593
rect 8389 20553 8401 20587
rect 8435 20553 8447 20587
rect 20990 20584 20996 20596
rect 20951 20556 20996 20584
rect 8389 20547 8447 20553
rect 3602 20516 3608 20528
rect 3563 20488 3608 20516
rect 3602 20476 3608 20488
rect 3660 20476 3666 20528
rect 7469 20519 7527 20525
rect 7469 20485 7481 20519
rect 7515 20516 7527 20519
rect 7742 20516 7748 20528
rect 7515 20488 7748 20516
rect 7515 20485 7527 20488
rect 7469 20479 7527 20485
rect 7742 20476 7748 20488
rect 7800 20516 7806 20528
rect 8404 20516 8432 20547
rect 20990 20544 20996 20556
rect 21048 20544 21054 20596
rect 21634 20544 21640 20596
rect 21692 20584 21698 20596
rect 22189 20587 22247 20593
rect 22189 20584 22201 20587
rect 21692 20556 22201 20584
rect 21692 20544 21698 20556
rect 22189 20553 22201 20556
rect 22235 20584 22247 20587
rect 22278 20584 22284 20596
rect 22235 20556 22284 20584
rect 22235 20553 22247 20556
rect 22189 20547 22247 20553
rect 22278 20544 22284 20556
rect 22336 20584 22342 20596
rect 24670 20584 24676 20596
rect 22336 20556 24676 20584
rect 22336 20544 22342 20556
rect 24670 20544 24676 20556
rect 24728 20584 24734 20596
rect 25958 20584 25964 20596
rect 24728 20556 25964 20584
rect 24728 20544 24734 20556
rect 25958 20544 25964 20556
rect 26016 20544 26022 20596
rect 31570 20584 31576 20596
rect 31531 20556 31576 20584
rect 31570 20544 31576 20556
rect 31628 20544 31634 20596
rect 32582 20584 32588 20596
rect 32543 20556 32588 20584
rect 32582 20544 32588 20556
rect 32640 20544 32646 20596
rect 14274 20516 14280 20528
rect 7800 20488 8432 20516
rect 13464 20488 14280 20516
rect 7800 20476 7806 20488
rect 3142 20448 3148 20460
rect 3103 20420 3148 20448
rect 3142 20408 3148 20420
rect 3200 20408 3206 20460
rect 3237 20451 3295 20457
rect 3237 20417 3249 20451
rect 3283 20448 3295 20451
rect 3970 20448 3976 20460
rect 3283 20420 3976 20448
rect 3283 20417 3295 20420
rect 3237 20411 3295 20417
rect 3970 20408 3976 20420
rect 4028 20408 4034 20460
rect 4433 20451 4491 20457
rect 4433 20417 4445 20451
rect 4479 20417 4491 20451
rect 4433 20411 4491 20417
rect 3050 20340 3056 20392
rect 3108 20380 3114 20392
rect 3418 20380 3424 20392
rect 3108 20352 3424 20380
rect 3108 20340 3114 20352
rect 3418 20340 3424 20352
rect 3476 20380 3482 20392
rect 3513 20383 3571 20389
rect 3513 20380 3525 20383
rect 3476 20352 3525 20380
rect 3476 20340 3482 20352
rect 3513 20349 3525 20352
rect 3559 20349 3571 20383
rect 4062 20380 4068 20392
rect 4023 20352 4068 20380
rect 3513 20343 3571 20349
rect 4062 20340 4068 20352
rect 4120 20340 4126 20392
rect 4338 20380 4344 20392
rect 4299 20352 4344 20380
rect 4338 20340 4344 20352
rect 4396 20340 4402 20392
rect 1854 20272 1860 20324
rect 1912 20312 1918 20324
rect 4448 20312 4476 20411
rect 7282 20408 7288 20460
rect 7340 20448 7346 20460
rect 7377 20451 7435 20457
rect 7377 20448 7389 20451
rect 7340 20420 7389 20448
rect 7340 20408 7346 20420
rect 7377 20417 7389 20420
rect 7423 20417 7435 20451
rect 7377 20411 7435 20417
rect 7653 20451 7711 20457
rect 7653 20417 7665 20451
rect 7699 20448 7711 20451
rect 8018 20448 8024 20460
rect 7699 20420 8024 20448
rect 7699 20417 7711 20420
rect 7653 20411 7711 20417
rect 8018 20408 8024 20420
rect 8076 20408 8082 20460
rect 8297 20451 8355 20457
rect 8297 20417 8309 20451
rect 8343 20417 8355 20451
rect 8478 20448 8484 20460
rect 8439 20420 8484 20448
rect 8297 20411 8355 20417
rect 8312 20380 8340 20411
rect 8478 20408 8484 20420
rect 8536 20408 8542 20460
rect 8573 20451 8631 20457
rect 8573 20417 8585 20451
rect 8619 20448 8631 20451
rect 10226 20448 10232 20460
rect 8619 20420 10232 20448
rect 8619 20417 8631 20420
rect 8573 20411 8631 20417
rect 10226 20408 10232 20420
rect 10284 20408 10290 20460
rect 11054 20448 11060 20460
rect 11015 20420 11060 20448
rect 11054 20408 11060 20420
rect 11112 20408 11118 20460
rect 13464 20457 13492 20488
rect 14274 20476 14280 20488
rect 14332 20476 14338 20528
rect 16206 20516 16212 20528
rect 14384 20488 16212 20516
rect 13449 20451 13507 20457
rect 13449 20417 13461 20451
rect 13495 20417 13507 20451
rect 13449 20411 13507 20417
rect 13817 20451 13875 20457
rect 13817 20417 13829 20451
rect 13863 20417 13875 20451
rect 13817 20411 13875 20417
rect 14001 20451 14059 20457
rect 14001 20417 14013 20451
rect 14047 20448 14059 20451
rect 14384 20448 14412 20488
rect 16206 20476 16212 20488
rect 16264 20476 16270 20528
rect 19702 20476 19708 20528
rect 19760 20516 19766 20528
rect 20625 20519 20683 20525
rect 20625 20516 20637 20519
rect 19760 20488 20637 20516
rect 19760 20476 19766 20488
rect 20625 20485 20637 20488
rect 20671 20485 20683 20519
rect 20625 20479 20683 20485
rect 20714 20476 20720 20528
rect 20772 20516 20778 20528
rect 20772 20488 20817 20516
rect 20772 20476 20778 20488
rect 22370 20476 22376 20528
rect 22428 20516 22434 20528
rect 23201 20519 23259 20525
rect 23201 20516 23213 20519
rect 22428 20488 23213 20516
rect 22428 20476 22434 20488
rect 23201 20485 23213 20488
rect 23247 20485 23259 20519
rect 23201 20479 23259 20485
rect 15102 20448 15108 20460
rect 14047 20420 14412 20448
rect 15063 20420 15108 20448
rect 14047 20417 14059 20420
rect 14001 20411 14059 20417
rect 8938 20380 8944 20392
rect 8312 20352 8944 20380
rect 8938 20340 8944 20352
rect 8996 20340 9002 20392
rect 10410 20380 10416 20392
rect 10371 20352 10416 20380
rect 10410 20340 10416 20352
rect 10468 20340 10474 20392
rect 12805 20383 12863 20389
rect 12805 20380 12817 20383
rect 12406 20352 12817 20380
rect 5074 20312 5080 20324
rect 1912 20284 5080 20312
rect 1912 20272 1918 20284
rect 5074 20272 5080 20284
rect 5132 20272 5138 20324
rect 6914 20272 6920 20324
rect 6972 20312 6978 20324
rect 7834 20312 7840 20324
rect 6972 20284 7840 20312
rect 6972 20272 6978 20284
rect 7834 20272 7840 20284
rect 7892 20312 7898 20324
rect 12406 20312 12434 20352
rect 12805 20349 12817 20352
rect 12851 20349 12863 20383
rect 12805 20343 12863 20349
rect 13541 20383 13599 20389
rect 13541 20349 13553 20383
rect 13587 20380 13599 20383
rect 13722 20380 13728 20392
rect 13587 20352 13728 20380
rect 13587 20349 13599 20352
rect 13541 20343 13599 20349
rect 13722 20340 13728 20352
rect 13780 20340 13786 20392
rect 7892 20284 12434 20312
rect 7892 20272 7898 20284
rect 13170 20272 13176 20324
rect 13228 20312 13234 20324
rect 13832 20312 13860 20411
rect 13228 20284 13860 20312
rect 13228 20272 13234 20284
rect 2774 20204 2780 20256
rect 2832 20244 2838 20256
rect 2961 20247 3019 20253
rect 2961 20244 2973 20247
rect 2832 20216 2973 20244
rect 2832 20204 2838 20216
rect 2961 20213 2973 20216
rect 3007 20213 3019 20247
rect 2961 20207 3019 20213
rect 12894 20204 12900 20256
rect 12952 20244 12958 20256
rect 14016 20244 14044 20411
rect 15102 20408 15108 20420
rect 15160 20408 15166 20460
rect 15378 20408 15384 20460
rect 15436 20448 15442 20460
rect 15657 20451 15715 20457
rect 15657 20448 15669 20451
rect 15436 20420 15669 20448
rect 15436 20408 15442 20420
rect 15657 20417 15669 20420
rect 15703 20417 15715 20451
rect 15657 20411 15715 20417
rect 15746 20408 15752 20460
rect 15804 20448 15810 20460
rect 15841 20451 15899 20457
rect 15841 20448 15853 20451
rect 15804 20420 15853 20448
rect 15804 20408 15810 20420
rect 15841 20417 15853 20420
rect 15887 20417 15899 20451
rect 15841 20411 15899 20417
rect 19981 20451 20039 20457
rect 19981 20417 19993 20451
rect 20027 20448 20039 20451
rect 20346 20448 20352 20460
rect 20027 20420 20352 20448
rect 20027 20417 20039 20420
rect 19981 20411 20039 20417
rect 20346 20408 20352 20420
rect 20404 20408 20410 20460
rect 20441 20451 20499 20457
rect 20441 20417 20453 20451
rect 20487 20417 20499 20451
rect 20441 20411 20499 20417
rect 14737 20383 14795 20389
rect 14737 20349 14749 20383
rect 14783 20349 14795 20383
rect 14737 20343 14795 20349
rect 16025 20383 16083 20389
rect 16025 20349 16037 20383
rect 16071 20380 16083 20383
rect 16942 20380 16948 20392
rect 16071 20352 16948 20380
rect 16071 20349 16083 20352
rect 16025 20343 16083 20349
rect 14090 20272 14096 20324
rect 14148 20312 14154 20324
rect 14752 20312 14780 20343
rect 16942 20340 16948 20352
rect 17000 20380 17006 20392
rect 17218 20380 17224 20392
rect 17000 20352 17224 20380
rect 17000 20340 17006 20352
rect 17218 20340 17224 20352
rect 17276 20340 17282 20392
rect 17310 20340 17316 20392
rect 17368 20380 17374 20392
rect 20456 20380 20484 20411
rect 20530 20408 20536 20460
rect 20588 20448 20594 20460
rect 20809 20451 20867 20457
rect 20809 20448 20821 20451
rect 20588 20420 20821 20448
rect 20588 20408 20594 20420
rect 20809 20417 20821 20420
rect 20855 20417 20867 20451
rect 20809 20411 20867 20417
rect 20990 20408 20996 20460
rect 21048 20448 21054 20460
rect 22097 20451 22155 20457
rect 22097 20448 22109 20451
rect 21048 20420 22109 20448
rect 21048 20408 21054 20420
rect 22097 20417 22109 20420
rect 22143 20417 22155 20451
rect 27982 20448 27988 20460
rect 27943 20420 27988 20448
rect 22097 20411 22155 20417
rect 27982 20408 27988 20420
rect 28040 20408 28046 20460
rect 31573 20451 31631 20457
rect 31573 20417 31585 20451
rect 31619 20417 31631 20451
rect 31573 20411 31631 20417
rect 31757 20451 31815 20457
rect 31757 20417 31769 20451
rect 31803 20448 31815 20451
rect 32582 20448 32588 20460
rect 31803 20420 32588 20448
rect 31803 20417 31815 20420
rect 31757 20411 31815 20417
rect 27890 20380 27896 20392
rect 17368 20352 20484 20380
rect 27851 20352 27896 20380
rect 17368 20340 17374 20352
rect 27890 20340 27896 20352
rect 27948 20340 27954 20392
rect 31588 20380 31616 20411
rect 32582 20408 32588 20420
rect 32640 20408 32646 20460
rect 32766 20448 32772 20460
rect 32727 20420 32772 20448
rect 32766 20408 32772 20420
rect 32824 20408 32830 20460
rect 33042 20448 33048 20460
rect 33003 20420 33048 20448
rect 33042 20408 33048 20420
rect 33100 20408 33106 20460
rect 31938 20380 31944 20392
rect 31588 20352 31944 20380
rect 31938 20340 31944 20352
rect 31996 20340 32002 20392
rect 14148 20284 14780 20312
rect 14148 20272 14154 20284
rect 12952 20216 14044 20244
rect 14752 20244 14780 20284
rect 14826 20272 14832 20324
rect 14884 20312 14890 20324
rect 14884 20284 18828 20312
rect 14884 20272 14890 20284
rect 17402 20244 17408 20256
rect 14752 20216 17408 20244
rect 12952 20204 12958 20216
rect 17402 20204 17408 20216
rect 17460 20204 17466 20256
rect 18690 20244 18696 20256
rect 18651 20216 18696 20244
rect 18690 20204 18696 20216
rect 18748 20204 18754 20256
rect 18800 20244 18828 20284
rect 20806 20272 20812 20324
rect 20864 20312 20870 20324
rect 24489 20315 24547 20321
rect 24489 20312 24501 20315
rect 20864 20284 24501 20312
rect 20864 20272 20870 20284
rect 24489 20281 24501 20284
rect 24535 20281 24547 20315
rect 24489 20275 24547 20281
rect 32306 20272 32312 20324
rect 32364 20312 32370 20324
rect 32950 20312 32956 20324
rect 32364 20284 32956 20312
rect 32364 20272 32370 20284
rect 32950 20272 32956 20284
rect 33008 20272 33014 20324
rect 27617 20247 27675 20253
rect 27617 20244 27629 20247
rect 18800 20216 27629 20244
rect 27617 20213 27629 20216
rect 27663 20213 27675 20247
rect 27617 20207 27675 20213
rect 27985 20247 28043 20253
rect 27985 20213 27997 20247
rect 28031 20244 28043 20247
rect 28074 20244 28080 20256
rect 28031 20216 28080 20244
rect 28031 20213 28043 20216
rect 27985 20207 28043 20213
rect 28074 20204 28080 20216
rect 28132 20204 28138 20256
rect 1104 20154 34868 20176
rect 1104 20102 5170 20154
rect 5222 20102 5234 20154
rect 5286 20102 5298 20154
rect 5350 20102 5362 20154
rect 5414 20102 5426 20154
rect 5478 20102 13611 20154
rect 13663 20102 13675 20154
rect 13727 20102 13739 20154
rect 13791 20102 13803 20154
rect 13855 20102 13867 20154
rect 13919 20102 22052 20154
rect 22104 20102 22116 20154
rect 22168 20102 22180 20154
rect 22232 20102 22244 20154
rect 22296 20102 22308 20154
rect 22360 20102 30493 20154
rect 30545 20102 30557 20154
rect 30609 20102 30621 20154
rect 30673 20102 30685 20154
rect 30737 20102 30749 20154
rect 30801 20102 34868 20154
rect 1104 20080 34868 20102
rect 3970 20040 3976 20052
rect 3931 20012 3976 20040
rect 3970 20000 3976 20012
rect 4028 20000 4034 20052
rect 4706 20000 4712 20052
rect 4764 20040 4770 20052
rect 5074 20040 5080 20052
rect 4764 20012 5080 20040
rect 4764 20000 4770 20012
rect 5074 20000 5080 20012
rect 5132 20000 5138 20052
rect 7561 20043 7619 20049
rect 7561 20009 7573 20043
rect 7607 20040 7619 20043
rect 7650 20040 7656 20052
rect 7607 20012 7656 20040
rect 7607 20009 7619 20012
rect 7561 20003 7619 20009
rect 3786 19932 3792 19984
rect 3844 19972 3850 19984
rect 6638 19972 6644 19984
rect 3844 19944 6644 19972
rect 3844 19932 3850 19944
rect 2409 19907 2467 19913
rect 2409 19904 2421 19907
rect 1688 19876 2421 19904
rect 1688 19845 1716 19876
rect 2409 19873 2421 19876
rect 2455 19904 2467 19907
rect 4338 19904 4344 19916
rect 2455 19876 4344 19904
rect 2455 19873 2467 19876
rect 2409 19867 2467 19873
rect 4338 19864 4344 19876
rect 4396 19864 4402 19916
rect 4448 19876 4844 19904
rect 1673 19839 1731 19845
rect 1673 19805 1685 19839
rect 1719 19805 1731 19839
rect 1854 19836 1860 19848
rect 1815 19808 1860 19836
rect 1673 19799 1731 19805
rect 1854 19796 1860 19808
rect 1912 19796 1918 19848
rect 2869 19839 2927 19845
rect 2869 19805 2881 19839
rect 2915 19805 2927 19839
rect 2869 19799 2927 19805
rect 3145 19839 3203 19845
rect 3145 19805 3157 19839
rect 3191 19836 3203 19839
rect 3191 19808 4108 19836
rect 3191 19805 3203 19808
rect 3145 19799 3203 19805
rect 2884 19768 2912 19799
rect 3234 19768 3240 19780
rect 2884 19740 3240 19768
rect 3234 19728 3240 19740
rect 3292 19768 3298 19780
rect 3970 19768 3976 19780
rect 3292 19740 3976 19768
rect 3292 19728 3298 19740
rect 3970 19728 3976 19740
rect 4028 19728 4034 19780
rect 1857 19703 1915 19709
rect 1857 19669 1869 19703
rect 1903 19700 1915 19703
rect 3326 19700 3332 19712
rect 1903 19672 3332 19700
rect 1903 19669 1915 19672
rect 1857 19663 1915 19669
rect 3326 19660 3332 19672
rect 3384 19660 3390 19712
rect 4080 19700 4108 19808
rect 4154 19796 4160 19848
rect 4212 19836 4218 19848
rect 4212 19808 4257 19836
rect 4212 19796 4218 19808
rect 4246 19768 4252 19780
rect 4207 19740 4252 19768
rect 4246 19728 4252 19740
rect 4304 19728 4310 19780
rect 4341 19771 4399 19777
rect 4341 19737 4353 19771
rect 4387 19768 4399 19771
rect 4448 19768 4476 19876
rect 4525 19839 4583 19845
rect 4525 19805 4537 19839
rect 4571 19805 4583 19839
rect 4525 19799 4583 19805
rect 4387 19740 4476 19768
rect 4387 19737 4399 19740
rect 4341 19731 4399 19737
rect 4430 19700 4436 19712
rect 4080 19672 4436 19700
rect 4430 19660 4436 19672
rect 4488 19660 4494 19712
rect 4540 19700 4568 19799
rect 4614 19796 4620 19848
rect 4672 19836 4678 19848
rect 4672 19808 4717 19836
rect 4672 19796 4678 19808
rect 4816 19768 4844 19876
rect 5276 19845 5304 19944
rect 6638 19932 6644 19944
rect 6696 19932 6702 19984
rect 7098 19972 7104 19984
rect 7059 19944 7104 19972
rect 7098 19932 7104 19944
rect 7156 19932 7162 19984
rect 7576 19904 7604 20003
rect 7650 20000 7656 20012
rect 7708 20000 7714 20052
rect 14553 20043 14611 20049
rect 14553 20009 14565 20043
rect 14599 20040 14611 20043
rect 15286 20040 15292 20052
rect 14599 20012 15292 20040
rect 14599 20009 14611 20012
rect 14553 20003 14611 20009
rect 15286 20000 15292 20012
rect 15344 20000 15350 20052
rect 20073 20043 20131 20049
rect 20073 20009 20085 20043
rect 20119 20040 20131 20043
rect 24762 20040 24768 20052
rect 20119 20012 24768 20040
rect 20119 20009 20131 20012
rect 20073 20003 20131 20009
rect 24762 20000 24768 20012
rect 24820 20000 24826 20052
rect 7742 19972 7748 19984
rect 7703 19944 7748 19972
rect 7742 19932 7748 19944
rect 7800 19932 7806 19984
rect 9125 19975 9183 19981
rect 9125 19941 9137 19975
rect 9171 19941 9183 19975
rect 20990 19972 20996 19984
rect 9125 19935 9183 19941
rect 18248 19944 20996 19972
rect 9140 19904 9168 19935
rect 10505 19907 10563 19913
rect 10505 19904 10517 19907
rect 6932 19876 7604 19904
rect 8312 19876 9168 19904
rect 9416 19876 10517 19904
rect 5261 19839 5319 19845
rect 5261 19805 5273 19839
rect 5307 19805 5319 19839
rect 5442 19836 5448 19848
rect 5403 19808 5448 19836
rect 5261 19799 5319 19805
rect 5442 19796 5448 19808
rect 5500 19796 5506 19848
rect 6932 19845 6960 19876
rect 6825 19839 6883 19845
rect 6825 19805 6837 19839
rect 6871 19805 6883 19839
rect 6825 19799 6883 19805
rect 6917 19839 6975 19845
rect 6917 19805 6929 19839
rect 6963 19805 6975 19839
rect 6917 19799 6975 19805
rect 7101 19839 7159 19845
rect 7101 19805 7113 19839
rect 7147 19836 7159 19839
rect 7374 19836 7380 19848
rect 7147 19808 7380 19836
rect 7147 19805 7159 19808
rect 7101 19799 7159 19805
rect 6546 19768 6552 19780
rect 4816 19740 6552 19768
rect 6546 19728 6552 19740
rect 6604 19728 6610 19780
rect 6840 19768 6868 19799
rect 7374 19796 7380 19808
rect 7432 19796 7438 19848
rect 8018 19836 8024 19848
rect 7931 19808 8024 19836
rect 8018 19796 8024 19808
rect 8076 19836 8082 19848
rect 8312 19836 8340 19876
rect 8076 19808 8340 19836
rect 8076 19796 8082 19808
rect 8478 19796 8484 19848
rect 8536 19836 8542 19848
rect 9416 19845 9444 19876
rect 10505 19873 10517 19876
rect 10551 19873 10563 19907
rect 11882 19904 11888 19916
rect 10505 19867 10563 19873
rect 10796 19876 11888 19904
rect 9401 19839 9459 19845
rect 9401 19836 9413 19839
rect 8536 19808 9413 19836
rect 8536 19796 8542 19808
rect 9401 19805 9413 19808
rect 9447 19805 9459 19839
rect 9401 19799 9459 19805
rect 9950 19796 9956 19848
rect 10008 19836 10014 19848
rect 10410 19836 10416 19848
rect 10008 19808 10416 19836
rect 10008 19796 10014 19808
rect 10410 19796 10416 19808
rect 10468 19796 10474 19848
rect 10796 19845 10824 19876
rect 11882 19864 11888 19876
rect 11940 19864 11946 19916
rect 13725 19907 13783 19913
rect 13725 19873 13737 19907
rect 13771 19904 13783 19907
rect 15102 19904 15108 19916
rect 13771 19876 15108 19904
rect 13771 19873 13783 19876
rect 13725 19867 13783 19873
rect 15102 19864 15108 19876
rect 15160 19864 15166 19916
rect 17034 19904 17040 19916
rect 15396 19876 17040 19904
rect 10781 19839 10839 19845
rect 10781 19805 10793 19839
rect 10827 19805 10839 19839
rect 10781 19799 10839 19805
rect 10870 19796 10876 19848
rect 10928 19836 10934 19848
rect 11701 19839 11759 19845
rect 11701 19836 11713 19839
rect 10928 19808 11713 19836
rect 10928 19796 10934 19808
rect 11701 19805 11713 19808
rect 11747 19805 11759 19839
rect 11701 19799 11759 19805
rect 12710 19796 12716 19848
rect 12768 19836 12774 19848
rect 13170 19836 13176 19848
rect 12768 19808 13176 19836
rect 12768 19796 12774 19808
rect 13170 19796 13176 19808
rect 13228 19836 13234 19848
rect 13357 19839 13415 19845
rect 13357 19836 13369 19839
rect 13228 19808 13369 19836
rect 13228 19796 13234 19808
rect 13357 19805 13369 19808
rect 13403 19805 13415 19839
rect 13357 19799 13415 19805
rect 13446 19796 13452 19848
rect 13504 19836 13510 19848
rect 13541 19839 13599 19845
rect 13541 19836 13553 19839
rect 13504 19808 13553 19836
rect 13504 19796 13510 19808
rect 13541 19805 13553 19808
rect 13587 19805 13599 19839
rect 14458 19836 14464 19848
rect 14419 19808 14464 19836
rect 13541 19799 13599 19805
rect 14458 19796 14464 19808
rect 14516 19796 14522 19848
rect 15396 19845 15424 19876
rect 17034 19864 17040 19876
rect 17092 19904 17098 19916
rect 17405 19907 17463 19913
rect 17405 19904 17417 19907
rect 17092 19876 17417 19904
rect 17092 19864 17098 19876
rect 17405 19873 17417 19876
rect 17451 19873 17463 19907
rect 17405 19867 17463 19873
rect 18248 19848 18276 19944
rect 20990 19932 20996 19944
rect 21048 19932 21054 19984
rect 32306 19972 32312 19984
rect 32267 19944 32312 19972
rect 32306 19932 32312 19944
rect 32364 19932 32370 19984
rect 19334 19864 19340 19916
rect 19392 19904 19398 19916
rect 20530 19904 20536 19916
rect 19392 19876 20536 19904
rect 19392 19864 19398 19876
rect 15381 19839 15439 19845
rect 15381 19805 15393 19839
rect 15427 19805 15439 19839
rect 15381 19799 15439 19805
rect 15657 19839 15715 19845
rect 15657 19805 15669 19839
rect 15703 19836 15715 19839
rect 15746 19836 15752 19848
rect 15703 19808 15752 19836
rect 15703 19805 15715 19808
rect 15657 19799 15715 19805
rect 7282 19768 7288 19780
rect 6840 19740 7288 19768
rect 7282 19728 7288 19740
rect 7340 19728 7346 19780
rect 8938 19728 8944 19780
rect 8996 19768 9002 19780
rect 9125 19771 9183 19777
rect 9125 19768 9137 19771
rect 8996 19740 9137 19768
rect 8996 19728 9002 19740
rect 9125 19737 9137 19740
rect 9171 19737 9183 19771
rect 9125 19731 9183 19737
rect 9309 19771 9367 19777
rect 9309 19737 9321 19771
rect 9355 19768 9367 19771
rect 9766 19768 9772 19780
rect 9355 19740 9772 19768
rect 9355 19737 9367 19740
rect 9309 19731 9367 19737
rect 9766 19728 9772 19740
rect 9824 19768 9830 19780
rect 10226 19768 10232 19780
rect 9824 19740 10232 19768
rect 9824 19728 9830 19740
rect 10226 19728 10232 19740
rect 10284 19728 10290 19780
rect 12434 19728 12440 19780
rect 12492 19768 12498 19780
rect 15672 19768 15700 19799
rect 15746 19796 15752 19808
rect 15804 19796 15810 19848
rect 15838 19796 15844 19848
rect 15896 19836 15902 19848
rect 16209 19839 16267 19845
rect 16209 19836 16221 19839
rect 15896 19808 16221 19836
rect 15896 19796 15902 19808
rect 16209 19805 16221 19808
rect 16255 19805 16267 19839
rect 17126 19836 17132 19848
rect 16209 19799 16267 19805
rect 16592 19808 17132 19836
rect 16592 19768 16620 19808
rect 17126 19796 17132 19808
rect 17184 19796 17190 19848
rect 17957 19839 18015 19845
rect 17957 19805 17969 19839
rect 18003 19836 18015 19839
rect 18230 19836 18236 19848
rect 18003 19808 18236 19836
rect 18003 19805 18015 19808
rect 17957 19799 18015 19805
rect 18230 19796 18236 19808
rect 18288 19796 18294 19848
rect 19426 19836 19432 19848
rect 19387 19808 19432 19836
rect 19426 19796 19432 19808
rect 19484 19796 19490 19848
rect 19518 19796 19524 19848
rect 19576 19836 19582 19848
rect 19794 19836 19800 19848
rect 19576 19808 19621 19836
rect 19755 19808 19800 19836
rect 19576 19796 19582 19808
rect 19794 19796 19800 19808
rect 19852 19796 19858 19848
rect 19904 19845 19932 19876
rect 20530 19864 20536 19876
rect 20588 19864 20594 19916
rect 22557 19907 22615 19913
rect 22557 19873 22569 19907
rect 22603 19904 22615 19907
rect 23198 19904 23204 19916
rect 22603 19876 23204 19904
rect 22603 19873 22615 19876
rect 22557 19867 22615 19873
rect 23198 19864 23204 19876
rect 23256 19864 23262 19916
rect 19894 19839 19952 19845
rect 19894 19805 19906 19839
rect 19940 19805 19952 19839
rect 19894 19799 19952 19805
rect 28537 19839 28595 19845
rect 28537 19805 28549 19839
rect 28583 19805 28595 19839
rect 28810 19836 28816 19848
rect 28771 19808 28816 19836
rect 28537 19799 28595 19805
rect 16758 19768 16764 19780
rect 12492 19740 16620 19768
rect 16719 19740 16764 19768
rect 12492 19728 12498 19740
rect 16758 19728 16764 19740
rect 16816 19728 16822 19780
rect 17678 19728 17684 19780
rect 17736 19768 17742 19780
rect 19702 19768 19708 19780
rect 17736 19740 19708 19768
rect 17736 19728 17742 19740
rect 19702 19728 19708 19740
rect 19760 19728 19766 19780
rect 20806 19768 20812 19780
rect 20767 19740 20812 19768
rect 20806 19728 20812 19740
rect 20864 19728 20870 19780
rect 28552 19768 28580 19799
rect 28810 19796 28816 19808
rect 28868 19796 28874 19848
rect 28902 19796 28908 19848
rect 28960 19836 28966 19848
rect 28997 19839 29055 19845
rect 28997 19836 29009 19839
rect 28960 19808 29009 19836
rect 28960 19796 28966 19808
rect 28997 19805 29009 19808
rect 29043 19836 29055 19839
rect 31754 19836 31760 19848
rect 29043 19808 31760 19836
rect 29043 19805 29055 19808
rect 28997 19799 29055 19805
rect 31754 19796 31760 19808
rect 31812 19796 31818 19848
rect 31938 19836 31944 19848
rect 31899 19808 31944 19836
rect 31938 19796 31944 19808
rect 31996 19796 32002 19848
rect 32214 19836 32220 19848
rect 32175 19808 32220 19836
rect 32214 19796 32220 19808
rect 32272 19796 32278 19848
rect 32398 19836 32404 19848
rect 32359 19808 32404 19836
rect 32398 19796 32404 19808
rect 32456 19796 32462 19848
rect 32582 19836 32588 19848
rect 32543 19808 32588 19836
rect 32582 19796 32588 19808
rect 32640 19796 32646 19848
rect 28718 19768 28724 19780
rect 28552 19740 28724 19768
rect 28718 19728 28724 19740
rect 28776 19728 28782 19780
rect 7466 19700 7472 19712
rect 4540 19672 7472 19700
rect 7466 19660 7472 19672
rect 7524 19660 7530 19712
rect 11514 19700 11520 19712
rect 11475 19672 11520 19700
rect 11514 19660 11520 19672
rect 11572 19660 11578 19712
rect 15197 19703 15255 19709
rect 15197 19669 15209 19703
rect 15243 19700 15255 19703
rect 15286 19700 15292 19712
rect 15243 19672 15292 19700
rect 15243 19669 15255 19672
rect 15197 19663 15255 19669
rect 15286 19660 15292 19672
rect 15344 19660 15350 19712
rect 15565 19703 15623 19709
rect 15565 19669 15577 19703
rect 15611 19700 15623 19703
rect 17310 19700 17316 19712
rect 15611 19672 17316 19700
rect 15611 19669 15623 19672
rect 15565 19663 15623 19669
rect 17310 19660 17316 19672
rect 17368 19660 17374 19712
rect 19426 19660 19432 19712
rect 19484 19700 19490 19712
rect 20254 19700 20260 19712
rect 19484 19672 20260 19700
rect 19484 19660 19490 19672
rect 20254 19660 20260 19672
rect 20312 19660 20318 19712
rect 28166 19660 28172 19712
rect 28224 19700 28230 19712
rect 28353 19703 28411 19709
rect 28353 19700 28365 19703
rect 28224 19672 28365 19700
rect 28224 19660 28230 19672
rect 28353 19669 28365 19672
rect 28399 19669 28411 19703
rect 28353 19663 28411 19669
rect 1104 19610 35027 19632
rect 1104 19558 9390 19610
rect 9442 19558 9454 19610
rect 9506 19558 9518 19610
rect 9570 19558 9582 19610
rect 9634 19558 9646 19610
rect 9698 19558 17831 19610
rect 17883 19558 17895 19610
rect 17947 19558 17959 19610
rect 18011 19558 18023 19610
rect 18075 19558 18087 19610
rect 18139 19558 26272 19610
rect 26324 19558 26336 19610
rect 26388 19558 26400 19610
rect 26452 19558 26464 19610
rect 26516 19558 26528 19610
rect 26580 19558 34713 19610
rect 34765 19558 34777 19610
rect 34829 19558 34841 19610
rect 34893 19558 34905 19610
rect 34957 19558 34969 19610
rect 35021 19558 35027 19610
rect 1104 19536 35027 19558
rect 4062 19456 4068 19508
rect 4120 19496 4126 19508
rect 4890 19496 4896 19508
rect 4120 19468 4896 19496
rect 4120 19456 4126 19468
rect 4890 19456 4896 19468
rect 4948 19496 4954 19508
rect 6914 19496 6920 19508
rect 4948 19468 6920 19496
rect 4948 19456 4954 19468
rect 6914 19456 6920 19468
rect 6972 19456 6978 19508
rect 16301 19499 16359 19505
rect 16301 19465 16313 19499
rect 16347 19496 16359 19499
rect 17221 19499 17279 19505
rect 17221 19496 17233 19499
rect 16347 19468 17233 19496
rect 16347 19465 16359 19468
rect 16301 19459 16359 19465
rect 17221 19465 17233 19468
rect 17267 19496 17279 19499
rect 19518 19496 19524 19508
rect 17267 19468 19524 19496
rect 17267 19465 17279 19468
rect 17221 19459 17279 19465
rect 19518 19456 19524 19468
rect 19576 19456 19582 19508
rect 20714 19456 20720 19508
rect 20772 19496 20778 19508
rect 20809 19499 20867 19505
rect 20809 19496 20821 19499
rect 20772 19468 20821 19496
rect 20772 19456 20778 19468
rect 20809 19465 20821 19468
rect 20855 19496 20867 19499
rect 22097 19499 22155 19505
rect 22097 19496 22109 19499
rect 20855 19468 22109 19496
rect 20855 19465 20867 19468
rect 20809 19459 20867 19465
rect 22097 19465 22109 19468
rect 22143 19465 22155 19499
rect 23014 19496 23020 19508
rect 22097 19459 22155 19465
rect 22204 19468 23020 19496
rect 4706 19428 4712 19440
rect 4632 19400 4712 19428
rect 2501 19363 2559 19369
rect 2501 19329 2513 19363
rect 2547 19360 2559 19363
rect 2547 19332 2636 19360
rect 2547 19329 2559 19332
rect 2501 19323 2559 19329
rect 2608 19292 2636 19332
rect 2774 19320 2780 19372
rect 2832 19360 2838 19372
rect 3510 19360 3516 19372
rect 2832 19332 2877 19360
rect 2976 19332 3516 19360
rect 2832 19320 2838 19332
rect 2976 19292 3004 19332
rect 3510 19320 3516 19332
rect 3568 19360 3574 19372
rect 3878 19360 3884 19372
rect 3568 19332 3884 19360
rect 3568 19320 3574 19332
rect 3878 19320 3884 19332
rect 3936 19360 3942 19372
rect 4632 19369 4660 19400
rect 4706 19388 4712 19400
rect 4764 19388 4770 19440
rect 16758 19388 16764 19440
rect 16816 19428 16822 19440
rect 22204 19428 22232 19468
rect 23014 19456 23020 19468
rect 23072 19456 23078 19508
rect 32214 19456 32220 19508
rect 32272 19496 32278 19508
rect 32677 19499 32735 19505
rect 32677 19496 32689 19499
rect 32272 19468 32689 19496
rect 32272 19456 32278 19468
rect 32677 19465 32689 19468
rect 32723 19465 32735 19499
rect 32677 19459 32735 19465
rect 32861 19499 32919 19505
rect 32861 19465 32873 19499
rect 32907 19496 32919 19499
rect 33042 19496 33048 19508
rect 32907 19468 33048 19496
rect 32907 19465 32919 19468
rect 32861 19459 32919 19465
rect 33042 19456 33048 19468
rect 33100 19456 33106 19508
rect 16816 19400 22232 19428
rect 24765 19431 24823 19437
rect 16816 19388 16822 19400
rect 4617 19363 4675 19369
rect 3936 19332 4568 19360
rect 3936 19320 3942 19332
rect 2608 19264 3004 19292
rect 4540 19292 4568 19332
rect 4617 19329 4629 19363
rect 4663 19329 4675 19363
rect 4798 19360 4804 19372
rect 4759 19332 4804 19360
rect 4617 19323 4675 19329
rect 4798 19320 4804 19332
rect 4856 19320 4862 19372
rect 4890 19320 4896 19372
rect 4948 19360 4954 19372
rect 7101 19363 7159 19369
rect 7101 19360 7113 19363
rect 4948 19332 4993 19360
rect 5092 19332 7113 19360
rect 4948 19320 4954 19332
rect 5092 19292 5120 19332
rect 7101 19329 7113 19332
rect 7147 19329 7159 19363
rect 7101 19323 7159 19329
rect 7368 19363 7426 19369
rect 7368 19329 7380 19363
rect 7414 19360 7426 19363
rect 7650 19360 7656 19372
rect 7414 19332 7656 19360
rect 7414 19329 7426 19332
rect 7368 19323 7426 19329
rect 7650 19320 7656 19332
rect 7708 19320 7714 19372
rect 8938 19320 8944 19372
rect 8996 19360 9002 19372
rect 9033 19363 9091 19369
rect 9033 19360 9045 19363
rect 8996 19332 9045 19360
rect 8996 19320 9002 19332
rect 9033 19329 9045 19332
rect 9079 19329 9091 19363
rect 9033 19323 9091 19329
rect 9217 19363 9275 19369
rect 9217 19329 9229 19363
rect 9263 19360 9275 19363
rect 9766 19360 9772 19372
rect 9263 19332 9772 19360
rect 9263 19329 9275 19332
rect 9217 19323 9275 19329
rect 9766 19320 9772 19332
rect 9824 19320 9830 19372
rect 10318 19320 10324 19372
rect 10376 19360 10382 19372
rect 10781 19363 10839 19369
rect 10781 19360 10793 19363
rect 10376 19332 10793 19360
rect 10376 19320 10382 19332
rect 10781 19329 10793 19332
rect 10827 19329 10839 19363
rect 12434 19360 12440 19372
rect 12395 19332 12440 19360
rect 10781 19323 10839 19329
rect 12434 19320 12440 19332
rect 12492 19320 12498 19372
rect 12713 19363 12771 19369
rect 12713 19329 12725 19363
rect 12759 19360 12771 19363
rect 13262 19360 13268 19372
rect 12759 19332 13268 19360
rect 12759 19329 12771 19332
rect 12713 19323 12771 19329
rect 13262 19320 13268 19332
rect 13320 19320 13326 19372
rect 17052 19369 17080 19400
rect 24765 19397 24777 19431
rect 24811 19428 24823 19431
rect 24946 19428 24952 19440
rect 24811 19400 24952 19428
rect 24811 19397 24823 19400
rect 24765 19391 24823 19397
rect 24946 19388 24952 19400
rect 25004 19428 25010 19440
rect 31938 19428 31944 19440
rect 25004 19400 31944 19428
rect 25004 19388 25010 19400
rect 15188 19363 15246 19369
rect 15188 19329 15200 19363
rect 15234 19360 15246 19363
rect 16853 19363 16911 19369
rect 16853 19360 16865 19363
rect 15234 19332 16865 19360
rect 15234 19329 15246 19332
rect 15188 19323 15246 19329
rect 16853 19329 16865 19332
rect 16899 19329 16911 19363
rect 16853 19323 16911 19329
rect 17037 19363 17095 19369
rect 17037 19329 17049 19363
rect 17083 19329 17095 19363
rect 17037 19323 17095 19329
rect 17126 19320 17132 19372
rect 17184 19360 17190 19372
rect 17313 19363 17371 19369
rect 17313 19360 17325 19363
rect 17184 19332 17325 19360
rect 17184 19320 17190 19332
rect 17313 19329 17325 19332
rect 17359 19329 17371 19363
rect 17313 19323 17371 19329
rect 18690 19320 18696 19372
rect 18748 19360 18754 19372
rect 19429 19363 19487 19369
rect 19429 19360 19441 19363
rect 18748 19332 19441 19360
rect 18748 19320 18754 19332
rect 19429 19329 19441 19332
rect 19475 19329 19487 19363
rect 19429 19323 19487 19329
rect 19696 19363 19754 19369
rect 19696 19329 19708 19363
rect 19742 19360 19754 19363
rect 19742 19332 20944 19360
rect 19742 19329 19754 19332
rect 19696 19323 19754 19329
rect 4540 19264 5120 19292
rect 10505 19295 10563 19301
rect 10505 19261 10517 19295
rect 10551 19292 10563 19295
rect 11054 19292 11060 19304
rect 10551 19264 11060 19292
rect 10551 19261 10563 19264
rect 10505 19255 10563 19261
rect 11054 19252 11060 19264
rect 11112 19292 11118 19304
rect 11514 19292 11520 19304
rect 11112 19264 11520 19292
rect 11112 19252 11118 19264
rect 11514 19252 11520 19264
rect 11572 19252 11578 19304
rect 14734 19252 14740 19304
rect 14792 19292 14798 19304
rect 14921 19295 14979 19301
rect 14921 19292 14933 19295
rect 14792 19264 14933 19292
rect 14792 19252 14798 19264
rect 14921 19261 14933 19264
rect 14967 19261 14979 19295
rect 20916 19292 20944 19332
rect 20990 19320 20996 19372
rect 21048 19360 21054 19372
rect 22005 19363 22063 19369
rect 22005 19360 22017 19363
rect 21048 19332 22017 19360
rect 21048 19320 21054 19332
rect 22005 19329 22017 19332
rect 22051 19329 22063 19363
rect 22005 19323 22063 19329
rect 22281 19363 22339 19369
rect 22281 19329 22293 19363
rect 22327 19360 22339 19363
rect 22370 19360 22376 19372
rect 22327 19332 22376 19360
rect 22327 19329 22339 19332
rect 22281 19323 22339 19329
rect 22370 19320 22376 19332
rect 22428 19320 22434 19372
rect 23109 19363 23167 19369
rect 23109 19329 23121 19363
rect 23155 19360 23167 19363
rect 23198 19360 23204 19372
rect 23155 19332 23204 19360
rect 23155 19329 23167 19332
rect 23109 19323 23167 19329
rect 23198 19320 23204 19332
rect 23256 19320 23262 19372
rect 27249 19363 27307 19369
rect 27249 19329 27261 19363
rect 27295 19360 27307 19363
rect 27338 19360 27344 19372
rect 27295 19332 27344 19360
rect 27295 19329 27307 19332
rect 27249 19323 27307 19329
rect 27338 19320 27344 19332
rect 27396 19320 27402 19372
rect 27430 19320 27436 19372
rect 27488 19360 27494 19372
rect 28813 19363 28871 19369
rect 27488 19332 27533 19360
rect 27488 19320 27494 19332
rect 28813 19329 28825 19363
rect 28859 19360 28871 19363
rect 29086 19360 29092 19372
rect 28859 19332 28948 19360
rect 29047 19332 29092 19360
rect 28859 19329 28871 19332
rect 28813 19323 28871 19329
rect 22465 19295 22523 19301
rect 22465 19292 22477 19295
rect 20916 19264 22477 19292
rect 14921 19255 14979 19261
rect 22465 19261 22477 19264
rect 22511 19261 22523 19295
rect 23382 19292 23388 19304
rect 23343 19264 23388 19292
rect 22465 19255 22523 19261
rect 23382 19252 23388 19264
rect 23440 19252 23446 19304
rect 28718 19292 28724 19304
rect 28679 19264 28724 19292
rect 28718 19252 28724 19264
rect 28776 19252 28782 19304
rect 28920 19292 28948 19332
rect 29086 19320 29092 19332
rect 29144 19320 29150 19372
rect 29380 19369 29408 19400
rect 29365 19363 29423 19369
rect 29365 19329 29377 19363
rect 29411 19329 29423 19363
rect 29730 19360 29736 19372
rect 29691 19332 29736 19360
rect 29365 19323 29423 19329
rect 29730 19320 29736 19332
rect 29788 19320 29794 19372
rect 31202 19360 31208 19372
rect 29840 19332 31208 19360
rect 29840 19292 29868 19332
rect 31202 19320 31208 19332
rect 31260 19320 31266 19372
rect 31312 19369 31340 19400
rect 31938 19388 31944 19400
rect 31996 19428 32002 19440
rect 32309 19431 32367 19437
rect 32309 19428 32321 19431
rect 31996 19400 32321 19428
rect 31996 19388 32002 19400
rect 32309 19397 32321 19400
rect 32355 19397 32367 19431
rect 32309 19391 32367 19397
rect 32398 19388 32404 19440
rect 32456 19428 32462 19440
rect 32493 19431 32551 19437
rect 32493 19428 32505 19431
rect 32456 19400 32505 19428
rect 32456 19388 32462 19400
rect 32493 19397 32505 19400
rect 32539 19397 32551 19431
rect 32493 19391 32551 19397
rect 31297 19363 31355 19369
rect 31297 19329 31309 19363
rect 31343 19329 31355 19363
rect 31297 19323 31355 19329
rect 32582 19320 32588 19372
rect 32640 19360 32646 19372
rect 32640 19332 32685 19360
rect 32640 19320 32646 19332
rect 28920 19264 29868 19292
rect 31481 19295 31539 19301
rect 31481 19261 31493 19295
rect 31527 19261 31539 19295
rect 31754 19292 31760 19304
rect 31667 19264 31760 19292
rect 31481 19255 31539 19261
rect 4614 19224 4620 19236
rect 4575 19196 4620 19224
rect 4614 19184 4620 19196
rect 4672 19184 4678 19236
rect 9766 19224 9772 19236
rect 8036 19196 9772 19224
rect 4065 19159 4123 19165
rect 4065 19125 4077 19159
rect 4111 19156 4123 19159
rect 4246 19156 4252 19168
rect 4111 19128 4252 19156
rect 4111 19125 4123 19128
rect 4065 19119 4123 19125
rect 4246 19116 4252 19128
rect 4304 19156 4310 19168
rect 5442 19156 5448 19168
rect 4304 19128 5448 19156
rect 4304 19116 4310 19128
rect 5442 19116 5448 19128
rect 5500 19156 5506 19168
rect 8036 19156 8064 19196
rect 9766 19184 9772 19196
rect 9824 19184 9830 19236
rect 31496 19224 31524 19255
rect 31726 19252 31760 19264
rect 31812 19292 31818 19304
rect 32674 19292 32680 19304
rect 31812 19264 32680 19292
rect 31812 19252 31818 19264
rect 32674 19252 32680 19264
rect 32732 19252 32738 19304
rect 31726 19224 31754 19252
rect 31496 19196 31754 19224
rect 5500 19128 8064 19156
rect 5500 19116 5506 19128
rect 8202 19116 8208 19168
rect 8260 19156 8266 19168
rect 8481 19159 8539 19165
rect 8481 19156 8493 19159
rect 8260 19128 8493 19156
rect 8260 19116 8266 19128
rect 8481 19125 8493 19128
rect 8527 19125 8539 19159
rect 9122 19156 9128 19168
rect 9083 19128 9128 19156
rect 8481 19119 8539 19125
rect 9122 19116 9128 19128
rect 9180 19116 9186 19168
rect 10226 19156 10232 19168
rect 10187 19128 10232 19156
rect 10226 19116 10232 19128
rect 10284 19116 10290 19168
rect 10686 19156 10692 19168
rect 10647 19128 10692 19156
rect 10686 19116 10692 19128
rect 10744 19116 10750 19168
rect 26418 19116 26424 19168
rect 26476 19156 26482 19168
rect 27341 19159 27399 19165
rect 27341 19156 27353 19159
rect 26476 19128 27353 19156
rect 26476 19116 26482 19128
rect 27341 19125 27353 19128
rect 27387 19125 27399 19159
rect 27341 19119 27399 19125
rect 1104 19066 34868 19088
rect 1104 19014 5170 19066
rect 5222 19014 5234 19066
rect 5286 19014 5298 19066
rect 5350 19014 5362 19066
rect 5414 19014 5426 19066
rect 5478 19014 13611 19066
rect 13663 19014 13675 19066
rect 13727 19014 13739 19066
rect 13791 19014 13803 19066
rect 13855 19014 13867 19066
rect 13919 19014 22052 19066
rect 22104 19014 22116 19066
rect 22168 19014 22180 19066
rect 22232 19014 22244 19066
rect 22296 19014 22308 19066
rect 22360 19014 30493 19066
rect 30545 19014 30557 19066
rect 30609 19014 30621 19066
rect 30673 19014 30685 19066
rect 30737 19014 30749 19066
rect 30801 19014 34868 19066
rect 1104 18992 34868 19014
rect 7650 18952 7656 18964
rect 7611 18924 7656 18952
rect 7650 18912 7656 18924
rect 7708 18912 7714 18964
rect 16577 18955 16635 18961
rect 16577 18921 16589 18955
rect 16623 18952 16635 18955
rect 17310 18952 17316 18964
rect 16623 18924 17316 18952
rect 16623 18921 16635 18924
rect 16577 18915 16635 18921
rect 17310 18912 17316 18924
rect 17368 18912 17374 18964
rect 17402 18912 17408 18964
rect 17460 18952 17466 18964
rect 18601 18955 18659 18961
rect 18601 18952 18613 18955
rect 17460 18924 18613 18952
rect 17460 18912 17466 18924
rect 18601 18921 18613 18924
rect 18647 18921 18659 18955
rect 25866 18952 25872 18964
rect 25827 18924 25872 18952
rect 18601 18915 18659 18921
rect 25866 18912 25872 18924
rect 25924 18912 25930 18964
rect 28258 18952 28264 18964
rect 28219 18924 28264 18952
rect 28258 18912 28264 18924
rect 28316 18912 28322 18964
rect 33137 18955 33195 18961
rect 33137 18921 33149 18955
rect 33183 18952 33195 18955
rect 33318 18952 33324 18964
rect 33183 18924 33324 18952
rect 33183 18921 33195 18924
rect 33137 18915 33195 18921
rect 33318 18912 33324 18924
rect 33376 18912 33382 18964
rect 2958 18844 2964 18896
rect 3016 18884 3022 18896
rect 3145 18887 3203 18893
rect 3145 18884 3157 18887
rect 3016 18856 3157 18884
rect 3016 18844 3022 18856
rect 3145 18853 3157 18856
rect 3191 18853 3203 18887
rect 8478 18884 8484 18896
rect 3145 18847 3203 18853
rect 7944 18856 8484 18884
rect 7098 18776 7104 18828
rect 7156 18816 7162 18828
rect 7944 18825 7972 18856
rect 8478 18844 8484 18856
rect 8536 18844 8542 18896
rect 27798 18884 27804 18896
rect 26068 18856 27804 18884
rect 7837 18819 7895 18825
rect 7837 18816 7849 18819
rect 7156 18788 7849 18816
rect 7156 18776 7162 18788
rect 7837 18785 7849 18788
rect 7883 18785 7895 18819
rect 7837 18779 7895 18785
rect 7929 18819 7987 18825
rect 7929 18785 7941 18819
rect 7975 18785 7987 18819
rect 7929 18779 7987 18785
rect 8205 18819 8263 18825
rect 8205 18785 8217 18819
rect 8251 18816 8263 18819
rect 9122 18816 9128 18828
rect 8251 18788 9128 18816
rect 8251 18785 8263 18788
rect 8205 18779 8263 18785
rect 9122 18776 9128 18788
rect 9180 18776 9186 18828
rect 26068 18825 26096 18856
rect 27798 18844 27804 18856
rect 27856 18844 27862 18896
rect 26053 18819 26111 18825
rect 24044 18788 25084 18816
rect 3326 18748 3332 18760
rect 3287 18720 3332 18748
rect 3326 18708 3332 18720
rect 3384 18708 3390 18760
rect 3418 18708 3424 18760
rect 3476 18748 3482 18760
rect 8297 18751 8355 18757
rect 3476 18720 3521 18748
rect 3476 18708 3482 18720
rect 8297 18717 8309 18751
rect 8343 18748 8355 18751
rect 10226 18748 10232 18760
rect 8343 18720 10232 18748
rect 8343 18717 8355 18720
rect 8297 18711 8355 18717
rect 10226 18708 10232 18720
rect 10284 18708 10290 18760
rect 10413 18751 10471 18757
rect 10413 18717 10425 18751
rect 10459 18717 10471 18751
rect 10413 18711 10471 18717
rect 10505 18751 10563 18757
rect 10505 18717 10517 18751
rect 10551 18748 10563 18751
rect 10686 18748 10692 18760
rect 10551 18720 10692 18748
rect 10551 18717 10563 18720
rect 10505 18711 10563 18717
rect 3145 18683 3203 18689
rect 3145 18649 3157 18683
rect 3191 18680 3203 18683
rect 3234 18680 3240 18692
rect 3191 18652 3240 18680
rect 3191 18649 3203 18652
rect 3145 18643 3203 18649
rect 3234 18640 3240 18652
rect 3292 18680 3298 18692
rect 7190 18680 7196 18692
rect 3292 18652 7196 18680
rect 3292 18640 3298 18652
rect 7190 18640 7196 18652
rect 7248 18680 7254 18692
rect 7248 18652 8064 18680
rect 7248 18640 7254 18652
rect 8036 18621 8064 18652
rect 8202 18640 8208 18692
rect 8260 18680 8266 18692
rect 10428 18680 10456 18711
rect 10686 18708 10692 18720
rect 10744 18748 10750 18760
rect 11977 18751 12035 18757
rect 11977 18748 11989 18751
rect 10744 18720 11989 18748
rect 10744 18708 10750 18720
rect 11977 18717 11989 18720
rect 12023 18717 12035 18751
rect 11977 18711 12035 18717
rect 12253 18751 12311 18757
rect 12253 18717 12265 18751
rect 12299 18748 12311 18751
rect 12434 18748 12440 18760
rect 12299 18720 12440 18748
rect 12299 18717 12311 18720
rect 12253 18711 12311 18717
rect 12434 18708 12440 18720
rect 12492 18708 12498 18760
rect 14734 18708 14740 18760
rect 14792 18748 14798 18760
rect 15197 18751 15255 18757
rect 15197 18748 15209 18751
rect 14792 18720 15209 18748
rect 14792 18708 14798 18720
rect 15197 18717 15209 18720
rect 15243 18717 15255 18751
rect 15197 18711 15255 18717
rect 15286 18708 15292 18760
rect 15344 18748 15350 18760
rect 15453 18751 15511 18757
rect 15453 18748 15465 18751
rect 15344 18720 15465 18748
rect 15344 18708 15350 18720
rect 15453 18717 15465 18720
rect 15499 18717 15511 18751
rect 15453 18711 15511 18717
rect 18877 18751 18935 18757
rect 18877 18717 18889 18751
rect 18923 18748 18935 18751
rect 19429 18751 19487 18757
rect 19429 18748 19441 18751
rect 18923 18720 19441 18748
rect 18923 18717 18935 18720
rect 18877 18711 18935 18717
rect 19429 18717 19441 18720
rect 19475 18717 19487 18751
rect 19429 18711 19487 18717
rect 21726 18708 21732 18760
rect 21784 18748 21790 18760
rect 24044 18757 24072 18788
rect 23753 18751 23811 18757
rect 23753 18748 23765 18751
rect 21784 18720 23765 18748
rect 21784 18708 21790 18720
rect 23753 18717 23765 18720
rect 23799 18717 23811 18751
rect 23753 18711 23811 18717
rect 24029 18751 24087 18757
rect 24029 18717 24041 18751
rect 24075 18717 24087 18751
rect 24029 18711 24087 18717
rect 24486 18708 24492 18760
rect 24544 18748 24550 18760
rect 25056 18757 25084 18788
rect 26053 18785 26065 18819
rect 26099 18785 26111 18819
rect 26053 18779 26111 18785
rect 26145 18819 26203 18825
rect 26145 18785 26157 18819
rect 26191 18816 26203 18819
rect 26418 18816 26424 18828
rect 26191 18788 26424 18816
rect 26191 18785 26203 18788
rect 26145 18779 26203 18785
rect 26418 18776 26424 18788
rect 26476 18776 26482 18828
rect 28718 18816 28724 18828
rect 28679 18788 28724 18816
rect 28718 18776 28724 18788
rect 28776 18776 28782 18828
rect 28902 18816 28908 18828
rect 28863 18788 28908 18816
rect 28902 18776 28908 18788
rect 28960 18776 28966 18828
rect 29086 18776 29092 18828
rect 29144 18816 29150 18828
rect 31849 18819 31907 18825
rect 29144 18788 30052 18816
rect 29144 18776 29150 18788
rect 24765 18751 24823 18757
rect 24765 18748 24777 18751
rect 24544 18720 24777 18748
rect 24544 18708 24550 18720
rect 24765 18717 24777 18720
rect 24811 18717 24823 18751
rect 24765 18711 24823 18717
rect 25041 18751 25099 18757
rect 25041 18717 25053 18751
rect 25087 18748 25099 18751
rect 25222 18748 25228 18760
rect 25087 18720 25228 18748
rect 25087 18717 25099 18720
rect 25041 18711 25099 18717
rect 25222 18708 25228 18720
rect 25280 18748 25286 18760
rect 25498 18748 25504 18760
rect 25280 18720 25504 18748
rect 25280 18708 25286 18720
rect 25498 18708 25504 18720
rect 25556 18708 25562 18760
rect 26234 18748 26240 18760
rect 26195 18720 26240 18748
rect 26234 18708 26240 18720
rect 26292 18708 26298 18760
rect 26330 18751 26388 18757
rect 26330 18717 26342 18751
rect 26376 18717 26388 18751
rect 27338 18748 27344 18760
rect 27299 18720 27344 18748
rect 26330 18711 26388 18717
rect 8260 18652 10456 18680
rect 12345 18683 12403 18689
rect 8260 18640 8266 18652
rect 12345 18649 12357 18683
rect 12391 18680 12403 18683
rect 16206 18680 16212 18692
rect 12391 18652 16212 18680
rect 12391 18649 12403 18652
rect 12345 18643 12403 18649
rect 16206 18640 16212 18652
rect 16264 18640 16270 18692
rect 17310 18640 17316 18692
rect 17368 18680 17374 18692
rect 18417 18683 18475 18689
rect 18417 18680 18429 18683
rect 17368 18652 18429 18680
rect 17368 18640 17374 18652
rect 18417 18649 18429 18652
rect 18463 18680 18475 18683
rect 19518 18680 19524 18692
rect 18463 18652 19524 18680
rect 18463 18649 18475 18652
rect 18417 18643 18475 18649
rect 19518 18640 19524 18652
rect 19576 18680 19582 18692
rect 20898 18680 20904 18692
rect 19576 18652 20904 18680
rect 19576 18640 19582 18652
rect 20898 18640 20904 18652
rect 20956 18640 20962 18692
rect 25682 18640 25688 18692
rect 25740 18680 25746 18692
rect 26344 18680 26372 18711
rect 27338 18708 27344 18720
rect 27396 18708 27402 18760
rect 27430 18708 27436 18760
rect 27488 18748 27494 18760
rect 27525 18751 27583 18757
rect 27525 18748 27537 18751
rect 27488 18720 27537 18748
rect 27488 18708 27494 18720
rect 27525 18717 27537 18720
rect 27571 18748 27583 18751
rect 27614 18748 27620 18760
rect 27571 18720 27620 18748
rect 27571 18717 27583 18720
rect 27525 18711 27583 18717
rect 27614 18708 27620 18720
rect 27672 18708 27678 18760
rect 28629 18751 28687 18757
rect 28629 18717 28641 18751
rect 28675 18717 28687 18751
rect 28629 18711 28687 18717
rect 25740 18652 26372 18680
rect 28644 18680 28672 18711
rect 28810 18708 28816 18760
rect 28868 18748 28874 18760
rect 28997 18751 29055 18757
rect 28997 18748 29009 18751
rect 28868 18720 29009 18748
rect 28868 18708 28874 18720
rect 28997 18717 29009 18720
rect 29043 18748 29055 18751
rect 29733 18751 29791 18757
rect 29733 18748 29745 18751
rect 29043 18720 29745 18748
rect 29043 18717 29055 18720
rect 28997 18711 29055 18717
rect 29733 18717 29745 18720
rect 29779 18717 29791 18751
rect 29733 18711 29791 18717
rect 29822 18708 29828 18760
rect 29880 18748 29886 18760
rect 30024 18757 30052 18788
rect 31849 18785 31861 18819
rect 31895 18816 31907 18819
rect 32490 18816 32496 18828
rect 31895 18788 32496 18816
rect 31895 18785 31907 18788
rect 31849 18779 31907 18785
rect 32490 18776 32496 18788
rect 32548 18776 32554 18828
rect 32582 18776 32588 18828
rect 32640 18816 32646 18828
rect 32769 18819 32827 18825
rect 32769 18816 32781 18819
rect 32640 18788 32781 18816
rect 32640 18776 32646 18788
rect 32769 18785 32781 18788
rect 32815 18785 32827 18819
rect 32769 18779 32827 18785
rect 30009 18751 30067 18757
rect 29880 18720 29925 18748
rect 29880 18708 29886 18720
rect 30009 18717 30021 18751
rect 30055 18717 30067 18751
rect 30009 18711 30067 18717
rect 32033 18751 32091 18757
rect 32033 18717 32045 18751
rect 32079 18717 32091 18751
rect 32033 18711 32091 18717
rect 32217 18751 32275 18757
rect 32217 18717 32229 18751
rect 32263 18748 32275 18751
rect 32677 18751 32735 18757
rect 32677 18748 32689 18751
rect 32263 18720 32689 18748
rect 32263 18717 32275 18720
rect 32217 18711 32275 18717
rect 32677 18717 32689 18720
rect 32723 18717 32735 18751
rect 32677 18711 32735 18717
rect 29454 18680 29460 18692
rect 28644 18652 29460 18680
rect 25740 18640 25746 18652
rect 29454 18640 29460 18652
rect 29512 18640 29518 18692
rect 32048 18680 32076 18711
rect 32858 18708 32864 18760
rect 32916 18748 32922 18760
rect 32953 18751 33011 18757
rect 32953 18748 32965 18751
rect 32916 18720 32965 18748
rect 32916 18708 32922 18720
rect 32953 18717 32965 18720
rect 32999 18717 33011 18751
rect 32953 18711 33011 18717
rect 32398 18680 32404 18692
rect 32048 18652 32404 18680
rect 32398 18640 32404 18652
rect 32456 18640 32462 18692
rect 8021 18615 8079 18621
rect 8021 18581 8033 18615
rect 8067 18581 8079 18615
rect 8021 18575 8079 18581
rect 18601 18615 18659 18621
rect 18601 18581 18613 18615
rect 18647 18612 18659 18615
rect 19334 18612 19340 18624
rect 18647 18584 19340 18612
rect 18647 18581 18659 18584
rect 18601 18575 18659 18581
rect 19334 18572 19340 18584
rect 19392 18572 19398 18624
rect 20346 18572 20352 18624
rect 20404 18612 20410 18624
rect 20717 18615 20775 18621
rect 20717 18612 20729 18615
rect 20404 18584 20729 18612
rect 20404 18572 20410 18584
rect 20717 18581 20729 18584
rect 20763 18581 20775 18615
rect 20717 18575 20775 18581
rect 23474 18572 23480 18624
rect 23532 18612 23538 18624
rect 23569 18615 23627 18621
rect 23569 18612 23581 18615
rect 23532 18584 23581 18612
rect 23532 18572 23538 18584
rect 23569 18581 23581 18584
rect 23615 18581 23627 18615
rect 23569 18575 23627 18581
rect 23937 18615 23995 18621
rect 23937 18581 23949 18615
rect 23983 18612 23995 18615
rect 24210 18612 24216 18624
rect 23983 18584 24216 18612
rect 23983 18581 23995 18584
rect 23937 18575 23995 18581
rect 24210 18572 24216 18584
rect 24268 18572 24274 18624
rect 24578 18612 24584 18624
rect 24539 18584 24584 18612
rect 24578 18572 24584 18584
rect 24636 18572 24642 18624
rect 24949 18615 25007 18621
rect 24949 18581 24961 18615
rect 24995 18612 25007 18615
rect 25130 18612 25136 18624
rect 24995 18584 25136 18612
rect 24995 18581 25007 18584
rect 24949 18575 25007 18581
rect 25130 18572 25136 18584
rect 25188 18572 25194 18624
rect 26234 18572 26240 18624
rect 26292 18612 26298 18624
rect 27062 18612 27068 18624
rect 26292 18584 27068 18612
rect 26292 18572 26298 18584
rect 27062 18572 27068 18584
rect 27120 18612 27126 18624
rect 27249 18615 27307 18621
rect 27249 18612 27261 18615
rect 27120 18584 27261 18612
rect 27120 18572 27126 18584
rect 27249 18581 27261 18584
rect 27295 18581 27307 18615
rect 27249 18575 27307 18581
rect 1104 18522 35027 18544
rect 1104 18470 9390 18522
rect 9442 18470 9454 18522
rect 9506 18470 9518 18522
rect 9570 18470 9582 18522
rect 9634 18470 9646 18522
rect 9698 18470 17831 18522
rect 17883 18470 17895 18522
rect 17947 18470 17959 18522
rect 18011 18470 18023 18522
rect 18075 18470 18087 18522
rect 18139 18470 26272 18522
rect 26324 18470 26336 18522
rect 26388 18470 26400 18522
rect 26452 18470 26464 18522
rect 26516 18470 26528 18522
rect 26580 18470 34713 18522
rect 34765 18470 34777 18522
rect 34829 18470 34841 18522
rect 34893 18470 34905 18522
rect 34957 18470 34969 18522
rect 35021 18470 35027 18522
rect 1104 18448 35027 18470
rect 8205 18411 8263 18417
rect 8205 18377 8217 18411
rect 8251 18408 8263 18411
rect 8938 18408 8944 18420
rect 8251 18380 8944 18408
rect 8251 18377 8263 18380
rect 8205 18371 8263 18377
rect 8938 18368 8944 18380
rect 8996 18368 9002 18420
rect 17129 18411 17187 18417
rect 17129 18377 17141 18411
rect 17175 18408 17187 18411
rect 17678 18408 17684 18420
rect 17175 18380 17684 18408
rect 17175 18377 17187 18380
rect 17129 18371 17187 18377
rect 17678 18368 17684 18380
rect 17736 18368 17742 18420
rect 19794 18368 19800 18420
rect 19852 18408 19858 18420
rect 20073 18411 20131 18417
rect 20073 18408 20085 18411
rect 19852 18380 20085 18408
rect 19852 18368 19858 18380
rect 20073 18377 20085 18380
rect 20119 18377 20131 18411
rect 20073 18371 20131 18377
rect 20901 18411 20959 18417
rect 20901 18377 20913 18411
rect 20947 18408 20959 18411
rect 21082 18408 21088 18420
rect 20947 18380 21088 18408
rect 20947 18377 20959 18380
rect 20901 18371 20959 18377
rect 21082 18368 21088 18380
rect 21140 18368 21146 18420
rect 24486 18408 24492 18420
rect 22066 18380 24492 18408
rect 6825 18343 6883 18349
rect 6825 18309 6837 18343
rect 6871 18340 6883 18343
rect 7190 18340 7196 18352
rect 6871 18312 7196 18340
rect 6871 18309 6883 18312
rect 6825 18303 6883 18309
rect 7190 18300 7196 18312
rect 7248 18300 7254 18352
rect 11974 18300 11980 18352
rect 12032 18340 12038 18352
rect 14734 18340 14740 18352
rect 12032 18312 12480 18340
rect 14695 18312 14740 18340
rect 12032 18300 12038 18312
rect 6638 18232 6644 18284
rect 6696 18272 6702 18284
rect 8021 18275 8079 18281
rect 8021 18272 8033 18275
rect 6696 18244 8033 18272
rect 6696 18232 6702 18244
rect 8021 18241 8033 18244
rect 8067 18241 8079 18275
rect 8202 18272 8208 18284
rect 8163 18244 8208 18272
rect 8021 18235 8079 18241
rect 8202 18232 8208 18244
rect 8260 18232 8266 18284
rect 10321 18275 10379 18281
rect 10321 18241 10333 18275
rect 10367 18272 10379 18275
rect 11054 18272 11060 18284
rect 10367 18244 11060 18272
rect 10367 18241 10379 18244
rect 10321 18235 10379 18241
rect 11054 18232 11060 18244
rect 11112 18232 11118 18284
rect 11790 18232 11796 18284
rect 11848 18272 11854 18284
rect 12342 18272 12348 18284
rect 11848 18244 12348 18272
rect 11848 18232 11854 18244
rect 12342 18232 12348 18244
rect 12400 18232 12406 18284
rect 12452 18281 12480 18312
rect 14734 18300 14740 18312
rect 14792 18300 14798 18352
rect 15286 18300 15292 18352
rect 15344 18340 15350 18352
rect 16209 18343 16267 18349
rect 15344 18312 16160 18340
rect 15344 18300 15350 18312
rect 12437 18275 12495 18281
rect 12437 18241 12449 18275
rect 12483 18241 12495 18275
rect 12986 18272 12992 18284
rect 12947 18244 12992 18272
rect 12437 18235 12495 18241
rect 12986 18232 12992 18244
rect 13044 18232 13050 18284
rect 16025 18275 16083 18281
rect 16025 18241 16037 18275
rect 16071 18241 16083 18275
rect 16132 18272 16160 18312
rect 16209 18309 16221 18343
rect 16255 18340 16267 18343
rect 16666 18340 16672 18352
rect 16255 18312 16672 18340
rect 16255 18309 16267 18312
rect 16209 18303 16267 18309
rect 16666 18300 16672 18312
rect 16724 18300 16730 18352
rect 17310 18340 17316 18352
rect 17271 18312 17316 18340
rect 17310 18300 17316 18312
rect 17368 18300 17374 18352
rect 18966 18349 18972 18352
rect 18960 18340 18972 18349
rect 18927 18312 18972 18340
rect 18960 18303 18972 18312
rect 18966 18300 18972 18303
rect 19024 18300 19030 18352
rect 22066 18340 22094 18380
rect 24486 18368 24492 18380
rect 24544 18368 24550 18420
rect 25682 18408 25688 18420
rect 25643 18380 25688 18408
rect 25682 18368 25688 18380
rect 25740 18368 25746 18420
rect 27614 18368 27620 18420
rect 27672 18408 27678 18420
rect 28813 18411 28871 18417
rect 28813 18408 28825 18411
rect 27672 18380 28825 18408
rect 27672 18368 27678 18380
rect 28813 18377 28825 18380
rect 28859 18377 28871 18411
rect 28813 18371 28871 18377
rect 32769 18411 32827 18417
rect 32769 18377 32781 18411
rect 32815 18408 32827 18411
rect 32858 18408 32864 18420
rect 32815 18380 32864 18408
rect 32815 18377 32827 18380
rect 32769 18371 32827 18377
rect 32858 18368 32864 18380
rect 32916 18368 32922 18420
rect 20732 18312 22094 18340
rect 16301 18275 16359 18281
rect 16301 18272 16313 18275
rect 16132 18244 16313 18272
rect 16025 18235 16083 18241
rect 16301 18241 16313 18244
rect 16347 18241 16359 18275
rect 18690 18272 18696 18284
rect 18651 18244 18696 18272
rect 16301 18235 16359 18241
rect 6730 18204 6736 18216
rect 6691 18176 6736 18204
rect 6730 18164 6736 18176
rect 6788 18164 6794 18216
rect 6914 18204 6920 18216
rect 6875 18176 6920 18204
rect 6914 18164 6920 18176
rect 6972 18164 6978 18216
rect 12158 18204 12164 18216
rect 12119 18176 12164 18204
rect 12158 18164 12164 18176
rect 12216 18164 12222 18216
rect 7282 18136 7288 18148
rect 7243 18108 7288 18136
rect 7282 18096 7288 18108
rect 7340 18096 7346 18148
rect 16040 18136 16068 18235
rect 18690 18232 18696 18244
rect 18748 18232 18754 18284
rect 20732 18281 20760 18312
rect 24210 18300 24216 18352
rect 24268 18340 24274 18352
rect 24857 18343 24915 18349
rect 24857 18340 24869 18343
rect 24268 18312 24869 18340
rect 24268 18300 24274 18312
rect 24857 18309 24869 18312
rect 24903 18340 24915 18343
rect 29086 18340 29092 18352
rect 24903 18312 29092 18340
rect 24903 18309 24915 18312
rect 24857 18303 24915 18309
rect 29086 18300 29092 18312
rect 29144 18300 29150 18352
rect 20717 18275 20775 18281
rect 20717 18241 20729 18275
rect 20763 18241 20775 18275
rect 20717 18235 20775 18241
rect 20898 18232 20904 18284
rect 20956 18272 20962 18284
rect 20993 18275 21051 18281
rect 20993 18272 21005 18275
rect 20956 18244 21005 18272
rect 20956 18232 20962 18244
rect 20993 18241 21005 18244
rect 21039 18241 21051 18275
rect 23474 18272 23480 18284
rect 23435 18244 23480 18272
rect 20993 18235 21051 18241
rect 23474 18232 23480 18244
rect 23532 18232 23538 18284
rect 25314 18272 25320 18284
rect 25275 18244 25320 18272
rect 25314 18232 25320 18244
rect 25372 18232 25378 18284
rect 28166 18272 28172 18284
rect 28127 18244 28172 18272
rect 28166 18232 28172 18244
rect 28224 18232 28230 18284
rect 28534 18232 28540 18284
rect 28592 18272 28598 18284
rect 28810 18272 28816 18284
rect 28592 18244 28816 18272
rect 28592 18232 28598 18244
rect 28810 18232 28816 18244
rect 28868 18272 28874 18284
rect 28997 18275 29055 18281
rect 28997 18272 29009 18275
rect 28868 18244 29009 18272
rect 28868 18232 28874 18244
rect 28997 18241 29009 18244
rect 29043 18241 29055 18275
rect 29178 18272 29184 18284
rect 29139 18244 29184 18272
rect 28997 18235 29055 18241
rect 29178 18232 29184 18244
rect 29236 18232 29242 18284
rect 29270 18232 29276 18284
rect 29328 18272 29334 18284
rect 32490 18272 32496 18284
rect 29328 18244 29373 18272
rect 32451 18244 32496 18272
rect 29328 18232 29334 18244
rect 32490 18232 32496 18244
rect 32548 18232 32554 18284
rect 23106 18164 23112 18216
rect 23164 18204 23170 18216
rect 23201 18207 23259 18213
rect 23201 18204 23213 18207
rect 23164 18176 23213 18204
rect 23164 18164 23170 18176
rect 23201 18173 23213 18176
rect 23247 18173 23259 18207
rect 25406 18204 25412 18216
rect 25367 18176 25412 18204
rect 23201 18167 23259 18173
rect 25406 18164 25412 18176
rect 25464 18164 25470 18216
rect 27338 18164 27344 18216
rect 27396 18204 27402 18216
rect 27801 18207 27859 18213
rect 27801 18204 27813 18207
rect 27396 18176 27813 18204
rect 27396 18164 27402 18176
rect 27801 18173 27813 18176
rect 27847 18173 27859 18207
rect 27801 18167 27859 18173
rect 28261 18207 28319 18213
rect 28261 18173 28273 18207
rect 28307 18204 28319 18207
rect 29454 18204 29460 18216
rect 28307 18176 29460 18204
rect 28307 18173 28319 18176
rect 28261 18167 28319 18173
rect 29454 18164 29460 18176
rect 29512 18164 29518 18216
rect 32306 18204 32312 18216
rect 32267 18176 32312 18204
rect 32306 18164 32312 18176
rect 32364 18164 32370 18216
rect 32858 18204 32864 18216
rect 32819 18176 32864 18204
rect 32858 18164 32864 18176
rect 32916 18164 32922 18216
rect 34330 18204 34336 18216
rect 34291 18176 34336 18204
rect 34330 18164 34336 18176
rect 34388 18164 34394 18216
rect 17310 18136 17316 18148
rect 16040 18108 17316 18136
rect 17310 18096 17316 18108
rect 17368 18096 17374 18148
rect 10226 18068 10232 18080
rect 10187 18040 10232 18068
rect 10226 18028 10232 18040
rect 10284 18028 10290 18080
rect 15838 18068 15844 18080
rect 15799 18040 15844 18068
rect 15838 18028 15844 18040
rect 15896 18028 15902 18080
rect 16942 18068 16948 18080
rect 16903 18040 16948 18068
rect 16942 18028 16948 18040
rect 17000 18028 17006 18080
rect 17129 18071 17187 18077
rect 17129 18037 17141 18071
rect 17175 18068 17187 18071
rect 17402 18068 17408 18080
rect 17175 18040 17408 18068
rect 17175 18037 17187 18040
rect 17129 18031 17187 18037
rect 17402 18028 17408 18040
rect 17460 18028 17466 18080
rect 20530 18068 20536 18080
rect 20491 18040 20536 18068
rect 20530 18028 20536 18040
rect 20588 18028 20594 18080
rect 24946 18028 24952 18080
rect 25004 18068 25010 18080
rect 25317 18071 25375 18077
rect 25317 18068 25329 18071
rect 25004 18040 25329 18068
rect 25004 18028 25010 18040
rect 25317 18037 25329 18040
rect 25363 18037 25375 18071
rect 25317 18031 25375 18037
rect 1104 17978 34868 18000
rect 1104 17926 5170 17978
rect 5222 17926 5234 17978
rect 5286 17926 5298 17978
rect 5350 17926 5362 17978
rect 5414 17926 5426 17978
rect 5478 17926 13611 17978
rect 13663 17926 13675 17978
rect 13727 17926 13739 17978
rect 13791 17926 13803 17978
rect 13855 17926 13867 17978
rect 13919 17926 22052 17978
rect 22104 17926 22116 17978
rect 22168 17926 22180 17978
rect 22232 17926 22244 17978
rect 22296 17926 22308 17978
rect 22360 17926 30493 17978
rect 30545 17926 30557 17978
rect 30609 17926 30621 17978
rect 30673 17926 30685 17978
rect 30737 17926 30749 17978
rect 30801 17926 34868 17978
rect 1104 17904 34868 17926
rect 6457 17867 6515 17873
rect 6457 17833 6469 17867
rect 6503 17864 6515 17867
rect 6730 17864 6736 17876
rect 6503 17836 6736 17864
rect 6503 17833 6515 17836
rect 6457 17827 6515 17833
rect 6730 17824 6736 17836
rect 6788 17824 6794 17876
rect 27982 17864 27988 17876
rect 27943 17836 27988 17864
rect 27982 17824 27988 17836
rect 28040 17824 28046 17876
rect 29270 17824 29276 17876
rect 29328 17864 29334 17876
rect 30745 17867 30803 17873
rect 30745 17864 30757 17867
rect 29328 17836 30757 17864
rect 29328 17824 29334 17836
rect 30745 17833 30757 17836
rect 30791 17833 30803 17867
rect 32677 17867 32735 17873
rect 32677 17864 32689 17867
rect 30745 17827 30803 17833
rect 30852 17836 32689 17864
rect 3421 17799 3479 17805
rect 3421 17765 3433 17799
rect 3467 17796 3479 17799
rect 3510 17796 3516 17808
rect 3467 17768 3516 17796
rect 3467 17765 3479 17768
rect 3421 17759 3479 17765
rect 3510 17756 3516 17768
rect 3568 17756 3574 17808
rect 28537 17799 28595 17805
rect 28537 17796 28549 17799
rect 27816 17768 28549 17796
rect 11330 17688 11336 17740
rect 11388 17728 11394 17740
rect 12066 17728 12072 17740
rect 11388 17700 12072 17728
rect 11388 17688 11394 17700
rect 12066 17688 12072 17700
rect 12124 17728 12130 17740
rect 27614 17728 27620 17740
rect 12124 17700 13124 17728
rect 27575 17700 27620 17728
rect 12124 17688 12130 17700
rect 3234 17660 3240 17672
rect 3195 17632 3240 17660
rect 3234 17620 3240 17632
rect 3292 17620 3298 17672
rect 6362 17660 6368 17672
rect 6323 17632 6368 17660
rect 6362 17620 6368 17632
rect 6420 17620 6426 17672
rect 6546 17660 6552 17672
rect 6507 17632 6552 17660
rect 6546 17620 6552 17632
rect 6604 17620 6610 17672
rect 13096 17669 13124 17700
rect 27614 17688 27620 17700
rect 27672 17688 27678 17740
rect 27816 17737 27844 17768
rect 28537 17765 28549 17768
rect 28583 17765 28595 17799
rect 28537 17759 28595 17765
rect 29454 17756 29460 17808
rect 29512 17796 29518 17808
rect 30852 17796 30880 17836
rect 32677 17833 32689 17836
rect 32723 17833 32735 17867
rect 32677 17827 32735 17833
rect 32306 17796 32312 17808
rect 29512 17768 30880 17796
rect 31772 17768 32312 17796
rect 29512 17756 29518 17768
rect 27801 17731 27859 17737
rect 27801 17697 27813 17731
rect 27847 17697 27859 17731
rect 27801 17691 27859 17697
rect 13081 17663 13139 17669
rect 13081 17629 13093 17663
rect 13127 17660 13139 17663
rect 13538 17660 13544 17672
rect 13127 17632 13544 17660
rect 13127 17629 13139 17632
rect 13081 17623 13139 17629
rect 13538 17620 13544 17632
rect 13596 17620 13602 17672
rect 16942 17660 16948 17672
rect 16903 17632 16948 17660
rect 16942 17620 16948 17632
rect 17000 17620 17006 17672
rect 18690 17620 18696 17672
rect 18748 17660 18754 17672
rect 19429 17663 19487 17669
rect 19429 17660 19441 17663
rect 18748 17632 19441 17660
rect 18748 17620 18754 17632
rect 19429 17629 19441 17632
rect 19475 17629 19487 17663
rect 19429 17623 19487 17629
rect 19696 17663 19754 17669
rect 19696 17629 19708 17663
rect 19742 17660 19754 17663
rect 20530 17660 20536 17672
rect 19742 17632 20536 17660
rect 19742 17629 19754 17632
rect 19696 17623 19754 17629
rect 20530 17620 20536 17632
rect 20588 17620 20594 17672
rect 25222 17660 25228 17672
rect 25135 17632 25228 17660
rect 25222 17620 25228 17632
rect 25280 17620 25286 17672
rect 25682 17620 25688 17672
rect 25740 17660 25746 17672
rect 27525 17663 27583 17669
rect 27525 17660 27537 17663
rect 25740 17632 27537 17660
rect 25740 17620 25746 17632
rect 27525 17629 27537 17632
rect 27571 17629 27583 17663
rect 27525 17623 27583 17629
rect 27709 17663 27767 17669
rect 27709 17629 27721 17663
rect 27755 17660 27767 17663
rect 28534 17660 28540 17672
rect 27755 17632 27844 17660
rect 28495 17632 28540 17660
rect 27755 17629 27767 17632
rect 27709 17623 27767 17629
rect 2682 17552 2688 17604
rect 2740 17592 2746 17604
rect 2869 17595 2927 17601
rect 2869 17592 2881 17595
rect 2740 17564 2881 17592
rect 2740 17552 2746 17564
rect 2869 17561 2881 17564
rect 2915 17561 2927 17595
rect 2869 17555 2927 17561
rect 12158 17552 12164 17604
rect 12216 17552 12222 17604
rect 12805 17595 12863 17601
rect 12805 17561 12817 17595
rect 12851 17592 12863 17595
rect 12894 17592 12900 17604
rect 12851 17564 12900 17592
rect 12851 17561 12863 17564
rect 12805 17555 12863 17561
rect 12894 17552 12900 17564
rect 12952 17552 12958 17604
rect 15197 17595 15255 17601
rect 15197 17561 15209 17595
rect 15243 17561 15255 17595
rect 15197 17555 15255 17561
rect 3050 17524 3056 17536
rect 3011 17496 3056 17524
rect 3050 17484 3056 17496
rect 3108 17484 3114 17536
rect 3142 17484 3148 17536
rect 3200 17524 3206 17536
rect 3200 17496 3245 17524
rect 3200 17484 3206 17496
rect 10962 17484 10968 17536
rect 11020 17524 11026 17536
rect 11333 17527 11391 17533
rect 11333 17524 11345 17527
rect 11020 17496 11345 17524
rect 11020 17484 11026 17496
rect 11333 17493 11345 17496
rect 11379 17493 11391 17527
rect 11333 17487 11391 17493
rect 12986 17484 12992 17536
rect 13044 17524 13050 17536
rect 15212 17524 15240 17555
rect 24486 17552 24492 17604
rect 24544 17592 24550 17604
rect 24949 17595 25007 17601
rect 24949 17592 24961 17595
rect 24544 17564 24961 17592
rect 24544 17552 24550 17564
rect 24949 17561 24961 17564
rect 24995 17561 25007 17595
rect 25240 17592 25268 17620
rect 27816 17604 27844 17632
rect 28534 17620 28540 17632
rect 28592 17620 28598 17672
rect 28813 17663 28871 17669
rect 28813 17629 28825 17663
rect 28859 17660 28871 17663
rect 29270 17660 29276 17672
rect 28859 17632 29276 17660
rect 28859 17629 28871 17632
rect 28813 17623 28871 17629
rect 29270 17620 29276 17632
rect 29328 17620 29334 17672
rect 30926 17660 30932 17672
rect 30839 17632 30932 17660
rect 30926 17620 30932 17632
rect 30984 17660 30990 17672
rect 31772 17669 31800 17768
rect 32306 17756 32312 17768
rect 32364 17796 32370 17808
rect 32364 17768 33640 17796
rect 32364 17756 32370 17768
rect 33612 17737 33640 17768
rect 33597 17731 33655 17737
rect 31956 17700 33456 17728
rect 31956 17669 31984 17700
rect 33428 17672 33456 17700
rect 33597 17697 33609 17731
rect 33643 17697 33655 17731
rect 33597 17691 33655 17697
rect 31757 17663 31815 17669
rect 31757 17660 31769 17663
rect 30984 17632 31769 17660
rect 30984 17620 30990 17632
rect 31757 17629 31769 17632
rect 31803 17629 31815 17663
rect 31757 17623 31815 17629
rect 31941 17663 31999 17669
rect 31941 17629 31953 17663
rect 31987 17629 31999 17663
rect 32582 17660 32588 17672
rect 32543 17632 32588 17660
rect 31941 17623 31999 17629
rect 32582 17620 32588 17632
rect 32640 17660 32646 17672
rect 33229 17663 33287 17669
rect 33229 17660 33241 17663
rect 32640 17632 33241 17660
rect 32640 17620 32646 17632
rect 33229 17629 33241 17632
rect 33275 17629 33287 17663
rect 33229 17623 33287 17629
rect 33410 17620 33416 17672
rect 33468 17660 33474 17672
rect 33468 17632 33561 17660
rect 33468 17620 33474 17632
rect 26142 17592 26148 17604
rect 25240 17564 26148 17592
rect 24949 17555 25007 17561
rect 26142 17552 26148 17564
rect 26200 17552 26206 17604
rect 27798 17552 27804 17604
rect 27856 17552 27862 17604
rect 28629 17595 28687 17601
rect 28629 17561 28641 17595
rect 28675 17592 28687 17595
rect 29178 17592 29184 17604
rect 28675 17564 29184 17592
rect 28675 17561 28687 17564
rect 28629 17555 28687 17561
rect 29178 17552 29184 17564
rect 29236 17592 29242 17604
rect 29822 17592 29828 17604
rect 29236 17564 29828 17592
rect 29236 17552 29242 17564
rect 29822 17552 29828 17564
rect 29880 17552 29886 17604
rect 31110 17592 31116 17604
rect 31071 17564 31116 17592
rect 31110 17552 31116 17564
rect 31168 17552 31174 17604
rect 31849 17595 31907 17601
rect 31849 17561 31861 17595
rect 31895 17592 31907 17595
rect 32401 17595 32459 17601
rect 32401 17592 32413 17595
rect 31895 17564 32413 17592
rect 31895 17561 31907 17564
rect 31849 17555 31907 17561
rect 32401 17561 32413 17564
rect 32447 17561 32459 17595
rect 32401 17555 32459 17561
rect 13044 17496 15240 17524
rect 20809 17527 20867 17533
rect 13044 17484 13050 17496
rect 20809 17493 20821 17527
rect 20855 17524 20867 17527
rect 21082 17524 21088 17536
rect 20855 17496 21088 17524
rect 20855 17493 20867 17496
rect 20809 17487 20867 17493
rect 21082 17484 21088 17496
rect 21140 17484 21146 17536
rect 1104 17434 35027 17456
rect 1104 17382 9390 17434
rect 9442 17382 9454 17434
rect 9506 17382 9518 17434
rect 9570 17382 9582 17434
rect 9634 17382 9646 17434
rect 9698 17382 17831 17434
rect 17883 17382 17895 17434
rect 17947 17382 17959 17434
rect 18011 17382 18023 17434
rect 18075 17382 18087 17434
rect 18139 17382 26272 17434
rect 26324 17382 26336 17434
rect 26388 17382 26400 17434
rect 26452 17382 26464 17434
rect 26516 17382 26528 17434
rect 26580 17382 34713 17434
rect 34765 17382 34777 17434
rect 34829 17382 34841 17434
rect 34893 17382 34905 17434
rect 34957 17382 34969 17434
rect 35021 17382 35027 17434
rect 1104 17360 35027 17382
rect 4433 17323 4491 17329
rect 4433 17289 4445 17323
rect 4479 17320 4491 17323
rect 6914 17320 6920 17332
rect 4479 17292 6920 17320
rect 4479 17289 4491 17292
rect 4433 17283 4491 17289
rect 6914 17280 6920 17292
rect 6972 17280 6978 17332
rect 10318 17320 10324 17332
rect 9600 17292 10324 17320
rect 2958 17252 2964 17264
rect 2919 17224 2964 17252
rect 2958 17212 2964 17224
rect 3016 17212 3022 17264
rect 6932 17252 6960 17280
rect 6932 17224 8248 17252
rect 4246 17184 4252 17196
rect 4094 17156 4252 17184
rect 4246 17144 4252 17156
rect 4304 17144 4310 17196
rect 6730 17184 6736 17196
rect 6691 17156 6736 17184
rect 6730 17144 6736 17156
rect 6788 17144 6794 17196
rect 6822 17144 6828 17196
rect 6880 17184 6886 17196
rect 7101 17187 7159 17193
rect 7101 17184 7113 17187
rect 6880 17156 7113 17184
rect 6880 17144 6886 17156
rect 7101 17153 7113 17156
rect 7147 17153 7159 17187
rect 7101 17147 7159 17153
rect 7466 17144 7472 17196
rect 7524 17184 7530 17196
rect 7561 17187 7619 17193
rect 7561 17184 7573 17187
rect 7524 17156 7573 17184
rect 7524 17144 7530 17156
rect 7561 17153 7573 17156
rect 7607 17153 7619 17187
rect 7561 17147 7619 17153
rect 7742 17144 7748 17196
rect 7800 17184 7806 17196
rect 8220 17193 8248 17224
rect 8846 17212 8852 17264
rect 8904 17252 8910 17264
rect 9600 17261 9628 17292
rect 10318 17280 10324 17292
rect 10376 17320 10382 17332
rect 14458 17320 14464 17332
rect 10376 17292 14464 17320
rect 10376 17280 10382 17292
rect 14458 17280 14464 17292
rect 14516 17280 14522 17332
rect 24489 17323 24547 17329
rect 24489 17289 24501 17323
rect 24535 17320 24547 17323
rect 25130 17320 25136 17332
rect 24535 17292 25136 17320
rect 24535 17289 24547 17292
rect 24489 17283 24547 17289
rect 25130 17280 25136 17292
rect 25188 17280 25194 17332
rect 25682 17320 25688 17332
rect 25643 17292 25688 17320
rect 25682 17280 25688 17292
rect 25740 17280 25746 17332
rect 29822 17320 29828 17332
rect 29783 17292 29828 17320
rect 29822 17280 29828 17292
rect 29880 17280 29886 17332
rect 30006 17280 30012 17332
rect 30064 17320 30070 17332
rect 30745 17323 30803 17329
rect 30745 17320 30757 17323
rect 30064 17292 30757 17320
rect 30064 17280 30070 17292
rect 30745 17289 30757 17292
rect 30791 17289 30803 17323
rect 30926 17320 30932 17332
rect 30887 17292 30932 17320
rect 30745 17283 30803 17289
rect 30926 17280 30932 17292
rect 30984 17280 30990 17332
rect 31662 17320 31668 17332
rect 31496 17292 31668 17320
rect 9585 17255 9643 17261
rect 9585 17252 9597 17255
rect 8904 17224 9597 17252
rect 8904 17212 8910 17224
rect 9585 17221 9597 17224
rect 9631 17221 9643 17255
rect 9585 17215 9643 17221
rect 12250 17212 12256 17264
rect 12308 17212 12314 17264
rect 13265 17255 13323 17261
rect 13265 17221 13277 17255
rect 13311 17252 13323 17255
rect 13354 17252 13360 17264
rect 13311 17224 13360 17252
rect 13311 17221 13323 17224
rect 13265 17215 13323 17221
rect 13354 17212 13360 17224
rect 13412 17212 13418 17264
rect 20809 17255 20867 17261
rect 20809 17252 20821 17255
rect 16224 17224 20821 17252
rect 16224 17196 16252 17224
rect 20809 17221 20821 17224
rect 20855 17221 20867 17255
rect 20809 17215 20867 17221
rect 21177 17255 21235 17261
rect 21177 17221 21189 17255
rect 21223 17252 21235 17255
rect 21726 17252 21732 17264
rect 21223 17224 21732 17252
rect 21223 17221 21235 17224
rect 21177 17215 21235 17221
rect 8021 17187 8079 17193
rect 8021 17184 8033 17187
rect 7800 17156 8033 17184
rect 7800 17144 7806 17156
rect 8021 17153 8033 17156
rect 8067 17153 8079 17187
rect 8021 17147 8079 17153
rect 8205 17187 8263 17193
rect 8205 17153 8217 17187
rect 8251 17153 8263 17187
rect 9858 17184 9864 17196
rect 9819 17156 9864 17184
rect 8205 17147 8263 17153
rect 9858 17144 9864 17156
rect 9916 17144 9922 17196
rect 13538 17144 13544 17196
rect 13596 17184 13602 17196
rect 16206 17184 16212 17196
rect 13596 17156 13641 17184
rect 16167 17156 16212 17184
rect 13596 17144 13602 17156
rect 16206 17144 16212 17156
rect 16264 17144 16270 17196
rect 19144 17187 19202 17193
rect 19144 17153 19156 17187
rect 19190 17184 19202 17187
rect 19426 17184 19432 17196
rect 19190 17156 19432 17184
rect 19190 17153 19202 17156
rect 19144 17147 19202 17153
rect 19426 17144 19432 17156
rect 19484 17144 19490 17196
rect 20714 17144 20720 17196
rect 20772 17184 20778 17196
rect 21192 17184 21220 17215
rect 21726 17212 21732 17224
rect 21784 17212 21790 17264
rect 23376 17255 23434 17261
rect 23376 17221 23388 17255
rect 23422 17252 23434 17255
rect 24578 17252 24584 17264
rect 23422 17224 24584 17252
rect 23422 17221 23434 17224
rect 23376 17215 23434 17221
rect 24578 17212 24584 17224
rect 24636 17212 24642 17264
rect 25317 17255 25375 17261
rect 25317 17252 25329 17255
rect 24688 17224 25329 17252
rect 20772 17156 21220 17184
rect 20772 17144 20778 17156
rect 23750 17144 23756 17196
rect 23808 17184 23814 17196
rect 24688 17184 24716 17224
rect 25317 17221 25329 17224
rect 25363 17221 25375 17255
rect 25317 17215 25375 17221
rect 25409 17255 25467 17261
rect 25409 17221 25421 17255
rect 25455 17252 25467 17255
rect 25958 17252 25964 17264
rect 25455 17224 25964 17252
rect 25455 17221 25467 17224
rect 25409 17215 25467 17221
rect 25958 17212 25964 17224
rect 26016 17212 26022 17264
rect 31496 17261 31524 17292
rect 31662 17280 31668 17292
rect 31720 17320 31726 17332
rect 32509 17323 32567 17329
rect 32509 17320 32521 17323
rect 31720 17292 32521 17320
rect 31720 17280 31726 17292
rect 32509 17289 32521 17292
rect 32555 17289 32567 17323
rect 32509 17283 32567 17289
rect 32677 17323 32735 17329
rect 32677 17289 32689 17323
rect 32723 17320 32735 17323
rect 32858 17320 32864 17332
rect 32723 17292 32864 17320
rect 32723 17289 32735 17292
rect 32677 17283 32735 17289
rect 32858 17280 32864 17292
rect 32916 17280 32922 17332
rect 33229 17323 33287 17329
rect 33229 17289 33241 17323
rect 33275 17320 33287 17323
rect 33410 17320 33416 17332
rect 33275 17292 33416 17320
rect 33275 17289 33287 17292
rect 33229 17283 33287 17289
rect 33410 17280 33416 17292
rect 33468 17280 33474 17332
rect 30837 17255 30895 17261
rect 30837 17252 30849 17255
rect 29932 17224 30849 17252
rect 25038 17184 25044 17196
rect 23808 17156 24716 17184
rect 24999 17156 25044 17184
rect 23808 17144 23814 17156
rect 25038 17144 25044 17156
rect 25096 17144 25102 17196
rect 25134 17187 25192 17193
rect 25134 17153 25146 17187
rect 25180 17153 25192 17187
rect 25134 17147 25192 17153
rect 2682 17116 2688 17128
rect 2643 17088 2688 17116
rect 2682 17076 2688 17088
rect 2740 17076 2746 17128
rect 6638 17116 6644 17128
rect 6599 17088 6644 17116
rect 6638 17076 6644 17088
rect 6696 17076 6702 17128
rect 9766 17116 9772 17128
rect 9727 17088 9772 17116
rect 9766 17076 9772 17088
rect 9824 17076 9830 17128
rect 15933 17119 15991 17125
rect 15933 17085 15945 17119
rect 15979 17116 15991 17119
rect 16298 17116 16304 17128
rect 15979 17088 16304 17116
rect 15979 17085 15991 17088
rect 15933 17079 15991 17085
rect 16298 17076 16304 17088
rect 16356 17076 16362 17128
rect 18690 17076 18696 17128
rect 18748 17116 18754 17128
rect 18877 17119 18935 17125
rect 18877 17116 18889 17119
rect 18748 17088 18889 17116
rect 18748 17076 18754 17088
rect 18877 17085 18889 17088
rect 18923 17085 18935 17119
rect 18877 17079 18935 17085
rect 22554 17076 22560 17128
rect 22612 17116 22618 17128
rect 23106 17116 23112 17128
rect 22612 17088 23112 17116
rect 22612 17076 22618 17088
rect 23106 17076 23112 17088
rect 23164 17076 23170 17128
rect 25148 17048 25176 17147
rect 25498 17144 25504 17196
rect 25556 17193 25562 17196
rect 29932 17193 29960 17224
rect 30837 17221 30849 17224
rect 30883 17252 30895 17255
rect 31481 17255 31539 17261
rect 31481 17252 31493 17255
rect 30883 17224 31493 17252
rect 30883 17221 30895 17224
rect 30837 17215 30895 17221
rect 31481 17221 31493 17224
rect 31527 17221 31539 17255
rect 32309 17255 32367 17261
rect 32309 17252 32321 17255
rect 31481 17215 31539 17221
rect 31680 17224 32321 17252
rect 25556 17184 25564 17193
rect 29733 17187 29791 17193
rect 25556 17156 25601 17184
rect 25556 17147 25564 17156
rect 29733 17153 29745 17187
rect 29779 17153 29791 17187
rect 29733 17147 29791 17153
rect 29917 17187 29975 17193
rect 29917 17153 29929 17187
rect 29963 17153 29975 17187
rect 29917 17147 29975 17153
rect 30469 17187 30527 17193
rect 30469 17153 30481 17187
rect 30515 17153 30527 17187
rect 30469 17147 30527 17153
rect 30613 17187 30671 17193
rect 30613 17153 30625 17187
rect 30659 17184 30671 17187
rect 31294 17184 31300 17196
rect 30659 17156 31300 17184
rect 30659 17153 30671 17156
rect 30613 17147 30671 17153
rect 25556 17144 25562 17147
rect 29748 17116 29776 17147
rect 30282 17116 30288 17128
rect 29748 17088 30288 17116
rect 30282 17076 30288 17088
rect 30340 17116 30346 17128
rect 30484 17116 30512 17147
rect 31294 17144 31300 17156
rect 31352 17144 31358 17196
rect 31680 17193 31708 17224
rect 32309 17221 32321 17224
rect 32355 17221 32367 17255
rect 32309 17215 32367 17221
rect 31665 17187 31723 17193
rect 31665 17184 31677 17187
rect 31404 17156 31677 17184
rect 30340 17088 30512 17116
rect 30340 17076 30346 17088
rect 24044 17020 25176 17048
rect 8202 16980 8208 16992
rect 8163 16952 8208 16980
rect 8202 16940 8208 16952
rect 8260 16940 8266 16992
rect 8294 16940 8300 16992
rect 8352 16980 8358 16992
rect 9677 16983 9735 16989
rect 9677 16980 9689 16983
rect 8352 16952 9689 16980
rect 8352 16940 8358 16952
rect 9677 16949 9689 16952
rect 9723 16949 9735 16983
rect 10042 16980 10048 16992
rect 10003 16952 10048 16980
rect 9677 16943 9735 16949
rect 10042 16940 10048 16952
rect 10100 16940 10106 16992
rect 11146 16940 11152 16992
rect 11204 16980 11210 16992
rect 11793 16983 11851 16989
rect 11793 16980 11805 16983
rect 11204 16952 11805 16980
rect 11204 16940 11210 16952
rect 11793 16949 11805 16952
rect 11839 16949 11851 16983
rect 11793 16943 11851 16949
rect 19794 16940 19800 16992
rect 19852 16980 19858 16992
rect 20257 16983 20315 16989
rect 20257 16980 20269 16983
rect 19852 16952 20269 16980
rect 19852 16940 19858 16952
rect 20257 16949 20269 16952
rect 20303 16949 20315 16983
rect 20257 16943 20315 16949
rect 22370 16940 22376 16992
rect 22428 16980 22434 16992
rect 23290 16980 23296 16992
rect 22428 16952 23296 16980
rect 22428 16940 22434 16952
rect 23290 16940 23296 16952
rect 23348 16980 23354 16992
rect 24044 16980 24072 17020
rect 30006 17008 30012 17060
rect 30064 17048 30070 17060
rect 31404 17048 31432 17156
rect 31665 17153 31677 17156
rect 31711 17153 31723 17187
rect 31665 17147 31723 17153
rect 31757 17187 31815 17193
rect 31757 17153 31769 17187
rect 31803 17184 31815 17187
rect 32582 17184 32588 17196
rect 31803 17156 32588 17184
rect 31803 17153 31815 17156
rect 31757 17147 31815 17153
rect 32582 17144 32588 17156
rect 32640 17144 32646 17196
rect 32876 17184 32904 17280
rect 33137 17187 33195 17193
rect 33137 17184 33149 17187
rect 32876 17156 33149 17184
rect 33137 17153 33149 17156
rect 33183 17153 33195 17187
rect 33137 17147 33195 17153
rect 33321 17187 33379 17193
rect 33321 17153 33333 17187
rect 33367 17153 33379 17187
rect 33321 17147 33379 17153
rect 33336 17116 33364 17147
rect 31726 17088 33364 17116
rect 30064 17020 31432 17048
rect 31481 17051 31539 17057
rect 30064 17008 30070 17020
rect 31481 17017 31493 17051
rect 31527 17048 31539 17051
rect 31726 17048 31754 17088
rect 31527 17020 31754 17048
rect 31527 17017 31539 17020
rect 31481 17011 31539 17017
rect 23348 16952 24072 16980
rect 32493 16983 32551 16989
rect 23348 16940 23354 16952
rect 32493 16949 32505 16983
rect 32539 16980 32551 16983
rect 32582 16980 32588 16992
rect 32539 16952 32588 16980
rect 32539 16949 32551 16952
rect 32493 16943 32551 16949
rect 32582 16940 32588 16952
rect 32640 16940 32646 16992
rect 1104 16890 34868 16912
rect 1104 16838 5170 16890
rect 5222 16838 5234 16890
rect 5286 16838 5298 16890
rect 5350 16838 5362 16890
rect 5414 16838 5426 16890
rect 5478 16838 13611 16890
rect 13663 16838 13675 16890
rect 13727 16838 13739 16890
rect 13791 16838 13803 16890
rect 13855 16838 13867 16890
rect 13919 16838 22052 16890
rect 22104 16838 22116 16890
rect 22168 16838 22180 16890
rect 22232 16838 22244 16890
rect 22296 16838 22308 16890
rect 22360 16838 30493 16890
rect 30545 16838 30557 16890
rect 30609 16838 30621 16890
rect 30673 16838 30685 16890
rect 30737 16838 30749 16890
rect 30801 16838 34868 16890
rect 1104 16816 34868 16838
rect 2682 16736 2688 16788
rect 2740 16776 2746 16788
rect 3053 16779 3111 16785
rect 3053 16776 3065 16779
rect 2740 16748 3065 16776
rect 2740 16736 2746 16748
rect 3053 16745 3065 16748
rect 3099 16745 3111 16779
rect 3234 16776 3240 16788
rect 3195 16748 3240 16776
rect 3053 16739 3111 16745
rect 3234 16736 3240 16748
rect 3292 16736 3298 16788
rect 4246 16776 4252 16788
rect 4207 16748 4252 16776
rect 4246 16736 4252 16748
rect 4304 16736 4310 16788
rect 6270 16776 6276 16788
rect 5920 16748 6276 16776
rect 5920 16717 5948 16748
rect 6270 16736 6276 16748
rect 6328 16776 6334 16788
rect 6914 16776 6920 16788
rect 6328 16748 6920 16776
rect 6328 16736 6334 16748
rect 6914 16736 6920 16748
rect 6972 16776 6978 16788
rect 7331 16779 7389 16785
rect 7331 16776 7343 16779
rect 6972 16748 7343 16776
rect 6972 16736 6978 16748
rect 7331 16745 7343 16748
rect 7377 16745 7389 16779
rect 7331 16739 7389 16745
rect 5905 16711 5963 16717
rect 5905 16677 5917 16711
rect 5951 16677 5963 16711
rect 7190 16708 7196 16720
rect 7151 16680 7196 16708
rect 5905 16671 5963 16677
rect 7190 16668 7196 16680
rect 7248 16668 7254 16720
rect 7346 16708 7374 16739
rect 8202 16736 8208 16788
rect 8260 16776 8266 16788
rect 9769 16779 9827 16785
rect 9769 16776 9781 16779
rect 8260 16748 9781 16776
rect 8260 16736 8266 16748
rect 9769 16745 9781 16748
rect 9815 16745 9827 16779
rect 12250 16776 12256 16788
rect 12211 16748 12256 16776
rect 9769 16739 9827 16745
rect 12250 16736 12256 16748
rect 12308 16736 12314 16788
rect 19426 16776 19432 16788
rect 19387 16748 19432 16776
rect 19426 16736 19432 16748
rect 19484 16736 19490 16788
rect 22097 16779 22155 16785
rect 19536 16748 21680 16776
rect 10962 16708 10968 16720
rect 7346 16680 10968 16708
rect 10962 16668 10968 16680
rect 11020 16668 11026 16720
rect 14829 16711 14887 16717
rect 14829 16677 14841 16711
rect 14875 16708 14887 16711
rect 15194 16708 15200 16720
rect 14875 16680 15200 16708
rect 14875 16677 14887 16680
rect 14829 16671 14887 16677
rect 15194 16668 15200 16680
rect 15252 16668 15258 16720
rect 16298 16668 16304 16720
rect 16356 16708 16362 16720
rect 19536 16708 19564 16748
rect 16356 16680 19564 16708
rect 21652 16708 21680 16748
rect 22097 16745 22109 16779
rect 22143 16776 22155 16779
rect 22370 16776 22376 16788
rect 22143 16748 22376 16776
rect 22143 16745 22155 16748
rect 22097 16739 22155 16745
rect 22370 16736 22376 16748
rect 22428 16736 22434 16788
rect 25774 16776 25780 16788
rect 24596 16748 25780 16776
rect 24596 16708 24624 16748
rect 25774 16736 25780 16748
rect 25832 16736 25838 16788
rect 31110 16736 31116 16788
rect 31168 16776 31174 16788
rect 31205 16779 31263 16785
rect 31205 16776 31217 16779
rect 31168 16748 31217 16776
rect 31168 16736 31174 16748
rect 31205 16745 31217 16748
rect 31251 16745 31263 16779
rect 31205 16739 31263 16745
rect 31662 16736 31668 16788
rect 31720 16776 31726 16788
rect 32217 16779 32275 16785
rect 32217 16776 32229 16779
rect 31720 16748 32229 16776
rect 31720 16736 31726 16748
rect 32217 16745 32229 16748
rect 32263 16745 32275 16779
rect 32217 16739 32275 16745
rect 21652 16680 24624 16708
rect 16356 16668 16362 16680
rect 6546 16600 6552 16652
rect 6604 16640 6610 16652
rect 6733 16643 6791 16649
rect 6733 16640 6745 16643
rect 6604 16612 6745 16640
rect 6604 16600 6610 16612
rect 6733 16609 6745 16612
rect 6779 16609 6791 16643
rect 6733 16603 6791 16609
rect 7101 16643 7159 16649
rect 7101 16609 7113 16643
rect 7147 16609 7159 16643
rect 7208 16640 7236 16668
rect 7208 16612 9904 16640
rect 7101 16603 7159 16609
rect 4062 16572 4068 16584
rect 4023 16544 4068 16572
rect 4062 16532 4068 16544
rect 4120 16532 4126 16584
rect 4338 16572 4344 16584
rect 4299 16544 4344 16572
rect 4338 16532 4344 16544
rect 4396 16532 4402 16584
rect 6454 16532 6460 16584
rect 6512 16572 6518 16584
rect 7116 16572 7144 16603
rect 9876 16581 9904 16612
rect 11974 16600 11980 16652
rect 12032 16640 12038 16652
rect 12032 16612 12204 16640
rect 12032 16600 12038 16612
rect 9950 16581 9956 16584
rect 9677 16575 9735 16581
rect 9677 16572 9689 16575
rect 6512 16544 9689 16572
rect 6512 16532 6518 16544
rect 9677 16541 9689 16544
rect 9723 16541 9735 16575
rect 9876 16575 9956 16581
rect 9876 16572 9905 16575
rect 9803 16544 9905 16572
rect 9677 16535 9735 16541
rect 9893 16541 9905 16544
rect 9939 16541 9956 16575
rect 9893 16535 9956 16541
rect 9950 16532 9956 16535
rect 10008 16532 10014 16584
rect 10042 16532 10048 16584
rect 10100 16572 10106 16584
rect 12176 16581 12204 16612
rect 14734 16600 14740 16652
rect 14792 16640 14798 16652
rect 15289 16643 15347 16649
rect 15289 16640 15301 16643
rect 14792 16612 15301 16640
rect 14792 16600 14798 16612
rect 15289 16609 15301 16612
rect 15335 16609 15347 16643
rect 15289 16603 15347 16609
rect 19978 16600 19984 16652
rect 20036 16640 20042 16652
rect 20717 16643 20775 16649
rect 20717 16640 20729 16643
rect 20036 16612 20729 16640
rect 20036 16600 20042 16612
rect 20717 16609 20729 16612
rect 20763 16609 20775 16643
rect 20717 16603 20775 16609
rect 30024 16612 31524 16640
rect 30024 16584 30052 16612
rect 12161 16575 12219 16581
rect 10100 16544 10145 16572
rect 10100 16532 10106 16544
rect 12161 16541 12173 16575
rect 12207 16541 12219 16575
rect 12161 16535 12219 16541
rect 12434 16532 12440 16584
rect 12492 16572 12498 16584
rect 14369 16575 14427 16581
rect 12492 16544 12537 16572
rect 12492 16532 12498 16544
rect 14369 16541 14381 16575
rect 14415 16541 14427 16575
rect 14369 16535 14427 16541
rect 14645 16575 14703 16581
rect 14645 16541 14657 16575
rect 14691 16572 14703 16575
rect 15556 16575 15614 16581
rect 14691 16544 15516 16572
rect 14691 16541 14703 16544
rect 14645 16535 14703 16541
rect 3050 16464 3056 16516
rect 3108 16504 3114 16516
rect 3421 16507 3479 16513
rect 3421 16504 3433 16507
rect 3108 16476 3433 16504
rect 3108 16464 3114 16476
rect 3421 16473 3433 16476
rect 3467 16473 3479 16507
rect 3421 16467 3479 16473
rect 5537 16507 5595 16513
rect 5537 16473 5549 16507
rect 5583 16504 5595 16507
rect 6546 16504 6552 16516
rect 5583 16476 6552 16504
rect 5583 16473 5595 16476
rect 5537 16467 5595 16473
rect 6546 16464 6552 16476
rect 6604 16504 6610 16516
rect 7469 16507 7527 16513
rect 7469 16504 7481 16507
rect 6604 16476 7481 16504
rect 6604 16464 6610 16476
rect 7469 16473 7481 16476
rect 7515 16504 7527 16507
rect 11146 16504 11152 16516
rect 7515 16476 11152 16504
rect 7515 16473 7527 16476
rect 7469 16467 7527 16473
rect 11146 16464 11152 16476
rect 11204 16464 11210 16516
rect 14384 16504 14412 16535
rect 15286 16504 15292 16516
rect 14384 16476 15292 16504
rect 15286 16464 15292 16476
rect 15344 16464 15350 16516
rect 15488 16504 15516 16544
rect 15556 16541 15568 16575
rect 15602 16572 15614 16575
rect 15838 16572 15844 16584
rect 15602 16544 15844 16572
rect 15602 16541 15614 16544
rect 15556 16535 15614 16541
rect 15838 16532 15844 16544
rect 15896 16532 15902 16584
rect 17218 16572 17224 16584
rect 17179 16544 17224 16572
rect 17218 16532 17224 16544
rect 17276 16532 17282 16584
rect 19613 16575 19671 16581
rect 19613 16541 19625 16575
rect 19659 16541 19671 16575
rect 19794 16572 19800 16584
rect 19755 16544 19800 16572
rect 19613 16535 19671 16541
rect 16114 16504 16120 16516
rect 15488 16476 16120 16504
rect 16114 16464 16120 16476
rect 16172 16504 16178 16516
rect 16298 16504 16304 16516
rect 16172 16476 16304 16504
rect 16172 16464 16178 16476
rect 16298 16464 16304 16476
rect 16356 16464 16362 16516
rect 17310 16464 17316 16516
rect 17368 16504 17374 16516
rect 17589 16507 17647 16513
rect 17589 16504 17601 16507
rect 17368 16476 17601 16504
rect 17368 16464 17374 16476
rect 17589 16473 17601 16476
rect 17635 16473 17647 16507
rect 19628 16504 19656 16535
rect 19794 16532 19800 16544
rect 19852 16532 19858 16584
rect 19886 16532 19892 16584
rect 19944 16572 19950 16584
rect 24578 16572 24584 16584
rect 19944 16544 19989 16572
rect 24539 16544 24584 16572
rect 19944 16532 19950 16544
rect 24578 16532 24584 16544
rect 24636 16532 24642 16584
rect 24670 16532 24676 16584
rect 24728 16572 24734 16584
rect 26421 16575 26479 16581
rect 26421 16572 26433 16575
rect 24728 16544 26433 16572
rect 24728 16532 24734 16544
rect 26421 16541 26433 16544
rect 26467 16541 26479 16575
rect 26421 16535 26479 16541
rect 29086 16532 29092 16584
rect 29144 16572 29150 16584
rect 30006 16572 30012 16584
rect 29144 16544 30012 16572
rect 29144 16532 29150 16544
rect 30006 16532 30012 16544
rect 30064 16532 30070 16584
rect 30098 16532 30104 16584
rect 30156 16572 30162 16584
rect 31496 16581 31524 16612
rect 32214 16600 32220 16652
rect 32272 16640 32278 16652
rect 32490 16640 32496 16652
rect 32272 16612 32496 16640
rect 32272 16600 32278 16612
rect 31389 16575 31447 16581
rect 31389 16572 31401 16575
rect 30156 16544 31401 16572
rect 30156 16532 30162 16544
rect 31389 16541 31401 16544
rect 31435 16541 31447 16575
rect 31389 16535 31447 16541
rect 31481 16575 31539 16581
rect 31481 16541 31493 16575
rect 31527 16541 31539 16575
rect 31481 16535 31539 16541
rect 31609 16575 31667 16581
rect 31609 16541 31621 16575
rect 31655 16572 31667 16575
rect 32324 16572 32352 16612
rect 32490 16600 32496 16612
rect 32548 16640 32554 16652
rect 32585 16643 32643 16649
rect 32585 16640 32597 16643
rect 32548 16612 32597 16640
rect 32548 16600 32554 16612
rect 32585 16609 32597 16612
rect 32631 16609 32643 16643
rect 32585 16603 32643 16609
rect 31655 16544 32352 16572
rect 31655 16541 31667 16544
rect 31609 16535 31667 16541
rect 20714 16504 20720 16516
rect 19628 16476 20720 16504
rect 17589 16467 17647 16473
rect 20714 16464 20720 16476
rect 20772 16464 20778 16516
rect 20990 16513 20996 16516
rect 20984 16467 20996 16513
rect 21048 16504 21054 16516
rect 24848 16507 24906 16513
rect 21048 16476 21084 16504
rect 20990 16464 20996 16467
rect 21048 16464 21054 16476
rect 24848 16473 24860 16507
rect 24894 16504 24906 16507
rect 25866 16504 25872 16516
rect 24894 16476 25872 16504
rect 24894 16473 24906 16476
rect 24848 16467 24906 16473
rect 25866 16464 25872 16476
rect 25924 16464 25930 16516
rect 26142 16464 26148 16516
rect 26200 16504 26206 16516
rect 26697 16507 26755 16513
rect 26697 16504 26709 16507
rect 26200 16476 26709 16504
rect 26200 16464 26206 16476
rect 26697 16473 26709 16476
rect 26743 16473 26755 16507
rect 29730 16504 29736 16516
rect 29691 16476 29736 16504
rect 26697 16467 26755 16473
rect 29730 16464 29736 16476
rect 29788 16464 29794 16516
rect 29917 16507 29975 16513
rect 29917 16473 29929 16507
rect 29963 16504 29975 16507
rect 30374 16504 30380 16516
rect 29963 16476 30380 16504
rect 29963 16473 29975 16476
rect 29917 16467 29975 16473
rect 30374 16464 30380 16476
rect 30432 16504 30438 16516
rect 31205 16507 31263 16513
rect 31205 16504 31217 16507
rect 30432 16476 31217 16504
rect 30432 16464 30438 16476
rect 31205 16473 31217 16476
rect 31251 16504 31263 16507
rect 31294 16504 31300 16516
rect 31251 16476 31300 16504
rect 31251 16473 31263 16476
rect 31205 16467 31263 16473
rect 31294 16464 31300 16476
rect 31352 16464 31358 16516
rect 3221 16439 3279 16445
rect 3221 16405 3233 16439
rect 3267 16436 3279 16439
rect 5997 16439 6055 16445
rect 5997 16436 6009 16439
rect 3267 16408 6009 16436
rect 3267 16405 3279 16408
rect 3221 16399 3279 16405
rect 5997 16405 6009 16408
rect 6043 16436 6055 16439
rect 6362 16436 6368 16448
rect 6043 16408 6368 16436
rect 6043 16405 6055 16408
rect 5997 16399 6055 16405
rect 6362 16396 6368 16408
rect 6420 16396 6426 16448
rect 10229 16439 10287 16445
rect 10229 16405 10241 16439
rect 10275 16436 10287 16439
rect 10410 16436 10416 16448
rect 10275 16408 10416 16436
rect 10275 16405 10287 16408
rect 10229 16399 10287 16405
rect 10410 16396 10416 16408
rect 10468 16396 10474 16448
rect 14458 16436 14464 16448
rect 14419 16408 14464 16436
rect 14458 16396 14464 16408
rect 14516 16396 14522 16448
rect 16666 16436 16672 16448
rect 16579 16408 16672 16436
rect 16666 16396 16672 16408
rect 16724 16436 16730 16448
rect 17494 16436 17500 16448
rect 16724 16408 17500 16436
rect 16724 16396 16730 16408
rect 17494 16396 17500 16408
rect 17552 16396 17558 16448
rect 19886 16396 19892 16448
rect 19944 16436 19950 16448
rect 20898 16436 20904 16448
rect 19944 16408 20904 16436
rect 19944 16396 19950 16408
rect 20898 16396 20904 16408
rect 20956 16396 20962 16448
rect 25961 16439 26019 16445
rect 25961 16405 25973 16439
rect 26007 16436 26019 16439
rect 26050 16436 26056 16448
rect 26007 16408 26056 16436
rect 26007 16405 26019 16408
rect 25961 16399 26019 16405
rect 26050 16396 26056 16408
rect 26108 16396 26114 16448
rect 30098 16396 30104 16448
rect 30156 16436 30162 16448
rect 30282 16436 30288 16448
rect 30156 16408 30201 16436
rect 30243 16408 30288 16436
rect 30156 16396 30162 16408
rect 30282 16396 30288 16408
rect 30340 16396 30346 16448
rect 31404 16436 31432 16535
rect 32398 16532 32404 16584
rect 32456 16572 32462 16584
rect 32456 16544 32549 16572
rect 32456 16532 32462 16544
rect 32416 16504 32444 16532
rect 31726 16476 32444 16504
rect 31726 16436 31754 16476
rect 31404 16408 31754 16436
rect 1104 16346 35027 16368
rect 1104 16294 9390 16346
rect 9442 16294 9454 16346
rect 9506 16294 9518 16346
rect 9570 16294 9582 16346
rect 9634 16294 9646 16346
rect 9698 16294 17831 16346
rect 17883 16294 17895 16346
rect 17947 16294 17959 16346
rect 18011 16294 18023 16346
rect 18075 16294 18087 16346
rect 18139 16294 26272 16346
rect 26324 16294 26336 16346
rect 26388 16294 26400 16346
rect 26452 16294 26464 16346
rect 26516 16294 26528 16346
rect 26580 16294 34713 16346
rect 34765 16294 34777 16346
rect 34829 16294 34841 16346
rect 34893 16294 34905 16346
rect 34957 16294 34969 16346
rect 35021 16294 35027 16346
rect 1104 16272 35027 16294
rect 6730 16232 6736 16244
rect 6691 16204 6736 16232
rect 6730 16192 6736 16204
rect 6788 16192 6794 16244
rect 10965 16235 11023 16241
rect 10965 16201 10977 16235
rect 11011 16232 11023 16235
rect 12342 16232 12348 16244
rect 11011 16204 12348 16232
rect 11011 16201 11023 16204
rect 10965 16195 11023 16201
rect 12342 16192 12348 16204
rect 12400 16192 12406 16244
rect 13262 16192 13268 16244
rect 13320 16232 13326 16244
rect 13541 16235 13599 16241
rect 13541 16232 13553 16235
rect 13320 16204 13553 16232
rect 13320 16192 13326 16204
rect 13541 16201 13553 16204
rect 13587 16232 13599 16235
rect 18690 16232 18696 16244
rect 13587 16204 17724 16232
rect 18651 16204 18696 16232
rect 13587 16201 13599 16204
rect 13541 16195 13599 16201
rect 5718 16164 5724 16176
rect 5631 16136 5724 16164
rect 5718 16124 5724 16136
rect 5776 16164 5782 16176
rect 6822 16164 6828 16176
rect 5776 16136 6828 16164
rect 5776 16124 5782 16136
rect 6822 16124 6828 16136
rect 6880 16124 6886 16176
rect 8941 16167 8999 16173
rect 8941 16133 8953 16167
rect 8987 16164 8999 16167
rect 11330 16164 11336 16176
rect 8987 16136 11336 16164
rect 8987 16133 8999 16136
rect 8941 16127 8999 16133
rect 11330 16124 11336 16136
rect 11388 16124 11394 16176
rect 13446 16124 13452 16176
rect 13504 16164 13510 16176
rect 15194 16173 15200 16176
rect 14093 16167 14151 16173
rect 14093 16164 14105 16167
rect 13504 16136 14105 16164
rect 13504 16124 13510 16136
rect 14093 16133 14105 16136
rect 14139 16133 14151 16167
rect 15188 16164 15200 16173
rect 15155 16136 15200 16164
rect 14093 16127 14151 16133
rect 15188 16127 15200 16136
rect 15194 16124 15200 16127
rect 15252 16124 15258 16176
rect 5537 16099 5595 16105
rect 5537 16065 5549 16099
rect 5583 16065 5595 16099
rect 6546 16096 6552 16108
rect 6507 16068 6552 16096
rect 5537 16059 5595 16065
rect 5353 16031 5411 16037
rect 5353 15997 5365 16031
rect 5399 15997 5411 16031
rect 5552 16028 5580 16059
rect 6546 16056 6552 16068
rect 6604 16056 6610 16108
rect 6733 16099 6791 16105
rect 6733 16065 6745 16099
rect 6779 16096 6791 16099
rect 6914 16096 6920 16108
rect 6779 16068 6920 16096
rect 6779 16065 6791 16068
rect 6733 16059 6791 16065
rect 6914 16056 6920 16068
rect 6972 16056 6978 16108
rect 7374 16096 7380 16108
rect 7335 16068 7380 16096
rect 7374 16056 7380 16068
rect 7432 16056 7438 16108
rect 7466 16056 7472 16108
rect 7524 16096 7530 16108
rect 8849 16099 8907 16105
rect 8849 16096 8861 16099
rect 7524 16068 8861 16096
rect 7524 16056 7530 16068
rect 8849 16065 8861 16068
rect 8895 16065 8907 16099
rect 10410 16096 10416 16108
rect 10371 16068 10416 16096
rect 8849 16059 8907 16065
rect 10410 16056 10416 16068
rect 10468 16056 10474 16108
rect 10962 16096 10968 16108
rect 10923 16068 10968 16096
rect 10962 16056 10968 16068
rect 11020 16056 11026 16108
rect 11146 16096 11152 16108
rect 11107 16068 11152 16096
rect 11146 16056 11152 16068
rect 11204 16056 11210 16108
rect 13357 16099 13415 16105
rect 13357 16096 13369 16099
rect 12406 16068 13369 16096
rect 7190 16028 7196 16040
rect 5552 16000 7196 16028
rect 5353 15991 5411 15997
rect 5368 15960 5396 15991
rect 7190 15988 7196 16000
rect 7248 15988 7254 16040
rect 7653 16031 7711 16037
rect 7653 15997 7665 16031
rect 7699 15997 7711 16031
rect 7653 15991 7711 15997
rect 5534 15960 5540 15972
rect 5368 15932 5540 15960
rect 5534 15920 5540 15932
rect 5592 15960 5598 15972
rect 6454 15960 6460 15972
rect 5592 15932 6460 15960
rect 5592 15920 5598 15932
rect 6454 15920 6460 15932
rect 6512 15960 6518 15972
rect 7668 15960 7696 15991
rect 6512 15932 7696 15960
rect 7929 15963 7987 15969
rect 6512 15920 6518 15932
rect 7929 15929 7941 15963
rect 7975 15960 7987 15963
rect 12406 15960 12434 16068
rect 13357 16065 13369 16068
rect 13403 16065 13415 16099
rect 14274 16096 14280 16108
rect 14235 16068 14280 16096
rect 13357 16059 13415 16065
rect 14274 16056 14280 16068
rect 14332 16056 14338 16108
rect 14461 16099 14519 16105
rect 14461 16065 14473 16099
rect 14507 16096 14519 16099
rect 16298 16096 16304 16108
rect 14507 16068 16304 16096
rect 14507 16065 14519 16068
rect 14461 16059 14519 16065
rect 16298 16056 16304 16068
rect 16356 16056 16362 16108
rect 17402 16096 17408 16108
rect 17363 16068 17408 16096
rect 17402 16056 17408 16068
rect 17460 16056 17466 16108
rect 17586 16096 17592 16108
rect 17547 16068 17592 16096
rect 17586 16056 17592 16068
rect 17644 16056 17650 16108
rect 17696 16096 17724 16204
rect 18690 16192 18696 16204
rect 18748 16192 18754 16244
rect 22646 16232 22652 16244
rect 19904 16204 20760 16232
rect 17773 16167 17831 16173
rect 17773 16133 17785 16167
rect 17819 16164 17831 16167
rect 19334 16164 19340 16176
rect 17819 16136 19340 16164
rect 17819 16133 17831 16136
rect 17773 16127 17831 16133
rect 19334 16124 19340 16136
rect 19392 16164 19398 16176
rect 19904 16164 19932 16204
rect 19392 16136 19932 16164
rect 19981 16167 20039 16173
rect 19392 16124 19398 16136
rect 19981 16133 19993 16167
rect 20027 16164 20039 16167
rect 20346 16164 20352 16176
rect 20027 16136 20352 16164
rect 20027 16133 20039 16136
rect 19981 16127 20039 16133
rect 20346 16124 20352 16136
rect 20404 16124 20410 16176
rect 20732 16173 20760 16204
rect 20824 16204 22508 16232
rect 22607 16204 22652 16232
rect 20824 16173 20852 16204
rect 20717 16167 20775 16173
rect 20717 16133 20729 16167
rect 20763 16133 20775 16167
rect 20717 16127 20775 16133
rect 20809 16167 20867 16173
rect 20809 16133 20821 16167
rect 20855 16133 20867 16167
rect 20809 16127 20867 16133
rect 20162 16096 20168 16108
rect 17696 16068 20168 16096
rect 20162 16056 20168 16068
rect 20220 16056 20226 16108
rect 20438 16096 20444 16108
rect 20399 16068 20444 16096
rect 20438 16056 20444 16068
rect 20496 16056 20502 16108
rect 20534 16099 20592 16105
rect 20534 16065 20546 16099
rect 20580 16065 20592 16099
rect 20534 16059 20592 16065
rect 14734 15988 14740 16040
rect 14792 16028 14798 16040
rect 14921 16031 14979 16037
rect 14921 16028 14933 16031
rect 14792 16000 14933 16028
rect 14792 15988 14798 16000
rect 14921 15997 14933 16000
rect 14967 15997 14979 16031
rect 14921 15991 14979 15997
rect 19794 15988 19800 16040
rect 19852 16028 19858 16040
rect 20548 16028 20576 16059
rect 19852 16000 20576 16028
rect 20732 16028 20760 16127
rect 21082 16124 21088 16176
rect 21140 16164 21146 16176
rect 22480 16164 22508 16204
rect 22646 16192 22652 16204
rect 22704 16192 22710 16244
rect 25866 16192 25872 16244
rect 25924 16232 25930 16244
rect 25961 16235 26019 16241
rect 25961 16232 25973 16235
rect 25924 16204 25973 16232
rect 25924 16192 25930 16204
rect 25961 16201 25973 16204
rect 26007 16201 26019 16235
rect 25961 16195 26019 16201
rect 28997 16235 29055 16241
rect 28997 16201 29009 16235
rect 29043 16201 29055 16235
rect 28997 16195 29055 16201
rect 26050 16164 26056 16176
rect 21140 16136 22140 16164
rect 22480 16136 26056 16164
rect 21140 16124 21146 16136
rect 20947 16099 21005 16105
rect 20947 16065 20959 16099
rect 20993 16096 21005 16099
rect 21634 16096 21640 16108
rect 20993 16068 21640 16096
rect 20993 16065 21005 16068
rect 20947 16059 21005 16065
rect 21634 16056 21640 16068
rect 21692 16056 21698 16108
rect 22002 16096 22008 16108
rect 21963 16068 22008 16096
rect 22002 16056 22008 16068
rect 22060 16056 22066 16108
rect 22112 16105 22140 16136
rect 26050 16124 26056 16136
rect 26108 16164 26114 16176
rect 26329 16167 26387 16173
rect 26329 16164 26341 16167
rect 26108 16136 26341 16164
rect 26108 16124 26114 16136
rect 26329 16133 26341 16136
rect 26375 16133 26387 16167
rect 29012 16164 29040 16195
rect 32490 16192 32496 16244
rect 32548 16232 32554 16244
rect 33042 16232 33048 16244
rect 32548 16204 33048 16232
rect 32548 16192 32554 16204
rect 33042 16192 33048 16204
rect 33100 16232 33106 16244
rect 33689 16235 33747 16241
rect 33689 16232 33701 16235
rect 33100 16204 33701 16232
rect 33100 16192 33106 16204
rect 33689 16201 33701 16204
rect 33735 16201 33747 16235
rect 33689 16195 33747 16201
rect 26329 16127 26387 16133
rect 28184 16136 29040 16164
rect 29273 16167 29331 16173
rect 22098 16099 22156 16105
rect 22098 16065 22110 16099
rect 22144 16065 22156 16099
rect 22098 16059 22156 16065
rect 22281 16099 22339 16105
rect 22281 16065 22293 16099
rect 22327 16065 22339 16099
rect 22281 16059 22339 16065
rect 20732 16000 21956 16028
rect 19852 15988 19858 16000
rect 7975 15932 12434 15960
rect 7975 15929 7987 15932
rect 7929 15923 7987 15929
rect 20622 15920 20628 15972
rect 20680 15960 20686 15972
rect 21085 15963 21143 15969
rect 21085 15960 21097 15963
rect 20680 15932 21097 15960
rect 20680 15920 20686 15932
rect 21085 15929 21097 15932
rect 21131 15929 21143 15963
rect 21928 15960 21956 16000
rect 22296 15960 22324 16059
rect 22370 16056 22376 16108
rect 22428 16096 22434 16108
rect 22511 16099 22569 16105
rect 22428 16068 22473 16096
rect 22428 16056 22434 16068
rect 22511 16065 22523 16099
rect 22557 16096 22569 16099
rect 22646 16096 22652 16108
rect 22557 16068 22652 16096
rect 22557 16065 22569 16068
rect 22511 16059 22569 16065
rect 22646 16056 22652 16068
rect 22704 16056 22710 16108
rect 25130 16096 25136 16108
rect 25091 16068 25136 16096
rect 25130 16056 25136 16068
rect 25188 16056 25194 16108
rect 25774 16056 25780 16108
rect 25832 16096 25838 16108
rect 28184 16105 28212 16136
rect 29273 16133 29285 16167
rect 29319 16164 29331 16167
rect 30374 16164 30380 16176
rect 29319 16136 30380 16164
rect 29319 16133 29331 16136
rect 29273 16127 29331 16133
rect 30374 16124 30380 16136
rect 30432 16124 30438 16176
rect 26145 16099 26203 16105
rect 26145 16096 26157 16099
rect 25832 16068 26157 16096
rect 25832 16056 25838 16068
rect 26145 16065 26157 16068
rect 26191 16065 26203 16099
rect 26145 16059 26203 16065
rect 26421 16099 26479 16105
rect 26421 16065 26433 16099
rect 26467 16065 26479 16099
rect 26421 16059 26479 16065
rect 28169 16099 28227 16105
rect 28169 16065 28181 16099
rect 28215 16065 28227 16099
rect 28442 16096 28448 16108
rect 28403 16068 28448 16096
rect 28169 16059 28227 16065
rect 24486 15988 24492 16040
rect 24544 16028 24550 16040
rect 26436 16028 26464 16059
rect 28442 16056 28448 16068
rect 28500 16056 28506 16108
rect 29086 16056 29092 16108
rect 29144 16096 29150 16108
rect 29181 16099 29239 16105
rect 29181 16096 29193 16099
rect 29144 16068 29193 16096
rect 29144 16056 29150 16068
rect 29181 16065 29193 16068
rect 29227 16065 29239 16099
rect 29365 16099 29423 16105
rect 29365 16096 29377 16099
rect 29181 16059 29239 16065
rect 29288 16068 29377 16096
rect 27706 16028 27712 16040
rect 24544 16000 27712 16028
rect 24544 15988 24550 16000
rect 27706 15988 27712 16000
rect 27764 15988 27770 16040
rect 27798 15988 27804 16040
rect 27856 16028 27862 16040
rect 28261 16031 28319 16037
rect 28261 16028 28273 16031
rect 27856 16000 28273 16028
rect 27856 15988 27862 16000
rect 28261 15997 28273 16000
rect 28307 15997 28319 16031
rect 28261 15991 28319 15997
rect 28350 15988 28356 16040
rect 28408 16028 28414 16040
rect 29288 16028 29316 16068
rect 29365 16065 29377 16068
rect 29411 16065 29423 16099
rect 29365 16059 29423 16065
rect 29549 16099 29607 16105
rect 29549 16065 29561 16099
rect 29595 16096 29607 16099
rect 29730 16096 29736 16108
rect 29595 16068 29736 16096
rect 29595 16065 29607 16068
rect 29549 16059 29607 16065
rect 29730 16056 29736 16068
rect 29788 16056 29794 16108
rect 32576 16099 32634 16105
rect 32576 16065 32588 16099
rect 32622 16096 32634 16099
rect 33870 16096 33876 16108
rect 32622 16068 33876 16096
rect 32622 16065 32634 16068
rect 32576 16059 32634 16065
rect 33870 16056 33876 16068
rect 33928 16056 33934 16108
rect 30098 16028 30104 16040
rect 28408 16000 28453 16028
rect 29288 16000 30104 16028
rect 28408 15988 28414 16000
rect 27985 15963 28043 15969
rect 27985 15960 27997 15963
rect 21928 15932 22324 15960
rect 23768 15932 27997 15960
rect 21085 15923 21143 15929
rect 7742 15892 7748 15904
rect 7703 15864 7748 15892
rect 7742 15852 7748 15864
rect 7800 15852 7806 15904
rect 14458 15852 14464 15904
rect 14516 15892 14522 15904
rect 16301 15895 16359 15901
rect 16301 15892 16313 15895
rect 14516 15864 16313 15892
rect 14516 15852 14522 15864
rect 16301 15861 16313 15864
rect 16347 15892 16359 15895
rect 20070 15892 20076 15904
rect 16347 15864 20076 15892
rect 16347 15861 16359 15864
rect 16301 15855 16359 15861
rect 20070 15852 20076 15864
rect 20128 15852 20134 15904
rect 22002 15852 22008 15904
rect 22060 15892 22066 15904
rect 23768 15892 23796 15932
rect 27985 15929 27997 15932
rect 28031 15929 28043 15963
rect 27985 15923 28043 15929
rect 22060 15864 23796 15892
rect 23845 15895 23903 15901
rect 22060 15852 22066 15864
rect 23845 15861 23857 15895
rect 23891 15892 23903 15895
rect 24578 15892 24584 15904
rect 23891 15864 24584 15892
rect 23891 15861 23903 15864
rect 23845 15855 23903 15861
rect 24578 15852 24584 15864
rect 24636 15852 24642 15904
rect 25222 15852 25228 15904
rect 25280 15892 25286 15904
rect 29288 15892 29316 16000
rect 30098 15988 30104 16000
rect 30156 15988 30162 16040
rect 32306 16028 32312 16040
rect 32267 16000 32312 16028
rect 32306 15988 32312 16000
rect 32364 15988 32370 16040
rect 25280 15864 29316 15892
rect 25280 15852 25286 15864
rect 1104 15802 34868 15824
rect 1104 15750 5170 15802
rect 5222 15750 5234 15802
rect 5286 15750 5298 15802
rect 5350 15750 5362 15802
rect 5414 15750 5426 15802
rect 5478 15750 13611 15802
rect 13663 15750 13675 15802
rect 13727 15750 13739 15802
rect 13791 15750 13803 15802
rect 13855 15750 13867 15802
rect 13919 15750 22052 15802
rect 22104 15750 22116 15802
rect 22168 15750 22180 15802
rect 22232 15750 22244 15802
rect 22296 15750 22308 15802
rect 22360 15750 30493 15802
rect 30545 15750 30557 15802
rect 30609 15750 30621 15802
rect 30673 15750 30685 15802
rect 30737 15750 30749 15802
rect 30801 15750 34868 15802
rect 1104 15728 34868 15750
rect 4798 15648 4804 15700
rect 4856 15688 4862 15700
rect 5261 15691 5319 15697
rect 5261 15688 5273 15691
rect 4856 15660 5273 15688
rect 4856 15648 4862 15660
rect 5261 15657 5273 15660
rect 5307 15688 5319 15691
rect 7742 15688 7748 15700
rect 5307 15660 7748 15688
rect 5307 15657 5319 15660
rect 5261 15651 5319 15657
rect 7742 15648 7748 15660
rect 7800 15648 7806 15700
rect 18049 15691 18107 15697
rect 18049 15657 18061 15691
rect 18095 15688 18107 15691
rect 19242 15688 19248 15700
rect 18095 15660 19248 15688
rect 18095 15657 18107 15660
rect 18049 15651 18107 15657
rect 19242 15648 19248 15660
rect 19300 15648 19306 15700
rect 19886 15688 19892 15700
rect 19847 15660 19892 15688
rect 19886 15648 19892 15660
rect 19944 15648 19950 15700
rect 25130 15648 25136 15700
rect 25188 15688 25194 15700
rect 26050 15688 26056 15700
rect 25188 15660 26056 15688
rect 25188 15648 25194 15660
rect 26050 15648 26056 15660
rect 26108 15688 26114 15700
rect 26513 15691 26571 15697
rect 26513 15688 26525 15691
rect 26108 15660 26525 15688
rect 26108 15648 26114 15660
rect 26513 15657 26525 15660
rect 26559 15657 26571 15691
rect 26513 15651 26571 15657
rect 28350 15648 28356 15700
rect 28408 15688 28414 15700
rect 29089 15691 29147 15697
rect 29089 15688 29101 15691
rect 28408 15660 29101 15688
rect 28408 15648 28414 15660
rect 29089 15657 29101 15660
rect 29135 15657 29147 15691
rect 29089 15651 29147 15657
rect 31665 15691 31723 15697
rect 31665 15657 31677 15691
rect 31711 15688 31723 15691
rect 31754 15688 31760 15700
rect 31711 15660 31760 15688
rect 31711 15657 31723 15660
rect 31665 15651 31723 15657
rect 31754 15648 31760 15660
rect 31812 15688 31818 15700
rect 32306 15688 32312 15700
rect 31812 15660 32312 15688
rect 31812 15648 31818 15660
rect 32306 15648 32312 15660
rect 32364 15648 32370 15700
rect 33870 15688 33876 15700
rect 33831 15660 33876 15688
rect 33870 15648 33876 15660
rect 33928 15648 33934 15700
rect 13633 15623 13691 15629
rect 13633 15589 13645 15623
rect 13679 15620 13691 15623
rect 18230 15620 18236 15632
rect 13679 15592 18236 15620
rect 13679 15589 13691 15592
rect 13633 15583 13691 15589
rect 18230 15580 18236 15592
rect 18288 15580 18294 15632
rect 22370 15580 22376 15632
rect 22428 15620 22434 15632
rect 32674 15620 32680 15632
rect 22428 15592 32680 15620
rect 22428 15580 22434 15592
rect 32674 15580 32680 15592
rect 32732 15580 32738 15632
rect 4338 15552 4344 15564
rect 2700 15524 4344 15552
rect 2700 15493 2728 15524
rect 4338 15512 4344 15524
rect 4396 15512 4402 15564
rect 6546 15552 6552 15564
rect 6104 15524 6552 15552
rect 6104 15496 6132 15524
rect 6546 15512 6552 15524
rect 6604 15512 6610 15564
rect 13262 15512 13268 15564
rect 13320 15552 13326 15564
rect 16574 15552 16580 15564
rect 13320 15524 14320 15552
rect 13320 15512 13326 15524
rect 2685 15487 2743 15493
rect 2685 15453 2697 15487
rect 2731 15453 2743 15487
rect 2685 15447 2743 15453
rect 2869 15487 2927 15493
rect 2869 15453 2881 15487
rect 2915 15484 2927 15487
rect 4062 15484 4068 15496
rect 2915 15456 4068 15484
rect 2915 15453 2927 15456
rect 2869 15447 2927 15453
rect 4062 15444 4068 15456
rect 4120 15444 4126 15496
rect 6086 15484 6092 15496
rect 5999 15456 6092 15484
rect 6086 15444 6092 15456
rect 6144 15444 6150 15496
rect 6270 15484 6276 15496
rect 6231 15456 6276 15484
rect 6270 15444 6276 15456
rect 6328 15444 6334 15496
rect 6730 15484 6736 15496
rect 6691 15456 6736 15484
rect 6730 15444 6736 15456
rect 6788 15444 6794 15496
rect 9766 15444 9772 15496
rect 9824 15484 9830 15496
rect 14292 15493 14320 15524
rect 16224 15524 16580 15552
rect 16224 15493 16252 15524
rect 16574 15512 16580 15524
rect 16632 15552 16638 15564
rect 17402 15552 17408 15564
rect 16632 15524 17408 15552
rect 16632 15512 16638 15524
rect 17402 15512 17408 15524
rect 17460 15512 17466 15564
rect 17494 15512 17500 15564
rect 17552 15552 17558 15564
rect 21174 15552 21180 15564
rect 17552 15524 21180 15552
rect 17552 15512 17558 15524
rect 21174 15512 21180 15524
rect 21232 15512 21238 15564
rect 22554 15552 22560 15564
rect 22515 15524 22560 15552
rect 22554 15512 22560 15524
rect 22612 15512 22618 15564
rect 29546 15512 29552 15564
rect 29604 15552 29610 15564
rect 29604 15524 33732 15552
rect 29604 15512 29610 15524
rect 12529 15487 12587 15493
rect 12529 15484 12541 15487
rect 9824 15456 12541 15484
rect 9824 15444 9830 15456
rect 12529 15453 12541 15456
rect 12575 15453 12587 15487
rect 12529 15447 12587 15453
rect 12621 15487 12679 15493
rect 12621 15453 12633 15487
rect 12667 15484 12679 15487
rect 13357 15487 13415 15493
rect 13357 15484 13369 15487
rect 12667 15456 13369 15484
rect 12667 15453 12679 15456
rect 12621 15447 12679 15453
rect 13357 15453 13369 15456
rect 13403 15453 13415 15487
rect 13357 15447 13415 15453
rect 13633 15487 13691 15493
rect 13633 15453 13645 15487
rect 13679 15453 13691 15487
rect 13633 15447 13691 15453
rect 14277 15487 14335 15493
rect 14277 15453 14289 15487
rect 14323 15453 14335 15487
rect 14277 15447 14335 15453
rect 16209 15487 16267 15493
rect 16209 15453 16221 15487
rect 16255 15453 16267 15487
rect 16209 15447 16267 15453
rect 2958 15416 2964 15428
rect 2919 15388 2964 15416
rect 2958 15376 2964 15388
rect 3016 15376 3022 15428
rect 5445 15419 5503 15425
rect 5445 15385 5457 15419
rect 5491 15416 5503 15419
rect 5534 15416 5540 15428
rect 5491 15388 5540 15416
rect 5491 15385 5503 15388
rect 5445 15379 5503 15385
rect 5534 15376 5540 15388
rect 5592 15376 5598 15428
rect 6181 15419 6239 15425
rect 6181 15385 6193 15419
rect 6227 15416 6239 15419
rect 7374 15416 7380 15428
rect 6227 15388 7380 15416
rect 6227 15385 6239 15388
rect 6181 15379 6239 15385
rect 4430 15308 4436 15360
rect 4488 15348 4494 15360
rect 5077 15351 5135 15357
rect 5077 15348 5089 15351
rect 4488 15320 5089 15348
rect 4488 15308 4494 15320
rect 5077 15317 5089 15320
rect 5123 15317 5135 15351
rect 5077 15311 5135 15317
rect 5245 15351 5303 15357
rect 5245 15317 5257 15351
rect 5291 15348 5303 15351
rect 6196 15348 6224 15379
rect 7374 15376 7380 15388
rect 7432 15376 7438 15428
rect 13648 15416 13676 15447
rect 16298 15444 16304 15496
rect 16356 15484 16362 15496
rect 16393 15487 16451 15493
rect 16393 15484 16405 15487
rect 16356 15456 16405 15484
rect 16356 15444 16362 15456
rect 16393 15453 16405 15456
rect 16439 15453 16451 15487
rect 16393 15447 16451 15453
rect 17957 15487 18015 15493
rect 17957 15453 17969 15487
rect 18003 15484 18015 15487
rect 18322 15484 18328 15496
rect 18003 15456 18328 15484
rect 18003 15453 18015 15456
rect 17957 15447 18015 15453
rect 18322 15444 18328 15456
rect 18380 15444 18386 15496
rect 20806 15484 20812 15496
rect 20767 15456 20812 15484
rect 20806 15444 20812 15456
rect 20864 15444 20870 15496
rect 23014 15444 23020 15496
rect 23072 15484 23078 15496
rect 23382 15484 23388 15496
rect 23072 15456 23388 15484
rect 23072 15444 23078 15456
rect 23382 15444 23388 15456
rect 23440 15444 23446 15496
rect 23661 15487 23719 15493
rect 23661 15453 23673 15487
rect 23707 15484 23719 15487
rect 24486 15484 24492 15496
rect 23707 15456 24492 15484
rect 23707 15453 23719 15456
rect 23661 15447 23719 15453
rect 24486 15444 24492 15456
rect 24544 15444 24550 15496
rect 29181 15487 29239 15493
rect 29181 15453 29193 15487
rect 29227 15484 29239 15487
rect 30282 15484 30288 15496
rect 29227 15456 30288 15484
rect 29227 15453 29239 15456
rect 29181 15447 29239 15453
rect 30282 15444 30288 15456
rect 30340 15444 30346 15496
rect 33410 15484 33416 15496
rect 33371 15456 33416 15484
rect 33410 15444 33416 15456
rect 33468 15444 33474 15496
rect 33704 15493 33732 15524
rect 33689 15487 33747 15493
rect 33689 15453 33701 15487
rect 33735 15453 33747 15487
rect 33689 15447 33747 15453
rect 14553 15419 14611 15425
rect 14553 15416 14565 15419
rect 13648 15388 14565 15416
rect 14553 15385 14565 15388
rect 14599 15416 14611 15419
rect 15286 15416 15292 15428
rect 14599 15388 15292 15416
rect 14599 15385 14611 15388
rect 14553 15379 14611 15385
rect 15286 15376 15292 15388
rect 15344 15416 15350 15428
rect 17126 15416 17132 15428
rect 15344 15388 17132 15416
rect 15344 15376 15350 15388
rect 17126 15376 17132 15388
rect 17184 15376 17190 15428
rect 17402 15376 17408 15428
rect 17460 15416 17466 15428
rect 17586 15416 17592 15428
rect 17460 15388 17592 15416
rect 17460 15376 17466 15388
rect 17586 15376 17592 15388
rect 17644 15416 17650 15428
rect 17773 15419 17831 15425
rect 17773 15416 17785 15419
rect 17644 15388 17785 15416
rect 17644 15376 17650 15388
rect 17773 15385 17785 15388
rect 17819 15385 17831 15419
rect 20162 15416 20168 15428
rect 20075 15388 20168 15416
rect 17773 15379 17831 15385
rect 20162 15376 20168 15388
rect 20220 15416 20226 15428
rect 20530 15416 20536 15428
rect 20220 15388 20536 15416
rect 20220 15376 20226 15388
rect 20530 15376 20536 15388
rect 20588 15416 20594 15428
rect 24670 15416 24676 15428
rect 20588 15388 24676 15416
rect 20588 15376 20594 15388
rect 24670 15376 24676 15388
rect 24728 15376 24734 15428
rect 25222 15416 25228 15428
rect 25183 15388 25228 15416
rect 25222 15376 25228 15388
rect 25280 15376 25286 15428
rect 25774 15376 25780 15428
rect 25832 15416 25838 15428
rect 28994 15416 29000 15428
rect 25832 15388 29000 15416
rect 25832 15376 25838 15388
rect 28994 15376 29000 15388
rect 29052 15376 29058 15428
rect 32953 15419 33011 15425
rect 32953 15385 32965 15419
rect 32999 15416 33011 15419
rect 33594 15416 33600 15428
rect 32999 15388 33600 15416
rect 32999 15385 33011 15388
rect 32953 15379 33011 15385
rect 33594 15376 33600 15388
rect 33652 15376 33658 15428
rect 6822 15348 6828 15360
rect 5291 15320 6224 15348
rect 6783 15320 6828 15348
rect 5291 15317 5303 15320
rect 5245 15311 5303 15317
rect 6822 15308 6828 15320
rect 6880 15308 6886 15360
rect 16390 15348 16396 15360
rect 16351 15320 16396 15348
rect 16390 15308 16396 15320
rect 16448 15308 16454 15360
rect 17310 15308 17316 15360
rect 17368 15348 17374 15360
rect 17494 15348 17500 15360
rect 17368 15320 17500 15348
rect 17368 15308 17374 15320
rect 17494 15308 17500 15320
rect 17552 15308 17558 15360
rect 20990 15308 20996 15360
rect 21048 15348 21054 15360
rect 22922 15348 22928 15360
rect 21048 15320 22928 15348
rect 21048 15308 21054 15320
rect 22922 15308 22928 15320
rect 22980 15308 22986 15360
rect 23201 15351 23259 15357
rect 23201 15317 23213 15351
rect 23247 15348 23259 15351
rect 23474 15348 23480 15360
rect 23247 15320 23480 15348
rect 23247 15317 23259 15320
rect 23201 15311 23259 15317
rect 23474 15308 23480 15320
rect 23532 15308 23538 15360
rect 23569 15351 23627 15357
rect 23569 15317 23581 15351
rect 23615 15348 23627 15351
rect 25958 15348 25964 15360
rect 23615 15320 25964 15348
rect 23615 15317 23627 15320
rect 23569 15311 23627 15317
rect 25958 15308 25964 15320
rect 26016 15308 26022 15360
rect 33042 15308 33048 15360
rect 33100 15348 33106 15360
rect 33505 15351 33563 15357
rect 33505 15348 33517 15351
rect 33100 15320 33517 15348
rect 33100 15308 33106 15320
rect 33505 15317 33517 15320
rect 33551 15317 33563 15351
rect 33505 15311 33563 15317
rect 1104 15258 35027 15280
rect 1104 15206 9390 15258
rect 9442 15206 9454 15258
rect 9506 15206 9518 15258
rect 9570 15206 9582 15258
rect 9634 15206 9646 15258
rect 9698 15206 17831 15258
rect 17883 15206 17895 15258
rect 17947 15206 17959 15258
rect 18011 15206 18023 15258
rect 18075 15206 18087 15258
rect 18139 15206 26272 15258
rect 26324 15206 26336 15258
rect 26388 15206 26400 15258
rect 26452 15206 26464 15258
rect 26516 15206 26528 15258
rect 26580 15206 34713 15258
rect 34765 15206 34777 15258
rect 34829 15206 34841 15258
rect 34893 15206 34905 15258
rect 34957 15206 34969 15258
rect 35021 15206 35027 15258
rect 1104 15184 35027 15206
rect 5436 15147 5494 15153
rect 5436 15113 5448 15147
rect 5482 15144 5494 15147
rect 5718 15144 5724 15156
rect 5482 15116 5724 15144
rect 5482 15113 5494 15116
rect 5436 15107 5494 15113
rect 5718 15104 5724 15116
rect 5776 15104 5782 15156
rect 16025 15147 16083 15153
rect 16025 15113 16037 15147
rect 16071 15144 16083 15147
rect 18414 15144 18420 15156
rect 16071 15116 18420 15144
rect 16071 15113 16083 15116
rect 16025 15107 16083 15113
rect 18414 15104 18420 15116
rect 18472 15104 18478 15156
rect 21818 15144 21824 15156
rect 19444 15116 21824 15144
rect 2958 15036 2964 15088
rect 3016 15036 3022 15088
rect 5813 15079 5871 15085
rect 5813 15045 5825 15079
rect 5859 15076 5871 15079
rect 6270 15076 6276 15088
rect 5859 15048 6276 15076
rect 5859 15045 5871 15048
rect 5813 15039 5871 15045
rect 6270 15036 6276 15048
rect 6328 15036 6334 15088
rect 9677 15079 9735 15085
rect 9677 15045 9689 15079
rect 9723 15076 9735 15079
rect 11790 15076 11796 15088
rect 9723 15048 11796 15076
rect 9723 15045 9735 15048
rect 9677 15039 9735 15045
rect 11790 15036 11796 15048
rect 11848 15036 11854 15088
rect 16853 15079 16911 15085
rect 16853 15045 16865 15079
rect 16899 15076 16911 15079
rect 16942 15076 16948 15088
rect 16899 15048 16948 15076
rect 16899 15045 16911 15048
rect 16853 15039 16911 15045
rect 16942 15036 16948 15048
rect 17000 15076 17006 15088
rect 17862 15076 17868 15088
rect 17000 15048 17868 15076
rect 17000 15036 17006 15048
rect 17862 15036 17868 15048
rect 17920 15036 17926 15088
rect 19444 15076 19472 15116
rect 21818 15104 21824 15116
rect 21876 15104 21882 15156
rect 22922 15144 22928 15156
rect 22883 15116 22928 15144
rect 22922 15104 22928 15116
rect 22980 15104 22986 15156
rect 23290 15144 23296 15156
rect 23251 15116 23296 15144
rect 23290 15104 23296 15116
rect 23348 15104 23354 15156
rect 23382 15104 23388 15156
rect 23440 15144 23446 15156
rect 25130 15144 25136 15156
rect 23440 15116 25136 15144
rect 23440 15104 23446 15116
rect 25130 15104 25136 15116
rect 25188 15144 25194 15156
rect 29546 15144 29552 15156
rect 25188 15116 29552 15144
rect 25188 15104 25194 15116
rect 29546 15104 29552 15116
rect 29604 15104 29610 15156
rect 33594 15144 33600 15156
rect 33555 15116 33600 15144
rect 33594 15104 33600 15116
rect 33652 15104 33658 15156
rect 19978 15076 19984 15088
rect 18064 15048 19472 15076
rect 19939 15048 19984 15076
rect 4157 15011 4215 15017
rect 4157 14977 4169 15011
rect 4203 15008 4215 15011
rect 4522 15008 4528 15020
rect 4203 14980 4528 15008
rect 4203 14977 4215 14980
rect 4157 14971 4215 14977
rect 1670 14940 1676 14952
rect 1631 14912 1676 14940
rect 1670 14900 1676 14912
rect 1728 14900 1734 14952
rect 1949 14943 2007 14949
rect 1949 14909 1961 14943
rect 1995 14940 2007 14943
rect 2682 14940 2688 14952
rect 1995 14912 2688 14940
rect 1995 14909 2007 14912
rect 1949 14903 2007 14909
rect 2682 14900 2688 14912
rect 2740 14940 2746 14952
rect 4065 14943 4123 14949
rect 4065 14940 4077 14943
rect 2740 14912 4077 14940
rect 2740 14900 2746 14912
rect 4065 14909 4077 14912
rect 4111 14909 4123 14943
rect 4065 14903 4123 14909
rect 3234 14832 3240 14884
rect 3292 14872 3298 14884
rect 3421 14875 3479 14881
rect 3421 14872 3433 14875
rect 3292 14844 3433 14872
rect 3292 14832 3298 14844
rect 3421 14841 3433 14844
rect 3467 14872 3479 14875
rect 4172 14872 4200 14971
rect 4522 14968 4528 14980
rect 4580 14968 4586 15020
rect 9030 15008 9036 15020
rect 8991 14980 9036 15008
rect 9030 14968 9036 14980
rect 9088 14968 9094 15020
rect 9217 15011 9275 15017
rect 9217 14977 9229 15011
rect 9263 15008 9275 15011
rect 9950 15008 9956 15020
rect 9263 14980 9956 15008
rect 9263 14977 9275 14980
rect 9217 14971 9275 14977
rect 9950 14968 9956 14980
rect 10008 14968 10014 15020
rect 10505 15011 10563 15017
rect 10505 14977 10517 15011
rect 10551 14977 10563 15011
rect 10686 15008 10692 15020
rect 10647 14980 10692 15008
rect 10505 14971 10563 14977
rect 8938 14940 8944 14952
rect 8851 14912 8944 14940
rect 8938 14900 8944 14912
rect 8996 14940 9002 14952
rect 9858 14940 9864 14952
rect 8996 14912 9864 14940
rect 8996 14900 9002 14912
rect 9858 14900 9864 14912
rect 9916 14900 9922 14952
rect 10318 14900 10324 14952
rect 10376 14940 10382 14952
rect 10413 14943 10471 14949
rect 10413 14940 10425 14943
rect 10376 14912 10425 14940
rect 10376 14900 10382 14912
rect 10413 14909 10425 14912
rect 10459 14909 10471 14943
rect 10520 14940 10548 14971
rect 10686 14968 10692 14980
rect 10744 14968 10750 15020
rect 12158 15008 12164 15020
rect 10796 14980 12164 15008
rect 10796 14940 10824 14980
rect 12158 14968 12164 14980
rect 12216 14968 12222 15020
rect 16117 15011 16175 15017
rect 16117 14977 16129 15011
rect 16163 15008 16175 15011
rect 16206 15008 16212 15020
rect 16163 14980 16212 15008
rect 16163 14977 16175 14980
rect 16117 14971 16175 14977
rect 16206 14968 16212 14980
rect 16264 14968 16270 15020
rect 16301 15011 16359 15017
rect 16301 14977 16313 15011
rect 16347 15008 16359 15011
rect 16666 15008 16672 15020
rect 16347 14980 16672 15008
rect 16347 14977 16359 14980
rect 16301 14971 16359 14977
rect 16666 14968 16672 14980
rect 16724 14968 16730 15020
rect 17037 15011 17095 15017
rect 17037 14977 17049 15011
rect 17083 14977 17095 15011
rect 17037 14971 17095 14977
rect 17405 15011 17463 15017
rect 17405 14977 17417 15011
rect 17451 15008 17463 15011
rect 18064 15008 18092 15048
rect 19978 15036 19984 15048
rect 20036 15036 20042 15088
rect 22480 15048 23428 15076
rect 22480 15020 22508 15048
rect 18230 15008 18236 15020
rect 17451 14980 18092 15008
rect 18191 14980 18236 15008
rect 17451 14977 17463 14980
rect 17405 14971 17463 14977
rect 10520 14912 10824 14940
rect 11149 14943 11207 14949
rect 10413 14903 10471 14909
rect 11149 14909 11161 14943
rect 11195 14940 11207 14943
rect 12066 14940 12072 14952
rect 11195 14912 12072 14940
rect 11195 14909 11207 14912
rect 11149 14903 11207 14909
rect 3467 14844 4200 14872
rect 10428 14872 10456 14903
rect 12066 14900 12072 14912
rect 12124 14900 12130 14952
rect 16224 14940 16252 14968
rect 17052 14940 17080 14971
rect 18230 14968 18236 14980
rect 18288 14968 18294 15020
rect 18506 14968 18512 15020
rect 18564 15008 18570 15020
rect 19794 15008 19800 15020
rect 18564 14980 19800 15008
rect 18564 14968 18570 14980
rect 19794 14968 19800 14980
rect 19852 14968 19858 15020
rect 20441 15011 20499 15017
rect 20441 15008 20453 15011
rect 20089 14980 20453 15008
rect 16224 14912 17080 14940
rect 17218 14900 17224 14952
rect 17276 14940 17282 14952
rect 19886 14940 19892 14952
rect 17276 14912 19892 14940
rect 17276 14900 17282 14912
rect 19886 14900 19892 14912
rect 19944 14900 19950 14952
rect 13446 14872 13452 14884
rect 10428 14844 13452 14872
rect 3467 14841 3479 14844
rect 3421 14835 3479 14841
rect 13446 14832 13452 14844
rect 13504 14832 13510 14884
rect 15102 14832 15108 14884
rect 15160 14872 15166 14884
rect 20089 14872 20117 14980
rect 20441 14977 20453 14980
rect 20487 14977 20499 15011
rect 22186 15008 22192 15020
rect 22147 14980 22192 15008
rect 20441 14971 20499 14977
rect 22186 14968 22192 14980
rect 22244 14968 22250 15020
rect 22370 15008 22376 15020
rect 22331 14980 22376 15008
rect 22370 14968 22376 14980
rect 22428 14968 22434 15020
rect 22462 14968 22468 15020
rect 22520 15008 22526 15020
rect 22520 14980 22565 15008
rect 22520 14968 22526 14980
rect 23014 14968 23020 15020
rect 23072 15008 23078 15020
rect 23400 15017 23428 15048
rect 26142 15036 26148 15088
rect 26200 15076 26206 15088
rect 29917 15079 29975 15085
rect 29917 15076 29929 15079
rect 26200 15048 29929 15076
rect 26200 15036 26206 15048
rect 29917 15045 29929 15048
rect 29963 15045 29975 15079
rect 29917 15039 29975 15045
rect 23109 15011 23167 15017
rect 23109 15008 23121 15011
rect 23072 14980 23121 15008
rect 23072 14968 23078 14980
rect 23109 14977 23121 14980
rect 23155 14977 23167 15011
rect 23109 14971 23167 14977
rect 23385 15011 23443 15017
rect 23385 14977 23397 15011
rect 23431 14977 23443 15011
rect 25038 15008 25044 15020
rect 25096 15017 25102 15020
rect 25008 14980 25044 15008
rect 23385 14971 23443 14977
rect 25038 14968 25044 14980
rect 25096 14971 25108 15017
rect 25096 14968 25102 14971
rect 30006 14968 30012 15020
rect 30064 15008 30070 15020
rect 32309 15011 32367 15017
rect 32309 15008 32321 15011
rect 30064 14980 32321 15008
rect 30064 14968 30070 14980
rect 32309 14977 32321 14980
rect 32355 14977 32367 15011
rect 32309 14971 32367 14977
rect 20714 14940 20720 14952
rect 20675 14912 20720 14940
rect 20714 14900 20720 14912
rect 20772 14940 20778 14952
rect 21910 14940 21916 14952
rect 20772 14912 21916 14940
rect 20772 14900 20778 14912
rect 21910 14900 21916 14912
rect 21968 14900 21974 14952
rect 25317 14943 25375 14949
rect 25317 14909 25329 14943
rect 25363 14940 25375 14943
rect 26418 14940 26424 14952
rect 25363 14912 26424 14940
rect 25363 14909 25375 14912
rect 25317 14903 25375 14909
rect 26418 14900 26424 14912
rect 26476 14900 26482 14952
rect 15160 14844 20117 14872
rect 15160 14832 15166 14844
rect 29638 14832 29644 14884
rect 29696 14872 29702 14884
rect 29733 14875 29791 14881
rect 29733 14872 29745 14875
rect 29696 14844 29745 14872
rect 29696 14832 29702 14844
rect 29733 14841 29745 14844
rect 29779 14841 29791 14875
rect 29733 14835 29791 14841
rect 2958 14764 2964 14816
rect 3016 14804 3022 14816
rect 5261 14807 5319 14813
rect 5261 14804 5273 14807
rect 3016 14776 5273 14804
rect 3016 14764 3022 14776
rect 5261 14773 5273 14776
rect 5307 14773 5319 14807
rect 5261 14767 5319 14773
rect 5445 14807 5503 14813
rect 5445 14773 5457 14807
rect 5491 14804 5503 14807
rect 6086 14804 6092 14816
rect 5491 14776 6092 14804
rect 5491 14773 5503 14776
rect 5445 14767 5503 14773
rect 6086 14764 6092 14776
rect 6144 14764 6150 14816
rect 9950 14764 9956 14816
rect 10008 14804 10014 14816
rect 10686 14804 10692 14816
rect 10008 14776 10692 14804
rect 10008 14764 10014 14776
rect 10686 14764 10692 14776
rect 10744 14764 10750 14816
rect 19886 14764 19892 14816
rect 19944 14804 19950 14816
rect 22005 14807 22063 14813
rect 22005 14804 22017 14807
rect 19944 14776 22017 14804
rect 19944 14764 19950 14776
rect 22005 14773 22017 14776
rect 22051 14773 22063 14807
rect 22005 14767 22063 14773
rect 23658 14764 23664 14816
rect 23716 14804 23722 14816
rect 23937 14807 23995 14813
rect 23937 14804 23949 14807
rect 23716 14776 23949 14804
rect 23716 14764 23722 14776
rect 23937 14773 23949 14776
rect 23983 14773 23995 14807
rect 23937 14767 23995 14773
rect 1104 14714 34868 14736
rect 1104 14662 5170 14714
rect 5222 14662 5234 14714
rect 5286 14662 5298 14714
rect 5350 14662 5362 14714
rect 5414 14662 5426 14714
rect 5478 14662 13611 14714
rect 13663 14662 13675 14714
rect 13727 14662 13739 14714
rect 13791 14662 13803 14714
rect 13855 14662 13867 14714
rect 13919 14662 22052 14714
rect 22104 14662 22116 14714
rect 22168 14662 22180 14714
rect 22232 14662 22244 14714
rect 22296 14662 22308 14714
rect 22360 14662 30493 14714
rect 30545 14662 30557 14714
rect 30609 14662 30621 14714
rect 30673 14662 30685 14714
rect 30737 14662 30749 14714
rect 30801 14662 34868 14714
rect 1104 14640 34868 14662
rect 6181 14603 6239 14609
rect 6181 14569 6193 14603
rect 6227 14600 6239 14603
rect 6822 14600 6828 14612
rect 6227 14572 6828 14600
rect 6227 14569 6239 14572
rect 6181 14563 6239 14569
rect 6822 14560 6828 14572
rect 6880 14560 6886 14612
rect 7193 14603 7251 14609
rect 7193 14569 7205 14603
rect 7239 14600 7251 14603
rect 7374 14600 7380 14612
rect 7239 14572 7380 14600
rect 7239 14569 7251 14572
rect 7193 14563 7251 14569
rect 2746 14504 6224 14532
rect 1394 14424 1400 14476
rect 1452 14464 1458 14476
rect 2746 14464 2774 14504
rect 1452 14436 2774 14464
rect 6196 14464 6224 14504
rect 6270 14492 6276 14544
rect 6328 14532 6334 14544
rect 7208 14532 7236 14563
rect 7374 14560 7380 14572
rect 7432 14560 7438 14612
rect 14366 14600 14372 14612
rect 14327 14572 14372 14600
rect 14366 14560 14372 14572
rect 14424 14560 14430 14612
rect 19978 14600 19984 14612
rect 19628 14572 19984 14600
rect 6328 14504 7236 14532
rect 8481 14535 8539 14541
rect 6328 14492 6334 14504
rect 8481 14501 8493 14535
rect 8527 14532 8539 14535
rect 8662 14532 8668 14544
rect 8527 14504 8668 14532
rect 8527 14501 8539 14504
rect 8481 14495 8539 14501
rect 8662 14492 8668 14504
rect 8720 14492 8726 14544
rect 9214 14532 9220 14544
rect 9175 14504 9220 14532
rect 9214 14492 9220 14504
rect 9272 14492 9278 14544
rect 12728 14504 15608 14532
rect 12728 14464 12756 14504
rect 6196 14436 12756 14464
rect 12820 14436 14320 14464
rect 1452 14424 1458 14436
rect 2682 14396 2688 14408
rect 2643 14368 2688 14396
rect 2682 14356 2688 14368
rect 2740 14356 2746 14408
rect 2869 14399 2927 14405
rect 2869 14365 2881 14399
rect 2915 14396 2927 14399
rect 3050 14396 3056 14408
rect 2915 14368 3056 14396
rect 2915 14365 2927 14368
rect 2869 14359 2927 14365
rect 3050 14356 3056 14368
rect 3108 14356 3114 14408
rect 6089 14399 6147 14405
rect 6089 14365 6101 14399
rect 6135 14396 6147 14399
rect 6270 14396 6276 14408
rect 6135 14368 6276 14396
rect 6135 14365 6147 14368
rect 6089 14359 6147 14365
rect 6270 14356 6276 14368
rect 6328 14356 6334 14408
rect 6365 14399 6423 14405
rect 6365 14365 6377 14399
rect 6411 14365 6423 14399
rect 9582 14396 9588 14408
rect 6365 14359 6423 14365
rect 8220 14368 9588 14396
rect 2961 14331 3019 14337
rect 2961 14297 2973 14331
rect 3007 14328 3019 14331
rect 3142 14328 3148 14340
rect 3007 14300 3148 14328
rect 3007 14297 3019 14300
rect 2961 14291 3019 14297
rect 3142 14288 3148 14300
rect 3200 14288 3206 14340
rect 5718 14288 5724 14340
rect 5776 14328 5782 14340
rect 6380 14328 6408 14359
rect 6454 14328 6460 14340
rect 5776 14300 6460 14328
rect 5776 14288 5782 14300
rect 6454 14288 6460 14300
rect 6512 14328 6518 14340
rect 7009 14331 7067 14337
rect 7009 14328 7021 14331
rect 6512 14300 7021 14328
rect 6512 14288 6518 14300
rect 7009 14297 7021 14300
rect 7055 14297 7067 14331
rect 7926 14328 7932 14340
rect 7887 14300 7932 14328
rect 7009 14291 7067 14297
rect 7926 14288 7932 14300
rect 7984 14328 7990 14340
rect 8220 14337 8248 14368
rect 9582 14356 9588 14368
rect 9640 14356 9646 14408
rect 10226 14396 10232 14408
rect 9692 14368 10232 14396
rect 8205 14331 8263 14337
rect 7984 14300 8156 14328
rect 7984 14288 7990 14300
rect 6549 14263 6607 14269
rect 6549 14229 6561 14263
rect 6595 14260 6607 14263
rect 6914 14260 6920 14272
rect 6595 14232 6920 14260
rect 6595 14229 6607 14232
rect 6549 14223 6607 14229
rect 6914 14220 6920 14232
rect 6972 14220 6978 14272
rect 7190 14220 7196 14272
rect 7248 14269 7254 14272
rect 7248 14263 7267 14269
rect 7255 14229 7267 14263
rect 7248 14223 7267 14229
rect 7377 14263 7435 14269
rect 7377 14229 7389 14263
rect 7423 14260 7435 14263
rect 7742 14260 7748 14272
rect 7423 14232 7748 14260
rect 7423 14229 7435 14232
rect 7377 14223 7435 14229
rect 7248 14220 7254 14223
rect 7742 14220 7748 14232
rect 7800 14220 7806 14272
rect 7834 14220 7840 14272
rect 7892 14260 7898 14272
rect 8021 14263 8079 14269
rect 8021 14260 8033 14263
rect 7892 14232 8033 14260
rect 7892 14220 7898 14232
rect 8021 14229 8033 14232
rect 8067 14229 8079 14263
rect 8128 14260 8156 14300
rect 8205 14297 8217 14331
rect 8251 14297 8263 14331
rect 8205 14291 8263 14297
rect 8294 14288 8300 14340
rect 8352 14328 8358 14340
rect 9692 14337 9720 14368
rect 10226 14356 10232 14368
rect 10284 14356 10290 14408
rect 11974 14356 11980 14408
rect 12032 14396 12038 14408
rect 12820 14405 12848 14436
rect 14292 14405 14320 14436
rect 15580 14405 15608 14504
rect 18506 14464 18512 14476
rect 18467 14436 18512 14464
rect 18506 14424 18512 14436
rect 18564 14424 18570 14476
rect 19628 14473 19656 14572
rect 19978 14560 19984 14572
rect 20036 14560 20042 14612
rect 21726 14560 21732 14612
rect 21784 14600 21790 14612
rect 23658 14600 23664 14612
rect 21784 14572 23664 14600
rect 21784 14560 21790 14572
rect 23658 14560 23664 14572
rect 23716 14560 23722 14612
rect 23753 14603 23811 14609
rect 23753 14569 23765 14603
rect 23799 14569 23811 14603
rect 23753 14563 23811 14569
rect 23937 14603 23995 14609
rect 23937 14569 23949 14603
rect 23983 14600 23995 14603
rect 25222 14600 25228 14612
rect 23983 14572 25228 14600
rect 23983 14569 23995 14572
rect 23937 14563 23995 14569
rect 20993 14535 21051 14541
rect 20993 14501 21005 14535
rect 21039 14532 21051 14535
rect 21039 14504 22048 14532
rect 21039 14501 21051 14504
rect 20993 14495 21051 14501
rect 19613 14467 19671 14473
rect 19613 14433 19625 14467
rect 19659 14433 19671 14467
rect 19613 14427 19671 14433
rect 12805 14399 12863 14405
rect 12805 14396 12817 14399
rect 12032 14368 12817 14396
rect 12032 14356 12038 14368
rect 12805 14365 12817 14368
rect 12851 14365 12863 14399
rect 12805 14359 12863 14365
rect 12897 14399 12955 14405
rect 12897 14365 12909 14399
rect 12943 14396 12955 14399
rect 14277 14399 14335 14405
rect 12943 14368 14044 14396
rect 12943 14365 12955 14368
rect 12897 14359 12955 14365
rect 9493 14331 9551 14337
rect 9493 14328 9505 14331
rect 8352 14300 9505 14328
rect 8352 14288 8358 14300
rect 9493 14297 9505 14300
rect 9539 14297 9551 14331
rect 9493 14291 9551 14297
rect 9677 14331 9735 14337
rect 9677 14297 9689 14331
rect 9723 14297 9735 14331
rect 9677 14291 9735 14297
rect 9769 14331 9827 14337
rect 9769 14297 9781 14331
rect 9815 14328 9827 14331
rect 9950 14328 9956 14340
rect 9815 14300 9956 14328
rect 9815 14297 9827 14300
rect 9769 14291 9827 14297
rect 9784 14260 9812 14291
rect 9950 14288 9956 14300
rect 10008 14288 10014 14340
rect 11698 14288 11704 14340
rect 11756 14328 11762 14340
rect 12434 14328 12440 14340
rect 11756 14300 12440 14328
rect 11756 14288 11762 14300
rect 12434 14288 12440 14300
rect 12492 14328 12498 14340
rect 12912 14328 12940 14359
rect 13078 14328 13084 14340
rect 12492 14300 12940 14328
rect 13039 14300 13084 14328
rect 12492 14288 12498 14300
rect 13078 14288 13084 14300
rect 13136 14288 13142 14340
rect 14016 14328 14044 14368
rect 14277 14365 14289 14399
rect 14323 14365 14335 14399
rect 14277 14359 14335 14365
rect 14461 14399 14519 14405
rect 14461 14365 14473 14399
rect 14507 14365 14519 14399
rect 14461 14359 14519 14365
rect 15565 14399 15623 14405
rect 15565 14365 15577 14399
rect 15611 14365 15623 14399
rect 15565 14359 15623 14365
rect 14476 14328 14504 14359
rect 17402 14356 17408 14408
rect 17460 14396 17466 14408
rect 17773 14399 17831 14405
rect 17773 14396 17785 14399
rect 17460 14368 17785 14396
rect 17460 14356 17466 14368
rect 17773 14365 17785 14368
rect 17819 14365 17831 14399
rect 17773 14359 17831 14365
rect 17862 14356 17868 14408
rect 17920 14396 17926 14408
rect 18233 14399 18291 14405
rect 18233 14396 18245 14399
rect 17920 14368 18245 14396
rect 17920 14356 17926 14368
rect 18233 14365 18245 14368
rect 18279 14365 18291 14399
rect 21634 14396 21640 14408
rect 21595 14368 21640 14396
rect 18233 14359 18291 14365
rect 21634 14356 21640 14368
rect 21692 14356 21698 14408
rect 21726 14356 21732 14408
rect 21784 14396 21790 14408
rect 22020 14405 22048 14504
rect 22094 14492 22100 14544
rect 22152 14532 22158 14544
rect 23768 14532 23796 14563
rect 25222 14560 25228 14572
rect 25280 14560 25286 14612
rect 25958 14600 25964 14612
rect 25919 14572 25964 14600
rect 25958 14560 25964 14572
rect 26016 14560 26022 14612
rect 26694 14560 26700 14612
rect 26752 14600 26758 14612
rect 28721 14603 28779 14609
rect 28721 14600 28733 14603
rect 26752 14572 28733 14600
rect 26752 14560 26758 14572
rect 28721 14569 28733 14572
rect 28767 14569 28779 14603
rect 32490 14600 32496 14612
rect 28721 14563 28779 14569
rect 29656 14572 32496 14600
rect 22152 14504 23796 14532
rect 22152 14492 22158 14504
rect 23750 14464 23756 14476
rect 22940 14436 23756 14464
rect 22005 14399 22063 14405
rect 21784 14368 21829 14396
rect 21784 14356 21790 14368
rect 22005 14365 22017 14399
rect 22051 14396 22063 14399
rect 22370 14396 22376 14408
rect 22051 14368 22376 14396
rect 22051 14365 22063 14368
rect 22005 14359 22063 14365
rect 22370 14356 22376 14368
rect 22428 14356 22434 14408
rect 19886 14337 19892 14340
rect 14016 14300 14504 14328
rect 17313 14331 17371 14337
rect 17313 14297 17325 14331
rect 17359 14328 17371 14331
rect 19880 14328 19892 14337
rect 17359 14300 18000 14328
rect 19847 14300 19892 14328
rect 17359 14297 17371 14300
rect 17313 14291 17371 14297
rect 8128 14232 9812 14260
rect 8021 14223 8079 14229
rect 9858 14220 9864 14272
rect 9916 14260 9922 14272
rect 17328 14260 17356 14291
rect 9916 14232 17356 14260
rect 17972 14260 18000 14300
rect 19880 14291 19892 14300
rect 19886 14288 19892 14291
rect 19944 14288 19950 14340
rect 20622 14288 20628 14340
rect 20680 14328 20686 14340
rect 21818 14328 21824 14340
rect 20680 14300 20944 14328
rect 21779 14300 21824 14328
rect 20680 14288 20686 14300
rect 20806 14260 20812 14272
rect 17972 14232 20812 14260
rect 9916 14220 9922 14232
rect 20806 14220 20812 14232
rect 20864 14220 20870 14272
rect 20916 14260 20944 14300
rect 21818 14288 21824 14300
rect 21876 14328 21882 14340
rect 22940 14328 22968 14436
rect 23750 14424 23756 14436
rect 23808 14424 23814 14476
rect 24578 14464 24584 14476
rect 24539 14436 24584 14464
rect 24578 14424 24584 14436
rect 24636 14424 24642 14476
rect 23474 14356 23480 14408
rect 23532 14396 23538 14408
rect 24837 14399 24895 14405
rect 24837 14396 24849 14399
rect 23532 14368 24849 14396
rect 23532 14356 23538 14368
rect 24837 14365 24849 14368
rect 24883 14365 24895 14399
rect 26418 14396 26424 14408
rect 26331 14368 26424 14396
rect 24837 14359 24895 14365
rect 26418 14356 26424 14368
rect 26476 14396 26482 14408
rect 26970 14396 26976 14408
rect 26476 14368 26976 14396
rect 26476 14356 26482 14368
rect 26970 14356 26976 14368
rect 27028 14356 27034 14408
rect 27706 14356 27712 14408
rect 27764 14396 27770 14408
rect 28261 14399 28319 14405
rect 28261 14396 28273 14399
rect 27764 14368 28273 14396
rect 27764 14356 27770 14368
rect 28261 14365 28273 14368
rect 28307 14365 28319 14399
rect 28261 14359 28319 14365
rect 28537 14399 28595 14405
rect 28537 14365 28549 14399
rect 28583 14396 28595 14399
rect 28626 14396 28632 14408
rect 28583 14368 28632 14396
rect 28583 14365 28595 14368
rect 28537 14359 28595 14365
rect 28626 14356 28632 14368
rect 28684 14396 28690 14408
rect 29656 14396 29684 14572
rect 32490 14560 32496 14572
rect 32548 14560 32554 14612
rect 31389 14467 31447 14473
rect 31389 14433 31401 14467
rect 31435 14464 31447 14467
rect 31754 14464 31760 14476
rect 31435 14436 31760 14464
rect 31435 14433 31447 14436
rect 31389 14427 31447 14433
rect 31754 14424 31760 14436
rect 31812 14424 31818 14476
rect 31849 14467 31907 14473
rect 31849 14433 31861 14467
rect 31895 14464 31907 14467
rect 32306 14464 32312 14476
rect 31895 14436 32312 14464
rect 31895 14433 31907 14436
rect 31849 14427 31907 14433
rect 32306 14424 32312 14436
rect 32364 14424 32370 14476
rect 28684 14368 29684 14396
rect 28684 14356 28690 14368
rect 30098 14356 30104 14408
rect 30156 14396 30162 14408
rect 31113 14399 31171 14405
rect 31113 14396 31125 14399
rect 30156 14368 31125 14396
rect 30156 14356 30162 14368
rect 31113 14365 31125 14368
rect 31159 14365 31171 14399
rect 32122 14396 32128 14408
rect 32083 14368 32128 14396
rect 31113 14359 31171 14365
rect 32122 14356 32128 14368
rect 32180 14356 32186 14408
rect 23566 14328 23572 14340
rect 21876 14300 22968 14328
rect 23527 14300 23572 14328
rect 21876 14288 21882 14300
rect 23566 14288 23572 14300
rect 23624 14288 23630 14340
rect 26694 14337 26700 14340
rect 26688 14328 26700 14337
rect 26655 14300 26700 14328
rect 26688 14291 26700 14300
rect 26694 14288 26700 14291
rect 26752 14288 26758 14340
rect 27614 14288 27620 14340
rect 27672 14328 27678 14340
rect 29086 14328 29092 14340
rect 27672 14300 29092 14328
rect 27672 14288 27678 14300
rect 29086 14288 29092 14300
rect 29144 14288 29150 14340
rect 29730 14328 29736 14340
rect 29691 14300 29736 14328
rect 29730 14288 29736 14300
rect 29788 14288 29794 14340
rect 21453 14263 21511 14269
rect 21453 14260 21465 14263
rect 20916 14232 21465 14260
rect 21453 14229 21465 14232
rect 21499 14229 21511 14263
rect 21453 14223 21511 14229
rect 23753 14263 23811 14269
rect 23753 14229 23765 14263
rect 23799 14260 23811 14263
rect 24026 14260 24032 14272
rect 23799 14232 24032 14260
rect 23799 14229 23811 14232
rect 23753 14223 23811 14229
rect 24026 14220 24032 14232
rect 24084 14220 24090 14272
rect 27706 14220 27712 14272
rect 27764 14260 27770 14272
rect 27801 14263 27859 14269
rect 27801 14260 27813 14263
rect 27764 14232 27813 14260
rect 27764 14220 27770 14232
rect 27801 14229 27813 14232
rect 27847 14260 27859 14263
rect 28353 14263 28411 14269
rect 28353 14260 28365 14263
rect 27847 14232 28365 14260
rect 27847 14229 27859 14232
rect 27801 14223 27859 14229
rect 28353 14229 28365 14232
rect 28399 14229 28411 14263
rect 28353 14223 28411 14229
rect 28994 14220 29000 14272
rect 29052 14260 29058 14272
rect 29914 14260 29920 14272
rect 29052 14232 29920 14260
rect 29052 14220 29058 14232
rect 29914 14220 29920 14232
rect 29972 14220 29978 14272
rect 31294 14220 31300 14272
rect 31352 14260 31358 14272
rect 33042 14260 33048 14272
rect 31352 14232 33048 14260
rect 31352 14220 31358 14232
rect 33042 14220 33048 14232
rect 33100 14260 33106 14272
rect 33229 14263 33287 14269
rect 33229 14260 33241 14263
rect 33100 14232 33241 14260
rect 33100 14220 33106 14232
rect 33229 14229 33241 14232
rect 33275 14229 33287 14263
rect 33229 14223 33287 14229
rect 1104 14170 35027 14192
rect 1104 14118 9390 14170
rect 9442 14118 9454 14170
rect 9506 14118 9518 14170
rect 9570 14118 9582 14170
rect 9634 14118 9646 14170
rect 9698 14118 17831 14170
rect 17883 14118 17895 14170
rect 17947 14118 17959 14170
rect 18011 14118 18023 14170
rect 18075 14118 18087 14170
rect 18139 14118 26272 14170
rect 26324 14118 26336 14170
rect 26388 14118 26400 14170
rect 26452 14118 26464 14170
rect 26516 14118 26528 14170
rect 26580 14118 34713 14170
rect 34765 14118 34777 14170
rect 34829 14118 34841 14170
rect 34893 14118 34905 14170
rect 34957 14118 34969 14170
rect 35021 14118 35027 14170
rect 1104 14096 35027 14118
rect 1670 14016 1676 14068
rect 1728 14056 1734 14068
rect 2593 14059 2651 14065
rect 2593 14056 2605 14059
rect 1728 14028 2605 14056
rect 1728 14016 1734 14028
rect 2593 14025 2605 14028
rect 2639 14025 2651 14059
rect 2593 14019 2651 14025
rect 3142 14016 3148 14068
rect 3200 14056 3206 14068
rect 5905 14059 5963 14065
rect 3200 14028 5764 14056
rect 3200 14016 3206 14028
rect 4430 13988 4436 14000
rect 4391 13960 4436 13988
rect 4430 13948 4436 13960
rect 4488 13948 4494 14000
rect 2685 13923 2743 13929
rect 2685 13889 2697 13923
rect 2731 13920 2743 13923
rect 3050 13920 3056 13932
rect 2731 13892 3056 13920
rect 2731 13889 2743 13892
rect 2685 13883 2743 13889
rect 3050 13880 3056 13892
rect 3108 13880 3114 13932
rect 5534 13880 5540 13932
rect 5592 13880 5598 13932
rect 5736 13920 5764 14028
rect 5905 14025 5917 14059
rect 5951 14056 5963 14059
rect 7926 14056 7932 14068
rect 5951 14028 7932 14056
rect 5951 14025 5963 14028
rect 5905 14019 5963 14025
rect 7926 14016 7932 14028
rect 7984 14016 7990 14068
rect 8294 14056 8300 14068
rect 8207 14028 8300 14056
rect 8294 14016 8300 14028
rect 8352 14056 8358 14068
rect 8352 14028 10180 14056
rect 8352 14016 8358 14028
rect 6454 13948 6460 14000
rect 6512 13988 6518 14000
rect 6549 13991 6607 13997
rect 6549 13988 6561 13991
rect 6512 13960 6561 13988
rect 6512 13948 6518 13960
rect 6549 13957 6561 13960
rect 6595 13957 6607 13991
rect 6549 13951 6607 13957
rect 6733 13991 6791 13997
rect 6733 13957 6745 13991
rect 6779 13988 6791 13991
rect 7190 13988 7196 14000
rect 6779 13960 7196 13988
rect 6779 13957 6791 13960
rect 6733 13951 6791 13957
rect 6748 13920 6776 13951
rect 7190 13948 7196 13960
rect 7248 13988 7254 14000
rect 7466 13988 7472 14000
rect 7248 13960 7472 13988
rect 7248 13948 7254 13960
rect 7466 13948 7472 13960
rect 7524 13948 7530 14000
rect 9306 13948 9312 14000
rect 9364 13988 9370 14000
rect 9585 13991 9643 13997
rect 9585 13988 9597 13991
rect 9364 13960 9597 13988
rect 9364 13948 9370 13960
rect 9585 13957 9597 13960
rect 9631 13988 9643 13991
rect 9858 13988 9864 14000
rect 9631 13960 9864 13988
rect 9631 13957 9643 13960
rect 9585 13951 9643 13957
rect 9858 13948 9864 13960
rect 9916 13948 9922 14000
rect 10152 13988 10180 14028
rect 11054 14016 11060 14068
rect 11112 14056 11118 14068
rect 11790 14056 11796 14068
rect 11112 14028 11796 14056
rect 11112 14016 11118 14028
rect 11790 14016 11796 14028
rect 11848 14056 11854 14068
rect 20717 14059 20775 14065
rect 11848 14028 12112 14056
rect 11848 14016 11854 14028
rect 11974 13988 11980 14000
rect 10152 13960 11980 13988
rect 5736 13892 6776 13920
rect 7009 13923 7067 13929
rect 7009 13889 7021 13923
rect 7055 13920 7067 13923
rect 8386 13920 8392 13932
rect 7055 13892 8392 13920
rect 7055 13889 7067 13892
rect 7009 13883 7067 13889
rect 8386 13880 8392 13892
rect 8444 13880 8450 13932
rect 10152 13929 10180 13960
rect 11974 13948 11980 13960
rect 12032 13948 12038 14000
rect 12084 13997 12112 14028
rect 20717 14025 20729 14059
rect 20763 14056 20775 14059
rect 22370 14056 22376 14068
rect 20763 14028 22376 14056
rect 20763 14025 20775 14028
rect 20717 14019 20775 14025
rect 22370 14016 22376 14028
rect 22428 14016 22434 14068
rect 23658 14016 23664 14068
rect 23716 14056 23722 14068
rect 24673 14059 24731 14065
rect 24673 14056 24685 14059
rect 23716 14028 24685 14056
rect 23716 14016 23722 14028
rect 24673 14025 24685 14028
rect 24719 14025 24731 14059
rect 25038 14056 25044 14068
rect 24999 14028 25044 14056
rect 24673 14019 24731 14025
rect 25038 14016 25044 14028
rect 25096 14016 25102 14068
rect 27798 14016 27804 14068
rect 27856 14056 27862 14068
rect 28905 14059 28963 14065
rect 28905 14056 28917 14059
rect 27856 14028 28917 14056
rect 27856 14016 27862 14028
rect 28905 14025 28917 14028
rect 28951 14025 28963 14059
rect 28905 14019 28963 14025
rect 29089 14059 29147 14065
rect 29089 14025 29101 14059
rect 29135 14056 29147 14059
rect 30006 14056 30012 14068
rect 29135 14028 30012 14056
rect 29135 14025 29147 14028
rect 29089 14019 29147 14025
rect 30006 14016 30012 14028
rect 30064 14016 30070 14068
rect 30098 14016 30104 14068
rect 30156 14056 30162 14068
rect 31389 14059 31447 14065
rect 30156 14028 30201 14056
rect 30156 14016 30162 14028
rect 31389 14025 31401 14059
rect 31435 14056 31447 14059
rect 32582 14056 32588 14068
rect 31435 14028 32588 14056
rect 31435 14025 31447 14028
rect 31389 14019 31447 14025
rect 32582 14016 32588 14028
rect 32640 14056 32646 14068
rect 33689 14059 33747 14065
rect 33689 14056 33701 14059
rect 32640 14028 33701 14056
rect 32640 14016 32646 14028
rect 33689 14025 33701 14028
rect 33735 14025 33747 14059
rect 33689 14019 33747 14025
rect 12069 13991 12127 13997
rect 12069 13957 12081 13991
rect 12115 13957 12127 13991
rect 12069 13951 12127 13957
rect 13078 13948 13084 14000
rect 13136 13948 13142 14000
rect 14645 13991 14703 13997
rect 14645 13957 14657 13991
rect 14691 13988 14703 13991
rect 16666 13988 16672 14000
rect 14691 13960 16672 13988
rect 14691 13957 14703 13960
rect 14645 13951 14703 13957
rect 16666 13948 16672 13960
rect 16724 13988 16730 14000
rect 17586 13988 17592 14000
rect 16724 13960 17592 13988
rect 16724 13948 16730 13960
rect 10137 13923 10195 13929
rect 10137 13889 10149 13923
rect 10183 13889 10195 13923
rect 10137 13883 10195 13889
rect 10229 13923 10287 13929
rect 10229 13889 10241 13923
rect 10275 13920 10287 13923
rect 11698 13920 11704 13932
rect 10275 13892 11704 13920
rect 10275 13889 10287 13892
rect 10229 13883 10287 13889
rect 4154 13852 4160 13864
rect 4115 13824 4160 13852
rect 4154 13812 4160 13824
rect 4212 13812 4218 13864
rect 5074 13852 5080 13864
rect 4264 13824 5080 13852
rect 4062 13744 4068 13796
rect 4120 13784 4126 13796
rect 4264 13784 4292 13824
rect 5074 13812 5080 13824
rect 5132 13852 5138 13864
rect 10244 13852 10272 13883
rect 11698 13880 11704 13892
rect 11756 13880 11762 13932
rect 13998 13880 14004 13932
rect 14056 13920 14062 13932
rect 14093 13923 14151 13929
rect 14093 13920 14105 13923
rect 14056 13892 14105 13920
rect 14056 13880 14062 13892
rect 14093 13889 14105 13892
rect 14139 13889 14151 13923
rect 14093 13883 14151 13889
rect 14277 13923 14335 13929
rect 14277 13889 14289 13923
rect 14323 13920 14335 13923
rect 14550 13920 14556 13932
rect 14323 13892 14556 13920
rect 14323 13889 14335 13892
rect 14277 13883 14335 13889
rect 14550 13880 14556 13892
rect 14608 13880 14614 13932
rect 15194 13920 15200 13932
rect 15155 13892 15200 13920
rect 15194 13880 15200 13892
rect 15252 13880 15258 13932
rect 15562 13920 15568 13932
rect 15523 13892 15568 13920
rect 15562 13880 15568 13892
rect 15620 13880 15626 13932
rect 17144 13929 17172 13960
rect 17586 13948 17592 13960
rect 17644 13948 17650 14000
rect 19429 13991 19487 13997
rect 19429 13957 19441 13991
rect 19475 13988 19487 13991
rect 19518 13988 19524 14000
rect 19475 13960 19524 13988
rect 19475 13957 19487 13960
rect 19429 13951 19487 13957
rect 19518 13948 19524 13960
rect 19576 13948 19582 14000
rect 19610 13948 19616 14000
rect 19668 13988 19674 14000
rect 21818 13988 21824 14000
rect 19668 13960 21824 13988
rect 19668 13948 19674 13960
rect 21818 13948 21824 13960
rect 21876 13948 21882 14000
rect 27614 13948 27620 14000
rect 27672 13988 27678 14000
rect 28718 13988 28724 14000
rect 27672 13960 27717 13988
rect 28679 13960 28724 13988
rect 27672 13948 27678 13960
rect 28718 13948 28724 13960
rect 28776 13948 28782 14000
rect 29656 13960 31708 13988
rect 29656 13932 29684 13960
rect 17129 13923 17187 13929
rect 17129 13889 17141 13923
rect 17175 13889 17187 13923
rect 17310 13920 17316 13932
rect 17271 13892 17316 13920
rect 17129 13883 17187 13889
rect 17310 13880 17316 13892
rect 17368 13880 17374 13932
rect 20530 13920 20536 13932
rect 20491 13892 20536 13920
rect 20530 13880 20536 13892
rect 20588 13880 20594 13932
rect 21634 13880 21640 13932
rect 21692 13920 21698 13932
rect 24026 13920 24032 13932
rect 21692 13892 24032 13920
rect 21692 13880 21698 13892
rect 24026 13880 24032 13892
rect 24084 13880 24090 13932
rect 24486 13880 24492 13932
rect 24544 13920 24550 13932
rect 24581 13923 24639 13929
rect 24581 13920 24593 13923
rect 24544 13892 24593 13920
rect 24544 13880 24550 13892
rect 24581 13889 24593 13892
rect 24627 13889 24639 13923
rect 24581 13883 24639 13889
rect 24857 13923 24915 13929
rect 24857 13889 24869 13923
rect 24903 13889 24915 13923
rect 24857 13883 24915 13889
rect 11790 13852 11796 13864
rect 5132 13824 10272 13852
rect 11751 13824 11796 13852
rect 5132 13812 5138 13824
rect 11790 13812 11796 13824
rect 11848 13812 11854 13864
rect 13541 13855 13599 13861
rect 13541 13821 13553 13855
rect 13587 13852 13599 13855
rect 14016 13852 14044 13880
rect 13587 13824 14044 13852
rect 17589 13855 17647 13861
rect 13587 13821 13599 13824
rect 13541 13815 13599 13821
rect 17589 13821 17601 13855
rect 17635 13852 17647 13855
rect 17678 13852 17684 13864
rect 17635 13824 17684 13852
rect 17635 13821 17647 13824
rect 17589 13815 17647 13821
rect 17678 13812 17684 13824
rect 17736 13812 17742 13864
rect 4120 13756 4292 13784
rect 15749 13787 15807 13793
rect 4120 13744 4126 13756
rect 15749 13753 15761 13787
rect 15795 13784 15807 13787
rect 16206 13784 16212 13796
rect 15795 13756 16212 13784
rect 15795 13753 15807 13756
rect 15749 13747 15807 13753
rect 16206 13744 16212 13756
rect 16264 13744 16270 13796
rect 20714 13784 20720 13796
rect 19628 13756 20720 13784
rect 6733 13719 6791 13725
rect 6733 13685 6745 13719
rect 6779 13716 6791 13719
rect 6822 13716 6828 13728
rect 6779 13688 6828 13716
rect 6779 13685 6791 13688
rect 6733 13679 6791 13685
rect 6822 13676 6828 13688
rect 6880 13676 6886 13728
rect 10134 13716 10140 13728
rect 10095 13688 10140 13716
rect 10134 13676 10140 13688
rect 10192 13676 10198 13728
rect 19518 13676 19524 13728
rect 19576 13716 19582 13728
rect 19628 13725 19656 13756
rect 20714 13744 20720 13756
rect 20772 13744 20778 13796
rect 24670 13744 24676 13796
rect 24728 13784 24734 13796
rect 24863 13784 24891 13883
rect 25038 13880 25044 13932
rect 25096 13920 25102 13932
rect 27387 13923 27445 13929
rect 27387 13920 27399 13923
rect 25096 13892 27399 13920
rect 25096 13880 25102 13892
rect 27387 13889 27399 13892
rect 27433 13889 27445 13923
rect 27387 13883 27445 13889
rect 27525 13923 27583 13929
rect 27525 13889 27537 13923
rect 27571 13889 27583 13923
rect 27525 13883 27583 13889
rect 27709 13923 27767 13929
rect 27709 13889 27721 13923
rect 27755 13920 27767 13923
rect 27798 13920 27804 13932
rect 27755 13892 27804 13920
rect 27755 13889 27767 13892
rect 27709 13883 27767 13889
rect 26694 13812 26700 13864
rect 26752 13852 26758 13864
rect 27249 13855 27307 13861
rect 27249 13852 27261 13855
rect 26752 13824 27261 13852
rect 26752 13812 26758 13824
rect 27249 13821 27261 13824
rect 27295 13821 27307 13855
rect 27540 13852 27568 13883
rect 27798 13880 27804 13892
rect 27856 13880 27862 13932
rect 29638 13920 29644 13932
rect 27908 13892 29500 13920
rect 29599 13892 29644 13920
rect 27908 13852 27936 13892
rect 29472 13852 29500 13892
rect 29638 13880 29644 13892
rect 29696 13880 29702 13932
rect 29730 13880 29736 13932
rect 29788 13920 29794 13932
rect 29788 13892 29881 13920
rect 29788 13880 29794 13892
rect 29914 13880 29920 13932
rect 29972 13920 29978 13932
rect 31312 13929 31340 13960
rect 31297 13923 31355 13929
rect 29972 13892 30017 13920
rect 29972 13880 29978 13892
rect 31297 13889 31309 13923
rect 31343 13889 31355 13923
rect 31297 13883 31355 13889
rect 31573 13923 31631 13929
rect 31573 13889 31585 13923
rect 31619 13889 31631 13923
rect 31573 13883 31631 13889
rect 29748 13852 29776 13880
rect 30282 13852 30288 13864
rect 27540 13824 27936 13852
rect 28966 13824 29408 13852
rect 29472 13824 29776 13852
rect 29840 13824 30288 13852
rect 27249 13815 27307 13821
rect 28966 13784 28994 13824
rect 24728 13756 28994 13784
rect 29380 13784 29408 13824
rect 29840 13784 29868 13824
rect 30282 13812 30288 13824
rect 30340 13852 30346 13864
rect 31588 13852 31616 13883
rect 30340 13824 31616 13852
rect 30340 13812 30346 13824
rect 29380 13756 29868 13784
rect 24728 13744 24734 13756
rect 19613 13719 19671 13725
rect 19613 13716 19625 13719
rect 19576 13688 19625 13716
rect 19576 13676 19582 13688
rect 19613 13685 19625 13688
rect 19659 13685 19671 13719
rect 19794 13716 19800 13728
rect 19755 13688 19800 13716
rect 19613 13679 19671 13685
rect 19794 13676 19800 13688
rect 19852 13676 19858 13728
rect 27893 13719 27951 13725
rect 27893 13685 27905 13719
rect 27939 13716 27951 13719
rect 28534 13716 28540 13728
rect 27939 13688 28540 13716
rect 27939 13685 27951 13688
rect 27893 13679 27951 13685
rect 28534 13676 28540 13688
rect 28592 13676 28598 13728
rect 28905 13719 28963 13725
rect 28905 13685 28917 13719
rect 28951 13716 28963 13719
rect 29454 13716 29460 13728
rect 28951 13688 29460 13716
rect 28951 13685 28963 13688
rect 28905 13679 28963 13685
rect 29454 13676 29460 13688
rect 29512 13676 29518 13728
rect 31680 13716 31708 13960
rect 31757 13923 31815 13929
rect 31757 13889 31769 13923
rect 31803 13920 31815 13923
rect 32585 13923 32643 13929
rect 32585 13920 32597 13923
rect 31803 13892 32597 13920
rect 31803 13889 31815 13892
rect 31757 13883 31815 13889
rect 32585 13889 32597 13892
rect 32631 13889 32643 13923
rect 32585 13883 32643 13889
rect 32306 13852 32312 13864
rect 32267 13824 32312 13852
rect 32306 13812 32312 13824
rect 32364 13812 32370 13864
rect 33410 13716 33416 13728
rect 31680 13688 33416 13716
rect 33410 13676 33416 13688
rect 33468 13676 33474 13728
rect 1104 13626 34868 13648
rect 1104 13574 5170 13626
rect 5222 13574 5234 13626
rect 5286 13574 5298 13626
rect 5350 13574 5362 13626
rect 5414 13574 5426 13626
rect 5478 13574 13611 13626
rect 13663 13574 13675 13626
rect 13727 13574 13739 13626
rect 13791 13574 13803 13626
rect 13855 13574 13867 13626
rect 13919 13574 22052 13626
rect 22104 13574 22116 13626
rect 22168 13574 22180 13626
rect 22232 13574 22244 13626
rect 22296 13574 22308 13626
rect 22360 13574 30493 13626
rect 30545 13574 30557 13626
rect 30609 13574 30621 13626
rect 30673 13574 30685 13626
rect 30737 13574 30749 13626
rect 30801 13574 34868 13626
rect 1104 13552 34868 13574
rect 3421 13515 3479 13521
rect 3421 13481 3433 13515
rect 3467 13512 3479 13515
rect 4154 13512 4160 13524
rect 3467 13484 4160 13512
rect 3467 13481 3479 13484
rect 3421 13475 3479 13481
rect 4154 13472 4160 13484
rect 4212 13472 4218 13524
rect 5445 13515 5503 13521
rect 5445 13481 5457 13515
rect 5491 13512 5503 13515
rect 5534 13512 5540 13524
rect 5491 13484 5540 13512
rect 5491 13481 5503 13484
rect 5445 13475 5503 13481
rect 5534 13472 5540 13484
rect 5592 13472 5598 13524
rect 12802 13512 12808 13524
rect 8496 13484 12808 13512
rect 8496 13444 8524 13484
rect 12802 13472 12808 13484
rect 12860 13512 12866 13524
rect 13262 13512 13268 13524
rect 12860 13484 13268 13512
rect 12860 13472 12866 13484
rect 13262 13472 13268 13484
rect 13320 13472 13326 13524
rect 14274 13472 14280 13524
rect 14332 13512 14338 13524
rect 14369 13515 14427 13521
rect 14369 13512 14381 13515
rect 14332 13484 14381 13512
rect 14332 13472 14338 13484
rect 14369 13481 14381 13484
rect 14415 13481 14427 13515
rect 14369 13475 14427 13481
rect 16301 13515 16359 13521
rect 16301 13481 16313 13515
rect 16347 13512 16359 13515
rect 17310 13512 17316 13524
rect 16347 13484 17316 13512
rect 16347 13481 16359 13484
rect 16301 13475 16359 13481
rect 4264 13416 8524 13444
rect 14384 13444 14412 13475
rect 17310 13472 17316 13484
rect 17368 13472 17374 13524
rect 26970 13472 26976 13524
rect 27028 13512 27034 13524
rect 27341 13515 27399 13521
rect 27341 13512 27353 13515
rect 27028 13484 27353 13512
rect 27028 13472 27034 13484
rect 27341 13481 27353 13484
rect 27387 13481 27399 13515
rect 27341 13475 27399 13481
rect 31665 13515 31723 13521
rect 31665 13481 31677 13515
rect 31711 13512 31723 13515
rect 32306 13512 32312 13524
rect 31711 13484 32312 13512
rect 31711 13481 31723 13484
rect 31665 13475 31723 13481
rect 32306 13472 32312 13484
rect 32364 13472 32370 13524
rect 18322 13444 18328 13456
rect 14384 13416 18328 13444
rect 2332 13348 3096 13376
rect 2332 13317 2360 13348
rect 2317 13311 2375 13317
rect 2317 13277 2329 13311
rect 2363 13277 2375 13311
rect 2317 13271 2375 13277
rect 2501 13311 2559 13317
rect 2501 13277 2513 13311
rect 2547 13308 2559 13311
rect 2958 13308 2964 13320
rect 2547 13280 2964 13308
rect 2547 13277 2559 13280
rect 2501 13271 2559 13277
rect 2958 13268 2964 13280
rect 3016 13268 3022 13320
rect 3068 13317 3096 13348
rect 3053 13311 3111 13317
rect 3053 13277 3065 13311
rect 3099 13308 3111 13311
rect 3237 13311 3295 13317
rect 3099 13280 3188 13308
rect 3099 13277 3111 13280
rect 3053 13271 3111 13277
rect 2406 13172 2412 13184
rect 2367 13144 2412 13172
rect 2406 13132 2412 13144
rect 2464 13132 2470 13184
rect 3160 13172 3188 13280
rect 3237 13277 3249 13311
rect 3283 13308 3295 13311
rect 3878 13308 3884 13320
rect 3283 13280 3884 13308
rect 3283 13277 3295 13280
rect 3237 13271 3295 13277
rect 3878 13268 3884 13280
rect 3936 13268 3942 13320
rect 4264 13308 4292 13416
rect 4338 13336 4344 13388
rect 4396 13376 4402 13388
rect 4396 13348 5488 13376
rect 4396 13336 4402 13348
rect 4617 13311 4675 13317
rect 4617 13308 4629 13311
rect 4264 13280 4629 13308
rect 4617 13277 4629 13280
rect 4663 13277 4675 13311
rect 4617 13271 4675 13277
rect 5074 13268 5080 13320
rect 5132 13308 5138 13320
rect 5460 13317 5488 13348
rect 7742 13336 7748 13388
rect 7800 13376 7806 13388
rect 9122 13376 9128 13388
rect 7800 13348 9128 13376
rect 7800 13336 7806 13348
rect 9122 13336 9128 13348
rect 9180 13376 9186 13388
rect 11790 13376 11796 13388
rect 9180 13348 11796 13376
rect 9180 13336 9186 13348
rect 11790 13336 11796 13348
rect 11848 13336 11854 13388
rect 12066 13376 12072 13388
rect 12027 13348 12072 13376
rect 12066 13336 12072 13348
rect 12124 13336 12130 13388
rect 12802 13336 12808 13388
rect 12860 13376 12866 13388
rect 15562 13376 15568 13388
rect 12860 13348 15568 13376
rect 12860 13336 12866 13348
rect 15562 13336 15568 13348
rect 15620 13376 15626 13388
rect 15620 13348 15700 13376
rect 15620 13336 15626 13348
rect 5261 13311 5319 13317
rect 5261 13308 5273 13311
rect 5132 13280 5273 13308
rect 5132 13268 5138 13280
rect 5261 13277 5273 13280
rect 5307 13277 5319 13311
rect 5261 13271 5319 13277
rect 5445 13311 5503 13317
rect 5445 13277 5457 13311
rect 5491 13308 5503 13311
rect 8294 13308 8300 13320
rect 5491 13280 8300 13308
rect 5491 13277 5503 13280
rect 5445 13271 5503 13277
rect 8294 13268 8300 13280
rect 8352 13268 8358 13320
rect 8389 13311 8447 13317
rect 8389 13277 8401 13311
rect 8435 13277 8447 13311
rect 8389 13271 8447 13277
rect 3418 13200 3424 13252
rect 3476 13240 3482 13252
rect 4249 13243 4307 13249
rect 4249 13240 4261 13243
rect 3476 13212 4261 13240
rect 3476 13200 3482 13212
rect 4249 13209 4261 13212
rect 4295 13240 4307 13243
rect 8404 13240 8432 13271
rect 13998 13268 14004 13320
rect 14056 13308 14062 13320
rect 15672 13317 15700 13348
rect 14277 13311 14335 13317
rect 14277 13308 14289 13311
rect 14056 13280 14289 13308
rect 14056 13268 14062 13280
rect 14277 13277 14289 13280
rect 14323 13277 14335 13311
rect 14277 13271 14335 13277
rect 14829 13311 14887 13317
rect 14829 13277 14841 13311
rect 14875 13277 14887 13311
rect 14829 13271 14887 13277
rect 15657 13311 15715 13317
rect 15657 13277 15669 13311
rect 15703 13308 15715 13311
rect 15746 13308 15752 13320
rect 15703 13280 15752 13308
rect 15703 13277 15715 13280
rect 15657 13271 15715 13277
rect 4295 13212 8432 13240
rect 4295 13209 4307 13212
rect 4249 13203 4307 13209
rect 8478 13200 8484 13252
rect 8536 13240 8542 13252
rect 8573 13243 8631 13249
rect 8573 13240 8585 13243
rect 8536 13212 8585 13240
rect 8536 13200 8542 13212
rect 8573 13209 8585 13212
rect 8619 13209 8631 13243
rect 8573 13203 8631 13209
rect 8662 13200 8668 13252
rect 8720 13240 8726 13252
rect 9401 13243 9459 13249
rect 9401 13240 9413 13243
rect 8720 13212 9413 13240
rect 8720 13200 8726 13212
rect 9401 13209 9413 13212
rect 9447 13209 9459 13243
rect 9401 13203 9459 13209
rect 10134 13200 10140 13252
rect 10192 13200 10198 13252
rect 14366 13240 14372 13252
rect 13294 13212 14372 13240
rect 14366 13200 14372 13212
rect 14424 13200 14430 13252
rect 14550 13200 14556 13252
rect 14608 13240 14614 13252
rect 14844 13240 14872 13271
rect 15746 13268 15752 13280
rect 15804 13268 15810 13320
rect 17972 13317 18000 13416
rect 18322 13404 18328 13416
rect 18380 13404 18386 13456
rect 18601 13379 18659 13385
rect 18601 13345 18613 13379
rect 18647 13376 18659 13379
rect 21634 13376 21640 13388
rect 18647 13348 21640 13376
rect 18647 13345 18659 13348
rect 18601 13339 18659 13345
rect 21634 13336 21640 13348
rect 21692 13336 21698 13388
rect 16577 13311 16635 13317
rect 16577 13277 16589 13311
rect 16623 13277 16635 13311
rect 16577 13271 16635 13277
rect 17957 13311 18015 13317
rect 17957 13277 17969 13311
rect 18003 13277 18015 13311
rect 18322 13308 18328 13320
rect 18283 13280 18328 13308
rect 17957 13271 18015 13277
rect 16592 13240 16620 13271
rect 18322 13268 18328 13280
rect 18380 13268 18386 13320
rect 19794 13268 19800 13320
rect 19852 13308 19858 13320
rect 20625 13311 20683 13317
rect 20625 13308 20637 13311
rect 19852 13280 20637 13308
rect 19852 13268 19858 13280
rect 20625 13277 20637 13280
rect 20671 13277 20683 13311
rect 26050 13308 26056 13320
rect 26011 13280 26056 13308
rect 20625 13271 20683 13277
rect 26050 13268 26056 13280
rect 26108 13268 26114 13320
rect 32953 13311 33011 13317
rect 32953 13277 32965 13311
rect 32999 13308 33011 13311
rect 33594 13308 33600 13320
rect 32999 13280 33600 13308
rect 32999 13277 33011 13280
rect 32953 13271 33011 13277
rect 33594 13268 33600 13280
rect 33652 13268 33658 13320
rect 14608 13212 14872 13240
rect 15212 13212 16620 13240
rect 14608 13200 14614 13212
rect 4430 13172 4436 13184
rect 3160 13144 4436 13172
rect 4430 13132 4436 13144
rect 4488 13132 4494 13184
rect 7374 13132 7380 13184
rect 7432 13172 7438 13184
rect 8680 13172 8708 13200
rect 15212 13184 15240 13212
rect 7432 13144 8708 13172
rect 7432 13132 7438 13144
rect 9030 13132 9036 13184
rect 9088 13172 9094 13184
rect 10873 13175 10931 13181
rect 10873 13172 10885 13175
rect 9088 13144 10885 13172
rect 9088 13132 9094 13144
rect 10873 13141 10885 13144
rect 10919 13172 10931 13175
rect 12802 13172 12808 13184
rect 10919 13144 12808 13172
rect 10919 13141 10931 13144
rect 10873 13135 10931 13141
rect 12802 13132 12808 13144
rect 12860 13132 12866 13184
rect 13078 13132 13084 13184
rect 13136 13172 13142 13184
rect 13541 13175 13599 13181
rect 13541 13172 13553 13175
rect 13136 13144 13553 13172
rect 13136 13132 13142 13144
rect 13541 13141 13553 13144
rect 13587 13172 13599 13175
rect 15194 13172 15200 13184
rect 13587 13144 15200 13172
rect 13587 13141 13599 13144
rect 13541 13135 13599 13141
rect 15194 13132 15200 13144
rect 15252 13132 15258 13184
rect 18230 13132 18236 13184
rect 18288 13172 18294 13184
rect 21913 13175 21971 13181
rect 21913 13172 21925 13175
rect 18288 13144 21925 13172
rect 18288 13132 18294 13144
rect 21913 13141 21925 13144
rect 21959 13141 21971 13175
rect 21913 13135 21971 13141
rect 1104 13082 35027 13104
rect 1104 13030 9390 13082
rect 9442 13030 9454 13082
rect 9506 13030 9518 13082
rect 9570 13030 9582 13082
rect 9634 13030 9646 13082
rect 9698 13030 17831 13082
rect 17883 13030 17895 13082
rect 17947 13030 17959 13082
rect 18011 13030 18023 13082
rect 18075 13030 18087 13082
rect 18139 13030 26272 13082
rect 26324 13030 26336 13082
rect 26388 13030 26400 13082
rect 26452 13030 26464 13082
rect 26516 13030 26528 13082
rect 26580 13030 34713 13082
rect 34765 13030 34777 13082
rect 34829 13030 34841 13082
rect 34893 13030 34905 13082
rect 34957 13030 34969 13082
rect 35021 13030 35027 13082
rect 1104 13008 35027 13030
rect 4338 12968 4344 12980
rect 2148 12940 4344 12968
rect 2148 12841 2176 12940
rect 4338 12928 4344 12940
rect 4396 12928 4402 12980
rect 4430 12928 4436 12980
rect 4488 12968 4494 12980
rect 20438 12968 20444 12980
rect 4488 12940 4533 12968
rect 20399 12940 20444 12968
rect 4488 12928 4494 12940
rect 20438 12928 20444 12940
rect 20496 12928 20502 12980
rect 27706 12968 27712 12980
rect 27448 12940 27712 12968
rect 2406 12900 2412 12912
rect 2367 12872 2412 12900
rect 2406 12860 2412 12872
rect 2464 12860 2470 12912
rect 3142 12860 3148 12912
rect 3200 12860 3206 12912
rect 8478 12860 8484 12912
rect 8536 12860 8542 12912
rect 9214 12860 9220 12912
rect 9272 12900 9278 12912
rect 9493 12903 9551 12909
rect 9493 12900 9505 12903
rect 9272 12872 9505 12900
rect 9272 12860 9278 12872
rect 9493 12869 9505 12872
rect 9539 12869 9551 12903
rect 12986 12900 12992 12912
rect 12947 12872 12992 12900
rect 9493 12863 9551 12869
rect 12986 12860 12992 12872
rect 13044 12860 13050 12912
rect 14734 12900 14740 12912
rect 14695 12872 14740 12900
rect 14734 12860 14740 12872
rect 14792 12860 14798 12912
rect 18417 12903 18475 12909
rect 17144 12872 18276 12900
rect 2133 12835 2191 12841
rect 2133 12801 2145 12835
rect 2179 12801 2191 12835
rect 3970 12832 3976 12844
rect 2133 12795 2191 12801
rect 3620 12804 3976 12832
rect 3050 12724 3056 12776
rect 3108 12764 3114 12776
rect 3620 12764 3648 12804
rect 3970 12792 3976 12804
rect 4028 12832 4034 12844
rect 4341 12835 4399 12841
rect 4341 12832 4353 12835
rect 4028 12804 4353 12832
rect 4028 12792 4034 12804
rect 4341 12801 4353 12804
rect 4387 12801 4399 12835
rect 4522 12832 4528 12844
rect 4483 12804 4528 12832
rect 4341 12795 4399 12801
rect 4522 12792 4528 12804
rect 4580 12792 4586 12844
rect 15102 12792 15108 12844
rect 15160 12832 15166 12844
rect 15381 12835 15439 12841
rect 15381 12832 15393 12835
rect 15160 12804 15393 12832
rect 15160 12792 15166 12804
rect 15381 12801 15393 12804
rect 15427 12801 15439 12835
rect 15381 12795 15439 12801
rect 16025 12835 16083 12841
rect 16025 12801 16037 12835
rect 16071 12801 16083 12835
rect 16942 12832 16948 12844
rect 16903 12804 16948 12832
rect 16025 12795 16083 12801
rect 3878 12764 3884 12776
rect 3108 12736 3648 12764
rect 3839 12736 3884 12764
rect 3108 12724 3114 12736
rect 3878 12724 3884 12736
rect 3936 12724 3942 12776
rect 9122 12724 9128 12776
rect 9180 12764 9186 12776
rect 9769 12767 9827 12773
rect 9769 12764 9781 12767
rect 9180 12736 9781 12764
rect 9180 12724 9186 12736
rect 9769 12733 9781 12736
rect 9815 12733 9827 12767
rect 9769 12727 9827 12733
rect 14550 12724 14556 12776
rect 14608 12764 14614 12776
rect 16040 12764 16068 12795
rect 16942 12792 16948 12804
rect 17000 12792 17006 12844
rect 17144 12841 17172 12872
rect 17129 12835 17187 12841
rect 17129 12801 17141 12835
rect 17175 12801 17187 12835
rect 17129 12795 17187 12801
rect 17402 12792 17408 12844
rect 17460 12832 17466 12844
rect 18248 12841 18276 12872
rect 18417 12869 18429 12903
rect 18463 12900 18475 12903
rect 22646 12900 22652 12912
rect 18463 12872 22652 12900
rect 18463 12869 18475 12872
rect 18417 12863 18475 12869
rect 22646 12860 22652 12872
rect 22704 12860 22710 12912
rect 17681 12835 17739 12841
rect 17681 12832 17693 12835
rect 17460 12804 17693 12832
rect 17460 12792 17466 12804
rect 17681 12801 17693 12804
rect 17727 12801 17739 12835
rect 17681 12795 17739 12801
rect 18233 12835 18291 12841
rect 18233 12801 18245 12835
rect 18279 12832 18291 12835
rect 18322 12832 18328 12844
rect 18279 12804 18328 12832
rect 18279 12801 18291 12804
rect 18233 12795 18291 12801
rect 18322 12792 18328 12804
rect 18380 12792 18386 12844
rect 20625 12835 20683 12841
rect 20625 12801 20637 12835
rect 20671 12801 20683 12835
rect 20625 12795 20683 12801
rect 14608 12736 16068 12764
rect 16117 12767 16175 12773
rect 14608 12724 14614 12736
rect 16117 12733 16129 12767
rect 16163 12764 16175 12767
rect 16574 12764 16580 12776
rect 16163 12736 16580 12764
rect 16163 12733 16175 12736
rect 16117 12727 16175 12733
rect 16574 12724 16580 12736
rect 16632 12724 16638 12776
rect 17221 12767 17279 12773
rect 17221 12733 17233 12767
rect 17267 12764 17279 12767
rect 19610 12764 19616 12776
rect 17267 12736 19616 12764
rect 17267 12733 17279 12736
rect 17221 12727 17279 12733
rect 19610 12724 19616 12736
rect 19668 12764 19674 12776
rect 20640 12764 20668 12795
rect 20714 12792 20720 12844
rect 20772 12832 20778 12844
rect 20898 12832 20904 12844
rect 20772 12804 20817 12832
rect 20859 12804 20904 12832
rect 20772 12792 20778 12804
rect 20898 12792 20904 12804
rect 20956 12792 20962 12844
rect 20990 12792 20996 12844
rect 21048 12832 21054 12844
rect 21048 12804 21093 12832
rect 21048 12792 21054 12804
rect 26602 12792 26608 12844
rect 26660 12832 26666 12844
rect 27448 12841 27476 12940
rect 27706 12928 27712 12940
rect 27764 12928 27770 12980
rect 27893 12971 27951 12977
rect 27893 12937 27905 12971
rect 27939 12968 27951 12971
rect 28350 12968 28356 12980
rect 27939 12940 28356 12968
rect 27939 12937 27951 12940
rect 27893 12931 27951 12937
rect 28350 12928 28356 12940
rect 28408 12928 28414 12980
rect 32122 12928 32128 12980
rect 32180 12968 32186 12980
rect 32309 12971 32367 12977
rect 32309 12968 32321 12971
rect 32180 12940 32321 12968
rect 32180 12928 32186 12940
rect 32309 12937 32321 12940
rect 32355 12937 32367 12971
rect 32309 12931 32367 12937
rect 32677 12971 32735 12977
rect 32677 12937 32689 12971
rect 32723 12968 32735 12971
rect 33042 12968 33048 12980
rect 32723 12940 33048 12968
rect 32723 12937 32735 12940
rect 32677 12931 32735 12937
rect 33042 12928 33048 12940
rect 33100 12928 33106 12980
rect 27617 12903 27675 12909
rect 27617 12869 27629 12903
rect 27663 12900 27675 12903
rect 27798 12900 27804 12912
rect 27663 12872 27804 12900
rect 27663 12869 27675 12872
rect 27617 12863 27675 12869
rect 27798 12860 27804 12872
rect 27856 12860 27862 12912
rect 28442 12860 28448 12912
rect 28500 12900 28506 12912
rect 28721 12903 28779 12909
rect 28721 12900 28733 12903
rect 28500 12872 28733 12900
rect 28500 12860 28506 12872
rect 28721 12869 28733 12872
rect 28767 12869 28779 12903
rect 28721 12863 28779 12869
rect 27249 12835 27307 12841
rect 27249 12832 27261 12835
rect 26660 12804 27261 12832
rect 26660 12792 26666 12804
rect 27249 12801 27261 12804
rect 27295 12801 27307 12835
rect 27249 12795 27307 12801
rect 27397 12835 27476 12841
rect 27397 12801 27409 12835
rect 27443 12804 27476 12835
rect 27525 12835 27583 12841
rect 27443 12801 27455 12804
rect 27397 12795 27455 12801
rect 27525 12801 27537 12835
rect 27571 12801 27583 12835
rect 27714 12835 27772 12841
rect 27714 12832 27726 12835
rect 27525 12795 27583 12801
rect 27623 12804 27726 12832
rect 19668 12736 20668 12764
rect 19668 12724 19674 12736
rect 24026 12724 24032 12776
rect 24084 12764 24090 12776
rect 25498 12764 25504 12776
rect 24084 12736 25504 12764
rect 24084 12724 24090 12736
rect 25498 12724 25504 12736
rect 25556 12764 25562 12776
rect 27540 12764 27568 12795
rect 25556 12736 27568 12764
rect 25556 12724 25562 12736
rect 16592 12696 16620 12724
rect 17402 12696 17408 12708
rect 16592 12668 17408 12696
rect 17402 12656 17408 12668
rect 17460 12656 17466 12708
rect 20530 12656 20536 12708
rect 20588 12696 20594 12708
rect 27623 12696 27651 12804
rect 27714 12801 27726 12804
rect 27760 12801 27772 12835
rect 27714 12795 27772 12801
rect 28537 12835 28595 12841
rect 28537 12801 28549 12835
rect 28583 12801 28595 12835
rect 28537 12795 28595 12801
rect 28813 12835 28871 12841
rect 28813 12801 28825 12835
rect 28859 12832 28871 12835
rect 28859 12804 29592 12832
rect 28859 12801 28871 12804
rect 28813 12795 28871 12801
rect 28552 12764 28580 12795
rect 28994 12764 29000 12776
rect 28552 12736 29000 12764
rect 28994 12724 29000 12736
rect 29052 12724 29058 12776
rect 29564 12773 29592 12804
rect 29638 12792 29644 12844
rect 29696 12832 29702 12844
rect 29733 12835 29791 12841
rect 29733 12832 29745 12835
rect 29696 12804 29745 12832
rect 29696 12792 29702 12804
rect 29733 12801 29745 12804
rect 29779 12801 29791 12835
rect 32490 12832 32496 12844
rect 32451 12804 32496 12832
rect 29733 12795 29791 12801
rect 32490 12792 32496 12804
rect 32548 12792 32554 12844
rect 32769 12835 32827 12841
rect 32769 12801 32781 12835
rect 32815 12832 32827 12835
rect 33410 12832 33416 12844
rect 32815 12804 33416 12832
rect 32815 12801 32827 12804
rect 32769 12795 32827 12801
rect 33410 12792 33416 12804
rect 33468 12792 33474 12844
rect 29549 12767 29607 12773
rect 29549 12733 29561 12767
rect 29595 12764 29607 12767
rect 30190 12764 30196 12776
rect 29595 12736 30196 12764
rect 29595 12733 29607 12736
rect 29549 12727 29607 12733
rect 30190 12724 30196 12736
rect 30248 12724 30254 12776
rect 27890 12696 27896 12708
rect 20588 12668 27896 12696
rect 20588 12656 20594 12668
rect 27890 12656 27896 12668
rect 27948 12656 27954 12708
rect 29012 12696 29040 12724
rect 30374 12696 30380 12708
rect 29012 12668 30380 12696
rect 30374 12656 30380 12668
rect 30432 12656 30438 12708
rect 7466 12588 7472 12640
rect 7524 12628 7530 12640
rect 8021 12631 8079 12637
rect 8021 12628 8033 12631
rect 7524 12600 8033 12628
rect 7524 12588 7530 12600
rect 8021 12597 8033 12600
rect 8067 12628 8079 12631
rect 14550 12628 14556 12640
rect 8067 12600 14556 12628
rect 8067 12597 8079 12600
rect 8021 12591 8079 12597
rect 14550 12588 14556 12600
rect 14608 12588 14614 12640
rect 17494 12588 17500 12640
rect 17552 12628 17558 12640
rect 21358 12628 21364 12640
rect 17552 12600 21364 12628
rect 17552 12588 17558 12600
rect 21358 12588 21364 12600
rect 21416 12588 21422 12640
rect 21450 12588 21456 12640
rect 21508 12628 21514 12640
rect 25038 12628 25044 12640
rect 21508 12600 25044 12628
rect 21508 12588 21514 12600
rect 25038 12588 25044 12600
rect 25096 12588 25102 12640
rect 28350 12628 28356 12640
rect 28311 12600 28356 12628
rect 28350 12588 28356 12600
rect 28408 12588 28414 12640
rect 1104 12538 34868 12560
rect 1104 12486 5170 12538
rect 5222 12486 5234 12538
rect 5286 12486 5298 12538
rect 5350 12486 5362 12538
rect 5414 12486 5426 12538
rect 5478 12486 13611 12538
rect 13663 12486 13675 12538
rect 13727 12486 13739 12538
rect 13791 12486 13803 12538
rect 13855 12486 13867 12538
rect 13919 12486 22052 12538
rect 22104 12486 22116 12538
rect 22168 12486 22180 12538
rect 22232 12486 22244 12538
rect 22296 12486 22308 12538
rect 22360 12486 30493 12538
rect 30545 12486 30557 12538
rect 30609 12486 30621 12538
rect 30673 12486 30685 12538
rect 30737 12486 30749 12538
rect 30801 12486 34868 12538
rect 1104 12464 34868 12486
rect 3142 12424 3148 12436
rect 3103 12396 3148 12424
rect 3142 12384 3148 12396
rect 3200 12384 3206 12436
rect 13998 12384 14004 12436
rect 14056 12424 14062 12436
rect 15102 12424 15108 12436
rect 14056 12396 15108 12424
rect 14056 12384 14062 12396
rect 15102 12384 15108 12396
rect 15160 12384 15166 12436
rect 16942 12356 16948 12368
rect 15304 12328 16948 12356
rect 4338 12288 4344 12300
rect 3160 12260 4344 12288
rect 3160 12229 3188 12260
rect 4338 12248 4344 12260
rect 4396 12248 4402 12300
rect 15304 12297 15332 12328
rect 16942 12316 16948 12328
rect 17000 12316 17006 12368
rect 20898 12316 20904 12368
rect 20956 12356 20962 12368
rect 27893 12359 27951 12365
rect 27893 12356 27905 12359
rect 20956 12328 27905 12356
rect 20956 12316 20962 12328
rect 27893 12325 27905 12328
rect 27939 12325 27951 12359
rect 27893 12319 27951 12325
rect 15289 12291 15347 12297
rect 15289 12257 15301 12291
rect 15335 12257 15347 12291
rect 15289 12251 15347 12257
rect 16669 12291 16727 12297
rect 16669 12257 16681 12291
rect 16715 12288 16727 12291
rect 18322 12288 18328 12300
rect 16715 12260 18328 12288
rect 16715 12257 16727 12260
rect 16669 12251 16727 12257
rect 3145 12223 3203 12229
rect 3145 12189 3157 12223
rect 3191 12189 3203 12223
rect 3145 12183 3203 12189
rect 3329 12223 3387 12229
rect 3329 12189 3341 12223
rect 3375 12220 3387 12223
rect 3418 12220 3424 12232
rect 3375 12192 3424 12220
rect 3375 12189 3387 12192
rect 3329 12183 3387 12189
rect 3418 12180 3424 12192
rect 3476 12180 3482 12232
rect 14550 12220 14556 12232
rect 14511 12192 14556 12220
rect 14550 12180 14556 12192
rect 14608 12180 14614 12232
rect 15102 12180 15108 12232
rect 15160 12220 15166 12232
rect 15197 12223 15255 12229
rect 15197 12220 15209 12223
rect 15160 12192 15209 12220
rect 15160 12180 15166 12192
rect 15197 12189 15209 12192
rect 15243 12189 15255 12223
rect 15197 12183 15255 12189
rect 15746 12180 15752 12232
rect 15804 12220 15810 12232
rect 15933 12223 15991 12229
rect 15933 12220 15945 12223
rect 15804 12192 15945 12220
rect 15804 12180 15810 12192
rect 15933 12189 15945 12192
rect 15979 12189 15991 12223
rect 15933 12183 15991 12189
rect 16298 12180 16304 12232
rect 16356 12220 16362 12232
rect 16577 12223 16635 12229
rect 16577 12220 16589 12223
rect 16356 12192 16589 12220
rect 16356 12180 16362 12192
rect 16577 12189 16589 12192
rect 16623 12189 16635 12223
rect 17586 12220 17592 12232
rect 17547 12192 17592 12220
rect 16577 12183 16635 12189
rect 17586 12180 17592 12192
rect 17644 12180 17650 12232
rect 17972 12229 18000 12260
rect 18322 12248 18328 12260
rect 18380 12248 18386 12300
rect 22554 12288 22560 12300
rect 22515 12260 22560 12288
rect 22554 12248 22560 12260
rect 22612 12248 22618 12300
rect 28626 12288 28632 12300
rect 24780 12260 28632 12288
rect 17957 12223 18015 12229
rect 17957 12189 17969 12223
rect 18003 12189 18015 12223
rect 17957 12183 18015 12189
rect 21358 12180 21364 12232
rect 21416 12220 21422 12232
rect 24780 12229 24808 12260
rect 28626 12248 28632 12260
rect 28684 12248 28690 12300
rect 28074 12229 28080 12232
rect 24765 12223 24823 12229
rect 24765 12220 24777 12223
rect 21416 12192 24777 12220
rect 21416 12180 21422 12192
rect 24765 12189 24777 12192
rect 24811 12189 24823 12223
rect 24765 12183 24823 12189
rect 25041 12223 25099 12229
rect 25041 12189 25053 12223
rect 25087 12189 25099 12223
rect 28072 12220 28080 12229
rect 28035 12192 28080 12220
rect 25041 12183 25099 12189
rect 28072 12183 28080 12192
rect 18233 12155 18291 12161
rect 18233 12121 18245 12155
rect 18279 12152 18291 12155
rect 19150 12152 19156 12164
rect 18279 12124 19156 12152
rect 18279 12121 18291 12124
rect 18233 12115 18291 12121
rect 19150 12112 19156 12124
rect 19208 12112 19214 12164
rect 20806 12152 20812 12164
rect 20767 12124 20812 12152
rect 20806 12112 20812 12124
rect 20864 12112 20870 12164
rect 23658 12112 23664 12164
rect 23716 12152 23722 12164
rect 24486 12152 24492 12164
rect 23716 12124 24492 12152
rect 23716 12112 23722 12124
rect 24486 12112 24492 12124
rect 24544 12152 24550 12164
rect 25056 12152 25084 12183
rect 28074 12180 28080 12183
rect 28132 12180 28138 12232
rect 28442 12220 28448 12232
rect 28403 12192 28448 12220
rect 28442 12180 28448 12192
rect 28500 12180 28506 12232
rect 28534 12180 28540 12232
rect 28592 12220 28598 12232
rect 28592 12192 28637 12220
rect 28592 12180 28598 12192
rect 24544 12124 25084 12152
rect 28169 12155 28227 12161
rect 24544 12112 24550 12124
rect 28169 12121 28181 12155
rect 28215 12121 28227 12155
rect 28169 12115 28227 12121
rect 28261 12155 28319 12161
rect 28261 12121 28273 12155
rect 28307 12152 28319 12155
rect 28626 12152 28632 12164
rect 28307 12124 28632 12152
rect 28307 12121 28319 12124
rect 28261 12115 28319 12121
rect 17126 12044 17132 12096
rect 17184 12084 17190 12096
rect 17310 12084 17316 12096
rect 17184 12056 17316 12084
rect 17184 12044 17190 12056
rect 17310 12044 17316 12056
rect 17368 12044 17374 12096
rect 24578 12084 24584 12096
rect 24539 12056 24584 12084
rect 24578 12044 24584 12056
rect 24636 12044 24642 12096
rect 24946 12084 24952 12096
rect 24907 12056 24952 12084
rect 24946 12044 24952 12056
rect 25004 12044 25010 12096
rect 28184 12084 28212 12115
rect 28626 12112 28632 12124
rect 28684 12112 28690 12164
rect 31294 12084 31300 12096
rect 28184 12056 31300 12084
rect 31294 12044 31300 12056
rect 31352 12044 31358 12096
rect 1104 11994 35027 12016
rect 1104 11942 9390 11994
rect 9442 11942 9454 11994
rect 9506 11942 9518 11994
rect 9570 11942 9582 11994
rect 9634 11942 9646 11994
rect 9698 11942 17831 11994
rect 17883 11942 17895 11994
rect 17947 11942 17959 11994
rect 18011 11942 18023 11994
rect 18075 11942 18087 11994
rect 18139 11942 26272 11994
rect 26324 11942 26336 11994
rect 26388 11942 26400 11994
rect 26452 11942 26464 11994
rect 26516 11942 26528 11994
rect 26580 11942 34713 11994
rect 34765 11942 34777 11994
rect 34829 11942 34841 11994
rect 34893 11942 34905 11994
rect 34957 11942 34969 11994
rect 35021 11942 35027 11994
rect 1104 11920 35027 11942
rect 20530 11880 20536 11892
rect 18524 11852 20536 11880
rect 15746 11812 15752 11824
rect 15707 11784 15752 11812
rect 15746 11772 15752 11784
rect 15804 11772 15810 11824
rect 18414 11812 18420 11824
rect 18064 11784 18420 11812
rect 15194 11704 15200 11756
rect 15252 11744 15258 11756
rect 15933 11747 15991 11753
rect 15933 11744 15945 11747
rect 15252 11716 15945 11744
rect 15252 11704 15258 11716
rect 15933 11713 15945 11716
rect 15979 11744 15991 11747
rect 16298 11744 16304 11756
rect 15979 11716 16304 11744
rect 15979 11713 15991 11716
rect 15933 11707 15991 11713
rect 16298 11704 16304 11716
rect 16356 11704 16362 11756
rect 16574 11704 16580 11756
rect 16632 11744 16638 11756
rect 18064 11753 18092 11784
rect 18414 11772 18420 11784
rect 18472 11772 18478 11824
rect 18524 11821 18552 11852
rect 20530 11840 20536 11852
rect 20588 11840 20594 11892
rect 20714 11840 20720 11892
rect 20772 11880 20778 11892
rect 21085 11883 21143 11889
rect 21085 11880 21097 11883
rect 20772 11852 21097 11880
rect 20772 11840 20778 11852
rect 21085 11849 21097 11852
rect 21131 11849 21143 11883
rect 21085 11843 21143 11849
rect 22462 11840 22468 11892
rect 22520 11880 22526 11892
rect 28166 11880 28172 11892
rect 22520 11852 28172 11880
rect 22520 11840 22526 11852
rect 28166 11840 28172 11852
rect 28224 11840 28230 11892
rect 28442 11840 28448 11892
rect 28500 11880 28506 11892
rect 28721 11883 28779 11889
rect 28721 11880 28733 11883
rect 28500 11852 28733 11880
rect 28500 11840 28506 11852
rect 28721 11849 28733 11852
rect 28767 11849 28779 11883
rect 31294 11880 31300 11892
rect 31255 11852 31300 11880
rect 28721 11843 28779 11849
rect 31294 11840 31300 11852
rect 31352 11840 31358 11892
rect 32674 11880 32680 11892
rect 32635 11852 32680 11880
rect 32674 11840 32680 11852
rect 32732 11880 32738 11892
rect 33686 11880 33692 11892
rect 32732 11852 33692 11880
rect 32732 11840 32738 11852
rect 33686 11840 33692 11852
rect 33744 11840 33750 11892
rect 18509 11815 18567 11821
rect 18509 11781 18521 11815
rect 18555 11781 18567 11815
rect 18509 11775 18567 11781
rect 19720 11784 20576 11812
rect 19720 11756 19748 11784
rect 16945 11747 17003 11753
rect 16945 11744 16957 11747
rect 16632 11716 16957 11744
rect 16632 11704 16638 11716
rect 16945 11713 16957 11716
rect 16991 11713 17003 11747
rect 16945 11707 17003 11713
rect 17129 11747 17187 11753
rect 17129 11713 17141 11747
rect 17175 11713 17187 11747
rect 17129 11707 17187 11713
rect 18049 11747 18107 11753
rect 18049 11713 18061 11747
rect 18095 11713 18107 11747
rect 18049 11707 18107 11713
rect 18233 11747 18291 11753
rect 18233 11713 18245 11747
rect 18279 11713 18291 11747
rect 19702 11744 19708 11756
rect 19615 11716 19708 11744
rect 18233 11707 18291 11713
rect 16209 11679 16267 11685
rect 16209 11645 16221 11679
rect 16255 11676 16267 11679
rect 16850 11676 16856 11688
rect 16255 11648 16856 11676
rect 16255 11645 16267 11648
rect 16209 11639 16267 11645
rect 16850 11636 16856 11648
rect 16908 11676 16914 11688
rect 17144 11676 17172 11707
rect 18248 11676 18276 11707
rect 19702 11704 19708 11716
rect 19760 11704 19766 11756
rect 19972 11747 20030 11753
rect 19972 11713 19984 11747
rect 20018 11744 20030 11747
rect 20438 11744 20444 11756
rect 20018 11716 20444 11744
rect 20018 11713 20030 11716
rect 19972 11707 20030 11713
rect 20438 11704 20444 11716
rect 20496 11704 20502 11756
rect 20548 11744 20576 11784
rect 22554 11772 22560 11824
rect 22612 11812 22618 11824
rect 22738 11812 22744 11824
rect 22612 11784 22744 11812
rect 22612 11772 22618 11784
rect 22738 11772 22744 11784
rect 22796 11812 22802 11824
rect 25685 11815 25743 11821
rect 25685 11812 25697 11815
rect 22796 11784 25697 11812
rect 22796 11772 22802 11784
rect 25685 11781 25697 11784
rect 25731 11781 25743 11815
rect 25685 11775 25743 11781
rect 25869 11815 25927 11821
rect 25869 11781 25881 11815
rect 25915 11781 25927 11815
rect 25869 11775 25927 11781
rect 27608 11815 27666 11821
rect 27608 11781 27620 11815
rect 27654 11812 27666 11815
rect 28350 11812 28356 11824
rect 27654 11784 28356 11812
rect 27654 11781 27666 11784
rect 27608 11775 27666 11781
rect 22005 11747 22063 11753
rect 22005 11744 22017 11747
rect 20548 11716 22017 11744
rect 22005 11713 22017 11716
rect 22051 11713 22063 11747
rect 22261 11747 22319 11753
rect 22261 11744 22273 11747
rect 22005 11707 22063 11713
rect 22112 11716 22273 11744
rect 16908 11648 18276 11676
rect 16908 11636 16914 11648
rect 21542 11636 21548 11688
rect 21600 11676 21606 11688
rect 22112 11676 22140 11716
rect 22261 11713 22273 11716
rect 22307 11713 22319 11747
rect 22261 11707 22319 11713
rect 24112 11747 24170 11753
rect 24112 11713 24124 11747
rect 24158 11744 24170 11747
rect 24578 11744 24584 11756
rect 24158 11716 24584 11744
rect 24158 11713 24170 11716
rect 24112 11707 24170 11713
rect 24578 11704 24584 11716
rect 24636 11704 24642 11756
rect 25314 11704 25320 11756
rect 25372 11744 25378 11756
rect 25884 11744 25912 11775
rect 28350 11772 28356 11784
rect 28408 11772 28414 11824
rect 30374 11772 30380 11824
rect 30432 11812 30438 11824
rect 30432 11784 31524 11812
rect 30432 11772 30438 11784
rect 28626 11744 28632 11756
rect 25372 11716 28632 11744
rect 25372 11704 25378 11716
rect 28626 11704 28632 11716
rect 28684 11704 28690 11756
rect 30190 11704 30196 11756
rect 30248 11744 30254 11756
rect 31496 11753 31524 11784
rect 31205 11747 31263 11753
rect 31205 11744 31217 11747
rect 30248 11716 31217 11744
rect 30248 11704 30254 11716
rect 31205 11713 31217 11716
rect 31251 11713 31263 11747
rect 31205 11707 31263 11713
rect 31481 11747 31539 11753
rect 31481 11713 31493 11747
rect 31527 11713 31539 11747
rect 31481 11707 31539 11713
rect 23842 11676 23848 11688
rect 21600 11648 22140 11676
rect 23803 11648 23848 11676
rect 21600 11636 21606 11648
rect 23842 11636 23848 11648
rect 23900 11636 23906 11688
rect 27338 11676 27344 11688
rect 27299 11648 27344 11676
rect 27338 11636 27344 11648
rect 27396 11636 27402 11688
rect 31220 11676 31248 11707
rect 31846 11704 31852 11756
rect 31904 11744 31910 11756
rect 32490 11744 32496 11756
rect 31904 11716 32496 11744
rect 31904 11704 31910 11716
rect 32490 11704 32496 11716
rect 32548 11704 32554 11756
rect 32769 11747 32827 11753
rect 32769 11713 32781 11747
rect 32815 11713 32827 11747
rect 32769 11707 32827 11713
rect 32784 11676 32812 11707
rect 33410 11676 33416 11688
rect 31220 11648 33416 11676
rect 33410 11636 33416 11648
rect 33468 11636 33474 11688
rect 17221 11611 17279 11617
rect 17221 11577 17233 11611
rect 17267 11577 17279 11611
rect 17221 11571 17279 11577
rect 21008 11580 21220 11608
rect 17236 11540 17264 11571
rect 21008 11540 21036 11580
rect 17236 11512 21036 11540
rect 21192 11540 21220 11580
rect 25884 11580 26188 11608
rect 22646 11540 22652 11552
rect 21192 11512 22652 11540
rect 22646 11500 22652 11512
rect 22704 11500 22710 11552
rect 22922 11500 22928 11552
rect 22980 11540 22986 11552
rect 23385 11543 23443 11549
rect 23385 11540 23397 11543
rect 22980 11512 23397 11540
rect 22980 11500 22986 11512
rect 23385 11509 23397 11512
rect 23431 11509 23443 11543
rect 23385 11503 23443 11509
rect 23474 11500 23480 11552
rect 23532 11540 23538 11552
rect 24946 11540 24952 11552
rect 23532 11512 24952 11540
rect 23532 11500 23538 11512
rect 24946 11500 24952 11512
rect 25004 11540 25010 11552
rect 25884 11549 25912 11580
rect 25225 11543 25283 11549
rect 25225 11540 25237 11543
rect 25004 11512 25237 11540
rect 25004 11500 25010 11512
rect 25225 11509 25237 11512
rect 25271 11509 25283 11543
rect 25225 11503 25283 11509
rect 25869 11543 25927 11549
rect 25869 11509 25881 11543
rect 25915 11509 25927 11543
rect 26050 11540 26056 11552
rect 26011 11512 26056 11540
rect 25869 11503 25927 11509
rect 26050 11500 26056 11512
rect 26108 11500 26114 11552
rect 26160 11540 26188 11580
rect 29362 11540 29368 11552
rect 26160 11512 29368 11540
rect 29362 11500 29368 11512
rect 29420 11500 29426 11552
rect 31662 11540 31668 11552
rect 31623 11512 31668 11540
rect 31662 11500 31668 11512
rect 31720 11500 31726 11552
rect 32309 11543 32367 11549
rect 32309 11509 32321 11543
rect 32355 11540 32367 11543
rect 32398 11540 32404 11552
rect 32355 11512 32404 11540
rect 32355 11509 32367 11512
rect 32309 11503 32367 11509
rect 32398 11500 32404 11512
rect 32456 11500 32462 11552
rect 1104 11450 34868 11472
rect 1104 11398 5170 11450
rect 5222 11398 5234 11450
rect 5286 11398 5298 11450
rect 5350 11398 5362 11450
rect 5414 11398 5426 11450
rect 5478 11398 13611 11450
rect 13663 11398 13675 11450
rect 13727 11398 13739 11450
rect 13791 11398 13803 11450
rect 13855 11398 13867 11450
rect 13919 11398 22052 11450
rect 22104 11398 22116 11450
rect 22168 11398 22180 11450
rect 22232 11398 22244 11450
rect 22296 11398 22308 11450
rect 22360 11398 30493 11450
rect 30545 11398 30557 11450
rect 30609 11398 30621 11450
rect 30673 11398 30685 11450
rect 30737 11398 30749 11450
rect 30801 11398 34868 11450
rect 1104 11376 34868 11398
rect 4157 11339 4215 11345
rect 4157 11305 4169 11339
rect 4203 11336 4215 11339
rect 4522 11336 4528 11348
rect 4203 11308 4528 11336
rect 4203 11305 4215 11308
rect 4157 11299 4215 11305
rect 4522 11296 4528 11308
rect 4580 11296 4586 11348
rect 17310 11296 17316 11348
rect 17368 11336 17374 11348
rect 21082 11336 21088 11348
rect 17368 11308 21088 11336
rect 17368 11296 17374 11308
rect 21082 11296 21088 11308
rect 21140 11296 21146 11348
rect 21542 11336 21548 11348
rect 21503 11308 21548 11336
rect 21542 11296 21548 11308
rect 21600 11296 21606 11348
rect 22462 11336 22468 11348
rect 22066 11308 22468 11336
rect 13633 11271 13691 11277
rect 13633 11237 13645 11271
rect 13679 11268 13691 11271
rect 15930 11268 15936 11280
rect 13679 11240 15936 11268
rect 13679 11237 13691 11240
rect 13633 11231 13691 11237
rect 15930 11228 15936 11240
rect 15988 11228 15994 11280
rect 22066 11268 22094 11308
rect 22462 11296 22468 11308
rect 22520 11296 22526 11348
rect 22830 11336 22836 11348
rect 22791 11308 22836 11336
rect 22830 11296 22836 11308
rect 22888 11296 22894 11348
rect 25314 11336 25320 11348
rect 23492 11308 25320 11336
rect 20364 11240 22094 11268
rect 12164 11212 12216 11218
rect 2958 11160 2964 11212
rect 3016 11200 3022 11212
rect 3326 11200 3332 11212
rect 3016 11172 3332 11200
rect 3016 11160 3022 11172
rect 3326 11160 3332 11172
rect 3384 11200 3390 11212
rect 3384 11172 3464 11200
rect 3384 11160 3390 11172
rect 3234 11132 3240 11144
rect 3195 11104 3240 11132
rect 3234 11092 3240 11104
rect 3292 11092 3298 11144
rect 3436 11141 3464 11172
rect 17678 11160 17684 11212
rect 17736 11200 17742 11212
rect 17736 11172 20300 11200
rect 17736 11160 17742 11172
rect 12164 11154 12216 11160
rect 3421 11135 3479 11141
rect 3421 11101 3433 11135
rect 3467 11132 3479 11135
rect 5537 11135 5595 11141
rect 3467 11104 4108 11132
rect 3467 11101 3479 11104
rect 3421 11095 3479 11101
rect 2498 11024 2504 11076
rect 2556 11064 2562 11076
rect 3970 11064 3976 11076
rect 2556 11036 3976 11064
rect 2556 11024 2562 11036
rect 3970 11024 3976 11036
rect 4028 11024 4034 11076
rect 4080 11064 4108 11104
rect 5537 11101 5549 11135
rect 5583 11132 5595 11135
rect 6086 11132 6092 11144
rect 5583 11104 6092 11132
rect 5583 11101 5595 11104
rect 5537 11095 5595 11101
rect 6086 11092 6092 11104
rect 6144 11092 6150 11144
rect 10321 11135 10379 11141
rect 10321 11101 10333 11135
rect 10367 11132 10379 11135
rect 10410 11132 10416 11144
rect 10367 11104 10416 11132
rect 10367 11101 10379 11104
rect 10321 11095 10379 11101
rect 10410 11092 10416 11104
rect 10468 11092 10474 11144
rect 10588 11135 10646 11141
rect 10588 11101 10600 11135
rect 10634 11132 10646 11135
rect 11054 11132 11060 11144
rect 10634 11104 11060 11132
rect 10634 11101 10646 11104
rect 10588 11095 10646 11101
rect 11054 11092 11060 11104
rect 11112 11092 11118 11144
rect 12526 11092 12532 11144
rect 12584 11132 12590 11144
rect 12713 11135 12771 11141
rect 12713 11132 12725 11135
rect 12584 11104 12725 11132
rect 12584 11092 12590 11104
rect 12713 11101 12725 11104
rect 12759 11132 12771 11135
rect 12894 11132 12900 11144
rect 12759 11104 12900 11132
rect 12759 11101 12771 11104
rect 12713 11095 12771 11101
rect 12894 11092 12900 11104
rect 12952 11092 12958 11144
rect 13078 11132 13084 11144
rect 13039 11104 13084 11132
rect 13078 11092 13084 11104
rect 13136 11092 13142 11144
rect 16850 11132 16856 11144
rect 16811 11104 16856 11132
rect 16850 11092 16856 11104
rect 16908 11092 16914 11144
rect 16942 11092 16948 11144
rect 17000 11132 17006 11144
rect 17037 11135 17095 11141
rect 17037 11132 17049 11135
rect 17000 11104 17049 11132
rect 17000 11092 17006 11104
rect 17037 11101 17049 11104
rect 17083 11101 17095 11135
rect 17586 11132 17592 11144
rect 17547 11104 17592 11132
rect 17037 11095 17095 11101
rect 17586 11092 17592 11104
rect 17644 11092 17650 11144
rect 18049 11135 18107 11141
rect 18049 11101 18061 11135
rect 18095 11101 18107 11135
rect 19978 11132 19984 11144
rect 19939 11104 19984 11132
rect 18049 11095 18107 11101
rect 4173 11067 4231 11073
rect 4173 11064 4185 11067
rect 4080 11036 4185 11064
rect 4173 11033 4185 11036
rect 4219 11033 4231 11067
rect 4173 11027 4231 11033
rect 5626 11024 5632 11076
rect 5684 11064 5690 11076
rect 5804 11067 5862 11073
rect 5804 11064 5816 11067
rect 5684 11036 5816 11064
rect 5684 11024 5690 11036
rect 5804 11033 5816 11036
rect 5850 11064 5862 11067
rect 9214 11064 9220 11076
rect 5850 11036 9220 11064
rect 5850 11033 5862 11036
rect 5804 11027 5862 11033
rect 9214 11024 9220 11036
rect 9272 11024 9278 11076
rect 12434 11064 12440 11076
rect 11716 11036 12440 11064
rect 3142 10956 3148 11008
rect 3200 10996 3206 11008
rect 3237 10999 3295 11005
rect 3237 10996 3249 10999
rect 3200 10968 3249 10996
rect 3200 10956 3206 10968
rect 3237 10965 3249 10968
rect 3283 10965 3295 10999
rect 4338 10996 4344 11008
rect 4299 10968 4344 10996
rect 3237 10959 3295 10965
rect 4338 10956 4344 10968
rect 4396 10956 4402 11008
rect 6914 10996 6920 11008
rect 6875 10968 6920 10996
rect 6914 10956 6920 10968
rect 6972 10956 6978 11008
rect 7098 10956 7104 11008
rect 7156 10996 7162 11008
rect 8846 10996 8852 11008
rect 7156 10968 8852 10996
rect 7156 10956 7162 10968
rect 8846 10956 8852 10968
rect 8904 10956 8910 11008
rect 8938 10956 8944 11008
rect 8996 10996 9002 11008
rect 9950 10996 9956 11008
rect 8996 10968 9956 10996
rect 8996 10956 9002 10968
rect 9950 10956 9956 10968
rect 10008 10956 10014 11008
rect 11716 11005 11744 11036
rect 12434 11024 12440 11036
rect 12492 11024 12498 11076
rect 12618 11064 12624 11076
rect 12579 11036 12624 11064
rect 12618 11024 12624 11036
rect 12676 11024 12682 11076
rect 13446 11064 13452 11076
rect 13407 11036 13452 11064
rect 13446 11024 13452 11036
rect 13504 11024 13510 11076
rect 16758 11064 16764 11076
rect 16719 11036 16764 11064
rect 16758 11024 16764 11036
rect 16816 11024 16822 11076
rect 16868 11064 16896 11092
rect 18064 11064 18092 11095
rect 19978 11092 19984 11104
rect 20036 11092 20042 11144
rect 20070 11092 20076 11144
rect 20128 11132 20134 11144
rect 20272 11141 20300 11172
rect 20364 11141 20392 11240
rect 20530 11141 20536 11144
rect 20257 11135 20315 11141
rect 20128 11104 20173 11132
rect 20128 11092 20134 11104
rect 20257 11101 20269 11135
rect 20303 11101 20315 11135
rect 20257 11095 20315 11101
rect 20349 11135 20407 11141
rect 20349 11101 20361 11135
rect 20395 11101 20407 11135
rect 20349 11095 20407 11101
rect 20487 11135 20536 11141
rect 20487 11101 20499 11135
rect 20533 11101 20536 11135
rect 20487 11095 20536 11101
rect 16868 11036 18092 11064
rect 18325 11067 18383 11073
rect 18325 11033 18337 11067
rect 18371 11064 18383 11067
rect 19886 11064 19892 11076
rect 18371 11036 19892 11064
rect 18371 11033 18383 11036
rect 18325 11027 18383 11033
rect 19886 11024 19892 11036
rect 19944 11024 19950 11076
rect 20272 11064 20300 11095
rect 20530 11092 20536 11095
rect 20588 11092 20594 11144
rect 21082 11132 21088 11144
rect 21043 11104 21088 11132
rect 21082 11092 21088 11104
rect 21140 11092 21146 11144
rect 21358 11132 21364 11144
rect 21319 11104 21364 11132
rect 21358 11092 21364 11104
rect 21416 11092 21422 11144
rect 22186 11132 22192 11144
rect 22147 11104 22192 11132
rect 22186 11092 22192 11104
rect 22244 11092 22250 11144
rect 22278 11092 22284 11144
rect 22336 11132 22342 11144
rect 22336 11104 22381 11132
rect 22336 11092 22342 11104
rect 22646 11092 22652 11144
rect 22704 11141 22710 11144
rect 22704 11135 22753 11141
rect 22704 11101 22707 11135
rect 22741 11132 22753 11135
rect 23492 11132 23520 11308
rect 25314 11296 25320 11308
rect 25372 11296 25378 11348
rect 31294 11296 31300 11348
rect 31352 11336 31358 11348
rect 31481 11339 31539 11345
rect 31481 11336 31493 11339
rect 31352 11308 31493 11336
rect 31352 11296 31358 11308
rect 31481 11305 31493 11308
rect 31527 11305 31539 11339
rect 31481 11299 31539 11305
rect 23934 11200 23940 11212
rect 23847 11172 23940 11200
rect 22741 11104 23520 11132
rect 22741 11101 22753 11104
rect 22704 11095 22753 11101
rect 22704 11092 22710 11095
rect 23566 11092 23572 11144
rect 23624 11132 23630 11144
rect 23860 11141 23888 11172
rect 23934 11160 23940 11172
rect 23992 11200 23998 11212
rect 24670 11200 24676 11212
rect 23992 11172 24676 11200
rect 23992 11160 23998 11172
rect 24670 11160 24676 11172
rect 24728 11160 24734 11212
rect 23845 11135 23903 11141
rect 23624 11104 23669 11132
rect 23624 11092 23630 11104
rect 23845 11101 23857 11135
rect 23891 11101 23903 11135
rect 25866 11132 25872 11144
rect 23845 11095 23903 11101
rect 23952 11104 25872 11132
rect 20272 11036 21128 11064
rect 11701 10999 11759 11005
rect 11701 10965 11713 10999
rect 11747 10965 11759 10999
rect 11701 10959 11759 10965
rect 12345 10999 12403 11005
rect 12345 10965 12357 10999
rect 12391 10996 12403 10999
rect 12710 10996 12716 11008
rect 12391 10968 12716 10996
rect 12391 10965 12403 10968
rect 12345 10959 12403 10965
rect 12710 10956 12716 10968
rect 12768 10956 12774 11008
rect 20625 10999 20683 11005
rect 20625 10965 20637 10999
rect 20671 10996 20683 10999
rect 20990 10996 20996 11008
rect 20671 10968 20996 10996
rect 20671 10965 20683 10968
rect 20625 10959 20683 10965
rect 20990 10956 20996 10968
rect 21048 10956 21054 11008
rect 21100 10996 21128 11036
rect 21174 11024 21180 11076
rect 21232 11064 21238 11076
rect 22465 11067 22523 11073
rect 22465 11064 22477 11067
rect 21232 11036 21277 11064
rect 22204 11036 22477 11064
rect 21232 11024 21238 11036
rect 22204 10996 22232 11036
rect 22465 11033 22477 11036
rect 22511 11033 22523 11067
rect 22465 11027 22523 11033
rect 22557 11067 22615 11073
rect 22557 11033 22569 11067
rect 22603 11064 22615 11067
rect 23474 11064 23480 11076
rect 22603 11036 23480 11064
rect 22603 11033 22615 11036
rect 22557 11027 22615 11033
rect 23474 11024 23480 11036
rect 23532 11024 23538 11076
rect 23661 11067 23719 11073
rect 23661 11033 23673 11067
rect 23707 11064 23719 11067
rect 23952 11064 23980 11104
rect 25866 11092 25872 11104
rect 25924 11092 25930 11144
rect 26050 11132 26056 11144
rect 26011 11104 26056 11132
rect 26050 11092 26056 11104
rect 26108 11092 26114 11144
rect 26602 11092 26608 11144
rect 26660 11132 26666 11144
rect 26786 11132 26792 11144
rect 26660 11104 26792 11132
rect 26660 11092 26666 11104
rect 26786 11092 26792 11104
rect 26844 11092 26850 11144
rect 29546 11092 29552 11144
rect 29604 11132 29610 11144
rect 29917 11135 29975 11141
rect 29917 11132 29929 11135
rect 29604 11104 29929 11132
rect 29604 11092 29610 11104
rect 29917 11101 29929 11104
rect 29963 11101 29975 11135
rect 30190 11132 30196 11144
rect 30151 11104 30196 11132
rect 29917 11095 29975 11101
rect 23707 11036 23980 11064
rect 24029 11067 24087 11073
rect 23707 11033 23719 11036
rect 23661 11027 23719 11033
rect 24029 11033 24041 11067
rect 24075 11064 24087 11067
rect 24854 11064 24860 11076
rect 24075 11036 24860 11064
rect 24075 11033 24087 11036
rect 24029 11027 24087 11033
rect 24854 11024 24860 11036
rect 24912 11024 24918 11076
rect 28074 11024 28080 11076
rect 28132 11064 28138 11076
rect 29454 11064 29460 11076
rect 28132 11036 29460 11064
rect 28132 11024 28138 11036
rect 29454 11024 29460 11036
rect 29512 11024 29518 11076
rect 29932 11064 29960 11095
rect 30190 11092 30196 11104
rect 30248 11092 30254 11144
rect 32306 11092 32312 11144
rect 32364 11132 32370 11144
rect 32861 11135 32919 11141
rect 32861 11132 32873 11135
rect 32364 11104 32873 11132
rect 32364 11092 32370 11104
rect 32861 11101 32873 11104
rect 32907 11101 32919 11135
rect 32861 11095 32919 11101
rect 30834 11064 30840 11076
rect 29932 11036 30840 11064
rect 30834 11024 30840 11036
rect 30892 11024 30898 11076
rect 31662 11024 31668 11076
rect 31720 11064 31726 11076
rect 32594 11067 32652 11073
rect 32594 11064 32606 11067
rect 31720 11036 32606 11064
rect 31720 11024 31726 11036
rect 32594 11033 32606 11036
rect 32640 11033 32652 11067
rect 32594 11027 32652 11033
rect 21100 10968 22232 10996
rect 26602 10956 26608 11008
rect 26660 10996 26666 11008
rect 27341 10999 27399 11005
rect 27341 10996 27353 10999
rect 26660 10968 27353 10996
rect 26660 10956 26666 10968
rect 27341 10965 27353 10968
rect 27387 10965 27399 10999
rect 29730 10996 29736 11008
rect 29691 10968 29736 10996
rect 27341 10959 27399 10965
rect 29730 10956 29736 10968
rect 29788 10956 29794 11008
rect 30098 10996 30104 11008
rect 30059 10968 30104 10996
rect 30098 10956 30104 10968
rect 30156 10956 30162 11008
rect 1104 10906 35027 10928
rect 1104 10854 9390 10906
rect 9442 10854 9454 10906
rect 9506 10854 9518 10906
rect 9570 10854 9582 10906
rect 9634 10854 9646 10906
rect 9698 10854 17831 10906
rect 17883 10854 17895 10906
rect 17947 10854 17959 10906
rect 18011 10854 18023 10906
rect 18075 10854 18087 10906
rect 18139 10854 26272 10906
rect 26324 10854 26336 10906
rect 26388 10854 26400 10906
rect 26452 10854 26464 10906
rect 26516 10854 26528 10906
rect 26580 10854 34713 10906
rect 34765 10854 34777 10906
rect 34829 10854 34841 10906
rect 34893 10854 34905 10906
rect 34957 10854 34969 10906
rect 35021 10854 35027 10906
rect 1104 10832 35027 10854
rect 4183 10795 4241 10801
rect 4183 10761 4195 10795
rect 4229 10792 4241 10795
rect 4338 10792 4344 10804
rect 4229 10764 4344 10792
rect 4229 10761 4241 10764
rect 4183 10755 4241 10761
rect 4338 10752 4344 10764
rect 4396 10752 4402 10804
rect 6638 10752 6644 10804
rect 6696 10792 6702 10804
rect 7837 10795 7895 10801
rect 6696 10764 7788 10792
rect 6696 10752 6702 10764
rect 3973 10727 4031 10733
rect 3973 10693 3985 10727
rect 4019 10693 4031 10727
rect 6730 10724 6736 10736
rect 6691 10696 6736 10724
rect 3973 10687 4031 10693
rect 2501 10659 2559 10665
rect 2501 10625 2513 10659
rect 2547 10656 2559 10659
rect 2682 10656 2688 10668
rect 2547 10628 2688 10656
rect 2547 10625 2559 10628
rect 2501 10619 2559 10625
rect 2682 10616 2688 10628
rect 2740 10616 2746 10668
rect 3142 10656 3148 10668
rect 3103 10628 3148 10656
rect 3142 10616 3148 10628
rect 3200 10616 3206 10668
rect 3329 10659 3387 10665
rect 3329 10625 3341 10659
rect 3375 10656 3387 10659
rect 3988 10656 4016 10687
rect 6730 10684 6736 10696
rect 6788 10684 6794 10736
rect 6914 10684 6920 10736
rect 6972 10724 6978 10736
rect 7009 10727 7067 10733
rect 7009 10724 7021 10727
rect 6972 10696 7021 10724
rect 6972 10684 6978 10696
rect 7009 10693 7021 10696
rect 7055 10693 7067 10727
rect 7466 10724 7472 10736
rect 7427 10696 7472 10724
rect 7009 10687 7067 10693
rect 7466 10684 7472 10696
rect 7524 10684 7530 10736
rect 7760 10724 7788 10764
rect 7837 10761 7849 10795
rect 7883 10792 7895 10795
rect 8202 10792 8208 10804
rect 7883 10764 8208 10792
rect 7883 10761 7895 10764
rect 7837 10755 7895 10761
rect 8202 10752 8208 10764
rect 8260 10752 8266 10804
rect 8478 10752 8484 10804
rect 8536 10792 8542 10804
rect 8757 10795 8815 10801
rect 8757 10792 8769 10795
rect 8536 10764 8769 10792
rect 8536 10752 8542 10764
rect 8757 10761 8769 10764
rect 8803 10761 8815 10795
rect 8757 10755 8815 10761
rect 8938 10752 8944 10804
rect 8996 10792 9002 10804
rect 8996 10764 9628 10792
rect 8996 10752 9002 10764
rect 9140 10733 9168 10764
rect 9125 10727 9183 10733
rect 7760 10696 8616 10724
rect 4246 10656 4252 10668
rect 3375 10628 4252 10656
rect 3375 10625 3387 10628
rect 3329 10619 3387 10625
rect 4246 10616 4252 10628
rect 4304 10616 4310 10668
rect 7098 10656 7104 10668
rect 7059 10628 7104 10656
rect 7098 10616 7104 10628
rect 7156 10616 7162 10668
rect 2409 10591 2467 10597
rect 2409 10557 2421 10591
rect 2455 10588 2467 10591
rect 2958 10588 2964 10600
rect 2455 10560 2964 10588
rect 2455 10557 2467 10560
rect 2409 10551 2467 10557
rect 2958 10548 2964 10560
rect 3016 10548 3022 10600
rect 3237 10591 3295 10597
rect 3237 10557 3249 10591
rect 3283 10557 3295 10591
rect 3418 10588 3424 10600
rect 3379 10560 3424 10588
rect 3237 10551 3295 10557
rect 2130 10480 2136 10532
rect 2188 10520 2194 10532
rect 3252 10520 3280 10551
rect 3418 10548 3424 10560
rect 3476 10548 3482 10600
rect 6638 10548 6644 10600
rect 6696 10548 6702 10600
rect 8588 10520 8616 10696
rect 9125 10693 9137 10727
rect 9171 10693 9183 10727
rect 9125 10687 9183 10693
rect 9214 10684 9220 10736
rect 9272 10724 9278 10736
rect 9493 10727 9551 10733
rect 9493 10724 9505 10727
rect 9272 10696 9505 10724
rect 9272 10684 9278 10696
rect 9493 10693 9505 10696
rect 9539 10693 9551 10727
rect 9600 10724 9628 10764
rect 9766 10752 9772 10804
rect 9824 10792 9830 10804
rect 9861 10795 9919 10801
rect 9861 10792 9873 10795
rect 9824 10764 9873 10792
rect 9824 10752 9830 10764
rect 9861 10761 9873 10764
rect 9907 10761 9919 10795
rect 9861 10755 9919 10761
rect 9950 10752 9956 10804
rect 10008 10792 10014 10804
rect 13633 10795 13691 10801
rect 13633 10792 13645 10795
rect 10008 10764 13645 10792
rect 10008 10752 10014 10764
rect 13633 10761 13645 10764
rect 13679 10761 13691 10795
rect 19702 10792 19708 10804
rect 19663 10764 19708 10792
rect 13633 10755 13691 10761
rect 19702 10752 19708 10764
rect 19760 10752 19766 10804
rect 20438 10792 20444 10804
rect 20399 10764 20444 10792
rect 20438 10752 20444 10764
rect 20496 10752 20502 10804
rect 20714 10752 20720 10804
rect 20772 10792 20778 10804
rect 20809 10795 20867 10801
rect 20809 10792 20821 10795
rect 20772 10764 20821 10792
rect 20772 10752 20778 10764
rect 20809 10761 20821 10764
rect 20855 10761 20867 10795
rect 20809 10755 20867 10761
rect 22186 10752 22192 10804
rect 22244 10792 22250 10804
rect 22373 10795 22431 10801
rect 22373 10792 22385 10795
rect 22244 10764 22385 10792
rect 22244 10752 22250 10764
rect 22373 10761 22385 10764
rect 22419 10761 22431 10795
rect 23566 10792 23572 10804
rect 22373 10755 22431 10761
rect 22572 10764 23572 10792
rect 11882 10724 11888 10736
rect 9600 10696 11888 10724
rect 9493 10687 9551 10693
rect 11882 10684 11888 10696
rect 11940 10724 11946 10736
rect 12342 10724 12348 10736
rect 11940 10696 12348 10724
rect 11940 10684 11946 10696
rect 12342 10684 12348 10696
rect 12400 10684 12406 10736
rect 12526 10724 12532 10736
rect 12487 10696 12532 10724
rect 12526 10684 12532 10696
rect 12584 10684 12590 10736
rect 12894 10724 12900 10736
rect 12855 10696 12900 10724
rect 12894 10684 12900 10696
rect 12952 10684 12958 10736
rect 13265 10727 13323 10733
rect 13265 10693 13277 10727
rect 13311 10724 13323 10727
rect 13998 10724 14004 10736
rect 13311 10696 14004 10724
rect 13311 10693 13323 10696
rect 13265 10687 13323 10693
rect 13998 10684 14004 10696
rect 14056 10684 14062 10736
rect 18230 10724 18236 10736
rect 18191 10696 18236 10724
rect 18230 10684 18236 10696
rect 18288 10684 18294 10736
rect 19886 10684 19892 10736
rect 19944 10724 19950 10736
rect 22572 10724 22600 10764
rect 23566 10752 23572 10764
rect 23624 10752 23630 10804
rect 25866 10752 25872 10804
rect 25924 10792 25930 10804
rect 25961 10795 26019 10801
rect 25961 10792 25973 10795
rect 25924 10764 25973 10792
rect 25924 10752 25930 10764
rect 25961 10761 25973 10764
rect 26007 10761 26019 10795
rect 25961 10755 26019 10761
rect 28721 10795 28779 10801
rect 28721 10761 28733 10795
rect 28767 10792 28779 10795
rect 28994 10792 29000 10804
rect 28767 10764 29000 10792
rect 28767 10761 28779 10764
rect 28721 10755 28779 10761
rect 28994 10752 29000 10764
rect 29052 10792 29058 10804
rect 30098 10792 30104 10804
rect 29052 10764 30104 10792
rect 29052 10752 29058 10764
rect 30098 10752 30104 10764
rect 30156 10752 30162 10804
rect 33686 10792 33692 10804
rect 33647 10764 33692 10792
rect 33686 10752 33692 10764
rect 33744 10752 33750 10804
rect 19944 10696 22600 10724
rect 19944 10684 19950 10696
rect 9030 10616 9036 10668
rect 9088 10656 9094 10668
rect 9088 10628 9133 10656
rect 9088 10616 9094 10628
rect 12434 10616 12440 10668
rect 12492 10656 12498 10668
rect 12805 10659 12863 10665
rect 12805 10656 12817 10659
rect 12492 10628 12817 10656
rect 12492 10616 12498 10628
rect 12805 10625 12817 10628
rect 12851 10625 12863 10659
rect 12805 10619 12863 10625
rect 19334 10616 19340 10668
rect 19392 10656 19398 10668
rect 20625 10659 20683 10665
rect 20625 10656 20637 10659
rect 19392 10628 20637 10656
rect 19392 10616 19398 10628
rect 20625 10625 20637 10628
rect 20671 10625 20683 10659
rect 20625 10619 20683 10625
rect 20901 10659 20959 10665
rect 20901 10625 20913 10659
rect 20947 10656 20959 10659
rect 22370 10656 22376 10668
rect 20947 10628 22376 10656
rect 20947 10625 20959 10628
rect 20901 10619 20959 10625
rect 11146 10548 11152 10600
rect 11204 10588 11210 10600
rect 12158 10588 12164 10600
rect 11204 10560 12164 10588
rect 11204 10548 11210 10560
rect 12158 10548 12164 10560
rect 12216 10588 12222 10600
rect 20640 10588 20668 10619
rect 22370 10616 22376 10628
rect 22428 10616 22434 10668
rect 22572 10665 22600 10696
rect 22741 10727 22799 10733
rect 22741 10693 22753 10727
rect 22787 10724 22799 10727
rect 23750 10724 23756 10736
rect 22787 10696 23756 10724
rect 22787 10693 22799 10696
rect 22741 10687 22799 10693
rect 23750 10684 23756 10696
rect 23808 10684 23814 10736
rect 24854 10733 24860 10736
rect 24848 10724 24860 10733
rect 24815 10696 24860 10724
rect 24848 10687 24860 10696
rect 24854 10684 24860 10687
rect 24912 10684 24918 10736
rect 28074 10684 28080 10736
rect 28132 10724 28138 10736
rect 29365 10727 29423 10733
rect 29365 10724 29377 10727
rect 28132 10696 29377 10724
rect 28132 10684 28138 10696
rect 29365 10693 29377 10696
rect 29411 10693 29423 10727
rect 29365 10687 29423 10693
rect 29454 10684 29460 10736
rect 29512 10724 29518 10736
rect 29549 10727 29607 10733
rect 29549 10724 29561 10727
rect 29512 10696 29561 10724
rect 29512 10684 29518 10696
rect 29549 10693 29561 10696
rect 29595 10693 29607 10727
rect 29549 10687 29607 10693
rect 22557 10659 22615 10665
rect 22557 10625 22569 10659
rect 22603 10625 22615 10659
rect 22557 10619 22615 10625
rect 22649 10659 22707 10665
rect 22649 10625 22661 10659
rect 22695 10625 22707 10659
rect 22922 10656 22928 10668
rect 22883 10628 22928 10656
rect 22649 10619 22707 10625
rect 22664 10588 22692 10619
rect 22922 10616 22928 10628
rect 22980 10616 22986 10668
rect 27608 10659 27666 10665
rect 27608 10625 27620 10659
rect 27654 10656 27666 10659
rect 29730 10656 29736 10668
rect 27654 10628 29736 10656
rect 27654 10625 27666 10628
rect 27608 10619 27666 10625
rect 29730 10616 29736 10628
rect 29788 10616 29794 10668
rect 32398 10616 32404 10668
rect 32456 10656 32462 10668
rect 32565 10659 32623 10665
rect 32565 10656 32577 10659
rect 32456 10628 32577 10656
rect 32456 10616 32462 10628
rect 32565 10625 32577 10628
rect 32611 10625 32623 10659
rect 32565 10619 32623 10625
rect 23474 10588 23480 10600
rect 12216 10560 12374 10588
rect 20640 10560 22094 10588
rect 22664 10560 23480 10588
rect 12216 10548 12222 10560
rect 8662 10520 8668 10532
rect 2188 10492 4108 10520
rect 8588 10492 8668 10520
rect 2188 10480 2194 10492
rect 4080 10464 4108 10492
rect 8662 10480 8668 10492
rect 8720 10480 8726 10532
rect 22066 10520 22094 10560
rect 23474 10548 23480 10560
rect 23532 10548 23538 10600
rect 24578 10588 24584 10600
rect 24539 10560 24584 10588
rect 24578 10548 24584 10560
rect 24636 10548 24642 10600
rect 27338 10588 27344 10600
rect 27299 10560 27344 10588
rect 27338 10548 27344 10560
rect 27396 10548 27402 10600
rect 32306 10588 32312 10600
rect 32267 10560 32312 10588
rect 32306 10548 32312 10560
rect 32364 10548 32370 10600
rect 22646 10520 22652 10532
rect 22066 10492 22652 10520
rect 22646 10480 22652 10492
rect 22704 10480 22710 10532
rect 2866 10412 2872 10464
rect 2924 10452 2930 10464
rect 2961 10455 3019 10461
rect 2961 10452 2973 10455
rect 2924 10424 2973 10452
rect 2924 10412 2930 10424
rect 2961 10421 2973 10424
rect 3007 10421 3019 10455
rect 2961 10415 3019 10421
rect 4062 10412 4068 10464
rect 4120 10452 4126 10464
rect 4157 10455 4215 10461
rect 4157 10452 4169 10455
rect 4120 10424 4169 10452
rect 4120 10412 4126 10424
rect 4157 10421 4169 10424
rect 4203 10421 4215 10455
rect 4157 10415 4215 10421
rect 4341 10455 4399 10461
rect 4341 10421 4353 10455
rect 4387 10452 4399 10455
rect 5534 10452 5540 10464
rect 4387 10424 5540 10452
rect 4387 10421 4399 10424
rect 4341 10415 4399 10421
rect 5534 10412 5540 10424
rect 5592 10412 5598 10464
rect 7926 10412 7932 10464
rect 7984 10452 7990 10464
rect 8021 10455 8079 10461
rect 8021 10452 8033 10455
rect 7984 10424 8033 10452
rect 7984 10412 7990 10424
rect 8021 10421 8033 10424
rect 8067 10421 8079 10455
rect 10042 10452 10048 10464
rect 10003 10424 10048 10452
rect 8021 10415 8079 10421
rect 10042 10412 10048 10424
rect 10100 10412 10106 10464
rect 13817 10455 13875 10461
rect 13817 10421 13829 10455
rect 13863 10452 13875 10455
rect 14366 10452 14372 10464
rect 13863 10424 14372 10452
rect 13863 10421 13875 10424
rect 13817 10415 13875 10421
rect 14366 10412 14372 10424
rect 14424 10412 14430 10464
rect 29362 10412 29368 10464
rect 29420 10452 29426 10464
rect 29549 10455 29607 10461
rect 29549 10452 29561 10455
rect 29420 10424 29561 10452
rect 29420 10412 29426 10424
rect 29549 10421 29561 10424
rect 29595 10421 29607 10455
rect 29549 10415 29607 10421
rect 29733 10455 29791 10461
rect 29733 10421 29745 10455
rect 29779 10452 29791 10455
rect 31018 10452 31024 10464
rect 29779 10424 31024 10452
rect 29779 10421 29791 10424
rect 29733 10415 29791 10421
rect 31018 10412 31024 10424
rect 31076 10412 31082 10464
rect 1104 10362 34868 10384
rect 1104 10310 5170 10362
rect 5222 10310 5234 10362
rect 5286 10310 5298 10362
rect 5350 10310 5362 10362
rect 5414 10310 5426 10362
rect 5478 10310 13611 10362
rect 13663 10310 13675 10362
rect 13727 10310 13739 10362
rect 13791 10310 13803 10362
rect 13855 10310 13867 10362
rect 13919 10310 22052 10362
rect 22104 10310 22116 10362
rect 22168 10310 22180 10362
rect 22232 10310 22244 10362
rect 22296 10310 22308 10362
rect 22360 10310 30493 10362
rect 30545 10310 30557 10362
rect 30609 10310 30621 10362
rect 30673 10310 30685 10362
rect 30737 10310 30749 10362
rect 30801 10310 34868 10362
rect 1104 10288 34868 10310
rect 2682 10248 2688 10260
rect 2643 10220 2688 10248
rect 2682 10208 2688 10220
rect 2740 10248 2746 10260
rect 3050 10248 3056 10260
rect 2740 10220 3056 10248
rect 2740 10208 2746 10220
rect 3050 10208 3056 10220
rect 3108 10208 3114 10260
rect 4154 10248 4160 10260
rect 4115 10220 4160 10248
rect 4154 10208 4160 10220
rect 4212 10208 4218 10260
rect 5534 10248 5540 10260
rect 5368 10220 5540 10248
rect 2866 10112 2872 10124
rect 2056 10084 2872 10112
rect 1762 10044 1768 10056
rect 1723 10016 1768 10044
rect 1762 10004 1768 10016
rect 1820 10004 1826 10056
rect 2056 10053 2084 10084
rect 2866 10072 2872 10084
rect 2924 10072 2930 10124
rect 3234 10112 3240 10124
rect 3195 10084 3240 10112
rect 3234 10072 3240 10084
rect 3292 10072 3298 10124
rect 3326 10072 3332 10124
rect 3384 10112 3390 10124
rect 5368 10121 5396 10220
rect 5534 10208 5540 10220
rect 5592 10208 5598 10260
rect 6730 10248 6736 10260
rect 6691 10220 6736 10248
rect 6730 10208 6736 10220
rect 6788 10208 6794 10260
rect 8573 10251 8631 10257
rect 8573 10217 8585 10251
rect 8619 10248 8631 10251
rect 9030 10248 9036 10260
rect 8619 10220 9036 10248
rect 8619 10217 8631 10220
rect 8573 10211 8631 10217
rect 9030 10208 9036 10220
rect 9088 10208 9094 10260
rect 12618 10248 12624 10260
rect 12579 10220 12624 10248
rect 12618 10208 12624 10220
rect 12676 10208 12682 10260
rect 21269 10251 21327 10257
rect 21269 10217 21281 10251
rect 21315 10248 21327 10251
rect 23842 10248 23848 10260
rect 21315 10220 23848 10248
rect 21315 10217 21327 10220
rect 21269 10211 21327 10217
rect 23842 10208 23848 10220
rect 23900 10248 23906 10260
rect 24578 10248 24584 10260
rect 23900 10220 24584 10248
rect 23900 10208 23906 10220
rect 24578 10208 24584 10220
rect 24636 10208 24642 10260
rect 24949 10251 25007 10257
rect 24949 10217 24961 10251
rect 24995 10248 25007 10251
rect 25406 10248 25412 10260
rect 24995 10220 25412 10248
rect 24995 10217 25007 10220
rect 24949 10211 25007 10217
rect 25406 10208 25412 10220
rect 25464 10208 25470 10260
rect 27338 10248 27344 10260
rect 27299 10220 27344 10248
rect 27338 10208 27344 10220
rect 27396 10208 27402 10260
rect 28258 10248 28264 10260
rect 28219 10220 28264 10248
rect 28258 10208 28264 10220
rect 28316 10208 28322 10260
rect 31665 10251 31723 10257
rect 31665 10217 31677 10251
rect 31711 10248 31723 10251
rect 32306 10248 32312 10260
rect 31711 10220 32312 10248
rect 31711 10217 31723 10220
rect 31665 10211 31723 10217
rect 32306 10208 32312 10220
rect 32364 10208 32370 10260
rect 8662 10140 8668 10192
rect 8720 10180 8726 10192
rect 11146 10180 11152 10192
rect 8720 10152 11152 10180
rect 8720 10140 8726 10152
rect 11146 10140 11152 10152
rect 11204 10140 11210 10192
rect 28459 10152 30052 10180
rect 5353 10115 5411 10121
rect 3384 10084 3429 10112
rect 3384 10072 3390 10084
rect 5353 10081 5365 10115
rect 5399 10081 5411 10115
rect 5353 10075 5411 10081
rect 10410 10072 10416 10124
rect 10468 10112 10474 10124
rect 11241 10115 11299 10121
rect 11241 10112 11253 10115
rect 10468 10084 11253 10112
rect 10468 10072 10474 10084
rect 11241 10081 11253 10084
rect 11287 10081 11299 10115
rect 11241 10075 11299 10081
rect 22572 10084 26096 10112
rect 2041 10047 2099 10053
rect 2041 10013 2053 10047
rect 2087 10013 2099 10047
rect 2041 10007 2099 10013
rect 2961 10047 3019 10053
rect 2961 10013 2973 10047
rect 3007 10013 3019 10047
rect 2961 10007 3019 10013
rect 1857 9979 1915 9985
rect 1857 9945 1869 9979
rect 1903 9976 1915 9979
rect 2976 9976 3004 10007
rect 4338 10004 4344 10056
rect 4396 10004 4402 10056
rect 4433 10047 4491 10053
rect 4433 10013 4445 10047
rect 4479 10044 4491 10047
rect 6086 10044 6092 10056
rect 4479 10016 6092 10044
rect 4479 10013 4491 10016
rect 4433 10007 4491 10013
rect 6086 10004 6092 10016
rect 6144 10044 6150 10056
rect 7466 10053 7472 10056
rect 7193 10047 7251 10053
rect 7193 10044 7205 10047
rect 6144 10016 7205 10044
rect 6144 10004 6150 10016
rect 7193 10013 7205 10016
rect 7239 10013 7251 10047
rect 7460 10044 7472 10053
rect 7427 10016 7472 10044
rect 7193 10007 7251 10013
rect 7460 10007 7472 10016
rect 3973 9979 4031 9985
rect 3973 9976 3985 9979
rect 1903 9948 2774 9976
rect 2976 9948 3985 9976
rect 1903 9945 1915 9948
rect 1857 9939 1915 9945
rect 2130 9868 2136 9920
rect 2188 9908 2194 9920
rect 2225 9911 2283 9917
rect 2225 9908 2237 9911
rect 2188 9880 2237 9908
rect 2188 9868 2194 9880
rect 2225 9877 2237 9880
rect 2271 9877 2283 9911
rect 2746 9908 2774 9948
rect 3973 9945 3985 9948
rect 4019 9945 4031 9979
rect 3973 9939 4031 9945
rect 4157 9979 4215 9985
rect 4157 9945 4169 9979
rect 4203 9976 4215 9979
rect 4356 9976 4384 10004
rect 5626 9985 5632 9988
rect 5620 9976 5632 9985
rect 4203 9948 4384 9976
rect 5587 9948 5632 9976
rect 4203 9945 4215 9948
rect 4157 9939 4215 9945
rect 5620 9939 5632 9948
rect 2958 9908 2964 9920
rect 2746 9880 2964 9908
rect 2225 9871 2283 9877
rect 2958 9868 2964 9880
rect 3016 9868 3022 9920
rect 3050 9868 3056 9920
rect 3108 9908 3114 9920
rect 3988 9908 4016 9939
rect 5626 9936 5632 9939
rect 5684 9936 5690 9988
rect 7208 9976 7236 10007
rect 7466 10004 7472 10007
rect 7524 10004 7530 10056
rect 10428 9976 10456 10072
rect 22572 10053 22600 10084
rect 22557 10047 22615 10053
rect 22557 10013 22569 10047
rect 22603 10013 22615 10047
rect 22557 10007 22615 10013
rect 24762 10004 24768 10056
rect 24820 10044 24826 10056
rect 25087 10047 25145 10053
rect 25087 10044 25099 10047
rect 24820 10016 25099 10044
rect 24820 10004 24826 10016
rect 25087 10013 25099 10016
rect 25133 10013 25145 10047
rect 25314 10044 25320 10056
rect 25275 10016 25320 10044
rect 25087 10007 25145 10013
rect 25314 10004 25320 10016
rect 25372 10004 25378 10056
rect 26068 10053 26096 10084
rect 25500 10047 25558 10053
rect 25500 10013 25512 10047
rect 25546 10013 25558 10047
rect 25500 10007 25558 10013
rect 25593 10047 25651 10053
rect 25593 10013 25605 10047
rect 25639 10044 25651 10047
rect 26053 10047 26111 10053
rect 25639 10016 26004 10044
rect 25639 10013 25651 10016
rect 25593 10007 25651 10013
rect 7208 9948 10456 9976
rect 11508 9979 11566 9985
rect 11508 9945 11520 9979
rect 11554 9976 11566 9979
rect 11790 9976 11796 9988
rect 11554 9948 11796 9976
rect 11554 9945 11566 9948
rect 11508 9939 11566 9945
rect 11790 9936 11796 9948
rect 11848 9976 11854 9988
rect 12066 9976 12072 9988
rect 11848 9948 12072 9976
rect 11848 9936 11854 9948
rect 12066 9936 12072 9948
rect 12124 9936 12130 9988
rect 25222 9976 25228 9988
rect 25183 9948 25228 9976
rect 25222 9936 25228 9948
rect 25280 9936 25286 9988
rect 25516 9976 25544 10007
rect 25866 9976 25872 9988
rect 25516 9948 25872 9976
rect 25866 9936 25872 9948
rect 25924 9936 25930 9988
rect 25976 9976 26004 10016
rect 26053 10013 26065 10047
rect 26099 10044 26111 10047
rect 26602 10044 26608 10056
rect 26099 10016 26608 10044
rect 26099 10013 26111 10016
rect 26053 10007 26111 10013
rect 26602 10004 26608 10016
rect 26660 10004 26666 10056
rect 28459 10053 28487 10152
rect 28994 10112 29000 10124
rect 28828 10084 29000 10112
rect 28401 10047 28487 10053
rect 28401 10013 28413 10047
rect 28447 10016 28487 10047
rect 28626 10044 28632 10056
rect 28587 10016 28632 10044
rect 28447 10013 28459 10016
rect 28401 10007 28459 10013
rect 25976 9948 26096 9976
rect 4246 9908 4252 9920
rect 3108 9880 3153 9908
rect 3988 9880 4252 9908
rect 3108 9868 3114 9880
rect 4246 9868 4252 9880
rect 4304 9868 4310 9920
rect 7834 9868 7840 9920
rect 7892 9908 7898 9920
rect 13354 9908 13360 9920
rect 7892 9880 13360 9908
rect 7892 9868 7898 9880
rect 13354 9868 13360 9880
rect 13412 9868 13418 9920
rect 26068 9908 26096 9948
rect 27890 9936 27896 9988
rect 27948 9976 27954 9988
rect 28258 9976 28264 9988
rect 27948 9948 28264 9976
rect 27948 9936 27954 9948
rect 28258 9936 28264 9948
rect 28316 9976 28322 9988
rect 28414 9976 28442 10007
rect 28626 10004 28632 10016
rect 28684 10004 28690 10056
rect 28828 10053 28856 10084
rect 28994 10072 29000 10084
rect 29052 10072 29058 10124
rect 28812 10047 28870 10053
rect 28812 10013 28824 10047
rect 28858 10013 28870 10047
rect 28812 10007 28870 10013
rect 28902 10004 28908 10056
rect 28960 10044 28966 10056
rect 28960 10016 29005 10044
rect 28960 10004 28966 10016
rect 29454 10004 29460 10056
rect 29512 10044 29518 10056
rect 29917 10047 29975 10053
rect 29917 10044 29929 10047
rect 29512 10016 29929 10044
rect 29512 10004 29518 10016
rect 29917 10013 29929 10016
rect 29963 10013 29975 10047
rect 30024 10044 30052 10152
rect 30101 10047 30159 10053
rect 30101 10044 30113 10047
rect 30024 10016 30113 10044
rect 29917 10007 29975 10013
rect 30101 10013 30113 10016
rect 30147 10013 30159 10047
rect 30282 10044 30288 10056
rect 30243 10016 30288 10044
rect 30101 10007 30159 10013
rect 30282 10004 30288 10016
rect 30340 10004 30346 10056
rect 33410 10044 33416 10056
rect 33371 10016 33416 10044
rect 33410 10004 33416 10016
rect 33468 10004 33474 10056
rect 33594 10004 33600 10056
rect 33652 10044 33658 10056
rect 33689 10047 33747 10053
rect 33689 10044 33701 10047
rect 33652 10016 33701 10044
rect 33652 10004 33658 10016
rect 33689 10013 33701 10016
rect 33735 10013 33747 10047
rect 33689 10007 33747 10013
rect 28534 9976 28540 9988
rect 28316 9948 28442 9976
rect 28495 9948 28540 9976
rect 28316 9936 28322 9948
rect 28534 9936 28540 9948
rect 28592 9936 28598 9988
rect 30009 9979 30067 9985
rect 30009 9945 30021 9979
rect 30055 9945 30067 9979
rect 30009 9939 30067 9945
rect 32953 9979 33011 9985
rect 32953 9945 32965 9979
rect 32999 9976 33011 9979
rect 32999 9948 33732 9976
rect 32999 9945 33011 9948
rect 32953 9939 33011 9945
rect 29733 9911 29791 9917
rect 29733 9908 29745 9911
rect 26068 9880 29745 9908
rect 29733 9877 29745 9880
rect 29779 9877 29791 9911
rect 30024 9908 30052 9939
rect 33704 9920 33732 9948
rect 32306 9908 32312 9920
rect 30024 9880 32312 9908
rect 29733 9871 29791 9877
rect 32306 9868 32312 9880
rect 32364 9908 32370 9920
rect 33505 9911 33563 9917
rect 33505 9908 33517 9911
rect 32364 9880 33517 9908
rect 32364 9868 32370 9880
rect 33505 9877 33517 9880
rect 33551 9877 33563 9911
rect 33505 9871 33563 9877
rect 33686 9868 33692 9920
rect 33744 9868 33750 9920
rect 33870 9908 33876 9920
rect 33831 9880 33876 9908
rect 33870 9868 33876 9880
rect 33928 9868 33934 9920
rect 1104 9818 35027 9840
rect 1104 9766 9390 9818
rect 9442 9766 9454 9818
rect 9506 9766 9518 9818
rect 9570 9766 9582 9818
rect 9634 9766 9646 9818
rect 9698 9766 17831 9818
rect 17883 9766 17895 9818
rect 17947 9766 17959 9818
rect 18011 9766 18023 9818
rect 18075 9766 18087 9818
rect 18139 9766 26272 9818
rect 26324 9766 26336 9818
rect 26388 9766 26400 9818
rect 26452 9766 26464 9818
rect 26516 9766 26528 9818
rect 26580 9766 34713 9818
rect 34765 9766 34777 9818
rect 34829 9766 34841 9818
rect 34893 9766 34905 9818
rect 34957 9766 34969 9818
rect 35021 9766 35027 9818
rect 1104 9744 35027 9766
rect 1762 9664 1768 9716
rect 1820 9704 1826 9716
rect 1949 9707 2007 9713
rect 1949 9704 1961 9707
rect 1820 9676 1961 9704
rect 1820 9664 1826 9676
rect 1949 9673 1961 9676
rect 1995 9673 2007 9707
rect 4154 9704 4160 9716
rect 4115 9676 4160 9704
rect 1949 9667 2007 9673
rect 4154 9664 4160 9676
rect 4212 9664 4218 9716
rect 4246 9664 4252 9716
rect 4304 9704 4310 9716
rect 4801 9707 4859 9713
rect 4801 9704 4813 9707
rect 4304 9676 4813 9704
rect 4304 9664 4310 9676
rect 4801 9673 4813 9676
rect 4847 9673 4859 9707
rect 8478 9704 8484 9716
rect 8439 9676 8484 9704
rect 4801 9667 4859 9673
rect 8478 9664 8484 9676
rect 8536 9664 8542 9716
rect 10042 9664 10048 9716
rect 10100 9704 10106 9716
rect 17034 9704 17040 9716
rect 10100 9676 17040 9704
rect 10100 9664 10106 9676
rect 17034 9664 17040 9676
rect 17092 9664 17098 9716
rect 27709 9707 27767 9713
rect 19628 9676 19840 9704
rect 2317 9639 2375 9645
rect 2317 9605 2329 9639
rect 2363 9636 2375 9639
rect 3237 9639 3295 9645
rect 2363 9608 2774 9636
rect 2363 9605 2375 9608
rect 2317 9599 2375 9605
rect 2130 9568 2136 9580
rect 2091 9540 2136 9568
rect 2130 9528 2136 9540
rect 2188 9528 2194 9580
rect 2409 9571 2467 9577
rect 2409 9537 2421 9571
rect 2455 9537 2467 9571
rect 2746 9568 2774 9608
rect 3237 9605 3249 9639
rect 3283 9636 3295 9639
rect 4172 9636 4200 9664
rect 3283 9608 4200 9636
rect 7368 9639 7426 9645
rect 3283 9605 3295 9608
rect 3237 9599 3295 9605
rect 7368 9605 7380 9639
rect 7414 9636 7426 9639
rect 7466 9636 7472 9648
rect 7414 9608 7472 9636
rect 7414 9605 7426 9608
rect 7368 9599 7426 9605
rect 7466 9596 7472 9608
rect 7524 9596 7530 9648
rect 16390 9596 16396 9648
rect 16448 9636 16454 9648
rect 17221 9639 17279 9645
rect 17221 9636 17233 9639
rect 16448 9608 17233 9636
rect 16448 9596 16454 9608
rect 17221 9605 17233 9608
rect 17267 9636 17279 9639
rect 19628 9636 19656 9676
rect 17267 9608 19656 9636
rect 19812 9636 19840 9676
rect 27709 9673 27721 9707
rect 27755 9704 27767 9707
rect 28902 9704 28908 9716
rect 27755 9676 28908 9704
rect 27755 9673 27767 9676
rect 27709 9667 27767 9673
rect 28902 9664 28908 9676
rect 28960 9664 28966 9716
rect 31386 9704 31392 9716
rect 30944 9676 31392 9704
rect 20993 9639 21051 9645
rect 19812 9608 20760 9636
rect 17267 9605 17279 9608
rect 17221 9599 17279 9605
rect 3329 9571 3387 9577
rect 3329 9568 3341 9571
rect 2746 9540 3341 9568
rect 2409 9531 2467 9537
rect 3329 9537 3341 9540
rect 3375 9568 3387 9571
rect 4062 9568 4068 9580
rect 3375 9540 3556 9568
rect 4023 9540 4068 9568
rect 3375 9537 3387 9540
rect 3329 9531 3387 9537
rect 2424 9500 2452 9531
rect 3142 9500 3148 9512
rect 2424 9472 3148 9500
rect 3142 9460 3148 9472
rect 3200 9500 3206 9512
rect 3421 9503 3479 9509
rect 3421 9500 3433 9503
rect 3200 9472 3433 9500
rect 3200 9460 3206 9472
rect 3421 9469 3433 9472
rect 3467 9469 3479 9503
rect 3528 9500 3556 9540
rect 4062 9528 4068 9540
rect 4120 9528 4126 9580
rect 4706 9568 4712 9580
rect 4667 9540 4712 9568
rect 4706 9528 4712 9540
rect 4764 9528 4770 9580
rect 5534 9528 5540 9580
rect 5592 9568 5598 9580
rect 6822 9568 6828 9580
rect 5592 9540 6828 9568
rect 5592 9528 5598 9540
rect 6822 9528 6828 9540
rect 6880 9568 6886 9580
rect 7101 9571 7159 9577
rect 7101 9568 7113 9571
rect 6880 9540 7113 9568
rect 6880 9528 6886 9540
rect 7101 9537 7113 9540
rect 7147 9537 7159 9571
rect 7101 9531 7159 9537
rect 11790 9528 11796 9580
rect 11848 9568 11854 9580
rect 11957 9571 12015 9577
rect 11957 9568 11969 9571
rect 11848 9540 11969 9568
rect 11848 9528 11854 9540
rect 11957 9537 11969 9540
rect 12003 9537 12015 9571
rect 11957 9531 12015 9537
rect 17037 9571 17095 9577
rect 17037 9537 17049 9571
rect 17083 9568 17095 9571
rect 17126 9568 17132 9580
rect 17083 9540 17132 9568
rect 17083 9537 17095 9540
rect 17037 9531 17095 9537
rect 17126 9528 17132 9540
rect 17184 9528 17190 9580
rect 17310 9568 17316 9580
rect 17271 9540 17316 9568
rect 17310 9528 17316 9540
rect 17368 9528 17374 9580
rect 17586 9528 17592 9580
rect 17644 9568 17650 9580
rect 18233 9571 18291 9577
rect 18233 9568 18245 9571
rect 17644 9540 18245 9568
rect 17644 9528 17650 9540
rect 18233 9537 18245 9540
rect 18279 9537 18291 9571
rect 18414 9568 18420 9580
rect 18327 9540 18420 9568
rect 18233 9531 18291 9537
rect 4724 9500 4752 9528
rect 3528 9472 4752 9500
rect 3421 9463 3479 9469
rect 10778 9460 10784 9512
rect 10836 9500 10842 9512
rect 11701 9503 11759 9509
rect 11701 9500 11713 9503
rect 10836 9472 11713 9500
rect 10836 9460 10842 9472
rect 11701 9469 11713 9472
rect 11747 9469 11759 9503
rect 11701 9463 11759 9469
rect 16758 9460 16764 9512
rect 16816 9500 16822 9512
rect 18340 9500 18368 9540
rect 18414 9528 18420 9540
rect 18472 9528 18478 9580
rect 18509 9571 18567 9577
rect 18509 9537 18521 9571
rect 18555 9537 18567 9571
rect 18509 9531 18567 9537
rect 18601 9571 18659 9577
rect 18601 9537 18613 9571
rect 18647 9568 18659 9571
rect 18708 9568 18828 9574
rect 18647 9546 19012 9568
rect 18647 9540 18736 9546
rect 18800 9540 19012 9546
rect 18647 9537 18659 9540
rect 18601 9531 18659 9537
rect 18524 9500 18552 9531
rect 16816 9472 18368 9500
rect 18432 9472 18552 9500
rect 18984 9500 19012 9540
rect 19058 9528 19064 9580
rect 19116 9568 19122 9580
rect 19429 9571 19487 9577
rect 19429 9568 19441 9571
rect 19116 9540 19441 9568
rect 19116 9528 19122 9540
rect 19429 9537 19441 9540
rect 19475 9537 19487 9571
rect 19613 9571 19671 9577
rect 19613 9568 19625 9571
rect 19429 9531 19487 9537
rect 19536 9540 19625 9568
rect 19150 9500 19156 9512
rect 18984 9472 19156 9500
rect 16816 9460 16822 9472
rect 12710 9392 12716 9444
rect 12768 9432 12774 9444
rect 13081 9435 13139 9441
rect 13081 9432 13093 9435
rect 12768 9404 13093 9432
rect 12768 9392 12774 9404
rect 13081 9401 13093 9404
rect 13127 9401 13139 9435
rect 13081 9395 13139 9401
rect 2866 9364 2872 9376
rect 2827 9336 2872 9364
rect 2866 9324 2872 9336
rect 2924 9324 2930 9376
rect 15286 9324 15292 9376
rect 15344 9364 15350 9376
rect 16853 9367 16911 9373
rect 16853 9364 16865 9367
rect 15344 9336 16865 9364
rect 15344 9324 15350 9336
rect 16853 9333 16865 9336
rect 16899 9333 16911 9367
rect 18432 9364 18460 9472
rect 19150 9460 19156 9472
rect 19208 9460 19214 9512
rect 19536 9500 19564 9540
rect 19613 9537 19625 9540
rect 19659 9537 19671 9571
rect 19613 9531 19671 9537
rect 19702 9528 19708 9580
rect 19760 9568 19766 9580
rect 19886 9577 19892 9580
rect 19843 9571 19892 9577
rect 19760 9540 19805 9568
rect 19760 9528 19766 9540
rect 19843 9537 19855 9571
rect 19889 9537 19892 9571
rect 19843 9531 19892 9537
rect 19886 9528 19892 9531
rect 19944 9528 19950 9580
rect 20622 9568 20628 9580
rect 20583 9540 20628 9568
rect 20622 9528 20628 9540
rect 20680 9528 20686 9580
rect 20732 9577 20760 9608
rect 20993 9605 21005 9639
rect 21039 9636 21051 9639
rect 21266 9636 21272 9648
rect 21039 9608 21272 9636
rect 21039 9605 21051 9608
rect 20993 9599 21051 9605
rect 21266 9596 21272 9608
rect 21324 9636 21330 9648
rect 22373 9639 22431 9645
rect 22373 9636 22385 9639
rect 21324 9608 22385 9636
rect 21324 9596 21330 9608
rect 22373 9605 22385 9608
rect 22419 9605 22431 9639
rect 22373 9599 22431 9605
rect 23566 9596 23572 9648
rect 23624 9636 23630 9648
rect 24762 9636 24768 9648
rect 23624 9608 24768 9636
rect 23624 9596 23630 9608
rect 24762 9596 24768 9608
rect 24820 9636 24826 9648
rect 27341 9639 27399 9645
rect 27341 9636 27353 9639
rect 24820 9608 27353 9636
rect 24820 9596 24826 9608
rect 27341 9605 27353 9608
rect 27387 9605 27399 9639
rect 30944 9636 30972 9676
rect 31386 9664 31392 9676
rect 31444 9664 31450 9716
rect 27341 9599 27399 9605
rect 27448 9608 30972 9636
rect 20718 9571 20776 9577
rect 20718 9537 20730 9571
rect 20764 9537 20776 9571
rect 20718 9531 20776 9537
rect 20901 9571 20959 9577
rect 20901 9537 20913 9571
rect 20947 9537 20959 9571
rect 20901 9531 20959 9537
rect 21131 9571 21189 9577
rect 21131 9537 21143 9571
rect 21177 9568 21189 9571
rect 21450 9568 21456 9580
rect 21177 9540 21456 9568
rect 21177 9537 21189 9540
rect 21131 9531 21189 9537
rect 20916 9500 20944 9531
rect 21450 9528 21456 9540
rect 21508 9528 21514 9580
rect 22189 9571 22247 9577
rect 22189 9537 22201 9571
rect 22235 9537 22247 9571
rect 22462 9568 22468 9580
rect 22423 9540 22468 9568
rect 22189 9531 22247 9537
rect 19444 9472 19564 9500
rect 19812 9472 20944 9500
rect 22204 9500 22232 9531
rect 22462 9528 22468 9540
rect 22520 9528 22526 9580
rect 25958 9528 25964 9580
rect 26016 9568 26022 9580
rect 27448 9577 27476 9608
rect 31018 9596 31024 9648
rect 31076 9636 31082 9648
rect 32309 9639 32367 9645
rect 32309 9636 32321 9639
rect 31076 9608 32321 9636
rect 31076 9596 31082 9608
rect 32309 9605 32321 9608
rect 32355 9605 32367 9639
rect 32309 9599 32367 9605
rect 27157 9571 27215 9577
rect 27157 9568 27169 9571
rect 26016 9540 27169 9568
rect 26016 9528 26022 9540
rect 27157 9537 27169 9540
rect 27203 9537 27215 9571
rect 27157 9531 27215 9537
rect 27433 9571 27491 9577
rect 27433 9537 27445 9571
rect 27479 9537 27491 9571
rect 27433 9531 27491 9537
rect 27525 9571 27583 9577
rect 27525 9537 27537 9571
rect 27571 9568 27583 9571
rect 27982 9568 27988 9580
rect 27571 9540 27988 9568
rect 27571 9537 27583 9540
rect 27525 9531 27583 9537
rect 27982 9528 27988 9540
rect 28040 9528 28046 9580
rect 30098 9528 30104 9580
rect 30156 9568 30162 9580
rect 31297 9571 31355 9577
rect 31297 9568 31309 9571
rect 30156 9540 31309 9568
rect 30156 9528 30162 9540
rect 31297 9537 31309 9540
rect 31343 9537 31355 9571
rect 31570 9568 31576 9580
rect 31531 9540 31576 9568
rect 31297 9531 31355 9537
rect 31570 9528 31576 9540
rect 31628 9528 31634 9580
rect 23934 9500 23940 9512
rect 22204 9472 23940 9500
rect 18782 9432 18788 9444
rect 18743 9404 18788 9432
rect 18782 9392 18788 9404
rect 18840 9392 18846 9444
rect 18874 9392 18880 9444
rect 18932 9432 18938 9444
rect 19444 9432 19472 9472
rect 19812 9432 19840 9472
rect 23934 9460 23940 9472
rect 23992 9460 23998 9512
rect 33594 9500 33600 9512
rect 31726 9472 33600 9500
rect 19978 9432 19984 9444
rect 18932 9404 19840 9432
rect 19939 9404 19984 9432
rect 18932 9392 18938 9404
rect 19978 9392 19984 9404
rect 20036 9392 20042 9444
rect 20714 9432 20720 9444
rect 20088 9404 20720 9432
rect 20088 9364 20116 9404
rect 20714 9392 20720 9404
rect 20772 9392 20778 9444
rect 21269 9435 21327 9441
rect 21269 9401 21281 9435
rect 21315 9432 21327 9435
rect 25038 9432 25044 9444
rect 21315 9404 25044 9432
rect 21315 9401 21327 9404
rect 21269 9395 21327 9401
rect 25038 9392 25044 9404
rect 25096 9392 25102 9444
rect 30190 9392 30196 9444
rect 30248 9432 30254 9444
rect 31726 9432 31754 9472
rect 33594 9460 33600 9472
rect 33652 9460 33658 9512
rect 30248 9404 31754 9432
rect 30248 9392 30254 9404
rect 18432 9336 20116 9364
rect 16853 9327 16911 9333
rect 20162 9324 20168 9376
rect 20220 9364 20226 9376
rect 22005 9367 22063 9373
rect 22005 9364 22017 9367
rect 20220 9336 22017 9364
rect 20220 9324 20226 9336
rect 22005 9333 22017 9336
rect 22051 9333 22063 9367
rect 22005 9327 22063 9333
rect 30834 9324 30840 9376
rect 30892 9364 30898 9376
rect 31570 9364 31576 9376
rect 30892 9336 31576 9364
rect 30892 9324 30898 9336
rect 31570 9324 31576 9336
rect 31628 9324 31634 9376
rect 31754 9364 31760 9376
rect 31715 9336 31760 9364
rect 31754 9324 31760 9336
rect 31812 9324 31818 9376
rect 33597 9367 33655 9373
rect 33597 9333 33609 9367
rect 33643 9364 33655 9367
rect 33686 9364 33692 9376
rect 33643 9336 33692 9364
rect 33643 9333 33655 9336
rect 33597 9327 33655 9333
rect 33686 9324 33692 9336
rect 33744 9324 33750 9376
rect 1104 9274 34868 9296
rect 1104 9222 5170 9274
rect 5222 9222 5234 9274
rect 5286 9222 5298 9274
rect 5350 9222 5362 9274
rect 5414 9222 5426 9274
rect 5478 9222 13611 9274
rect 13663 9222 13675 9274
rect 13727 9222 13739 9274
rect 13791 9222 13803 9274
rect 13855 9222 13867 9274
rect 13919 9222 22052 9274
rect 22104 9222 22116 9274
rect 22168 9222 22180 9274
rect 22232 9222 22244 9274
rect 22296 9222 22308 9274
rect 22360 9222 30493 9274
rect 30545 9222 30557 9274
rect 30609 9222 30621 9274
rect 30673 9222 30685 9274
rect 30737 9222 30749 9274
rect 30801 9222 34868 9274
rect 1104 9200 34868 9222
rect 2958 9160 2964 9172
rect 2919 9132 2964 9160
rect 2958 9120 2964 9132
rect 3016 9120 3022 9172
rect 12161 9163 12219 9169
rect 12161 9129 12173 9163
rect 12207 9160 12219 9163
rect 12526 9160 12532 9172
rect 12207 9132 12532 9160
rect 12207 9129 12219 9132
rect 12161 9123 12219 9129
rect 12526 9120 12532 9132
rect 12584 9120 12590 9172
rect 16390 9160 16396 9172
rect 16351 9132 16396 9160
rect 16390 9120 16396 9132
rect 16448 9120 16454 9172
rect 18782 9120 18788 9172
rect 18840 9160 18846 9172
rect 20254 9160 20260 9172
rect 18840 9132 20260 9160
rect 18840 9120 18846 9132
rect 20254 9120 20260 9132
rect 20312 9120 20318 9172
rect 21266 9160 21272 9172
rect 21227 9132 21272 9160
rect 21266 9120 21272 9132
rect 21324 9120 21330 9172
rect 22830 9120 22836 9172
rect 22888 9160 22894 9172
rect 26694 9160 26700 9172
rect 22888 9132 26700 9160
rect 22888 9120 22894 9132
rect 26694 9120 26700 9132
rect 26752 9120 26758 9172
rect 32306 9160 32312 9172
rect 32267 9132 32312 9160
rect 32306 9120 32312 9132
rect 32364 9120 32370 9172
rect 2777 9095 2835 9101
rect 2777 9061 2789 9095
rect 2823 9061 2835 9095
rect 2777 9055 2835 9061
rect 2792 9024 2820 9055
rect 21082 9052 21088 9104
rect 21140 9092 21146 9104
rect 21140 9064 22968 9092
rect 21140 9052 21146 9064
rect 3973 9027 4031 9033
rect 3973 9024 3985 9027
rect 2792 8996 3985 9024
rect 3973 8993 3985 8996
rect 4019 9024 4031 9027
rect 4706 9024 4712 9036
rect 4019 8996 4712 9024
rect 4019 8993 4031 8996
rect 3973 8987 4031 8993
rect 4706 8984 4712 8996
rect 4764 8984 4770 9036
rect 6822 8984 6828 9036
rect 6880 9024 6886 9036
rect 10778 9024 10784 9036
rect 6880 8996 10784 9024
rect 6880 8984 6886 8996
rect 10778 8984 10784 8996
rect 10836 8984 10842 9036
rect 4157 8959 4215 8965
rect 4157 8925 4169 8959
rect 4203 8956 4215 8959
rect 4338 8956 4344 8968
rect 4203 8928 4344 8956
rect 4203 8925 4215 8928
rect 4157 8919 4215 8925
rect 4338 8916 4344 8928
rect 4396 8916 4402 8968
rect 11054 8965 11060 8968
rect 11048 8956 11060 8965
rect 11015 8928 11060 8956
rect 11048 8919 11060 8928
rect 11054 8916 11060 8919
rect 11112 8916 11118 8968
rect 15013 8959 15071 8965
rect 15013 8925 15025 8959
rect 15059 8956 15071 8959
rect 15102 8956 15108 8968
rect 15059 8928 15108 8956
rect 15059 8925 15071 8928
rect 15013 8919 15071 8925
rect 15102 8916 15108 8928
rect 15160 8916 15166 8968
rect 15286 8965 15292 8968
rect 15280 8956 15292 8965
rect 15247 8928 15292 8956
rect 15280 8919 15292 8928
rect 15286 8916 15292 8919
rect 15344 8916 15350 8968
rect 16850 8956 16856 8968
rect 16763 8928 16856 8956
rect 16850 8916 16856 8928
rect 16908 8956 16914 8968
rect 19518 8956 19524 8968
rect 16908 8928 19524 8956
rect 16908 8916 16914 8928
rect 19518 8916 19524 8928
rect 19576 8916 19582 8968
rect 19886 8956 19892 8968
rect 19847 8928 19892 8956
rect 19886 8916 19892 8928
rect 19944 8916 19950 8968
rect 20162 8965 20168 8968
rect 20156 8956 20168 8965
rect 20123 8928 20168 8956
rect 20156 8919 20168 8928
rect 20162 8916 20168 8919
rect 20220 8916 20226 8968
rect 22646 8956 22652 8968
rect 22559 8928 22652 8956
rect 22646 8916 22652 8928
rect 22704 8916 22710 8968
rect 22830 8956 22836 8968
rect 22791 8928 22836 8956
rect 22830 8916 22836 8928
rect 22888 8916 22894 8968
rect 22940 8965 22968 9064
rect 23382 9052 23388 9104
rect 23440 9092 23446 9104
rect 26786 9092 26792 9104
rect 23440 9064 26792 9092
rect 23440 9052 23446 9064
rect 26786 9052 26792 9064
rect 26844 9052 26850 9104
rect 30190 9052 30196 9104
rect 30248 9052 30254 9104
rect 30208 9024 30236 9052
rect 24872 8996 29040 9024
rect 22925 8959 22983 8965
rect 22925 8925 22937 8959
rect 22971 8925 22983 8959
rect 22925 8919 22983 8925
rect 23658 8916 23664 8968
rect 23716 8956 23722 8968
rect 24578 8956 24584 8968
rect 23716 8928 24584 8956
rect 23716 8916 23722 8928
rect 24578 8916 24584 8928
rect 24636 8916 24642 8968
rect 24872 8965 24900 8996
rect 24857 8959 24915 8965
rect 24857 8925 24869 8959
rect 24903 8925 24915 8959
rect 24857 8919 24915 8925
rect 28721 8959 28779 8965
rect 28721 8925 28733 8959
rect 28767 8956 28779 8959
rect 28902 8956 28908 8968
rect 28767 8928 28908 8956
rect 28767 8925 28779 8928
rect 28721 8919 28779 8925
rect 2866 8848 2872 8900
rect 2924 8897 2930 8900
rect 2924 8891 2973 8897
rect 2924 8857 2927 8891
rect 2961 8857 2973 8891
rect 2924 8851 2973 8857
rect 2924 8848 2930 8851
rect 3050 8848 3056 8900
rect 3108 8888 3114 8900
rect 3329 8891 3387 8897
rect 3329 8888 3341 8891
rect 3108 8860 3341 8888
rect 3108 8848 3114 8860
rect 3329 8857 3341 8860
rect 3375 8888 3387 8891
rect 3418 8888 3424 8900
rect 3375 8860 3424 8888
rect 3375 8857 3387 8860
rect 3329 8851 3387 8857
rect 3418 8848 3424 8860
rect 3476 8848 3482 8900
rect 17120 8891 17178 8897
rect 17120 8857 17132 8891
rect 17166 8888 17178 8891
rect 17218 8888 17224 8900
rect 17166 8860 17224 8888
rect 17166 8857 17178 8860
rect 17120 8851 17178 8857
rect 17218 8848 17224 8860
rect 17276 8848 17282 8900
rect 19702 8848 19708 8900
rect 19760 8888 19766 8900
rect 22664 8888 22692 8916
rect 24872 8888 24900 8919
rect 28902 8916 28908 8928
rect 28960 8916 28966 8968
rect 29012 8965 29040 8996
rect 29932 8996 30236 9024
rect 29932 8965 29960 8996
rect 28997 8959 29055 8965
rect 28997 8925 29009 8959
rect 29043 8925 29055 8959
rect 28997 8919 29055 8925
rect 29917 8959 29975 8965
rect 29917 8925 29929 8959
rect 29963 8925 29975 8959
rect 30190 8956 30196 8968
rect 29917 8919 29975 8925
rect 30024 8928 30196 8956
rect 19760 8860 22600 8888
rect 22664 8860 24900 8888
rect 19760 8848 19766 8860
rect 4338 8820 4344 8832
rect 4299 8792 4344 8820
rect 4338 8780 4344 8792
rect 4396 8780 4402 8832
rect 18233 8823 18291 8829
rect 18233 8789 18245 8823
rect 18279 8820 18291 8823
rect 18782 8820 18788 8832
rect 18279 8792 18788 8820
rect 18279 8789 18291 8792
rect 18233 8783 18291 8789
rect 18782 8780 18788 8792
rect 18840 8780 18846 8832
rect 21910 8780 21916 8832
rect 21968 8820 21974 8832
rect 22465 8823 22523 8829
rect 22465 8820 22477 8823
rect 21968 8792 22477 8820
rect 21968 8780 21974 8792
rect 22465 8789 22477 8792
rect 22511 8789 22523 8823
rect 22572 8820 22600 8860
rect 28166 8848 28172 8900
rect 28224 8888 28230 8900
rect 28813 8891 28871 8897
rect 28813 8888 28825 8891
rect 28224 8860 28825 8888
rect 28224 8848 28230 8860
rect 28813 8857 28825 8860
rect 28859 8857 28871 8891
rect 28920 8888 28948 8916
rect 30024 8888 30052 8928
rect 30190 8916 30196 8928
rect 30248 8916 30254 8968
rect 32306 8916 32312 8968
rect 32364 8956 32370 8968
rect 33689 8959 33747 8965
rect 33689 8956 33701 8959
rect 32364 8928 33701 8956
rect 32364 8916 32370 8928
rect 33689 8925 33701 8928
rect 33735 8925 33747 8959
rect 33689 8919 33747 8925
rect 28920 8860 30052 8888
rect 30101 8891 30159 8897
rect 28813 8851 28871 8857
rect 30101 8857 30113 8891
rect 30147 8888 30159 8891
rect 30282 8888 30288 8900
rect 30147 8860 30288 8888
rect 30147 8857 30159 8860
rect 30101 8851 30159 8857
rect 30282 8848 30288 8860
rect 30340 8848 30346 8900
rect 33444 8891 33502 8897
rect 33444 8857 33456 8891
rect 33490 8888 33502 8891
rect 33870 8888 33876 8900
rect 33490 8860 33876 8888
rect 33490 8857 33502 8860
rect 33444 8851 33502 8857
rect 33870 8848 33876 8860
rect 33928 8848 33934 8900
rect 23658 8820 23664 8832
rect 22572 8792 23664 8820
rect 22465 8783 22523 8789
rect 23658 8780 23664 8792
rect 23716 8820 23722 8832
rect 24673 8823 24731 8829
rect 24673 8820 24685 8823
rect 23716 8792 24685 8820
rect 23716 8780 23722 8792
rect 24673 8789 24685 8792
rect 24719 8789 24731 8823
rect 25038 8820 25044 8832
rect 24999 8792 25044 8820
rect 24673 8783 24731 8789
rect 25038 8780 25044 8792
rect 25096 8780 25102 8832
rect 29178 8820 29184 8832
rect 29139 8792 29184 8820
rect 29178 8780 29184 8792
rect 29236 8780 29242 8832
rect 29730 8820 29736 8832
rect 29691 8792 29736 8820
rect 29730 8780 29736 8792
rect 29788 8780 29794 8832
rect 1104 8730 35027 8752
rect 1104 8678 9390 8730
rect 9442 8678 9454 8730
rect 9506 8678 9518 8730
rect 9570 8678 9582 8730
rect 9634 8678 9646 8730
rect 9698 8678 17831 8730
rect 17883 8678 17895 8730
rect 17947 8678 17959 8730
rect 18011 8678 18023 8730
rect 18075 8678 18087 8730
rect 18139 8678 26272 8730
rect 26324 8678 26336 8730
rect 26388 8678 26400 8730
rect 26452 8678 26464 8730
rect 26516 8678 26528 8730
rect 26580 8678 34713 8730
rect 34765 8678 34777 8730
rect 34829 8678 34841 8730
rect 34893 8678 34905 8730
rect 34957 8678 34969 8730
rect 35021 8678 35027 8730
rect 1104 8656 35027 8678
rect 16206 8576 16212 8628
rect 16264 8616 16270 8628
rect 16264 8588 17540 8616
rect 16264 8576 16270 8588
rect 9306 8508 9312 8560
rect 9364 8548 9370 8560
rect 9585 8551 9643 8557
rect 9585 8548 9597 8551
rect 9364 8520 9597 8548
rect 9364 8508 9370 8520
rect 9585 8517 9597 8520
rect 9631 8517 9643 8551
rect 9585 8511 9643 8517
rect 16056 8551 16114 8557
rect 16056 8517 16068 8551
rect 16102 8548 16114 8551
rect 16390 8548 16396 8560
rect 16102 8520 16396 8548
rect 16102 8517 16114 8520
rect 16056 8511 16114 8517
rect 16390 8508 16396 8520
rect 16448 8508 16454 8560
rect 16301 8483 16359 8489
rect 15304 8452 16252 8480
rect 8297 8347 8355 8353
rect 8297 8313 8309 8347
rect 8343 8344 8355 8347
rect 9858 8344 9864 8356
rect 8343 8316 9864 8344
rect 8343 8313 8355 8316
rect 8297 8307 8355 8313
rect 9858 8304 9864 8316
rect 9916 8304 9922 8356
rect 14921 8347 14979 8353
rect 14921 8313 14933 8347
rect 14967 8344 14979 8347
rect 15304 8344 15332 8452
rect 16224 8412 16252 8452
rect 16301 8449 16313 8483
rect 16347 8480 16359 8483
rect 16850 8480 16856 8492
rect 16347 8452 16856 8480
rect 16347 8449 16359 8452
rect 16301 8443 16359 8449
rect 16850 8440 16856 8452
rect 16908 8440 16914 8492
rect 17512 8489 17540 8588
rect 17678 8576 17684 8628
rect 17736 8616 17742 8628
rect 19058 8616 19064 8628
rect 17736 8588 19064 8616
rect 17736 8576 17742 8588
rect 19058 8576 19064 8588
rect 19116 8576 19122 8628
rect 19150 8576 19156 8628
rect 19208 8616 19214 8628
rect 20993 8619 21051 8625
rect 19208 8588 20944 8616
rect 19208 8576 19214 8588
rect 18874 8508 18880 8560
rect 18932 8548 18938 8560
rect 20625 8551 20683 8557
rect 20625 8548 20637 8551
rect 18932 8520 20637 8548
rect 18932 8508 18938 8520
rect 20625 8517 20637 8520
rect 20671 8517 20683 8551
rect 20625 8511 20683 8517
rect 20717 8551 20775 8557
rect 20717 8517 20729 8551
rect 20763 8517 20775 8551
rect 20717 8511 20775 8517
rect 17497 8483 17555 8489
rect 17497 8449 17509 8483
rect 17543 8449 17555 8483
rect 17497 8443 17555 8449
rect 17773 8483 17831 8489
rect 17773 8449 17785 8483
rect 17819 8449 17831 8483
rect 17773 8443 17831 8449
rect 18233 8483 18291 8489
rect 18233 8449 18245 8483
rect 18279 8480 18291 8483
rect 18690 8480 18696 8492
rect 18279 8452 18696 8480
rect 18279 8449 18291 8452
rect 18233 8443 18291 8449
rect 17586 8412 17592 8424
rect 16224 8384 17592 8412
rect 17586 8372 17592 8384
rect 17644 8372 17650 8424
rect 14967 8316 15332 8344
rect 14967 8313 14979 8316
rect 14921 8307 14979 8313
rect 16298 8304 16304 8356
rect 16356 8344 16362 8356
rect 17313 8347 17371 8353
rect 17313 8344 17325 8347
rect 16356 8316 17325 8344
rect 16356 8304 16362 8316
rect 17313 8313 17325 8316
rect 17359 8313 17371 8347
rect 17313 8307 17371 8313
rect 17126 8236 17132 8288
rect 17184 8276 17190 8288
rect 17788 8276 17816 8443
rect 18690 8440 18696 8452
rect 18748 8440 18754 8492
rect 18782 8440 18788 8492
rect 18840 8480 18846 8492
rect 20441 8483 20499 8489
rect 20441 8480 20453 8483
rect 18840 8452 20453 8480
rect 18840 8440 18846 8452
rect 20441 8449 20453 8452
rect 20487 8449 20499 8483
rect 20441 8443 20499 8449
rect 19886 8372 19892 8424
rect 19944 8412 19950 8424
rect 19981 8415 20039 8421
rect 19981 8412 19993 8415
rect 19944 8384 19993 8412
rect 19944 8372 19950 8384
rect 19981 8381 19993 8384
rect 20027 8412 20039 8415
rect 20530 8412 20536 8424
rect 20027 8384 20536 8412
rect 20027 8381 20039 8384
rect 19981 8375 20039 8381
rect 20530 8372 20536 8384
rect 20588 8372 20594 8424
rect 20732 8412 20760 8511
rect 20809 8483 20867 8489
rect 20809 8449 20821 8483
rect 20855 8480 20867 8483
rect 20916 8480 20944 8588
rect 20993 8585 21005 8619
rect 21039 8616 21051 8619
rect 23382 8616 23388 8628
rect 21039 8588 23388 8616
rect 21039 8585 21051 8588
rect 20993 8579 21051 8585
rect 23382 8576 23388 8588
rect 23440 8576 23446 8628
rect 23658 8616 23664 8628
rect 23619 8588 23664 8616
rect 23658 8576 23664 8588
rect 23716 8576 23722 8628
rect 23934 8576 23940 8628
rect 23992 8616 23998 8628
rect 23992 8588 25176 8616
rect 23992 8576 23998 8588
rect 22738 8548 22744 8560
rect 22699 8520 22744 8548
rect 22738 8508 22744 8520
rect 22796 8508 22802 8560
rect 22925 8551 22983 8557
rect 22925 8517 22937 8551
rect 22971 8548 22983 8551
rect 23566 8548 23572 8560
rect 22971 8520 23572 8548
rect 22971 8517 22983 8520
rect 22925 8511 22983 8517
rect 23566 8508 23572 8520
rect 23624 8508 23630 8560
rect 24796 8551 24854 8557
rect 24796 8517 24808 8551
rect 24842 8548 24854 8551
rect 25038 8548 25044 8560
rect 24842 8520 25044 8548
rect 24842 8517 24854 8520
rect 24796 8511 24854 8517
rect 25038 8508 25044 8520
rect 25096 8508 25102 8560
rect 25148 8548 25176 8588
rect 25222 8576 25228 8628
rect 25280 8616 25286 8628
rect 25866 8616 25872 8628
rect 25280 8588 25872 8616
rect 25280 8576 25286 8588
rect 25866 8576 25872 8588
rect 25924 8576 25930 8628
rect 28902 8576 28908 8628
rect 28960 8616 28966 8628
rect 30009 8619 30067 8625
rect 28960 8588 29224 8616
rect 28960 8576 28966 8588
rect 29086 8548 29092 8560
rect 25148 8520 25728 8548
rect 21450 8480 21456 8492
rect 20855 8452 21456 8480
rect 20855 8449 20867 8452
rect 20809 8443 20867 8449
rect 21450 8440 21456 8452
rect 21508 8440 21514 8492
rect 24946 8440 24952 8492
rect 25004 8480 25010 8492
rect 25700 8489 25728 8520
rect 28644 8520 29092 8548
rect 25501 8483 25559 8489
rect 25501 8480 25513 8483
rect 25004 8452 25513 8480
rect 25004 8440 25010 8452
rect 25501 8449 25513 8452
rect 25547 8449 25559 8483
rect 25501 8443 25559 8449
rect 25685 8483 25743 8489
rect 25685 8449 25697 8483
rect 25731 8449 25743 8483
rect 25685 8443 25743 8449
rect 25961 8483 26019 8489
rect 25961 8449 25973 8483
rect 26007 8480 26019 8483
rect 26050 8480 26056 8492
rect 26007 8452 26056 8480
rect 26007 8449 26019 8452
rect 25961 8443 26019 8449
rect 26050 8440 26056 8452
rect 26108 8440 26114 8492
rect 28644 8489 28672 8520
rect 29086 8508 29092 8520
rect 29144 8508 29150 8560
rect 29196 8548 29224 8588
rect 30009 8585 30021 8619
rect 30055 8616 30067 8619
rect 30282 8616 30288 8628
rect 30055 8588 30288 8616
rect 30055 8585 30067 8588
rect 30009 8579 30067 8585
rect 30282 8576 30288 8588
rect 30340 8576 30346 8628
rect 30837 8619 30895 8625
rect 30837 8585 30849 8619
rect 30883 8616 30895 8619
rect 30926 8616 30932 8628
rect 30883 8588 30932 8616
rect 30883 8585 30895 8588
rect 30837 8579 30895 8585
rect 30926 8576 30932 8588
rect 30984 8576 30990 8628
rect 31386 8576 31392 8628
rect 31444 8616 31450 8628
rect 33689 8619 33747 8625
rect 33689 8616 33701 8619
rect 31444 8588 33701 8616
rect 31444 8576 31450 8588
rect 33689 8585 33701 8588
rect 33735 8585 33747 8619
rect 33689 8579 33747 8585
rect 30469 8551 30527 8557
rect 30469 8548 30481 8551
rect 29196 8520 30481 8548
rect 30469 8517 30481 8520
rect 30515 8517 30527 8551
rect 30469 8511 30527 8517
rect 30576 8520 30972 8548
rect 28629 8483 28687 8489
rect 28629 8449 28641 8483
rect 28675 8449 28687 8483
rect 28629 8443 28687 8449
rect 28896 8483 28954 8489
rect 28896 8449 28908 8483
rect 28942 8480 28954 8483
rect 29730 8480 29736 8492
rect 28942 8452 29736 8480
rect 28942 8449 28954 8452
rect 28896 8443 28954 8449
rect 29730 8440 29736 8452
rect 29788 8440 29794 8492
rect 30190 8440 30196 8492
rect 30248 8480 30254 8492
rect 30576 8480 30604 8520
rect 30944 8489 30972 8520
rect 31754 8508 31760 8560
rect 31812 8548 31818 8560
rect 32554 8551 32612 8557
rect 32554 8548 32566 8551
rect 31812 8520 32566 8548
rect 31812 8508 31818 8520
rect 32554 8517 32566 8520
rect 32600 8517 32612 8551
rect 32554 8511 32612 8517
rect 30248 8452 30604 8480
rect 30653 8483 30711 8489
rect 30248 8440 30254 8452
rect 30653 8449 30665 8483
rect 30699 8449 30711 8483
rect 30653 8443 30711 8449
rect 30929 8483 30987 8489
rect 30929 8449 30941 8483
rect 30975 8449 30987 8483
rect 31846 8480 31852 8492
rect 30929 8443 30987 8449
rect 31726 8452 31852 8480
rect 20898 8412 20904 8424
rect 20732 8384 20904 8412
rect 20898 8372 20904 8384
rect 20956 8372 20962 8424
rect 25038 8412 25044 8424
rect 24999 8384 25044 8412
rect 25038 8372 25044 8384
rect 25096 8372 25102 8424
rect 30668 8412 30696 8443
rect 31726 8412 31754 8452
rect 31846 8440 31852 8452
rect 31904 8440 31910 8492
rect 32306 8480 32312 8492
rect 32267 8452 32312 8480
rect 32306 8440 32312 8452
rect 32364 8440 32370 8492
rect 30668 8384 31754 8412
rect 23109 8347 23167 8353
rect 23109 8313 23121 8347
rect 23155 8344 23167 8347
rect 24026 8344 24032 8356
rect 23155 8316 24032 8344
rect 23155 8313 23167 8316
rect 23109 8307 23167 8313
rect 24026 8304 24032 8316
rect 24084 8304 24090 8356
rect 17184 8248 17816 8276
rect 17184 8236 17190 8248
rect 19334 8236 19340 8288
rect 19392 8276 19398 8288
rect 22925 8279 22983 8285
rect 22925 8276 22937 8279
rect 19392 8248 22937 8276
rect 19392 8236 19398 8248
rect 22925 8245 22937 8248
rect 22971 8276 22983 8279
rect 29362 8276 29368 8288
rect 22971 8248 29368 8276
rect 22971 8245 22983 8248
rect 22925 8239 22983 8245
rect 29362 8236 29368 8248
rect 29420 8236 29426 8288
rect 1104 8186 34868 8208
rect 1104 8134 5170 8186
rect 5222 8134 5234 8186
rect 5286 8134 5298 8186
rect 5350 8134 5362 8186
rect 5414 8134 5426 8186
rect 5478 8134 13611 8186
rect 13663 8134 13675 8186
rect 13727 8134 13739 8186
rect 13791 8134 13803 8186
rect 13855 8134 13867 8186
rect 13919 8134 22052 8186
rect 22104 8134 22116 8186
rect 22168 8134 22180 8186
rect 22232 8134 22244 8186
rect 22296 8134 22308 8186
rect 22360 8134 30493 8186
rect 30545 8134 30557 8186
rect 30609 8134 30621 8186
rect 30673 8134 30685 8186
rect 30737 8134 30749 8186
rect 30801 8134 34868 8186
rect 1104 8112 34868 8134
rect 15654 8032 15660 8084
rect 15712 8072 15718 8084
rect 18601 8075 18659 8081
rect 18601 8072 18613 8075
rect 15712 8044 18613 8072
rect 15712 8032 15718 8044
rect 18601 8041 18613 8044
rect 18647 8041 18659 8075
rect 18601 8035 18659 8041
rect 18616 8004 18644 8035
rect 18690 8032 18696 8084
rect 18748 8072 18754 8084
rect 22925 8075 22983 8081
rect 22925 8072 22937 8075
rect 18748 8044 22937 8072
rect 18748 8032 18754 8044
rect 22925 8041 22937 8044
rect 22971 8041 22983 8075
rect 22925 8035 22983 8041
rect 28261 8075 28319 8081
rect 28261 8041 28273 8075
rect 28307 8072 28319 8075
rect 29362 8072 29368 8084
rect 28307 8044 29368 8072
rect 28307 8041 28319 8044
rect 28261 8035 28319 8041
rect 29362 8032 29368 8044
rect 29420 8032 29426 8084
rect 32306 8032 32312 8084
rect 32364 8072 32370 8084
rect 32401 8075 32459 8081
rect 32401 8072 32413 8075
rect 32364 8044 32413 8072
rect 32364 8032 32370 8044
rect 32401 8041 32413 8044
rect 32447 8041 32459 8075
rect 32401 8035 32459 8041
rect 19334 8004 19340 8016
rect 18616 7976 19340 8004
rect 19334 7964 19340 7976
rect 19392 7964 19398 8016
rect 7116 7908 9904 7936
rect 4062 7828 4068 7880
rect 4120 7868 4126 7880
rect 7116 7877 7144 7908
rect 9876 7880 9904 7908
rect 20622 7896 20628 7948
rect 20680 7936 20686 7948
rect 25130 7936 25136 7948
rect 20680 7908 25136 7936
rect 20680 7896 20686 7908
rect 25130 7896 25136 7908
rect 25188 7896 25194 7948
rect 7101 7871 7159 7877
rect 7101 7868 7113 7871
rect 4120 7840 7113 7868
rect 4120 7828 4126 7840
rect 7101 7837 7113 7840
rect 7147 7837 7159 7871
rect 7101 7831 7159 7837
rect 7285 7871 7343 7877
rect 7285 7837 7297 7871
rect 7331 7868 7343 7871
rect 9858 7868 9864 7880
rect 7331 7840 8248 7868
rect 9819 7840 9864 7868
rect 7331 7837 7343 7840
rect 7285 7831 7343 7837
rect 8220 7812 8248 7840
rect 9858 7828 9864 7840
rect 9916 7828 9922 7880
rect 10045 7871 10103 7877
rect 10045 7837 10057 7871
rect 10091 7837 10103 7871
rect 10045 7831 10103 7837
rect 18877 7871 18935 7877
rect 18877 7837 18889 7871
rect 18923 7868 18935 7871
rect 21637 7871 21695 7877
rect 21637 7868 21649 7871
rect 18923 7840 21649 7868
rect 18923 7837 18935 7840
rect 18877 7831 18935 7837
rect 21637 7837 21649 7840
rect 21683 7837 21695 7871
rect 21637 7831 21695 7837
rect 7374 7800 7380 7812
rect 7335 7772 7380 7800
rect 7374 7760 7380 7772
rect 7432 7760 7438 7812
rect 8202 7760 8208 7812
rect 8260 7800 8266 7812
rect 10060 7800 10088 7831
rect 24026 7828 24032 7880
rect 24084 7868 24090 7880
rect 24581 7871 24639 7877
rect 24581 7868 24593 7871
rect 24084 7840 24593 7868
rect 24084 7828 24090 7840
rect 24581 7837 24593 7840
rect 24627 7837 24639 7871
rect 24581 7831 24639 7837
rect 28537 7871 28595 7877
rect 28537 7837 28549 7871
rect 28583 7868 28595 7871
rect 29733 7871 29791 7877
rect 29733 7868 29745 7871
rect 28583 7840 29745 7868
rect 28583 7837 28595 7840
rect 28537 7831 28595 7837
rect 29733 7837 29745 7840
rect 29779 7837 29791 7871
rect 33686 7868 33692 7880
rect 33647 7840 33692 7868
rect 29733 7831 29791 7837
rect 33686 7828 33692 7840
rect 33744 7828 33750 7880
rect 10226 7800 10232 7812
rect 8260 7772 10088 7800
rect 10187 7772 10232 7800
rect 8260 7760 8266 7772
rect 10226 7760 10232 7772
rect 10284 7760 10290 7812
rect 15562 7760 15568 7812
rect 15620 7800 15626 7812
rect 16209 7803 16267 7809
rect 16209 7800 16221 7803
rect 15620 7772 16221 7800
rect 15620 7760 15626 7772
rect 16209 7769 16221 7772
rect 16255 7769 16267 7803
rect 16209 7763 16267 7769
rect 17310 7760 17316 7812
rect 17368 7800 17374 7812
rect 18417 7803 18475 7809
rect 18417 7800 18429 7803
rect 17368 7772 18429 7800
rect 17368 7760 17374 7772
rect 18417 7769 18429 7772
rect 18463 7800 18475 7803
rect 19429 7803 19487 7809
rect 18463 7772 19380 7800
rect 18463 7769 18475 7772
rect 18417 7763 18475 7769
rect 17494 7732 17500 7744
rect 17455 7704 17500 7732
rect 17494 7692 17500 7704
rect 17552 7692 17558 7744
rect 18601 7735 18659 7741
rect 18601 7701 18613 7735
rect 18647 7732 18659 7735
rect 19150 7732 19156 7744
rect 18647 7704 19156 7732
rect 18647 7701 18659 7704
rect 18601 7695 18659 7701
rect 19150 7692 19156 7704
rect 19208 7692 19214 7744
rect 19352 7732 19380 7772
rect 19429 7769 19441 7803
rect 19475 7800 19487 7803
rect 20806 7800 20812 7812
rect 19475 7772 20812 7800
rect 19475 7769 19487 7772
rect 19429 7763 19487 7769
rect 20806 7760 20812 7772
rect 20864 7760 20870 7812
rect 28074 7800 28080 7812
rect 28035 7772 28080 7800
rect 28074 7760 28080 7772
rect 28132 7800 28138 7812
rect 28442 7800 28448 7812
rect 28132 7772 28448 7800
rect 28132 7760 28138 7772
rect 28442 7760 28448 7772
rect 28500 7760 28506 7812
rect 20717 7735 20775 7741
rect 20717 7732 20729 7735
rect 19352 7704 20729 7732
rect 20717 7701 20729 7704
rect 20763 7701 20775 7735
rect 20717 7695 20775 7701
rect 23382 7692 23388 7744
rect 23440 7732 23446 7744
rect 25869 7735 25927 7741
rect 25869 7732 25881 7735
rect 23440 7704 25881 7732
rect 23440 7692 23446 7704
rect 25869 7701 25881 7704
rect 25915 7701 25927 7735
rect 28258 7732 28264 7744
rect 28219 7704 28264 7732
rect 25869 7695 25927 7701
rect 28258 7692 28264 7704
rect 28316 7692 28322 7744
rect 30374 7692 30380 7744
rect 30432 7732 30438 7744
rect 31021 7735 31079 7741
rect 31021 7732 31033 7735
rect 30432 7704 31033 7732
rect 30432 7692 30438 7704
rect 31021 7701 31033 7704
rect 31067 7701 31079 7735
rect 31021 7695 31079 7701
rect 1104 7642 35027 7664
rect 1104 7590 9390 7642
rect 9442 7590 9454 7642
rect 9506 7590 9518 7642
rect 9570 7590 9582 7642
rect 9634 7590 9646 7642
rect 9698 7590 17831 7642
rect 17883 7590 17895 7642
rect 17947 7590 17959 7642
rect 18011 7590 18023 7642
rect 18075 7590 18087 7642
rect 18139 7590 26272 7642
rect 26324 7590 26336 7642
rect 26388 7590 26400 7642
rect 26452 7590 26464 7642
rect 26516 7590 26528 7642
rect 26580 7590 34713 7642
rect 34765 7590 34777 7642
rect 34829 7590 34841 7642
rect 34893 7590 34905 7642
rect 34957 7590 34969 7642
rect 35021 7590 35027 7642
rect 1104 7568 35027 7590
rect 10686 7528 10692 7540
rect 10599 7500 10692 7528
rect 10686 7488 10692 7500
rect 10744 7528 10750 7540
rect 12161 7531 12219 7537
rect 12161 7528 12173 7531
rect 10744 7500 12173 7528
rect 10744 7488 10750 7500
rect 12161 7497 12173 7500
rect 12207 7497 12219 7531
rect 15562 7528 15568 7540
rect 15523 7500 15568 7528
rect 12161 7491 12219 7497
rect 15562 7488 15568 7500
rect 15620 7488 15626 7540
rect 15749 7531 15807 7537
rect 15749 7497 15761 7531
rect 15795 7528 15807 7531
rect 16758 7528 16764 7540
rect 15795 7500 16764 7528
rect 15795 7497 15807 7500
rect 15749 7491 15807 7497
rect 16758 7488 16764 7500
rect 16816 7488 16822 7540
rect 17494 7488 17500 7540
rect 17552 7488 17558 7540
rect 17681 7531 17739 7537
rect 17681 7497 17693 7531
rect 17727 7528 17739 7531
rect 18782 7528 18788 7540
rect 17727 7500 18788 7528
rect 17727 7497 17739 7500
rect 17681 7491 17739 7497
rect 18782 7488 18788 7500
rect 18840 7488 18846 7540
rect 19518 7528 19524 7540
rect 19479 7500 19524 7528
rect 19518 7488 19524 7500
rect 19576 7488 19582 7540
rect 20714 7488 20720 7540
rect 20772 7528 20778 7540
rect 20809 7531 20867 7537
rect 20809 7528 20821 7531
rect 20772 7500 20821 7528
rect 20772 7488 20778 7500
rect 20809 7497 20821 7500
rect 20855 7497 20867 7531
rect 20809 7491 20867 7497
rect 20898 7488 20904 7540
rect 20956 7528 20962 7540
rect 22373 7531 22431 7537
rect 22373 7528 22385 7531
rect 20956 7500 22385 7528
rect 20956 7488 20962 7500
rect 22373 7497 22385 7500
rect 22419 7497 22431 7531
rect 25958 7528 25964 7540
rect 25919 7500 25964 7528
rect 22373 7491 22431 7497
rect 25958 7488 25964 7500
rect 26016 7488 26022 7540
rect 29086 7528 29092 7540
rect 29047 7500 29092 7528
rect 29086 7488 29092 7500
rect 29144 7488 29150 7540
rect 5626 7420 5632 7472
rect 5684 7460 5690 7472
rect 6825 7463 6883 7469
rect 6825 7460 6837 7463
rect 5684 7432 6837 7460
rect 5684 7420 5690 7432
rect 6825 7429 6837 7432
rect 6871 7429 6883 7463
rect 6825 7423 6883 7429
rect 7374 7420 7380 7472
rect 7432 7420 7438 7472
rect 10226 7420 10232 7472
rect 10284 7420 10290 7472
rect 15933 7463 15991 7469
rect 15933 7429 15945 7463
rect 15979 7460 15991 7463
rect 17310 7460 17316 7472
rect 15979 7432 17316 7460
rect 15979 7429 15991 7432
rect 15933 7423 15991 7429
rect 17310 7420 17316 7432
rect 17368 7420 17374 7472
rect 17512 7460 17540 7488
rect 18233 7463 18291 7469
rect 18233 7460 18245 7463
rect 17420 7432 18245 7460
rect 2498 7392 2504 7404
rect 2459 7364 2504 7392
rect 2498 7352 2504 7364
rect 2556 7352 2562 7404
rect 8386 7352 8392 7404
rect 8444 7392 8450 7404
rect 8938 7392 8944 7404
rect 8444 7364 8944 7392
rect 8444 7352 8450 7364
rect 8938 7352 8944 7364
rect 8996 7352 9002 7404
rect 14737 7395 14795 7401
rect 14737 7361 14749 7395
rect 14783 7392 14795 7395
rect 17420 7392 17448 7432
rect 18233 7429 18245 7432
rect 18279 7429 18291 7463
rect 22278 7460 22284 7472
rect 18233 7423 18291 7429
rect 20916 7432 22284 7460
rect 14783 7364 17448 7392
rect 14783 7361 14795 7364
rect 14737 7355 14795 7361
rect 17494 7352 17500 7404
rect 17552 7392 17558 7404
rect 17773 7395 17831 7401
rect 17552 7364 17597 7392
rect 17552 7352 17558 7364
rect 17773 7361 17785 7395
rect 17819 7392 17831 7395
rect 17862 7392 17868 7404
rect 17819 7364 17868 7392
rect 17819 7361 17831 7364
rect 17773 7355 17831 7361
rect 17862 7352 17868 7364
rect 17920 7352 17926 7404
rect 19334 7352 19340 7404
rect 19392 7392 19398 7404
rect 20622 7392 20628 7404
rect 19392 7364 20628 7392
rect 19392 7352 19398 7364
rect 20622 7352 20628 7364
rect 20680 7352 20686 7404
rect 20916 7401 20944 7432
rect 22278 7420 22284 7432
rect 22336 7420 22342 7472
rect 23382 7460 23388 7472
rect 23343 7432 23388 7460
rect 23382 7420 23388 7432
rect 23440 7420 23446 7472
rect 25038 7460 25044 7472
rect 24999 7432 25044 7460
rect 25038 7420 25044 7432
rect 25096 7420 25102 7472
rect 20901 7395 20959 7401
rect 20901 7361 20913 7395
rect 20947 7361 20959 7395
rect 20901 7355 20959 7361
rect 22189 7395 22247 7401
rect 22189 7361 22201 7395
rect 22235 7361 22247 7395
rect 22296 7392 22324 7420
rect 22465 7395 22523 7401
rect 22465 7392 22477 7395
rect 22296 7364 22477 7392
rect 22189 7355 22247 7361
rect 22465 7361 22477 7364
rect 22511 7361 22523 7395
rect 22465 7355 22523 7361
rect 6549 7327 6607 7333
rect 6549 7293 6561 7327
rect 6595 7324 6607 7327
rect 8404 7324 8432 7352
rect 6595 7296 8432 7324
rect 9217 7327 9275 7333
rect 6595 7293 6607 7296
rect 6549 7287 6607 7293
rect 9217 7293 9229 7327
rect 9263 7324 9275 7327
rect 11054 7324 11060 7336
rect 9263 7296 11060 7324
rect 9263 7293 9275 7296
rect 9217 7287 9275 7293
rect 11054 7284 11060 7296
rect 11112 7284 11118 7336
rect 11146 7284 11152 7336
rect 11204 7324 11210 7336
rect 11882 7324 11888 7336
rect 11204 7296 11888 7324
rect 11204 7284 11210 7296
rect 11882 7284 11888 7296
rect 11940 7284 11946 7336
rect 12069 7327 12127 7333
rect 12069 7293 12081 7327
rect 12115 7324 12127 7327
rect 13078 7324 13084 7336
rect 12115 7296 13084 7324
rect 12115 7293 12127 7296
rect 12069 7287 12127 7293
rect 13078 7284 13084 7296
rect 13136 7284 13142 7336
rect 17218 7284 17224 7336
rect 17276 7324 17282 7336
rect 17313 7327 17371 7333
rect 17313 7324 17325 7327
rect 17276 7296 17325 7324
rect 17276 7284 17282 7296
rect 17313 7293 17325 7296
rect 17359 7293 17371 7327
rect 17512 7324 17540 7352
rect 22204 7324 22232 7355
rect 25130 7352 25136 7404
rect 25188 7392 25194 7404
rect 25777 7395 25835 7401
rect 25777 7392 25789 7395
rect 25188 7364 25789 7392
rect 25188 7352 25194 7364
rect 25777 7361 25789 7364
rect 25823 7361 25835 7395
rect 26050 7392 26056 7404
rect 25963 7364 26056 7392
rect 25777 7355 25835 7361
rect 26050 7352 26056 7364
rect 26108 7352 26114 7404
rect 30374 7392 30380 7404
rect 30335 7364 30380 7392
rect 30374 7352 30380 7364
rect 30432 7352 30438 7404
rect 23750 7324 23756 7336
rect 17512 7296 23756 7324
rect 17313 7287 17371 7293
rect 23750 7284 23756 7296
rect 23808 7284 23814 7336
rect 24026 7284 24032 7336
rect 24084 7324 24090 7336
rect 24578 7324 24584 7336
rect 24084 7296 24584 7324
rect 24084 7284 24090 7296
rect 24578 7284 24584 7296
rect 24636 7324 24642 7336
rect 26068 7324 26096 7352
rect 24636 7296 26096 7324
rect 24636 7284 24642 7296
rect 2590 7188 2596 7200
rect 2551 7160 2596 7188
rect 2590 7148 2596 7160
rect 2648 7148 2654 7200
rect 8294 7188 8300 7200
rect 8255 7160 8300 7188
rect 8294 7148 8300 7160
rect 8352 7148 8358 7200
rect 12526 7188 12532 7200
rect 12487 7160 12532 7188
rect 12526 7148 12532 7160
rect 12584 7148 12590 7200
rect 13449 7191 13507 7197
rect 13449 7157 13461 7191
rect 13495 7188 13507 7191
rect 15102 7188 15108 7200
rect 13495 7160 15108 7188
rect 13495 7157 13507 7160
rect 13449 7151 13507 7157
rect 15102 7148 15108 7160
rect 15160 7148 15166 7200
rect 15654 7148 15660 7200
rect 15712 7188 15718 7200
rect 15749 7191 15807 7197
rect 15749 7188 15761 7191
rect 15712 7160 15761 7188
rect 15712 7148 15718 7160
rect 15749 7157 15761 7160
rect 15795 7157 15807 7191
rect 20438 7188 20444 7200
rect 20399 7160 20444 7188
rect 15749 7151 15807 7157
rect 20438 7148 20444 7160
rect 20496 7148 20502 7200
rect 20714 7148 20720 7200
rect 20772 7188 20778 7200
rect 22005 7191 22063 7197
rect 22005 7188 22017 7191
rect 20772 7160 22017 7188
rect 20772 7148 20778 7160
rect 22005 7157 22017 7160
rect 22051 7157 22063 7191
rect 25590 7188 25596 7200
rect 25551 7160 25596 7188
rect 22005 7151 22063 7157
rect 25590 7148 25596 7160
rect 25648 7148 25654 7200
rect 1104 7098 34868 7120
rect 1104 7046 5170 7098
rect 5222 7046 5234 7098
rect 5286 7046 5298 7098
rect 5350 7046 5362 7098
rect 5414 7046 5426 7098
rect 5478 7046 13611 7098
rect 13663 7046 13675 7098
rect 13727 7046 13739 7098
rect 13791 7046 13803 7098
rect 13855 7046 13867 7098
rect 13919 7046 22052 7098
rect 22104 7046 22116 7098
rect 22168 7046 22180 7098
rect 22232 7046 22244 7098
rect 22296 7046 22308 7098
rect 22360 7046 30493 7098
rect 30545 7046 30557 7098
rect 30609 7046 30621 7098
rect 30673 7046 30685 7098
rect 30737 7046 30749 7098
rect 30801 7046 34868 7098
rect 1104 7024 34868 7046
rect 1673 6987 1731 6993
rect 1673 6953 1685 6987
rect 1719 6984 1731 6987
rect 2498 6984 2504 6996
rect 1719 6956 2504 6984
rect 1719 6953 1731 6956
rect 1673 6947 1731 6953
rect 2498 6944 2504 6956
rect 2556 6944 2562 6996
rect 2590 6944 2596 6996
rect 2648 6984 2654 6996
rect 3157 6987 3215 6993
rect 3157 6984 3169 6987
rect 2648 6956 3169 6984
rect 2648 6944 2654 6956
rect 3157 6953 3169 6956
rect 3203 6953 3215 6987
rect 13078 6984 13084 6996
rect 13039 6956 13084 6984
rect 3157 6947 3215 6953
rect 13078 6944 13084 6956
rect 13136 6944 13142 6996
rect 20806 6984 20812 6996
rect 20767 6956 20812 6984
rect 20806 6944 20812 6956
rect 20864 6944 20870 6996
rect 7852 6888 8340 6916
rect 4338 6808 4344 6860
rect 4396 6848 4402 6860
rect 5074 6848 5080 6860
rect 4396 6820 5080 6848
rect 4396 6808 4402 6820
rect 5074 6808 5080 6820
rect 5132 6848 5138 6860
rect 5445 6851 5503 6857
rect 5445 6848 5457 6851
rect 5132 6820 5457 6848
rect 5132 6808 5138 6820
rect 5445 6817 5457 6820
rect 5491 6817 5503 6851
rect 5445 6811 5503 6817
rect 3418 6740 3424 6792
rect 3476 6780 3482 6792
rect 4062 6780 4068 6792
rect 3476 6752 4068 6780
rect 3476 6740 3482 6752
rect 4062 6740 4068 6752
rect 4120 6740 4126 6792
rect 5718 6789 5724 6792
rect 5712 6780 5724 6789
rect 5679 6752 5724 6780
rect 5712 6743 5724 6752
rect 5718 6740 5724 6743
rect 5776 6740 5782 6792
rect 7653 6783 7711 6789
rect 7653 6749 7665 6783
rect 7699 6780 7711 6783
rect 7852 6780 7880 6888
rect 8312 6860 8340 6888
rect 17218 6876 17224 6928
rect 17276 6916 17282 6928
rect 17862 6916 17868 6928
rect 17276 6888 17868 6916
rect 17276 6876 17282 6888
rect 17862 6876 17868 6888
rect 17920 6876 17926 6928
rect 7929 6851 7987 6857
rect 7929 6817 7941 6851
rect 7975 6848 7987 6851
rect 7975 6820 8248 6848
rect 7975 6817 7987 6820
rect 7929 6811 7987 6817
rect 7699 6752 7880 6780
rect 7699 6749 7711 6752
rect 7653 6743 7711 6749
rect 2682 6672 2688 6724
rect 2740 6672 2746 6724
rect 7745 6715 7803 6721
rect 7745 6712 7757 6715
rect 6840 6684 7757 6712
rect 6840 6653 6868 6684
rect 7745 6681 7757 6684
rect 7791 6681 7803 6715
rect 7745 6675 7803 6681
rect 6825 6647 6883 6653
rect 6825 6613 6837 6647
rect 6871 6613 6883 6647
rect 6825 6607 6883 6613
rect 6914 6604 6920 6656
rect 6972 6644 6978 6656
rect 7285 6647 7343 6653
rect 7285 6644 7297 6647
rect 6972 6616 7297 6644
rect 6972 6604 6978 6616
rect 7285 6613 7297 6616
rect 7331 6613 7343 6647
rect 8220 6644 8248 6820
rect 8294 6808 8300 6860
rect 8352 6848 8358 6860
rect 10137 6851 10195 6857
rect 10137 6848 10149 6851
rect 8352 6820 10149 6848
rect 8352 6808 8358 6820
rect 10137 6817 10149 6820
rect 10183 6817 10195 6851
rect 10137 6811 10195 6817
rect 10318 6808 10324 6860
rect 10376 6848 10382 6860
rect 10689 6851 10747 6857
rect 10689 6848 10701 6851
rect 10376 6820 10701 6848
rect 10376 6808 10382 6820
rect 10689 6817 10701 6820
rect 10735 6817 10747 6851
rect 10689 6811 10747 6817
rect 15102 6808 15108 6860
rect 15160 6848 15166 6860
rect 15565 6851 15623 6857
rect 15565 6848 15577 6851
rect 15160 6820 15577 6848
rect 15160 6808 15166 6820
rect 15565 6817 15577 6820
rect 15611 6817 15623 6851
rect 19334 6848 19340 6860
rect 15565 6811 15623 6817
rect 17604 6820 19340 6848
rect 10229 6783 10287 6789
rect 10229 6749 10241 6783
rect 10275 6749 10287 6783
rect 10229 6743 10287 6749
rect 10244 6712 10272 6743
rect 10410 6740 10416 6792
rect 10468 6780 10474 6792
rect 10551 6783 10609 6789
rect 10551 6780 10563 6783
rect 10468 6752 10563 6780
rect 10468 6740 10474 6752
rect 10551 6749 10563 6752
rect 10597 6749 10609 6783
rect 11146 6780 11152 6792
rect 10551 6743 10609 6749
rect 10796 6752 11152 6780
rect 10686 6712 10692 6724
rect 10244 6684 10692 6712
rect 10686 6672 10692 6684
rect 10744 6672 10750 6724
rect 10796 6644 10824 6752
rect 11146 6740 11152 6752
rect 11204 6740 11210 6792
rect 11698 6780 11704 6792
rect 11659 6752 11704 6780
rect 11698 6740 11704 6752
rect 11756 6740 11762 6792
rect 13541 6783 13599 6789
rect 13541 6749 13553 6783
rect 13587 6749 13599 6783
rect 13541 6743 13599 6749
rect 13725 6783 13783 6789
rect 13725 6749 13737 6783
rect 13771 6780 13783 6783
rect 15654 6780 15660 6792
rect 13771 6752 15660 6780
rect 13771 6749 13783 6752
rect 13725 6743 13783 6749
rect 11054 6672 11060 6724
rect 11112 6712 11118 6724
rect 11946 6715 12004 6721
rect 11946 6712 11958 6715
rect 11112 6684 11958 6712
rect 11112 6672 11118 6684
rect 11946 6681 11958 6684
rect 11992 6681 12004 6715
rect 12802 6712 12808 6724
rect 11946 6675 12004 6681
rect 12406 6684 12808 6712
rect 8220 6616 10824 6644
rect 10965 6647 11023 6653
rect 7285 6607 7343 6613
rect 10965 6613 10977 6647
rect 11011 6644 11023 6647
rect 12406 6644 12434 6684
rect 12802 6672 12808 6684
rect 12860 6672 12866 6724
rect 13556 6712 13584 6743
rect 15654 6740 15660 6752
rect 15712 6740 15718 6792
rect 15832 6783 15890 6789
rect 15832 6749 15844 6783
rect 15878 6780 15890 6783
rect 16298 6780 16304 6792
rect 15878 6752 16304 6780
rect 15878 6749 15890 6752
rect 15832 6743 15890 6749
rect 16298 6740 16304 6752
rect 16356 6740 16362 6792
rect 16390 6740 16396 6792
rect 16448 6780 16454 6792
rect 17604 6789 17632 6820
rect 19334 6808 19340 6820
rect 19392 6808 19398 6860
rect 20530 6808 20536 6860
rect 20588 6848 20594 6860
rect 21269 6851 21327 6857
rect 21269 6848 21281 6851
rect 20588 6820 21281 6848
rect 20588 6808 20594 6820
rect 21269 6817 21281 6820
rect 21315 6817 21327 6851
rect 21269 6811 21327 6817
rect 17405 6783 17463 6789
rect 17405 6780 17417 6783
rect 16448 6752 17417 6780
rect 16448 6740 16454 6752
rect 17405 6749 17417 6752
rect 17451 6749 17463 6783
rect 17405 6743 17463 6749
rect 17589 6783 17647 6789
rect 17589 6749 17601 6783
rect 17635 6749 17647 6783
rect 17862 6780 17868 6792
rect 17823 6752 17868 6780
rect 17589 6743 17647 6749
rect 17862 6740 17868 6752
rect 17920 6740 17926 6792
rect 19429 6783 19487 6789
rect 19429 6749 19441 6783
rect 19475 6780 19487 6783
rect 19518 6780 19524 6792
rect 19475 6752 19524 6780
rect 19475 6749 19487 6752
rect 19429 6743 19487 6749
rect 19518 6740 19524 6752
rect 19576 6740 19582 6792
rect 19696 6783 19754 6789
rect 19696 6749 19708 6783
rect 19742 6780 19754 6783
rect 20438 6780 20444 6792
rect 19742 6752 20444 6780
rect 19742 6749 19754 6752
rect 19696 6743 19754 6749
rect 20438 6740 20444 6752
rect 20496 6740 20502 6792
rect 21536 6783 21594 6789
rect 21536 6749 21548 6783
rect 21582 6780 21594 6783
rect 21910 6780 21916 6792
rect 21582 6752 21916 6780
rect 21582 6749 21594 6752
rect 21536 6743 21594 6749
rect 21910 6740 21916 6752
rect 21968 6740 21974 6792
rect 23750 6780 23756 6792
rect 23711 6752 23756 6780
rect 23750 6740 23756 6752
rect 23808 6740 23814 6792
rect 24026 6780 24032 6792
rect 23987 6752 24032 6780
rect 24026 6740 24032 6752
rect 24084 6740 24090 6792
rect 24581 6783 24639 6789
rect 24581 6749 24593 6783
rect 24627 6780 24639 6783
rect 24627 6752 25084 6780
rect 24627 6749 24639 6752
rect 24581 6743 24639 6749
rect 25056 6724 25084 6752
rect 28902 6740 28908 6792
rect 28960 6789 28966 6792
rect 28960 6780 28972 6789
rect 28960 6752 29005 6780
rect 28960 6743 28972 6752
rect 28960 6740 28966 6743
rect 29086 6740 29092 6792
rect 29144 6780 29150 6792
rect 29181 6783 29239 6789
rect 29181 6780 29193 6783
rect 29144 6752 29193 6780
rect 29144 6740 29150 6752
rect 29181 6749 29193 6752
rect 29227 6749 29239 6783
rect 29181 6743 29239 6749
rect 29822 6740 29828 6792
rect 29880 6780 29886 6792
rect 30101 6783 30159 6789
rect 30101 6780 30113 6783
rect 29880 6752 30113 6780
rect 29880 6740 29886 6752
rect 30101 6749 30113 6752
rect 30147 6749 30159 6783
rect 30101 6743 30159 6749
rect 17218 6712 17224 6724
rect 13556 6684 17224 6712
rect 17218 6672 17224 6684
rect 17276 6672 17282 6724
rect 17494 6672 17500 6724
rect 17552 6712 17558 6724
rect 17773 6715 17831 6721
rect 17773 6712 17785 6715
rect 17552 6684 17785 6712
rect 17552 6672 17558 6684
rect 17773 6681 17785 6684
rect 17819 6681 17831 6715
rect 17773 6675 17831 6681
rect 23474 6672 23480 6724
rect 23532 6712 23538 6724
rect 23937 6715 23995 6721
rect 23937 6712 23949 6715
rect 23532 6684 23949 6712
rect 23532 6672 23538 6684
rect 23937 6681 23949 6684
rect 23983 6681 23995 6715
rect 23937 6675 23995 6681
rect 24848 6715 24906 6721
rect 24848 6681 24860 6715
rect 24894 6712 24906 6715
rect 24946 6712 24952 6724
rect 24894 6684 24952 6712
rect 24894 6681 24906 6684
rect 24848 6675 24906 6681
rect 24946 6672 24952 6684
rect 25004 6672 25010 6724
rect 25038 6672 25044 6724
rect 25096 6672 25102 6724
rect 29270 6672 29276 6724
rect 29328 6712 29334 6724
rect 30346 6715 30404 6721
rect 30346 6712 30358 6715
rect 29328 6684 30358 6712
rect 29328 6672 29334 6684
rect 30346 6681 30358 6684
rect 30392 6681 30404 6715
rect 30346 6675 30404 6681
rect 13630 6644 13636 6656
rect 11011 6616 12434 6644
rect 13591 6616 13636 6644
rect 11011 6613 11023 6616
rect 10965 6607 11023 6613
rect 13630 6604 13636 6616
rect 13688 6604 13694 6656
rect 16945 6647 17003 6653
rect 16945 6613 16957 6647
rect 16991 6644 17003 6647
rect 17678 6644 17684 6656
rect 16991 6616 17684 6644
rect 16991 6613 17003 6616
rect 16945 6607 17003 6613
rect 17678 6604 17684 6616
rect 17736 6604 17742 6656
rect 22649 6647 22707 6653
rect 22649 6613 22661 6647
rect 22695 6644 22707 6647
rect 22830 6644 22836 6656
rect 22695 6616 22836 6644
rect 22695 6613 22707 6616
rect 22649 6607 22707 6613
rect 22830 6604 22836 6616
rect 22888 6604 22894 6656
rect 23566 6644 23572 6656
rect 23527 6616 23572 6644
rect 23566 6604 23572 6616
rect 23624 6604 23630 6656
rect 25866 6604 25872 6656
rect 25924 6644 25930 6656
rect 25961 6647 26019 6653
rect 25961 6644 25973 6647
rect 25924 6616 25973 6644
rect 25924 6604 25930 6616
rect 25961 6613 25973 6616
rect 26007 6613 26019 6647
rect 27798 6644 27804 6656
rect 27759 6616 27804 6644
rect 25961 6607 26019 6613
rect 27798 6604 27804 6616
rect 27856 6604 27862 6656
rect 28534 6604 28540 6656
rect 28592 6644 28598 6656
rect 31481 6647 31539 6653
rect 31481 6644 31493 6647
rect 28592 6616 31493 6644
rect 28592 6604 28598 6616
rect 31481 6613 31493 6616
rect 31527 6613 31539 6647
rect 31481 6607 31539 6613
rect 1104 6554 35027 6576
rect 1104 6502 9390 6554
rect 9442 6502 9454 6554
rect 9506 6502 9518 6554
rect 9570 6502 9582 6554
rect 9634 6502 9646 6554
rect 9698 6502 17831 6554
rect 17883 6502 17895 6554
rect 17947 6502 17959 6554
rect 18011 6502 18023 6554
rect 18075 6502 18087 6554
rect 18139 6502 26272 6554
rect 26324 6502 26336 6554
rect 26388 6502 26400 6554
rect 26452 6502 26464 6554
rect 26516 6502 26528 6554
rect 26580 6502 34713 6554
rect 34765 6502 34777 6554
rect 34829 6502 34841 6554
rect 34893 6502 34905 6554
rect 34957 6502 34969 6554
rect 35021 6502 35027 6554
rect 1104 6480 35027 6502
rect 2498 6400 2504 6452
rect 2556 6440 2562 6452
rect 6914 6440 6920 6452
rect 2556 6412 3740 6440
rect 6875 6412 6920 6440
rect 2556 6400 2562 6412
rect 2682 6332 2688 6384
rect 2740 6372 2746 6384
rect 3712 6381 3740 6412
rect 6914 6400 6920 6412
rect 6972 6400 6978 6452
rect 12526 6400 12532 6452
rect 12584 6440 12590 6452
rect 12989 6443 13047 6449
rect 12989 6440 13001 6443
rect 12584 6412 13001 6440
rect 12584 6400 12590 6412
rect 12989 6409 13001 6412
rect 13035 6409 13047 6443
rect 20898 6440 20904 6452
rect 20859 6412 20904 6440
rect 12989 6403 13047 6409
rect 20898 6400 20904 6412
rect 20956 6400 20962 6452
rect 27798 6400 27804 6452
rect 27856 6440 27862 6452
rect 30926 6440 30932 6452
rect 27856 6412 30932 6440
rect 27856 6400 27862 6412
rect 30926 6400 30932 6412
rect 30984 6400 30990 6452
rect 2777 6375 2835 6381
rect 2777 6372 2789 6375
rect 2740 6344 2789 6372
rect 2740 6332 2746 6344
rect 2777 6341 2789 6344
rect 2823 6341 2835 6375
rect 2777 6335 2835 6341
rect 3697 6375 3755 6381
rect 3697 6341 3709 6375
rect 3743 6341 3755 6375
rect 3697 6335 3755 6341
rect 6825 6375 6883 6381
rect 6825 6341 6837 6375
rect 6871 6372 6883 6375
rect 7006 6372 7012 6384
rect 6871 6344 7012 6372
rect 6871 6341 6883 6344
rect 6825 6335 6883 6341
rect 7006 6332 7012 6344
rect 7064 6332 7070 6384
rect 12897 6375 12955 6381
rect 12897 6341 12909 6375
rect 12943 6372 12955 6375
rect 13630 6372 13636 6384
rect 12943 6344 13636 6372
rect 12943 6341 12955 6344
rect 12897 6335 12955 6341
rect 13630 6332 13636 6344
rect 13688 6332 13694 6384
rect 19788 6375 19846 6381
rect 19788 6341 19800 6375
rect 19834 6372 19846 6375
rect 20714 6372 20720 6384
rect 19834 6344 20720 6372
rect 19834 6341 19846 6344
rect 19788 6335 19846 6341
rect 20714 6332 20720 6344
rect 20772 6332 20778 6384
rect 23566 6332 23572 6384
rect 23624 6372 23630 6384
rect 24682 6375 24740 6381
rect 24682 6372 24694 6375
rect 23624 6344 24694 6372
rect 23624 6332 23630 6344
rect 24682 6341 24694 6344
rect 24728 6341 24740 6375
rect 24682 6335 24740 6341
rect 29178 6332 29184 6384
rect 29236 6372 29242 6384
rect 29558 6375 29616 6381
rect 29558 6372 29570 6375
rect 29236 6344 29570 6372
rect 29236 6332 29242 6344
rect 29558 6341 29570 6344
rect 29604 6341 29616 6375
rect 29558 6335 29616 6341
rect 2958 6304 2964 6316
rect 2919 6276 2964 6304
rect 2958 6264 2964 6276
rect 3016 6264 3022 6316
rect 3145 6307 3203 6313
rect 3145 6273 3157 6307
rect 3191 6304 3203 6307
rect 3418 6304 3424 6316
rect 3191 6276 3424 6304
rect 3191 6273 3203 6276
rect 3145 6267 3203 6273
rect 3418 6264 3424 6276
rect 3476 6264 3482 6316
rect 5718 6196 5724 6248
rect 5776 6236 5782 6248
rect 6641 6239 6699 6245
rect 6641 6236 6653 6239
rect 5776 6208 6653 6236
rect 5776 6196 5782 6208
rect 6641 6205 6653 6208
rect 6687 6236 6699 6239
rect 12342 6236 12348 6248
rect 6687 6208 12348 6236
rect 6687 6205 6699 6208
rect 6641 6199 6699 6205
rect 12342 6196 12348 6208
rect 12400 6236 12406 6248
rect 12713 6239 12771 6245
rect 12713 6236 12725 6239
rect 12400 6208 12725 6236
rect 12400 6196 12406 6208
rect 12713 6205 12725 6208
rect 12759 6205 12771 6239
rect 19518 6236 19524 6248
rect 19479 6208 19524 6236
rect 12713 6199 12771 6205
rect 19518 6196 19524 6208
rect 19576 6196 19582 6248
rect 24949 6239 25007 6245
rect 24949 6205 24961 6239
rect 24995 6205 25007 6239
rect 29822 6236 29828 6248
rect 29783 6208 29828 6236
rect 24949 6199 25007 6205
rect 7285 6171 7343 6177
rect 7285 6137 7297 6171
rect 7331 6168 7343 6171
rect 18414 6168 18420 6180
rect 7331 6140 18420 6168
rect 7331 6137 7343 6140
rect 7285 6131 7343 6137
rect 18414 6128 18420 6140
rect 18472 6128 18478 6180
rect 23474 6128 23480 6180
rect 23532 6168 23538 6180
rect 23569 6171 23627 6177
rect 23569 6168 23581 6171
rect 23532 6140 23581 6168
rect 23532 6128 23538 6140
rect 23569 6137 23581 6140
rect 23615 6137 23627 6171
rect 23569 6131 23627 6137
rect 3789 6103 3847 6109
rect 3789 6069 3801 6103
rect 3835 6100 3847 6103
rect 3970 6100 3976 6112
rect 3835 6072 3976 6100
rect 3835 6069 3847 6072
rect 3789 6063 3847 6069
rect 3970 6060 3976 6072
rect 4028 6060 4034 6112
rect 13357 6103 13415 6109
rect 13357 6069 13369 6103
rect 13403 6100 13415 6103
rect 20162 6100 20168 6112
rect 13403 6072 20168 6100
rect 13403 6069 13415 6072
rect 13357 6063 13415 6069
rect 20162 6060 20168 6072
rect 20220 6060 20226 6112
rect 24670 6060 24676 6112
rect 24728 6100 24734 6112
rect 24964 6100 24992 6199
rect 29822 6196 29828 6208
rect 29880 6196 29886 6248
rect 28166 6128 28172 6180
rect 28224 6168 28230 6180
rect 28445 6171 28503 6177
rect 28445 6168 28457 6171
rect 28224 6140 28457 6168
rect 28224 6128 28230 6140
rect 28445 6137 28457 6140
rect 28491 6137 28503 6171
rect 28445 6131 28503 6137
rect 24728 6072 24992 6100
rect 24728 6060 24734 6072
rect 1104 6010 34868 6032
rect 1104 5958 5170 6010
rect 5222 5958 5234 6010
rect 5286 5958 5298 6010
rect 5350 5958 5362 6010
rect 5414 5958 5426 6010
rect 5478 5958 13611 6010
rect 13663 5958 13675 6010
rect 13727 5958 13739 6010
rect 13791 5958 13803 6010
rect 13855 5958 13867 6010
rect 13919 5958 22052 6010
rect 22104 5958 22116 6010
rect 22168 5958 22180 6010
rect 22232 5958 22244 6010
rect 22296 5958 22308 6010
rect 22360 5958 30493 6010
rect 30545 5958 30557 6010
rect 30609 5958 30621 6010
rect 30673 5958 30685 6010
rect 30737 5958 30749 6010
rect 30801 5958 34868 6010
rect 1104 5936 34868 5958
rect 25958 5896 25964 5908
rect 25919 5868 25964 5896
rect 25958 5856 25964 5868
rect 26016 5856 26022 5908
rect 29181 5899 29239 5905
rect 29181 5865 29193 5899
rect 29227 5896 29239 5899
rect 29270 5896 29276 5908
rect 29227 5868 29276 5896
rect 29227 5865 29239 5868
rect 29181 5859 29239 5865
rect 29270 5856 29276 5868
rect 29328 5856 29334 5908
rect 28994 5828 29000 5840
rect 28736 5800 29000 5828
rect 3970 5760 3976 5772
rect 3931 5732 3976 5760
rect 3970 5720 3976 5732
rect 4028 5720 4034 5772
rect 4341 5763 4399 5769
rect 4341 5729 4353 5763
rect 4387 5760 4399 5763
rect 5534 5760 5540 5772
rect 4387 5732 5540 5760
rect 4387 5729 4399 5732
rect 4341 5723 4399 5729
rect 5534 5720 5540 5732
rect 5592 5720 5598 5772
rect 5718 5760 5724 5772
rect 5679 5732 5724 5760
rect 5718 5720 5724 5732
rect 5776 5720 5782 5772
rect 11882 5720 11888 5772
rect 11940 5760 11946 5772
rect 12897 5763 12955 5769
rect 12897 5760 12909 5763
rect 11940 5732 12909 5760
rect 11940 5720 11946 5732
rect 12897 5729 12909 5732
rect 12943 5729 12955 5763
rect 12897 5723 12955 5729
rect 12342 5652 12348 5704
rect 12400 5692 12406 5704
rect 12621 5695 12679 5701
rect 12621 5692 12633 5695
rect 12400 5664 12633 5692
rect 12400 5652 12406 5664
rect 12621 5661 12633 5664
rect 12667 5661 12679 5695
rect 12621 5655 12679 5661
rect 12710 5652 12716 5704
rect 12768 5692 12774 5704
rect 24581 5695 24639 5701
rect 12768 5664 12813 5692
rect 12768 5652 12774 5664
rect 24581 5661 24593 5695
rect 24627 5692 24639 5695
rect 24670 5692 24676 5704
rect 24627 5664 24676 5692
rect 24627 5661 24639 5664
rect 24581 5655 24639 5661
rect 24670 5652 24676 5664
rect 24728 5652 24734 5704
rect 24848 5695 24906 5701
rect 24848 5661 24860 5695
rect 24894 5692 24906 5695
rect 25590 5692 25596 5704
rect 24894 5664 25596 5692
rect 24894 5661 24906 5664
rect 24848 5655 24906 5661
rect 25590 5652 25596 5664
rect 25648 5652 25654 5704
rect 28736 5701 28764 5800
rect 28994 5788 29000 5800
rect 29052 5788 29058 5840
rect 28721 5695 28779 5701
rect 28721 5661 28733 5695
rect 28767 5661 28779 5695
rect 28721 5655 28779 5661
rect 28997 5695 29055 5701
rect 28997 5661 29009 5695
rect 29043 5692 29055 5695
rect 30834 5692 30840 5704
rect 29043 5664 30840 5692
rect 29043 5661 29055 5664
rect 28997 5655 29055 5661
rect 30834 5652 30840 5664
rect 30892 5652 30898 5704
rect 4706 5584 4712 5636
rect 4764 5584 4770 5636
rect 28534 5584 28540 5636
rect 28592 5624 28598 5636
rect 28813 5627 28871 5633
rect 28813 5624 28825 5627
rect 28592 5596 28825 5624
rect 28592 5584 28598 5596
rect 28813 5593 28825 5596
rect 28859 5593 28871 5627
rect 28813 5587 28871 5593
rect 12897 5559 12955 5565
rect 12897 5525 12909 5559
rect 12943 5556 12955 5559
rect 14274 5556 14280 5568
rect 12943 5528 14280 5556
rect 12943 5525 12955 5528
rect 12897 5519 12955 5525
rect 14274 5516 14280 5528
rect 14332 5516 14338 5568
rect 1104 5466 35027 5488
rect 1104 5414 9390 5466
rect 9442 5414 9454 5466
rect 9506 5414 9518 5466
rect 9570 5414 9582 5466
rect 9634 5414 9646 5466
rect 9698 5414 17831 5466
rect 17883 5414 17895 5466
rect 17947 5414 17959 5466
rect 18011 5414 18023 5466
rect 18075 5414 18087 5466
rect 18139 5414 26272 5466
rect 26324 5414 26336 5466
rect 26388 5414 26400 5466
rect 26452 5414 26464 5466
rect 26516 5414 26528 5466
rect 26580 5414 34713 5466
rect 34765 5414 34777 5466
rect 34829 5414 34841 5466
rect 34893 5414 34905 5466
rect 34957 5414 34969 5466
rect 35021 5414 35027 5466
rect 1104 5392 35027 5414
rect 5534 5312 5540 5364
rect 5592 5352 5598 5364
rect 5629 5355 5687 5361
rect 5629 5352 5641 5355
rect 5592 5324 5641 5352
rect 5592 5312 5598 5324
rect 5629 5321 5641 5324
rect 5675 5321 5687 5355
rect 5629 5315 5687 5321
rect 9493 5355 9551 5361
rect 9493 5321 9505 5355
rect 9539 5352 9551 5355
rect 10226 5352 10232 5364
rect 9539 5324 10232 5352
rect 9539 5321 9551 5324
rect 9493 5315 9551 5321
rect 4341 5287 4399 5293
rect 4341 5253 4353 5287
rect 4387 5284 4399 5287
rect 4706 5284 4712 5296
rect 4387 5256 4712 5284
rect 4387 5253 4399 5256
rect 4341 5247 4399 5253
rect 4706 5244 4712 5256
rect 4764 5244 4770 5296
rect 5644 5284 5672 5315
rect 10226 5312 10232 5324
rect 10284 5312 10290 5364
rect 10410 5352 10416 5364
rect 10371 5324 10416 5352
rect 10410 5312 10416 5324
rect 10468 5312 10474 5364
rect 12710 5312 12716 5364
rect 12768 5352 12774 5364
rect 13081 5355 13139 5361
rect 13081 5352 13093 5355
rect 12768 5324 13093 5352
rect 12768 5312 12774 5324
rect 13081 5321 13093 5324
rect 13127 5321 13139 5355
rect 19518 5352 19524 5364
rect 19479 5324 19524 5352
rect 13081 5315 13139 5321
rect 19518 5312 19524 5324
rect 19576 5312 19582 5364
rect 24670 5352 24676 5364
rect 24631 5324 24676 5352
rect 24670 5312 24676 5324
rect 24728 5312 24734 5364
rect 6638 5284 6644 5296
rect 5644 5256 6644 5284
rect 6638 5244 6644 5256
rect 6696 5284 6702 5296
rect 6696 5256 8340 5284
rect 6696 5244 6702 5256
rect 4062 5216 4068 5228
rect 4023 5188 4068 5216
rect 4062 5176 4068 5188
rect 4120 5176 4126 5228
rect 4249 5219 4307 5225
rect 4249 5185 4261 5219
rect 4295 5185 4307 5219
rect 5718 5216 5724 5228
rect 5679 5188 5724 5216
rect 4249 5179 4307 5185
rect 2958 5108 2964 5160
rect 3016 5148 3022 5160
rect 4264 5148 4292 5179
rect 5718 5176 5724 5188
rect 5776 5176 5782 5228
rect 8202 5148 8208 5160
rect 3016 5120 8208 5148
rect 3016 5108 3022 5120
rect 8202 5108 8208 5120
rect 8260 5108 8266 5160
rect 8312 5148 8340 5256
rect 9214 5244 9220 5296
rect 9272 5284 9278 5296
rect 18233 5287 18291 5293
rect 9272 5256 10364 5284
rect 9272 5244 9278 5256
rect 10336 5225 10364 5256
rect 18233 5253 18245 5287
rect 18279 5284 18291 5287
rect 18690 5284 18696 5296
rect 18279 5256 18696 5284
rect 18279 5253 18291 5256
rect 18233 5247 18291 5253
rect 18690 5244 18696 5256
rect 18748 5244 18754 5296
rect 23382 5284 23388 5296
rect 23343 5256 23388 5284
rect 23382 5244 23388 5256
rect 23440 5244 23446 5296
rect 25777 5287 25835 5293
rect 25777 5253 25789 5287
rect 25823 5284 25835 5287
rect 26050 5284 26056 5296
rect 25823 5256 26056 5284
rect 25823 5253 25835 5256
rect 25777 5247 25835 5253
rect 26050 5244 26056 5256
rect 26108 5244 26114 5296
rect 10321 5219 10379 5225
rect 10321 5185 10333 5219
rect 10367 5185 10379 5219
rect 10321 5179 10379 5185
rect 10505 5219 10563 5225
rect 10505 5185 10517 5219
rect 10551 5216 10563 5219
rect 10870 5216 10876 5228
rect 10551 5188 10876 5216
rect 10551 5185 10563 5188
rect 10505 5179 10563 5185
rect 10870 5176 10876 5188
rect 10928 5176 10934 5228
rect 11790 5176 11796 5228
rect 11848 5216 11854 5228
rect 11957 5219 12015 5225
rect 11957 5216 11969 5219
rect 11848 5188 11969 5216
rect 11848 5176 11854 5188
rect 11957 5185 11969 5188
rect 12003 5185 12015 5219
rect 15194 5216 15200 5228
rect 15155 5188 15200 5216
rect 11957 5179 12015 5185
rect 15194 5176 15200 5188
rect 15252 5176 15258 5228
rect 25961 5219 26019 5225
rect 25961 5185 25973 5219
rect 26007 5216 26019 5219
rect 26234 5216 26240 5228
rect 26007 5188 26240 5216
rect 26007 5185 26019 5188
rect 25961 5179 26019 5185
rect 26234 5176 26240 5188
rect 26292 5176 26298 5228
rect 9217 5151 9275 5157
rect 9217 5148 9229 5151
rect 8312 5120 9229 5148
rect 9217 5117 9229 5120
rect 9263 5117 9275 5151
rect 9217 5111 9275 5117
rect 9306 5108 9312 5160
rect 9364 5148 9370 5160
rect 9401 5151 9459 5157
rect 9401 5148 9413 5151
rect 9364 5120 9413 5148
rect 9364 5108 9370 5120
rect 9401 5117 9413 5120
rect 9447 5117 9459 5151
rect 11698 5148 11704 5160
rect 9401 5111 9459 5117
rect 9508 5120 11704 5148
rect 7190 5040 7196 5092
rect 7248 5080 7254 5092
rect 9508 5080 9536 5120
rect 11698 5108 11704 5120
rect 11756 5108 11762 5160
rect 7248 5052 9536 5080
rect 9861 5083 9919 5089
rect 7248 5040 7254 5052
rect 9861 5049 9873 5083
rect 9907 5080 9919 5083
rect 9907 5052 11192 5080
rect 9907 5049 9919 5052
rect 9861 5043 9919 5049
rect 11164 5012 11192 5052
rect 14826 5012 14832 5024
rect 11164 4984 14832 5012
rect 14826 4972 14832 4984
rect 14884 4972 14890 5024
rect 14918 4972 14924 5024
rect 14976 5012 14982 5024
rect 15105 5015 15163 5021
rect 15105 5012 15117 5015
rect 14976 4984 15117 5012
rect 14976 4972 14982 4984
rect 15105 4981 15117 4984
rect 15151 4981 15163 5015
rect 25590 5012 25596 5024
rect 25551 4984 25596 5012
rect 15105 4975 15163 4981
rect 25590 4972 25596 4984
rect 25648 4972 25654 5024
rect 1104 4922 34868 4944
rect 1104 4870 5170 4922
rect 5222 4870 5234 4922
rect 5286 4870 5298 4922
rect 5350 4870 5362 4922
rect 5414 4870 5426 4922
rect 5478 4870 13611 4922
rect 13663 4870 13675 4922
rect 13727 4870 13739 4922
rect 13791 4870 13803 4922
rect 13855 4870 13867 4922
rect 13919 4870 22052 4922
rect 22104 4870 22116 4922
rect 22168 4870 22180 4922
rect 22232 4870 22244 4922
rect 22296 4870 22308 4922
rect 22360 4870 30493 4922
rect 30545 4870 30557 4922
rect 30609 4870 30621 4922
rect 30673 4870 30685 4922
rect 30737 4870 30749 4922
rect 30801 4870 34868 4922
rect 1104 4848 34868 4870
rect 10870 4808 10876 4820
rect 10831 4780 10876 4808
rect 10870 4768 10876 4780
rect 10928 4768 10934 4820
rect 11882 4768 11888 4820
rect 11940 4808 11946 4820
rect 11977 4811 12035 4817
rect 11977 4808 11989 4811
rect 11940 4780 11989 4808
rect 11940 4768 11946 4780
rect 11977 4777 11989 4780
rect 12023 4777 12035 4811
rect 11977 4771 12035 4777
rect 13262 4768 13268 4820
rect 13320 4808 13326 4820
rect 26234 4808 26240 4820
rect 13320 4780 22094 4808
rect 13320 4768 13326 4780
rect 5074 4632 5080 4684
rect 5132 4672 5138 4684
rect 7190 4672 7196 4684
rect 5132 4644 7196 4672
rect 5132 4632 5138 4644
rect 7190 4632 7196 4644
rect 7248 4632 7254 4684
rect 8938 4632 8944 4684
rect 8996 4672 9002 4684
rect 9125 4675 9183 4681
rect 9125 4672 9137 4675
rect 8996 4644 9137 4672
rect 8996 4632 9002 4644
rect 9125 4641 9137 4644
rect 9171 4641 9183 4675
rect 9125 4635 9183 4641
rect 7466 4613 7472 4616
rect 7460 4604 7472 4613
rect 7427 4576 7472 4604
rect 7460 4567 7472 4576
rect 7466 4564 7472 4567
rect 7524 4564 7530 4616
rect 10888 4604 10916 4768
rect 14553 4743 14611 4749
rect 14553 4709 14565 4743
rect 14599 4740 14611 4743
rect 20714 4740 20720 4752
rect 14599 4712 20720 4740
rect 14599 4709 14611 4712
rect 14553 4703 14611 4709
rect 20714 4700 20720 4712
rect 20772 4700 20778 4752
rect 14182 4632 14188 4684
rect 14240 4672 14246 4684
rect 16209 4675 16267 4681
rect 16209 4672 16221 4675
rect 14240 4644 16221 4672
rect 14240 4632 14246 4644
rect 11885 4607 11943 4613
rect 11885 4604 11897 4607
rect 10888 4576 11897 4604
rect 11885 4573 11897 4576
rect 11931 4573 11943 4607
rect 11885 4567 11943 4573
rect 12253 4607 12311 4613
rect 12253 4573 12265 4607
rect 12299 4604 12311 4607
rect 12342 4604 12348 4616
rect 12299 4576 12348 4604
rect 12299 4573 12311 4576
rect 12253 4567 12311 4573
rect 12342 4564 12348 4576
rect 12400 4564 12406 4616
rect 14274 4604 14280 4616
rect 14235 4576 14280 4604
rect 14274 4564 14280 4576
rect 14332 4564 14338 4616
rect 14568 4613 14596 4644
rect 16209 4641 16221 4644
rect 16255 4672 16267 4675
rect 18693 4675 18751 4681
rect 18693 4672 18705 4675
rect 16255 4644 18705 4672
rect 16255 4641 16267 4644
rect 16209 4635 16267 4641
rect 18693 4641 18705 4644
rect 18739 4672 18751 4675
rect 20438 4672 20444 4684
rect 18739 4644 20444 4672
rect 18739 4641 18751 4644
rect 18693 4635 18751 4641
rect 20438 4632 20444 4644
rect 20496 4632 20502 4684
rect 22066 4672 22094 4780
rect 24596 4780 26240 4808
rect 24596 4681 24624 4780
rect 26234 4768 26240 4780
rect 26292 4808 26298 4820
rect 26602 4808 26608 4820
rect 26292 4780 26608 4808
rect 26292 4768 26298 4780
rect 26602 4768 26608 4780
rect 26660 4768 26666 4820
rect 24946 4740 24952 4752
rect 24907 4712 24952 4740
rect 24946 4700 24952 4712
rect 25004 4700 25010 4752
rect 24581 4675 24639 4681
rect 24581 4672 24593 4675
rect 22066 4644 24593 4672
rect 24581 4641 24593 4644
rect 24627 4641 24639 4675
rect 24581 4635 24639 4641
rect 14553 4607 14611 4613
rect 14553 4573 14565 4607
rect 14599 4573 14611 4607
rect 15930 4604 15936 4616
rect 15891 4576 15936 4604
rect 14553 4567 14611 4573
rect 15930 4564 15936 4576
rect 15988 4564 15994 4616
rect 17310 4564 17316 4616
rect 17368 4604 17374 4616
rect 17405 4607 17463 4613
rect 17405 4604 17417 4607
rect 17368 4576 17417 4604
rect 17368 4564 17374 4576
rect 17405 4573 17417 4576
rect 17451 4573 17463 4607
rect 18414 4604 18420 4616
rect 18375 4576 18420 4604
rect 17405 4567 17463 4573
rect 18414 4564 18420 4576
rect 18472 4564 18478 4616
rect 20162 4604 20168 4616
rect 20123 4576 20168 4604
rect 20162 4564 20168 4576
rect 20220 4564 20226 4616
rect 20898 4564 20904 4616
rect 20956 4604 20962 4616
rect 21637 4607 21695 4613
rect 21637 4604 21649 4607
rect 20956 4576 21649 4604
rect 20956 4564 20962 4576
rect 21637 4573 21649 4576
rect 21683 4604 21695 4607
rect 22281 4607 22339 4613
rect 22281 4604 22293 4607
rect 21683 4576 22293 4604
rect 21683 4573 21695 4576
rect 21637 4567 21695 4573
rect 22281 4573 22293 4576
rect 22327 4573 22339 4607
rect 25866 4604 25872 4616
rect 25827 4576 25872 4604
rect 22281 4567 22339 4573
rect 25866 4564 25872 4576
rect 25924 4564 25930 4616
rect 9401 4539 9459 4545
rect 9401 4505 9413 4539
rect 9447 4505 9459 4539
rect 9401 4499 9459 4505
rect 8570 4468 8576 4480
rect 8531 4440 8576 4468
rect 8570 4428 8576 4440
rect 8628 4428 8634 4480
rect 9416 4468 9444 4499
rect 10410 4496 10416 4548
rect 10468 4496 10474 4548
rect 26142 4545 26148 4548
rect 26136 4499 26148 4545
rect 26200 4536 26206 4548
rect 26200 4508 26236 4536
rect 26142 4496 26148 4499
rect 26200 4496 26206 4508
rect 11790 4468 11796 4480
rect 9416 4440 11796 4468
rect 11790 4428 11796 4440
rect 11848 4428 11854 4480
rect 12437 4471 12495 4477
rect 12437 4437 12449 4471
rect 12483 4468 12495 4471
rect 14369 4471 14427 4477
rect 14369 4468 14381 4471
rect 12483 4440 14381 4468
rect 12483 4437 12495 4440
rect 12437 4431 12495 4437
rect 14369 4437 14381 4440
rect 14415 4437 14427 4471
rect 15562 4468 15568 4480
rect 15523 4440 15568 4468
rect 14369 4431 14427 4437
rect 15562 4428 15568 4440
rect 15620 4428 15626 4480
rect 16025 4471 16083 4477
rect 16025 4437 16037 4471
rect 16071 4468 16083 4471
rect 16298 4468 16304 4480
rect 16071 4440 16304 4468
rect 16071 4437 16083 4440
rect 16025 4431 16083 4437
rect 16298 4428 16304 4440
rect 16356 4428 16362 4480
rect 17494 4468 17500 4480
rect 17455 4440 17500 4468
rect 17494 4428 17500 4440
rect 17552 4428 17558 4480
rect 18049 4471 18107 4477
rect 18049 4437 18061 4471
rect 18095 4468 18107 4471
rect 18230 4468 18236 4480
rect 18095 4440 18236 4468
rect 18095 4437 18107 4440
rect 18049 4431 18107 4437
rect 18230 4428 18236 4440
rect 18288 4428 18294 4480
rect 18509 4471 18567 4477
rect 18509 4437 18521 4471
rect 18555 4468 18567 4471
rect 19058 4468 19064 4480
rect 18555 4440 19064 4468
rect 18555 4437 18567 4440
rect 18509 4431 18567 4437
rect 19058 4428 19064 4440
rect 19116 4428 19122 4480
rect 19794 4468 19800 4480
rect 19755 4440 19800 4468
rect 19794 4428 19800 4440
rect 19852 4428 19858 4480
rect 20257 4471 20315 4477
rect 20257 4437 20269 4471
rect 20303 4468 20315 4471
rect 20806 4468 20812 4480
rect 20303 4440 20812 4468
rect 20303 4437 20315 4440
rect 20257 4431 20315 4437
rect 20806 4428 20812 4440
rect 20864 4428 20870 4480
rect 21542 4468 21548 4480
rect 21503 4440 21548 4468
rect 21542 4428 21548 4440
rect 21600 4428 21606 4480
rect 22094 4428 22100 4480
rect 22152 4468 22158 4480
rect 22189 4471 22247 4477
rect 22189 4468 22201 4471
rect 22152 4440 22201 4468
rect 22152 4428 22158 4440
rect 22189 4437 22201 4440
rect 22235 4437 22247 4471
rect 25038 4468 25044 4480
rect 24999 4440 25044 4468
rect 22189 4431 22247 4437
rect 25038 4428 25044 4440
rect 25096 4428 25102 4480
rect 27246 4468 27252 4480
rect 27207 4440 27252 4468
rect 27246 4428 27252 4440
rect 27304 4428 27310 4480
rect 1104 4378 35027 4400
rect 1104 4326 9390 4378
rect 9442 4326 9454 4378
rect 9506 4326 9518 4378
rect 9570 4326 9582 4378
rect 9634 4326 9646 4378
rect 9698 4326 17831 4378
rect 17883 4326 17895 4378
rect 17947 4326 17959 4378
rect 18011 4326 18023 4378
rect 18075 4326 18087 4378
rect 18139 4326 26272 4378
rect 26324 4326 26336 4378
rect 26388 4326 26400 4378
rect 26452 4326 26464 4378
rect 26516 4326 26528 4378
rect 26580 4326 34713 4378
rect 34765 4326 34777 4378
rect 34829 4326 34841 4378
rect 34893 4326 34905 4378
rect 34957 4326 34969 4378
rect 35021 4326 35027 4378
rect 1104 4304 35027 4326
rect 7466 4224 7472 4276
rect 7524 4224 7530 4276
rect 8570 4224 8576 4276
rect 8628 4264 8634 4276
rect 9677 4267 9735 4273
rect 9677 4264 9689 4267
rect 8628 4236 9689 4264
rect 8628 4224 8634 4236
rect 9677 4233 9689 4236
rect 9723 4233 9735 4267
rect 13354 4264 13360 4276
rect 13315 4236 13360 4264
rect 9677 4227 9735 4233
rect 13354 4224 13360 4236
rect 13412 4224 13418 4276
rect 14826 4224 14832 4276
rect 14884 4264 14890 4276
rect 22462 4264 22468 4276
rect 14884 4236 22468 4264
rect 14884 4224 14890 4236
rect 22462 4224 22468 4236
rect 22520 4224 22526 4276
rect 26142 4264 26148 4276
rect 26103 4236 26148 4264
rect 26142 4224 26148 4236
rect 26200 4224 26206 4276
rect 7285 4199 7343 4205
rect 7285 4165 7297 4199
rect 7331 4196 7343 4199
rect 7484 4196 7512 4224
rect 7331 4168 7512 4196
rect 7331 4165 7343 4168
rect 7285 4159 7343 4165
rect 7926 4156 7932 4208
rect 7984 4156 7990 4208
rect 9214 4156 9220 4208
rect 9272 4196 9278 4208
rect 9585 4199 9643 4205
rect 9585 4196 9597 4199
rect 9272 4168 9597 4196
rect 9272 4156 9278 4168
rect 9585 4165 9597 4168
rect 9631 4165 9643 4199
rect 9585 4159 9643 4165
rect 15188 4199 15246 4205
rect 15188 4165 15200 4199
rect 15234 4196 15246 4199
rect 15562 4196 15568 4208
rect 15234 4168 15568 4196
rect 15234 4165 15246 4168
rect 15188 4159 15246 4165
rect 15562 4156 15568 4168
rect 15620 4156 15626 4208
rect 25440 4199 25498 4205
rect 17328 4168 18092 4196
rect 8938 4128 8944 4140
rect 8496 4100 8944 4128
rect 7009 4063 7067 4069
rect 7009 4029 7021 4063
rect 7055 4060 7067 4063
rect 8496 4060 8524 4100
rect 8938 4088 8944 4100
rect 8996 4088 9002 4140
rect 7055 4032 8524 4060
rect 8757 4063 8815 4069
rect 7055 4029 7067 4032
rect 7009 4023 7067 4029
rect 8757 4029 8769 4063
rect 8803 4060 8815 4063
rect 9232 4060 9260 4156
rect 17328 4140 17356 4168
rect 10410 4128 10416 4140
rect 10371 4100 10416 4128
rect 10410 4088 10416 4100
rect 10468 4088 10474 4140
rect 10502 4088 10508 4140
rect 10560 4128 10566 4140
rect 10778 4128 10784 4140
rect 10560 4100 10605 4128
rect 10739 4100 10784 4128
rect 10560 4088 10566 4100
rect 10778 4088 10784 4100
rect 10836 4088 10842 4140
rect 13449 4131 13507 4137
rect 13449 4097 13461 4131
rect 13495 4128 13507 4131
rect 13998 4128 14004 4140
rect 13495 4100 14004 4128
rect 13495 4097 13507 4100
rect 13449 4091 13507 4097
rect 13998 4088 14004 4100
rect 14056 4088 14062 4140
rect 14918 4128 14924 4140
rect 14879 4100 14924 4128
rect 14918 4088 14924 4100
rect 14976 4088 14982 4140
rect 17037 4131 17095 4137
rect 17037 4097 17049 4131
rect 17083 4128 17095 4131
rect 17310 4128 17316 4140
rect 17083 4100 17316 4128
rect 17083 4097 17095 4100
rect 17037 4091 17095 4097
rect 17310 4088 17316 4100
rect 17368 4088 17374 4140
rect 17494 4088 17500 4140
rect 17552 4128 17558 4140
rect 17954 4137 17960 4140
rect 17681 4131 17739 4137
rect 17681 4128 17693 4131
rect 17552 4100 17693 4128
rect 17552 4088 17558 4100
rect 17681 4097 17693 4100
rect 17727 4097 17739 4131
rect 17948 4128 17960 4137
rect 17915 4100 17960 4128
rect 17681 4091 17739 4097
rect 17948 4091 17960 4100
rect 17954 4088 17960 4091
rect 18012 4088 18018 4140
rect 18064 4128 18092 4168
rect 25440 4165 25452 4199
rect 25486 4196 25498 4199
rect 25590 4196 25596 4208
rect 25486 4168 25596 4196
rect 25486 4165 25498 4168
rect 25440 4159 25498 4165
rect 25590 4156 25596 4168
rect 25648 4156 25654 4208
rect 28184 4168 28488 4196
rect 20898 4128 20904 4140
rect 18064 4100 20904 4128
rect 20898 4088 20904 4100
rect 20956 4088 20962 4140
rect 21174 4128 21180 4140
rect 21232 4137 21238 4140
rect 21144 4100 21180 4128
rect 21174 4088 21180 4100
rect 21232 4091 21244 4137
rect 21453 4131 21511 4137
rect 21453 4097 21465 4131
rect 21499 4128 21511 4131
rect 21542 4128 21548 4140
rect 21499 4100 21548 4128
rect 21499 4097 21511 4100
rect 21453 4091 21511 4097
rect 21232 4088 21238 4091
rect 21542 4088 21548 4100
rect 21600 4088 21606 4140
rect 22005 4131 22063 4137
rect 22005 4097 22017 4131
rect 22051 4128 22063 4131
rect 22094 4128 22100 4140
rect 22051 4100 22100 4128
rect 22051 4097 22063 4100
rect 22005 4091 22063 4097
rect 22094 4088 22100 4100
rect 22152 4088 22158 4140
rect 22278 4137 22284 4140
rect 22272 4091 22284 4137
rect 22336 4128 22342 4140
rect 25685 4131 25743 4137
rect 22336 4100 22372 4128
rect 22278 4088 22284 4091
rect 22336 4088 22342 4100
rect 25685 4097 25697 4131
rect 25731 4128 25743 4131
rect 25866 4128 25872 4140
rect 25731 4100 25872 4128
rect 25731 4097 25743 4100
rect 25685 4091 25743 4097
rect 25866 4088 25872 4100
rect 25924 4128 25930 4140
rect 28184 4128 28212 4168
rect 28460 4140 28488 4168
rect 25924 4100 28212 4128
rect 25924 4088 25930 4100
rect 28258 4088 28264 4140
rect 28316 4137 28322 4140
rect 28316 4128 28328 4137
rect 28316 4100 28361 4128
rect 28316 4091 28328 4100
rect 28316 4088 28322 4091
rect 28442 4088 28448 4140
rect 28500 4128 28506 4140
rect 28537 4131 28595 4137
rect 28537 4128 28549 4131
rect 28500 4100 28549 4128
rect 28500 4088 28506 4100
rect 28537 4097 28549 4100
rect 28583 4097 28595 4131
rect 28537 4091 28595 4097
rect 8803 4032 9260 4060
rect 9861 4063 9919 4069
rect 8803 4029 8815 4032
rect 8757 4023 8815 4029
rect 9861 4029 9873 4063
rect 9907 4060 9919 4063
rect 11882 4060 11888 4072
rect 9907 4032 11888 4060
rect 9907 4029 9919 4032
rect 9861 4023 9919 4029
rect 11882 4020 11888 4032
rect 11940 4020 11946 4072
rect 13633 4063 13691 4069
rect 13633 4029 13645 4063
rect 13679 4060 13691 4063
rect 14182 4060 14188 4072
rect 13679 4032 14188 4060
rect 13679 4029 13691 4032
rect 13633 4023 13691 4029
rect 14182 4020 14188 4032
rect 14240 4020 14246 4072
rect 26602 4060 26608 4072
rect 26563 4032 26608 4060
rect 26602 4020 26608 4032
rect 26660 4020 26666 4072
rect 9217 3995 9275 4001
rect 9217 3961 9229 3995
rect 9263 3992 9275 3995
rect 9306 3992 9312 4004
rect 9263 3964 9312 3992
rect 9263 3961 9275 3964
rect 9217 3955 9275 3961
rect 9306 3952 9312 3964
rect 9364 3952 9370 4004
rect 26234 3992 26240 4004
rect 26195 3964 26240 3992
rect 26234 3952 26240 3964
rect 26292 3952 26298 4004
rect 12986 3924 12992 3936
rect 12947 3896 12992 3924
rect 12986 3884 12992 3896
rect 13044 3884 13050 3936
rect 16298 3924 16304 3936
rect 16259 3896 16304 3924
rect 16298 3884 16304 3896
rect 16356 3884 16362 3936
rect 16666 3884 16672 3936
rect 16724 3924 16730 3936
rect 16945 3927 17003 3933
rect 16945 3924 16957 3927
rect 16724 3896 16957 3924
rect 16724 3884 16730 3896
rect 16945 3893 16957 3896
rect 16991 3893 17003 3927
rect 19058 3924 19064 3936
rect 19019 3896 19064 3924
rect 16945 3887 17003 3893
rect 19058 3884 19064 3896
rect 19116 3884 19122 3936
rect 20073 3927 20131 3933
rect 20073 3893 20085 3927
rect 20119 3924 20131 3927
rect 21082 3924 21088 3936
rect 20119 3896 21088 3924
rect 20119 3893 20131 3896
rect 20073 3887 20131 3893
rect 21082 3884 21088 3896
rect 21140 3884 21146 3936
rect 23382 3924 23388 3936
rect 23343 3896 23388 3924
rect 23382 3884 23388 3896
rect 23440 3884 23446 3936
rect 24305 3927 24363 3933
rect 24305 3893 24317 3927
rect 24351 3924 24363 3927
rect 24946 3924 24952 3936
rect 24351 3896 24952 3924
rect 24351 3893 24363 3896
rect 24305 3887 24363 3893
rect 24946 3884 24952 3896
rect 25004 3884 25010 3936
rect 27157 3927 27215 3933
rect 27157 3893 27169 3927
rect 27203 3924 27215 3927
rect 27614 3924 27620 3936
rect 27203 3896 27620 3924
rect 27203 3893 27215 3896
rect 27157 3887 27215 3893
rect 27614 3884 27620 3896
rect 27672 3884 27678 3936
rect 1104 3834 34868 3856
rect 1104 3782 5170 3834
rect 5222 3782 5234 3834
rect 5286 3782 5298 3834
rect 5350 3782 5362 3834
rect 5414 3782 5426 3834
rect 5478 3782 13611 3834
rect 13663 3782 13675 3834
rect 13727 3782 13739 3834
rect 13791 3782 13803 3834
rect 13855 3782 13867 3834
rect 13919 3782 22052 3834
rect 22104 3782 22116 3834
rect 22168 3782 22180 3834
rect 22232 3782 22244 3834
rect 22296 3782 22308 3834
rect 22360 3782 30493 3834
rect 30545 3782 30557 3834
rect 30609 3782 30621 3834
rect 30673 3782 30685 3834
rect 30737 3782 30749 3834
rect 30801 3782 34868 3834
rect 1104 3760 34868 3782
rect 7926 3720 7932 3732
rect 7887 3692 7932 3720
rect 7926 3680 7932 3692
rect 7984 3680 7990 3732
rect 13725 3723 13783 3729
rect 13725 3689 13737 3723
rect 13771 3720 13783 3723
rect 13998 3720 14004 3732
rect 13771 3692 14004 3720
rect 13771 3689 13783 3692
rect 13725 3683 13783 3689
rect 13998 3680 14004 3692
rect 14056 3680 14062 3732
rect 20806 3680 20812 3732
rect 20864 3720 20870 3732
rect 20901 3723 20959 3729
rect 20901 3720 20913 3723
rect 20864 3692 20913 3720
rect 20864 3680 20870 3692
rect 20901 3689 20913 3692
rect 20947 3689 20959 3723
rect 20901 3683 20959 3689
rect 22097 3723 22155 3729
rect 22097 3689 22109 3723
rect 22143 3720 22155 3723
rect 22370 3720 22376 3732
rect 22143 3692 22376 3720
rect 22143 3689 22155 3692
rect 22097 3683 22155 3689
rect 22370 3680 22376 3692
rect 22428 3680 22434 3732
rect 26786 3720 26792 3732
rect 26699 3692 26792 3720
rect 26786 3680 26792 3692
rect 26844 3720 26850 3732
rect 27801 3723 27859 3729
rect 26844 3692 27200 3720
rect 26844 3680 26850 3692
rect 22066 3624 24624 3652
rect 9858 3584 9864 3596
rect 7944 3556 9864 3584
rect 7944 3525 7972 3556
rect 9858 3544 9864 3556
rect 9916 3584 9922 3596
rect 10778 3584 10784 3596
rect 9916 3556 10784 3584
rect 9916 3544 9922 3556
rect 10778 3544 10784 3556
rect 10836 3544 10842 3596
rect 16666 3584 16672 3596
rect 16627 3556 16672 3584
rect 16666 3544 16672 3556
rect 16724 3544 16730 3596
rect 7929 3519 7987 3525
rect 7929 3485 7941 3519
rect 7975 3485 7987 3519
rect 7929 3479 7987 3485
rect 8113 3519 8171 3525
rect 8113 3485 8125 3519
rect 8159 3516 8171 3519
rect 8202 3516 8208 3528
rect 8159 3488 8208 3516
rect 8159 3485 8171 3488
rect 8113 3479 8171 3485
rect 8202 3476 8208 3488
rect 8260 3516 8266 3528
rect 10502 3516 10508 3528
rect 8260 3488 10508 3516
rect 8260 3476 8266 3488
rect 10502 3476 10508 3488
rect 10560 3476 10566 3528
rect 12342 3516 12348 3528
rect 12303 3488 12348 3516
rect 12342 3476 12348 3488
rect 12400 3476 12406 3528
rect 12612 3519 12670 3525
rect 12612 3485 12624 3519
rect 12658 3516 12670 3519
rect 12986 3516 12992 3528
rect 12658 3488 12992 3516
rect 12658 3485 12670 3488
rect 12612 3479 12670 3485
rect 12986 3476 12992 3488
rect 13044 3476 13050 3528
rect 15654 3516 15660 3528
rect 15615 3488 15660 3516
rect 15654 3476 15660 3488
rect 15712 3476 15718 3528
rect 16758 3476 16764 3528
rect 16816 3516 16822 3528
rect 19518 3516 19524 3528
rect 16816 3488 17172 3516
rect 19479 3488 19524 3516
rect 16816 3476 16822 3488
rect 14734 3408 14740 3460
rect 14792 3448 14798 3460
rect 16942 3457 16948 3460
rect 15390 3451 15448 3457
rect 15390 3448 15402 3451
rect 14792 3420 15402 3448
rect 14792 3408 14798 3420
rect 15390 3417 15402 3420
rect 15436 3417 15448 3451
rect 15390 3411 15448 3417
rect 16936 3411 16948 3457
rect 17000 3448 17006 3460
rect 17144 3448 17172 3488
rect 19518 3476 19524 3488
rect 19576 3476 19582 3528
rect 19794 3525 19800 3528
rect 19788 3516 19800 3525
rect 19755 3488 19800 3516
rect 19788 3479 19800 3488
rect 19794 3476 19800 3479
rect 19852 3476 19858 3528
rect 20898 3476 20904 3528
rect 20956 3516 20962 3528
rect 22066 3516 22094 3624
rect 22738 3584 22744 3596
rect 22699 3556 22744 3584
rect 22738 3544 22744 3556
rect 22796 3544 22802 3596
rect 20956 3488 22094 3516
rect 20956 3476 20962 3488
rect 22462 3476 22468 3528
rect 22520 3516 22526 3528
rect 24596 3525 24624 3624
rect 25590 3612 25596 3664
rect 25648 3652 25654 3664
rect 26421 3655 26479 3661
rect 26421 3652 26433 3655
rect 25648 3624 26433 3652
rect 25648 3612 25654 3624
rect 26421 3621 26433 3624
rect 26467 3621 26479 3655
rect 26421 3615 26479 3621
rect 26881 3655 26939 3661
rect 26881 3621 26893 3655
rect 26927 3652 26939 3655
rect 27172 3652 27200 3692
rect 27801 3689 27813 3723
rect 27847 3720 27859 3723
rect 28258 3720 28264 3732
rect 27847 3692 28264 3720
rect 27847 3689 27859 3692
rect 27801 3683 27859 3689
rect 28258 3680 28264 3692
rect 28316 3680 28322 3732
rect 27246 3652 27252 3664
rect 26927 3624 27108 3652
rect 27159 3624 27252 3652
rect 26927 3621 26939 3624
rect 26881 3615 26939 3621
rect 26234 3544 26240 3596
rect 26292 3584 26298 3596
rect 26973 3587 27031 3593
rect 26973 3584 26985 3587
rect 26292 3556 26985 3584
rect 26292 3544 26298 3556
rect 26973 3553 26985 3556
rect 27019 3553 27031 3587
rect 26973 3547 27031 3553
rect 27080 3584 27108 3624
rect 27246 3612 27252 3624
rect 27304 3652 27310 3664
rect 27890 3652 27896 3664
rect 27304 3624 27896 3652
rect 27304 3612 27310 3624
rect 27890 3612 27896 3624
rect 27948 3612 27954 3664
rect 27614 3584 27620 3596
rect 27080 3556 27620 3584
rect 24581 3519 24639 3525
rect 22520 3488 22565 3516
rect 22520 3476 22526 3488
rect 24581 3485 24593 3519
rect 24627 3516 24639 3519
rect 25866 3516 25872 3528
rect 24627 3488 25872 3516
rect 24627 3485 24639 3488
rect 24581 3479 24639 3485
rect 25866 3476 25872 3488
rect 25924 3476 25930 3528
rect 26050 3476 26056 3528
rect 26108 3516 26114 3528
rect 27080 3516 27108 3556
rect 27614 3544 27620 3556
rect 27672 3584 27678 3596
rect 28350 3584 28356 3596
rect 27672 3556 28356 3584
rect 27672 3544 27678 3556
rect 28350 3544 28356 3556
rect 28408 3544 28414 3596
rect 26108 3488 27108 3516
rect 26108 3476 26114 3488
rect 22557 3451 22615 3457
rect 17000 3420 17036 3448
rect 17144 3420 22094 3448
rect 16942 3408 16948 3411
rect 17000 3408 17006 3420
rect 14274 3380 14280 3392
rect 14235 3352 14280 3380
rect 14274 3340 14280 3352
rect 14332 3340 14338 3392
rect 18049 3383 18107 3389
rect 18049 3349 18061 3383
rect 18095 3380 18107 3383
rect 18230 3380 18236 3392
rect 18095 3352 18236 3380
rect 18095 3349 18107 3352
rect 18049 3343 18107 3349
rect 18230 3340 18236 3352
rect 18288 3340 18294 3392
rect 22066 3380 22094 3420
rect 22557 3417 22569 3451
rect 22603 3448 22615 3451
rect 23382 3448 23388 3460
rect 22603 3420 23388 3448
rect 22603 3417 22615 3420
rect 22557 3411 22615 3417
rect 23382 3408 23388 3420
rect 23440 3408 23446 3460
rect 24848 3451 24906 3457
rect 24848 3417 24860 3451
rect 24894 3448 24906 3451
rect 25038 3448 25044 3460
rect 24894 3420 25044 3448
rect 24894 3417 24906 3420
rect 24848 3411 24906 3417
rect 25038 3408 25044 3420
rect 25096 3408 25102 3460
rect 27341 3451 27399 3457
rect 27341 3448 27353 3451
rect 25148 3420 27353 3448
rect 25148 3380 25176 3420
rect 27341 3417 27353 3420
rect 27387 3417 27399 3451
rect 27341 3411 27399 3417
rect 28261 3451 28319 3457
rect 28261 3417 28273 3451
rect 28307 3417 28319 3451
rect 28261 3411 28319 3417
rect 25958 3380 25964 3392
rect 22066 3352 25176 3380
rect 25919 3352 25964 3380
rect 25958 3340 25964 3352
rect 26016 3380 26022 3392
rect 26234 3380 26240 3392
rect 26016 3352 26240 3380
rect 26016 3340 26022 3352
rect 26234 3340 26240 3352
rect 26292 3340 26298 3392
rect 26602 3340 26608 3392
rect 26660 3380 26666 3392
rect 28276 3380 28304 3411
rect 26660 3352 28304 3380
rect 26660 3340 26666 3352
rect 1104 3290 35027 3312
rect 1104 3238 9390 3290
rect 9442 3238 9454 3290
rect 9506 3238 9518 3290
rect 9570 3238 9582 3290
rect 9634 3238 9646 3290
rect 9698 3238 17831 3290
rect 17883 3238 17895 3290
rect 17947 3238 17959 3290
rect 18011 3238 18023 3290
rect 18075 3238 18087 3290
rect 18139 3238 26272 3290
rect 26324 3238 26336 3290
rect 26388 3238 26400 3290
rect 26452 3238 26464 3290
rect 26516 3238 26528 3290
rect 26580 3238 34713 3290
rect 34765 3238 34777 3290
rect 34829 3238 34841 3290
rect 34893 3238 34905 3290
rect 34957 3238 34969 3290
rect 35021 3238 35027 3290
rect 1104 3216 35027 3238
rect 12342 3136 12348 3188
rect 12400 3176 12406 3188
rect 12529 3179 12587 3185
rect 12529 3176 12541 3179
rect 12400 3148 12541 3176
rect 12400 3136 12406 3148
rect 12529 3145 12541 3148
rect 12575 3145 12587 3179
rect 14366 3176 14372 3188
rect 14327 3148 14372 3176
rect 12529 3139 12587 3145
rect 14366 3136 14372 3148
rect 14424 3136 14430 3188
rect 14734 3176 14740 3188
rect 14695 3148 14740 3176
rect 14734 3136 14740 3148
rect 14792 3136 14798 3188
rect 15289 3179 15347 3185
rect 15289 3145 15301 3179
rect 15335 3176 15347 3179
rect 15654 3176 15660 3188
rect 15335 3148 15660 3176
rect 15335 3145 15347 3148
rect 15289 3139 15347 3145
rect 15654 3136 15660 3148
rect 15712 3136 15718 3188
rect 16942 3176 16948 3188
rect 16903 3148 16948 3176
rect 16942 3136 16948 3148
rect 17000 3136 17006 3188
rect 17034 3136 17040 3188
rect 17092 3176 17098 3188
rect 17313 3179 17371 3185
rect 17313 3176 17325 3179
rect 17092 3148 17325 3176
rect 17092 3136 17098 3148
rect 17313 3145 17325 3148
rect 17359 3145 17371 3179
rect 17313 3139 17371 3145
rect 17405 3179 17463 3185
rect 17405 3145 17417 3179
rect 17451 3176 17463 3179
rect 18230 3176 18236 3188
rect 17451 3148 18236 3176
rect 17451 3145 17463 3148
rect 17405 3139 17463 3145
rect 18230 3136 18236 3148
rect 18288 3136 18294 3188
rect 19518 3136 19524 3188
rect 19576 3176 19582 3188
rect 19705 3179 19763 3185
rect 19705 3176 19717 3179
rect 19576 3148 19717 3176
rect 19576 3136 19582 3148
rect 19705 3145 19717 3148
rect 19751 3145 19763 3179
rect 19705 3139 19763 3145
rect 20898 3136 20904 3188
rect 20956 3136 20962 3188
rect 21082 3176 21088 3188
rect 21043 3148 21088 3176
rect 21082 3136 21088 3148
rect 21140 3136 21146 3188
rect 29089 3179 29147 3185
rect 29089 3145 29101 3179
rect 29135 3176 29147 3179
rect 29822 3176 29828 3188
rect 29135 3148 29828 3176
rect 29135 3145 29147 3148
rect 29089 3139 29147 3145
rect 29822 3136 29828 3148
rect 29880 3136 29886 3188
rect 20916 3108 20944 3136
rect 30374 3108 30380 3120
rect 12636 3080 15240 3108
rect 10778 3000 10784 3052
rect 10836 3040 10842 3052
rect 12636 3049 12664 3080
rect 15212 3052 15240 3080
rect 19812 3080 20944 3108
rect 30335 3080 30380 3108
rect 12621 3043 12679 3049
rect 12621 3040 12633 3043
rect 10836 3012 12633 3040
rect 10836 3000 10842 3012
rect 12621 3009 12633 3012
rect 12667 3009 12679 3043
rect 15194 3040 15200 3052
rect 15155 3012 15200 3040
rect 12621 3003 12679 3009
rect 15194 3000 15200 3012
rect 15252 3000 15258 3052
rect 19812 3049 19840 3080
rect 30374 3068 30380 3080
rect 30432 3068 30438 3120
rect 19797 3043 19855 3049
rect 19797 3009 19809 3043
rect 19843 3009 19855 3043
rect 19797 3003 19855 3009
rect 20714 3000 20720 3052
rect 20772 3040 20778 3052
rect 20901 3043 20959 3049
rect 20901 3040 20913 3043
rect 20772 3012 20913 3040
rect 20772 3000 20778 3012
rect 20901 3009 20913 3012
rect 20947 3009 20959 3043
rect 20901 3003 20959 3009
rect 21177 3043 21235 3049
rect 21177 3009 21189 3043
rect 21223 3040 21235 3043
rect 22738 3040 22744 3052
rect 21223 3012 22744 3040
rect 21223 3009 21235 3012
rect 21177 3003 21235 3009
rect 14182 2972 14188 2984
rect 14143 2944 14188 2972
rect 14182 2932 14188 2944
rect 14240 2932 14246 2984
rect 14274 2932 14280 2984
rect 14332 2972 14338 2984
rect 15470 2972 15476 2984
rect 14332 2944 15476 2972
rect 14332 2932 14338 2944
rect 15470 2932 15476 2944
rect 15528 2932 15534 2984
rect 17589 2975 17647 2981
rect 17589 2941 17601 2975
rect 17635 2972 17647 2975
rect 20438 2972 20444 2984
rect 17635 2944 20444 2972
rect 17635 2941 17647 2944
rect 17589 2935 17647 2941
rect 20438 2932 20444 2944
rect 20496 2972 20502 2984
rect 21192 2972 21220 3003
rect 22738 3000 22744 3012
rect 22796 3040 22802 3052
rect 25133 3043 25191 3049
rect 25133 3040 25145 3043
rect 22796 3012 25145 3040
rect 22796 3000 22802 3012
rect 25133 3009 25145 3012
rect 25179 3009 25191 3043
rect 25133 3003 25191 3009
rect 26053 3043 26111 3049
rect 26053 3009 26065 3043
rect 26099 3040 26111 3043
rect 26786 3040 26792 3052
rect 26099 3012 26792 3040
rect 26099 3009 26111 3012
rect 26053 3003 26111 3009
rect 26786 3000 26792 3012
rect 26844 3000 26850 3052
rect 20496 2944 21220 2972
rect 25501 2975 25559 2981
rect 20496 2932 20502 2944
rect 25501 2941 25513 2975
rect 25547 2972 25559 2975
rect 25958 2972 25964 2984
rect 25547 2944 25964 2972
rect 25547 2941 25559 2944
rect 25501 2935 25559 2941
rect 25958 2932 25964 2944
rect 26016 2972 26022 2984
rect 26234 2972 26240 2984
rect 26016 2944 26240 2972
rect 26016 2932 26022 2944
rect 26234 2932 26240 2944
rect 26292 2932 26298 2984
rect 20717 2907 20775 2913
rect 20717 2873 20729 2907
rect 20763 2904 20775 2907
rect 21174 2904 21180 2916
rect 20763 2876 21180 2904
rect 20763 2873 20775 2876
rect 20717 2867 20775 2873
rect 21174 2864 21180 2876
rect 21232 2864 21238 2916
rect 24946 2864 24952 2916
rect 25004 2904 25010 2916
rect 25590 2904 25596 2916
rect 25004 2876 25596 2904
rect 25004 2864 25010 2876
rect 25590 2864 25596 2876
rect 25648 2864 25654 2916
rect 25685 2907 25743 2913
rect 25685 2873 25697 2907
rect 25731 2904 25743 2907
rect 26050 2904 26056 2916
rect 25731 2876 26056 2904
rect 25731 2873 25743 2876
rect 25685 2867 25743 2873
rect 26050 2864 26056 2876
rect 26108 2864 26114 2916
rect 1104 2746 34868 2768
rect 1104 2694 5170 2746
rect 5222 2694 5234 2746
rect 5286 2694 5298 2746
rect 5350 2694 5362 2746
rect 5414 2694 5426 2746
rect 5478 2694 13611 2746
rect 13663 2694 13675 2746
rect 13727 2694 13739 2746
rect 13791 2694 13803 2746
rect 13855 2694 13867 2746
rect 13919 2694 22052 2746
rect 22104 2694 22116 2746
rect 22168 2694 22180 2746
rect 22232 2694 22244 2746
rect 22296 2694 22308 2746
rect 22360 2694 30493 2746
rect 30545 2694 30557 2746
rect 30609 2694 30621 2746
rect 30673 2694 30685 2746
rect 30737 2694 30749 2746
rect 30801 2694 34868 2746
rect 1104 2672 34868 2694
rect 15930 2632 15936 2644
rect 4448 2604 15936 2632
rect 2056 2468 4384 2496
rect 2056 2437 2084 2468
rect 2041 2431 2099 2437
rect 2041 2397 2053 2431
rect 2087 2397 2099 2431
rect 2041 2391 2099 2397
rect 3053 2431 3111 2437
rect 3053 2397 3065 2431
rect 3099 2397 3111 2431
rect 3053 2391 3111 2397
rect 1210 2320 1216 2372
rect 1268 2360 1274 2372
rect 1765 2363 1823 2369
rect 1765 2360 1777 2363
rect 1268 2332 1777 2360
rect 1268 2320 1274 2332
rect 1765 2329 1777 2332
rect 1811 2329 1823 2363
rect 1765 2323 1823 2329
rect 2498 2320 2504 2372
rect 2556 2360 2562 2372
rect 2777 2363 2835 2369
rect 2777 2360 2789 2363
rect 2556 2332 2789 2360
rect 2556 2320 2562 2332
rect 2777 2329 2789 2332
rect 2823 2329 2835 2363
rect 2777 2323 2835 2329
rect 3068 2292 3096 2391
rect 3786 2320 3792 2372
rect 3844 2360 3850 2372
rect 4157 2363 4215 2369
rect 4157 2360 4169 2363
rect 3844 2332 4169 2360
rect 3844 2320 3850 2332
rect 4157 2329 4169 2332
rect 4203 2329 4215 2363
rect 4356 2360 4384 2468
rect 4448 2437 4476 2604
rect 15930 2592 15936 2604
rect 15988 2592 15994 2644
rect 10042 2564 10048 2576
rect 5644 2536 10048 2564
rect 5644 2437 5672 2536
rect 10042 2524 10048 2536
rect 10100 2524 10106 2576
rect 18230 2496 18236 2508
rect 18064 2468 18236 2496
rect 4433 2431 4491 2437
rect 4433 2397 4445 2431
rect 4479 2397 4491 2431
rect 5629 2431 5687 2437
rect 4433 2391 4491 2397
rect 5000 2400 5488 2428
rect 5000 2360 5028 2400
rect 4356 2332 5028 2360
rect 4157 2323 4215 2329
rect 5074 2320 5080 2372
rect 5132 2360 5138 2372
rect 5353 2363 5411 2369
rect 5353 2360 5365 2363
rect 5132 2332 5365 2360
rect 5132 2320 5138 2332
rect 5353 2329 5365 2332
rect 5399 2329 5411 2363
rect 5460 2360 5488 2400
rect 5629 2397 5641 2431
rect 5675 2397 5687 2431
rect 5629 2391 5687 2397
rect 6362 2388 6368 2440
rect 6420 2428 6426 2440
rect 6549 2431 6607 2437
rect 6549 2428 6561 2431
rect 6420 2400 6561 2428
rect 6420 2388 6426 2400
rect 6549 2397 6561 2400
rect 6595 2397 6607 2431
rect 6549 2391 6607 2397
rect 7650 2388 7656 2440
rect 7708 2428 7714 2440
rect 7745 2431 7803 2437
rect 7745 2428 7757 2431
rect 7708 2400 7757 2428
rect 7708 2388 7714 2400
rect 7745 2397 7757 2400
rect 7791 2397 7803 2431
rect 7745 2391 7803 2397
rect 8938 2388 8944 2440
rect 8996 2428 9002 2440
rect 9125 2431 9183 2437
rect 9125 2428 9137 2431
rect 8996 2400 9137 2428
rect 8996 2388 9002 2400
rect 9125 2397 9137 2400
rect 9171 2397 9183 2431
rect 9125 2391 9183 2397
rect 10226 2388 10232 2440
rect 10284 2428 10290 2440
rect 10321 2431 10379 2437
rect 10321 2428 10333 2431
rect 10284 2400 10333 2428
rect 10284 2388 10290 2400
rect 10321 2397 10333 2400
rect 10367 2397 10379 2431
rect 10321 2391 10379 2397
rect 11514 2388 11520 2440
rect 11572 2428 11578 2440
rect 11701 2431 11759 2437
rect 11701 2428 11713 2431
rect 11572 2400 11713 2428
rect 11572 2388 11578 2400
rect 11701 2397 11713 2400
rect 11747 2397 11759 2431
rect 11701 2391 11759 2397
rect 12802 2388 12808 2440
rect 12860 2428 12866 2440
rect 12897 2431 12955 2437
rect 12897 2428 12909 2431
rect 12860 2400 12909 2428
rect 12860 2388 12866 2400
rect 12897 2397 12909 2400
rect 12943 2397 12955 2431
rect 12897 2391 12955 2397
rect 13998 2388 14004 2440
rect 14056 2428 14062 2440
rect 14277 2431 14335 2437
rect 14277 2428 14289 2431
rect 14056 2400 14289 2428
rect 14056 2388 14062 2400
rect 14277 2397 14289 2400
rect 14323 2397 14335 2431
rect 15470 2428 15476 2440
rect 15431 2400 15476 2428
rect 14277 2391 14335 2397
rect 15470 2388 15476 2400
rect 15528 2388 15534 2440
rect 16298 2388 16304 2440
rect 16356 2428 16362 2440
rect 18064 2437 18092 2468
rect 18230 2456 18236 2468
rect 18288 2456 18294 2508
rect 20898 2456 20904 2508
rect 20956 2456 20962 2508
rect 16853 2431 16911 2437
rect 16853 2428 16865 2431
rect 16356 2400 16865 2428
rect 16356 2388 16362 2400
rect 16853 2397 16865 2400
rect 16899 2397 16911 2431
rect 16853 2391 16911 2397
rect 18049 2431 18107 2437
rect 18049 2397 18061 2431
rect 18095 2397 18107 2431
rect 18049 2391 18107 2397
rect 19058 2388 19064 2440
rect 19116 2428 19122 2440
rect 19429 2431 19487 2437
rect 19429 2428 19441 2431
rect 19116 2400 19441 2428
rect 19116 2388 19122 2400
rect 19429 2397 19441 2400
rect 19475 2397 19487 2431
rect 19429 2391 19487 2397
rect 20625 2431 20683 2437
rect 20625 2397 20637 2431
rect 20671 2428 20683 2431
rect 20916 2428 20944 2456
rect 20671 2400 20944 2428
rect 20671 2397 20683 2400
rect 20625 2391 20683 2397
rect 21082 2388 21088 2440
rect 21140 2428 21146 2440
rect 22005 2431 22063 2437
rect 22005 2428 22017 2431
rect 21140 2400 22017 2428
rect 21140 2388 21146 2400
rect 22005 2397 22017 2400
rect 22051 2397 22063 2431
rect 22005 2391 22063 2397
rect 23201 2431 23259 2437
rect 23201 2397 23213 2431
rect 23247 2428 23259 2431
rect 23382 2428 23388 2440
rect 23247 2400 23388 2428
rect 23247 2397 23259 2400
rect 23201 2391 23259 2397
rect 23382 2388 23388 2400
rect 23440 2388 23446 2440
rect 25041 2431 25099 2437
rect 25041 2397 25053 2431
rect 25087 2428 25099 2431
rect 25590 2428 25596 2440
rect 25087 2400 25596 2428
rect 25087 2397 25099 2400
rect 25041 2391 25099 2397
rect 25590 2388 25596 2400
rect 25648 2388 25654 2440
rect 26234 2388 26240 2440
rect 26292 2428 26298 2440
rect 27617 2431 27675 2437
rect 26292 2400 26337 2428
rect 26292 2388 26298 2400
rect 27617 2397 27629 2431
rect 27663 2428 27675 2431
rect 27890 2428 27896 2440
rect 27663 2400 27896 2428
rect 27663 2397 27675 2400
rect 27617 2391 27675 2397
rect 27890 2388 27896 2400
rect 27948 2388 27954 2440
rect 28350 2428 28356 2440
rect 28311 2400 28356 2428
rect 28350 2388 28356 2400
rect 28408 2388 28414 2440
rect 29546 2388 29552 2440
rect 29604 2428 29610 2440
rect 29733 2431 29791 2437
rect 29733 2428 29745 2431
rect 29604 2400 29745 2428
rect 29604 2388 29610 2400
rect 29733 2397 29745 2400
rect 29779 2397 29791 2431
rect 29733 2391 29791 2397
rect 30834 2388 30840 2440
rect 30892 2428 30898 2440
rect 30929 2431 30987 2437
rect 30929 2428 30941 2431
rect 30892 2400 30941 2428
rect 30892 2388 30898 2400
rect 30929 2397 30941 2400
rect 30975 2397 30987 2431
rect 30929 2391 30987 2397
rect 32122 2388 32128 2440
rect 32180 2428 32186 2440
rect 32309 2431 32367 2437
rect 32309 2428 32321 2431
rect 32180 2400 32321 2428
rect 32180 2388 32186 2400
rect 32309 2397 32321 2400
rect 32355 2397 32367 2431
rect 32309 2391 32367 2397
rect 33410 2388 33416 2440
rect 33468 2428 33474 2440
rect 33505 2431 33563 2437
rect 33505 2428 33517 2431
rect 33468 2400 33517 2428
rect 33468 2388 33474 2400
rect 33505 2397 33517 2400
rect 33551 2397 33563 2431
rect 33505 2391 33563 2397
rect 7834 2360 7840 2372
rect 5460 2332 7840 2360
rect 5353 2323 5411 2329
rect 7834 2320 7840 2332
rect 7892 2320 7898 2372
rect 14090 2320 14096 2372
rect 14148 2360 14154 2372
rect 14553 2363 14611 2369
rect 14553 2360 14565 2363
rect 14148 2332 14565 2360
rect 14148 2320 14154 2332
rect 14553 2329 14565 2332
rect 14599 2329 14611 2363
rect 14553 2323 14611 2329
rect 15378 2320 15384 2372
rect 15436 2360 15442 2372
rect 15749 2363 15807 2369
rect 15749 2360 15761 2363
rect 15436 2332 15761 2360
rect 15436 2320 15442 2332
rect 15749 2329 15761 2332
rect 15795 2329 15807 2363
rect 15749 2323 15807 2329
rect 16666 2320 16672 2372
rect 16724 2360 16730 2372
rect 17129 2363 17187 2369
rect 17129 2360 17141 2363
rect 16724 2332 17141 2360
rect 16724 2320 16730 2332
rect 17129 2329 17141 2332
rect 17175 2329 17187 2363
rect 17129 2323 17187 2329
rect 18230 2320 18236 2372
rect 18288 2360 18294 2372
rect 18325 2363 18383 2369
rect 18325 2360 18337 2363
rect 18288 2332 18337 2360
rect 18288 2320 18294 2332
rect 18325 2329 18337 2332
rect 18371 2329 18383 2363
rect 18325 2323 18383 2329
rect 19242 2320 19248 2372
rect 19300 2360 19306 2372
rect 19705 2363 19763 2369
rect 19705 2360 19717 2363
rect 19300 2332 19717 2360
rect 19300 2320 19306 2332
rect 19705 2329 19717 2332
rect 19751 2329 19763 2363
rect 19705 2323 19763 2329
rect 20530 2320 20536 2372
rect 20588 2360 20594 2372
rect 20901 2363 20959 2369
rect 20901 2360 20913 2363
rect 20588 2332 20913 2360
rect 20588 2320 20594 2332
rect 20901 2329 20913 2332
rect 20947 2329 20959 2363
rect 20901 2323 20959 2329
rect 21818 2320 21824 2372
rect 21876 2360 21882 2372
rect 22281 2363 22339 2369
rect 22281 2360 22293 2363
rect 21876 2332 22293 2360
rect 21876 2320 21882 2332
rect 22281 2329 22293 2332
rect 22327 2329 22339 2363
rect 22281 2323 22339 2329
rect 23106 2320 23112 2372
rect 23164 2360 23170 2372
rect 23477 2363 23535 2369
rect 23477 2360 23489 2363
rect 23164 2332 23489 2360
rect 23164 2320 23170 2332
rect 23477 2329 23489 2332
rect 23523 2329 23535 2363
rect 23477 2323 23535 2329
rect 24394 2320 24400 2372
rect 24452 2360 24458 2372
rect 24765 2363 24823 2369
rect 24765 2360 24777 2363
rect 24452 2332 24777 2360
rect 24452 2320 24458 2332
rect 24765 2329 24777 2332
rect 24811 2329 24823 2363
rect 24765 2323 24823 2329
rect 25682 2320 25688 2372
rect 25740 2360 25746 2372
rect 25961 2363 26019 2369
rect 25961 2360 25973 2363
rect 25740 2332 25973 2360
rect 25740 2320 25746 2332
rect 25961 2329 25973 2332
rect 26007 2329 26019 2363
rect 25961 2323 26019 2329
rect 26970 2320 26976 2372
rect 27028 2360 27034 2372
rect 27341 2363 27399 2369
rect 27341 2360 27353 2363
rect 27028 2332 27353 2360
rect 27028 2320 27034 2332
rect 27341 2329 27353 2332
rect 27387 2329 27399 2363
rect 27341 2323 27399 2329
rect 28258 2320 28264 2372
rect 28316 2360 28322 2372
rect 28629 2363 28687 2369
rect 28629 2360 28641 2363
rect 28316 2332 28641 2360
rect 28316 2320 28322 2332
rect 28629 2329 28641 2332
rect 28675 2329 28687 2363
rect 28629 2323 28687 2329
rect 14366 2292 14372 2304
rect 3068 2264 14372 2292
rect 14366 2252 14372 2264
rect 14424 2252 14430 2304
rect 34333 2295 34391 2301
rect 34333 2261 34345 2295
rect 34379 2292 34391 2295
rect 34606 2292 34612 2304
rect 34379 2264 34612 2292
rect 34379 2261 34391 2264
rect 34333 2255 34391 2261
rect 34606 2252 34612 2264
rect 34664 2252 34670 2304
rect 1104 2202 35027 2224
rect 1104 2150 9390 2202
rect 9442 2150 9454 2202
rect 9506 2150 9518 2202
rect 9570 2150 9582 2202
rect 9634 2150 9646 2202
rect 9698 2150 17831 2202
rect 17883 2150 17895 2202
rect 17947 2150 17959 2202
rect 18011 2150 18023 2202
rect 18075 2150 18087 2202
rect 18139 2150 26272 2202
rect 26324 2150 26336 2202
rect 26388 2150 26400 2202
rect 26452 2150 26464 2202
rect 26516 2150 26528 2202
rect 26580 2150 34713 2202
rect 34765 2150 34777 2202
rect 34829 2150 34841 2202
rect 34893 2150 34905 2202
rect 34957 2150 34969 2202
rect 35021 2150 35027 2202
rect 1104 2128 35027 2150
<< via1 >>
rect 9390 33702 9442 33754
rect 9454 33702 9506 33754
rect 9518 33702 9570 33754
rect 9582 33702 9634 33754
rect 9646 33702 9698 33754
rect 17831 33702 17883 33754
rect 17895 33702 17947 33754
rect 17959 33702 18011 33754
rect 18023 33702 18075 33754
rect 18087 33702 18139 33754
rect 26272 33702 26324 33754
rect 26336 33702 26388 33754
rect 26400 33702 26452 33754
rect 26464 33702 26516 33754
rect 26528 33702 26580 33754
rect 34713 33702 34765 33754
rect 34777 33702 34829 33754
rect 34841 33702 34893 33754
rect 34905 33702 34957 33754
rect 34969 33702 35021 33754
rect 4896 33575 4948 33584
rect 4896 33541 4905 33575
rect 4905 33541 4939 33575
rect 4939 33541 4948 33575
rect 4896 33532 4948 33541
rect 7840 33575 7892 33584
rect 7840 33541 7849 33575
rect 7849 33541 7883 33575
rect 7883 33541 7892 33575
rect 7840 33532 7892 33541
rect 10600 33532 10652 33584
rect 13820 33532 13872 33584
rect 16580 33532 16632 33584
rect 19432 33532 19484 33584
rect 22652 33575 22704 33584
rect 22652 33541 22661 33575
rect 22661 33541 22695 33575
rect 22695 33541 22704 33575
rect 22652 33532 22704 33541
rect 25596 33575 25648 33584
rect 25596 33541 25605 33575
rect 25605 33541 25639 33575
rect 25639 33541 25648 33575
rect 25596 33532 25648 33541
rect 28264 33532 28316 33584
rect 31484 33575 31536 33584
rect 31484 33541 31493 33575
rect 31493 33541 31527 33575
rect 31527 33541 31536 33575
rect 31484 33532 31536 33541
rect 34244 33575 34296 33584
rect 34244 33541 34253 33575
rect 34253 33541 34287 33575
rect 34287 33541 34296 33575
rect 34244 33532 34296 33541
rect 8024 33371 8076 33380
rect 8024 33337 8033 33371
rect 8033 33337 8067 33371
rect 8067 33337 8076 33371
rect 8024 33328 8076 33337
rect 12256 33328 12308 33380
rect 14280 33371 14332 33380
rect 14280 33337 14289 33371
rect 14289 33337 14323 33371
rect 14323 33337 14332 33371
rect 14280 33328 14332 33337
rect 16856 33371 16908 33380
rect 16856 33337 16865 33371
rect 16865 33337 16899 33371
rect 16899 33337 16908 33371
rect 16856 33328 16908 33337
rect 19524 33371 19576 33380
rect 19524 33337 19533 33371
rect 19533 33337 19567 33371
rect 19567 33337 19576 33371
rect 19524 33328 19576 33337
rect 22468 33371 22520 33380
rect 22468 33337 22477 33371
rect 22477 33337 22511 33371
rect 22511 33337 22520 33371
rect 22468 33328 22520 33337
rect 25412 33371 25464 33380
rect 25412 33337 25421 33371
rect 25421 33337 25455 33371
rect 25455 33337 25464 33371
rect 25412 33328 25464 33337
rect 28356 33371 28408 33380
rect 28356 33337 28365 33371
rect 28365 33337 28399 33371
rect 28399 33337 28408 33371
rect 28356 33328 28408 33337
rect 31300 33371 31352 33380
rect 31300 33337 31309 33371
rect 31309 33337 31343 33371
rect 31343 33337 31352 33371
rect 31300 33328 31352 33337
rect 33416 33328 33468 33380
rect 4988 33303 5040 33312
rect 4988 33269 4997 33303
rect 4997 33269 5031 33303
rect 5031 33269 5040 33303
rect 4988 33260 5040 33269
rect 5170 33158 5222 33210
rect 5234 33158 5286 33210
rect 5298 33158 5350 33210
rect 5362 33158 5414 33210
rect 5426 33158 5478 33210
rect 13611 33158 13663 33210
rect 13675 33158 13727 33210
rect 13739 33158 13791 33210
rect 13803 33158 13855 33210
rect 13867 33158 13919 33210
rect 22052 33158 22104 33210
rect 22116 33158 22168 33210
rect 22180 33158 22232 33210
rect 22244 33158 22296 33210
rect 22308 33158 22360 33210
rect 30493 33158 30545 33210
rect 30557 33158 30609 33210
rect 30621 33158 30673 33210
rect 30685 33158 30737 33210
rect 30749 33158 30801 33210
rect 10508 32852 10560 32904
rect 16856 32920 16908 32972
rect 20628 32963 20680 32972
rect 20628 32929 20637 32963
rect 20637 32929 20671 32963
rect 20671 32929 20680 32963
rect 20628 32920 20680 32929
rect 16212 32784 16264 32836
rect 16764 32784 16816 32836
rect 20536 32895 20588 32904
rect 20536 32861 20545 32895
rect 20545 32861 20579 32895
rect 20579 32861 20588 32895
rect 24584 32988 24636 33040
rect 20812 32920 20864 32972
rect 25412 32920 25464 32972
rect 20536 32852 20588 32861
rect 22928 32852 22980 32904
rect 28356 32784 28408 32836
rect 10140 32759 10192 32768
rect 10140 32725 10149 32759
rect 10149 32725 10183 32759
rect 10183 32725 10192 32759
rect 10140 32716 10192 32725
rect 13268 32716 13320 32768
rect 20812 32716 20864 32768
rect 21272 32716 21324 32768
rect 22008 32716 22060 32768
rect 9390 32614 9442 32666
rect 9454 32614 9506 32666
rect 9518 32614 9570 32666
rect 9582 32614 9634 32666
rect 9646 32614 9698 32666
rect 17831 32614 17883 32666
rect 17895 32614 17947 32666
rect 17959 32614 18011 32666
rect 18023 32614 18075 32666
rect 18087 32614 18139 32666
rect 26272 32614 26324 32666
rect 26336 32614 26388 32666
rect 26400 32614 26452 32666
rect 26464 32614 26516 32666
rect 26528 32614 26580 32666
rect 34713 32614 34765 32666
rect 34777 32614 34829 32666
rect 34841 32614 34893 32666
rect 34905 32614 34957 32666
rect 34969 32614 35021 32666
rect 12256 32555 12308 32564
rect 12256 32521 12265 32555
rect 12265 32521 12299 32555
rect 12299 32521 12308 32555
rect 12256 32512 12308 32521
rect 14280 32512 14332 32564
rect 10692 32444 10744 32496
rect 13268 32487 13320 32496
rect 13268 32453 13277 32487
rect 13277 32453 13311 32487
rect 13311 32453 13320 32487
rect 13268 32444 13320 32453
rect 22468 32512 22520 32564
rect 10508 32419 10560 32428
rect 10508 32385 10517 32419
rect 10517 32385 10551 32419
rect 10551 32385 10560 32419
rect 10508 32376 10560 32385
rect 17868 32376 17920 32428
rect 18236 32419 18288 32428
rect 18236 32385 18245 32419
rect 18245 32385 18279 32419
rect 18279 32385 18288 32419
rect 18236 32376 18288 32385
rect 12348 32351 12400 32360
rect 8576 32240 8628 32292
rect 12348 32317 12357 32351
rect 12357 32317 12391 32351
rect 12391 32317 12400 32351
rect 12348 32308 12400 32317
rect 13452 32240 13504 32292
rect 10048 32172 10100 32224
rect 10600 32215 10652 32224
rect 10600 32181 10609 32215
rect 10609 32181 10643 32215
rect 10643 32181 10652 32215
rect 10600 32172 10652 32181
rect 11980 32172 12032 32224
rect 13176 32172 13228 32224
rect 14004 32308 14056 32360
rect 17408 32351 17460 32360
rect 13636 32240 13688 32292
rect 17408 32317 17417 32351
rect 17417 32317 17451 32351
rect 17451 32317 17460 32351
rect 17408 32308 17460 32317
rect 19524 32240 19576 32292
rect 22008 32419 22060 32428
rect 22008 32385 22017 32419
rect 22017 32385 22051 32419
rect 22051 32385 22060 32419
rect 22008 32376 22060 32385
rect 22560 32376 22612 32428
rect 23296 32419 23348 32428
rect 21272 32351 21324 32360
rect 21272 32317 21281 32351
rect 21281 32317 21315 32351
rect 21315 32317 21324 32351
rect 21272 32308 21324 32317
rect 23296 32385 23305 32419
rect 23305 32385 23339 32419
rect 23339 32385 23348 32419
rect 23296 32376 23348 32385
rect 23388 32308 23440 32360
rect 24584 32376 24636 32428
rect 27712 32419 27764 32428
rect 27712 32385 27721 32419
rect 27721 32385 27755 32419
rect 27755 32385 27764 32419
rect 27712 32376 27764 32385
rect 28632 32419 28684 32428
rect 28632 32385 28641 32419
rect 28641 32385 28675 32419
rect 28675 32385 28684 32419
rect 28632 32376 28684 32385
rect 31300 32376 31352 32428
rect 33416 32419 33468 32428
rect 33416 32385 33425 32419
rect 33425 32385 33459 32419
rect 33459 32385 33468 32419
rect 33416 32376 33468 32385
rect 24768 32308 24820 32360
rect 21180 32240 21232 32292
rect 16764 32172 16816 32224
rect 18512 32172 18564 32224
rect 22744 32172 22796 32224
rect 22928 32172 22980 32224
rect 25044 32172 25096 32224
rect 30196 32172 30248 32224
rect 33232 32215 33284 32224
rect 33232 32181 33241 32215
rect 33241 32181 33275 32215
rect 33275 32181 33284 32215
rect 33232 32172 33284 32181
rect 5170 32070 5222 32122
rect 5234 32070 5286 32122
rect 5298 32070 5350 32122
rect 5362 32070 5414 32122
rect 5426 32070 5478 32122
rect 13611 32070 13663 32122
rect 13675 32070 13727 32122
rect 13739 32070 13791 32122
rect 13803 32070 13855 32122
rect 13867 32070 13919 32122
rect 22052 32070 22104 32122
rect 22116 32070 22168 32122
rect 22180 32070 22232 32122
rect 22244 32070 22296 32122
rect 22308 32070 22360 32122
rect 30493 32070 30545 32122
rect 30557 32070 30609 32122
rect 30621 32070 30673 32122
rect 30685 32070 30737 32122
rect 30749 32070 30801 32122
rect 8576 31900 8628 31952
rect 8760 31900 8812 31952
rect 10508 31968 10560 32020
rect 11704 31900 11756 31952
rect 9864 31875 9916 31884
rect 9864 31841 9873 31875
rect 9873 31841 9907 31875
rect 9907 31841 9916 31875
rect 9864 31832 9916 31841
rect 10140 31764 10192 31816
rect 12348 31764 12400 31816
rect 16120 31968 16172 32020
rect 18236 31968 18288 32020
rect 20628 31968 20680 32020
rect 23296 31968 23348 32020
rect 14004 31900 14056 31952
rect 16672 31900 16724 31952
rect 14004 31764 14056 31816
rect 14280 31807 14332 31816
rect 14280 31773 14289 31807
rect 14289 31773 14323 31807
rect 14323 31773 14332 31807
rect 14280 31764 14332 31773
rect 14648 31764 14700 31816
rect 20536 31900 20588 31952
rect 17132 31875 17184 31884
rect 17132 31841 17141 31875
rect 17141 31841 17175 31875
rect 17175 31841 17184 31875
rect 17132 31832 17184 31841
rect 22560 31900 22612 31952
rect 17316 31807 17368 31816
rect 17316 31773 17325 31807
rect 17325 31773 17359 31807
rect 17359 31773 17368 31807
rect 17316 31764 17368 31773
rect 17868 31764 17920 31816
rect 18512 31807 18564 31816
rect 18512 31773 18521 31807
rect 18521 31773 18555 31807
rect 18555 31773 18564 31807
rect 18512 31764 18564 31773
rect 22744 31832 22796 31884
rect 25044 31875 25096 31884
rect 25044 31841 25053 31875
rect 25053 31841 25087 31875
rect 25087 31841 25096 31875
rect 25044 31832 25096 31841
rect 25136 31875 25188 31884
rect 25136 31841 25145 31875
rect 25145 31841 25179 31875
rect 25179 31841 25188 31875
rect 25136 31832 25188 31841
rect 20812 31764 20864 31816
rect 21088 31764 21140 31816
rect 21180 31764 21232 31816
rect 22928 31807 22980 31816
rect 22928 31773 22937 31807
rect 22937 31773 22971 31807
rect 22971 31773 22980 31807
rect 22928 31764 22980 31773
rect 23756 31807 23808 31816
rect 23756 31773 23765 31807
rect 23765 31773 23799 31807
rect 23799 31773 23808 31807
rect 23756 31764 23808 31773
rect 26608 31807 26660 31816
rect 10048 31696 10100 31748
rect 15568 31739 15620 31748
rect 15568 31705 15577 31739
rect 15577 31705 15611 31739
rect 15611 31705 15620 31739
rect 15568 31696 15620 31705
rect 16120 31696 16172 31748
rect 8024 31628 8076 31680
rect 15752 31671 15804 31680
rect 15752 31637 15777 31671
rect 15777 31637 15804 31671
rect 15752 31628 15804 31637
rect 21272 31739 21324 31748
rect 21272 31705 21281 31739
rect 21281 31705 21315 31739
rect 21315 31705 21324 31739
rect 21272 31696 21324 31705
rect 22652 31696 22704 31748
rect 23388 31696 23440 31748
rect 26608 31773 26617 31807
rect 26617 31773 26651 31807
rect 26651 31773 26660 31807
rect 26608 31764 26660 31773
rect 27344 31807 27396 31816
rect 27344 31773 27353 31807
rect 27353 31773 27387 31807
rect 27387 31773 27396 31807
rect 27344 31764 27396 31773
rect 27712 31696 27764 31748
rect 23572 31671 23624 31680
rect 23572 31637 23581 31671
rect 23581 31637 23615 31671
rect 23615 31637 23624 31671
rect 23572 31628 23624 31637
rect 24584 31628 24636 31680
rect 24768 31628 24820 31680
rect 9390 31526 9442 31578
rect 9454 31526 9506 31578
rect 9518 31526 9570 31578
rect 9582 31526 9634 31578
rect 9646 31526 9698 31578
rect 17831 31526 17883 31578
rect 17895 31526 17947 31578
rect 17959 31526 18011 31578
rect 18023 31526 18075 31578
rect 18087 31526 18139 31578
rect 26272 31526 26324 31578
rect 26336 31526 26388 31578
rect 26400 31526 26452 31578
rect 26464 31526 26516 31578
rect 26528 31526 26580 31578
rect 34713 31526 34765 31578
rect 34777 31526 34829 31578
rect 34841 31526 34893 31578
rect 34905 31526 34957 31578
rect 34969 31526 35021 31578
rect 9864 31424 9916 31476
rect 14280 31424 14332 31476
rect 16120 31467 16172 31476
rect 16120 31433 16129 31467
rect 16129 31433 16163 31467
rect 16163 31433 16172 31467
rect 16120 31424 16172 31433
rect 17316 31424 17368 31476
rect 20812 31467 20864 31476
rect 20812 31433 20846 31467
rect 20846 31433 20864 31467
rect 20812 31424 20864 31433
rect 25136 31424 25188 31476
rect 26608 31424 26660 31476
rect 28632 31424 28684 31476
rect 10048 31356 10100 31408
rect 10600 31356 10652 31408
rect 9864 31288 9916 31340
rect 10232 31331 10284 31340
rect 10232 31297 10241 31331
rect 10241 31297 10275 31331
rect 10275 31297 10284 31331
rect 10232 31288 10284 31297
rect 9404 31220 9456 31272
rect 10048 31220 10100 31272
rect 13084 31288 13136 31340
rect 15568 31356 15620 31408
rect 20444 31356 20496 31408
rect 14096 31331 14148 31340
rect 14096 31297 14105 31331
rect 14105 31297 14139 31331
rect 14139 31297 14148 31331
rect 14096 31288 14148 31297
rect 14832 31331 14884 31340
rect 14832 31297 14841 31331
rect 14841 31297 14875 31331
rect 14875 31297 14884 31331
rect 14832 31288 14884 31297
rect 10416 31263 10468 31272
rect 10416 31229 10425 31263
rect 10425 31229 10459 31263
rect 10459 31229 10468 31263
rect 13268 31263 13320 31272
rect 10416 31220 10468 31229
rect 13268 31229 13277 31263
rect 13277 31229 13311 31263
rect 13311 31229 13320 31263
rect 13268 31220 13320 31229
rect 10968 31195 11020 31204
rect 10968 31161 10977 31195
rect 10977 31161 11011 31195
rect 11011 31161 11020 31195
rect 10968 31152 11020 31161
rect 10692 31084 10744 31136
rect 14280 31127 14332 31136
rect 14280 31093 14289 31127
rect 14289 31093 14323 31127
rect 14323 31093 14332 31127
rect 14280 31084 14332 31093
rect 14648 31220 14700 31272
rect 15476 31288 15528 31340
rect 16304 31331 16356 31340
rect 16304 31297 16313 31331
rect 16313 31297 16347 31331
rect 16347 31297 16356 31331
rect 16304 31288 16356 31297
rect 17132 31331 17184 31340
rect 17132 31297 17141 31331
rect 17141 31297 17175 31331
rect 17175 31297 17184 31331
rect 17132 31288 17184 31297
rect 15752 31220 15804 31272
rect 17684 31288 17736 31340
rect 20168 31288 20220 31340
rect 20996 31288 21048 31340
rect 22652 31331 22704 31340
rect 22652 31297 22661 31331
rect 22661 31297 22695 31331
rect 22695 31297 22704 31331
rect 22652 31288 22704 31297
rect 22744 31331 22796 31340
rect 22744 31297 22753 31331
rect 22753 31297 22787 31331
rect 22787 31297 22796 31331
rect 23020 31331 23072 31340
rect 22744 31288 22796 31297
rect 23020 31297 23029 31331
rect 23029 31297 23063 31331
rect 23063 31297 23072 31331
rect 23020 31288 23072 31297
rect 23572 31331 23624 31340
rect 20536 31263 20588 31272
rect 20536 31229 20545 31263
rect 20545 31229 20579 31263
rect 20579 31229 20588 31263
rect 20536 31220 20588 31229
rect 20904 31152 20956 31204
rect 21272 31152 21324 31204
rect 21456 31220 21508 31272
rect 23572 31297 23581 31331
rect 23581 31297 23615 31331
rect 23615 31297 23624 31331
rect 23572 31288 23624 31297
rect 24492 31288 24544 31340
rect 25044 31288 25096 31340
rect 25320 31288 25372 31340
rect 26056 31288 26108 31340
rect 27344 31331 27396 31340
rect 27344 31297 27353 31331
rect 27353 31297 27387 31331
rect 27387 31297 27396 31331
rect 27344 31288 27396 31297
rect 27528 31288 27580 31340
rect 27712 31288 27764 31340
rect 28540 31288 28592 31340
rect 25780 31220 25832 31272
rect 21732 31152 21784 31204
rect 22744 31152 22796 31204
rect 23572 31152 23624 31204
rect 28448 31195 28500 31204
rect 17040 31084 17092 31136
rect 28448 31161 28457 31195
rect 28457 31161 28491 31195
rect 28491 31161 28500 31195
rect 28448 31152 28500 31161
rect 25596 31084 25648 31136
rect 5170 30982 5222 31034
rect 5234 30982 5286 31034
rect 5298 30982 5350 31034
rect 5362 30982 5414 31034
rect 5426 30982 5478 31034
rect 13611 30982 13663 31034
rect 13675 30982 13727 31034
rect 13739 30982 13791 31034
rect 13803 30982 13855 31034
rect 13867 30982 13919 31034
rect 22052 30982 22104 31034
rect 22116 30982 22168 31034
rect 22180 30982 22232 31034
rect 22244 30982 22296 31034
rect 22308 30982 22360 31034
rect 30493 30982 30545 31034
rect 30557 30982 30609 31034
rect 30621 30982 30673 31034
rect 30685 30982 30737 31034
rect 30749 30982 30801 31034
rect 9404 30923 9456 30932
rect 9404 30889 9413 30923
rect 9413 30889 9447 30923
rect 9447 30889 9456 30923
rect 9404 30880 9456 30889
rect 10048 30923 10100 30932
rect 10048 30889 10057 30923
rect 10057 30889 10091 30923
rect 10091 30889 10100 30923
rect 10048 30880 10100 30889
rect 10232 30880 10284 30932
rect 13268 30880 13320 30932
rect 17408 30880 17460 30932
rect 20996 30923 21048 30932
rect 20996 30889 21005 30923
rect 21005 30889 21039 30923
rect 21039 30889 21048 30923
rect 20996 30880 21048 30889
rect 23020 30880 23072 30932
rect 14832 30812 14884 30864
rect 24952 30855 25004 30864
rect 10508 30744 10560 30796
rect 9956 30719 10008 30728
rect 9956 30685 9965 30719
rect 9965 30685 9999 30719
rect 9999 30685 10008 30719
rect 9956 30676 10008 30685
rect 10692 30676 10744 30728
rect 15752 30787 15804 30796
rect 15752 30753 15761 30787
rect 15761 30753 15795 30787
rect 15795 30753 15804 30787
rect 15752 30744 15804 30753
rect 10416 30608 10468 30660
rect 10508 30608 10560 30660
rect 14096 30676 14148 30728
rect 14556 30719 14608 30728
rect 14556 30685 14565 30719
rect 14565 30685 14599 30719
rect 14599 30685 14608 30719
rect 14556 30676 14608 30685
rect 14924 30719 14976 30728
rect 14924 30685 14933 30719
rect 14933 30685 14967 30719
rect 14967 30685 14976 30719
rect 14924 30676 14976 30685
rect 15476 30719 15528 30728
rect 15476 30685 15485 30719
rect 15485 30685 15519 30719
rect 15519 30685 15528 30719
rect 15476 30676 15528 30685
rect 24952 30821 24961 30855
rect 24961 30821 24995 30855
rect 24995 30821 25004 30855
rect 24952 30812 25004 30821
rect 16672 30676 16724 30728
rect 17040 30719 17092 30728
rect 17040 30685 17049 30719
rect 17049 30685 17083 30719
rect 17083 30685 17092 30719
rect 17040 30676 17092 30685
rect 21456 30676 21508 30728
rect 23388 30744 23440 30796
rect 23296 30719 23348 30728
rect 14004 30540 14056 30592
rect 16304 30608 16356 30660
rect 18788 30608 18840 30660
rect 23296 30685 23305 30719
rect 23305 30685 23339 30719
rect 23339 30685 23348 30719
rect 23296 30676 23348 30685
rect 25320 30676 25372 30728
rect 25596 30719 25648 30728
rect 25596 30685 25605 30719
rect 25605 30685 25639 30719
rect 25639 30685 25648 30719
rect 25596 30676 25648 30685
rect 25780 30719 25832 30728
rect 25780 30685 25789 30719
rect 25789 30685 25823 30719
rect 25823 30685 25832 30719
rect 25780 30676 25832 30685
rect 26056 30676 26108 30728
rect 27712 30676 27764 30728
rect 28080 30719 28132 30728
rect 28080 30685 28089 30719
rect 28089 30685 28123 30719
rect 28123 30685 28132 30719
rect 28080 30676 28132 30685
rect 28632 30719 28684 30728
rect 23756 30608 23808 30660
rect 25044 30608 25096 30660
rect 28632 30685 28641 30719
rect 28641 30685 28675 30719
rect 28675 30685 28684 30719
rect 28632 30676 28684 30685
rect 28540 30608 28592 30660
rect 9390 30438 9442 30490
rect 9454 30438 9506 30490
rect 9518 30438 9570 30490
rect 9582 30438 9634 30490
rect 9646 30438 9698 30490
rect 17831 30438 17883 30490
rect 17895 30438 17947 30490
rect 17959 30438 18011 30490
rect 18023 30438 18075 30490
rect 18087 30438 18139 30490
rect 26272 30438 26324 30490
rect 26336 30438 26388 30490
rect 26400 30438 26452 30490
rect 26464 30438 26516 30490
rect 26528 30438 26580 30490
rect 34713 30438 34765 30490
rect 34777 30438 34829 30490
rect 34841 30438 34893 30490
rect 34905 30438 34957 30490
rect 34969 30438 35021 30490
rect 25044 30336 25096 30388
rect 18788 30268 18840 30320
rect 14280 30243 14332 30252
rect 14280 30209 14289 30243
rect 14289 30209 14323 30243
rect 14323 30209 14332 30243
rect 14280 30200 14332 30209
rect 14924 30243 14976 30252
rect 14924 30209 14933 30243
rect 14933 30209 14967 30243
rect 14967 30209 14976 30243
rect 14924 30200 14976 30209
rect 21548 30268 21600 30320
rect 20260 30200 20312 30252
rect 21272 30200 21324 30252
rect 24676 30243 24728 30252
rect 24676 30209 24685 30243
rect 24685 30209 24719 30243
rect 24719 30209 24728 30243
rect 24676 30200 24728 30209
rect 25320 30243 25372 30252
rect 25320 30209 25329 30243
rect 25329 30209 25363 30243
rect 25363 30209 25372 30243
rect 25320 30200 25372 30209
rect 25596 30200 25648 30252
rect 25412 30132 25464 30184
rect 25780 30200 25832 30252
rect 26056 30243 26108 30252
rect 26056 30209 26065 30243
rect 26065 30209 26099 30243
rect 26099 30209 26108 30243
rect 26056 30200 26108 30209
rect 27160 30336 27212 30388
rect 27344 30336 27396 30388
rect 28448 30336 28500 30388
rect 28080 30268 28132 30320
rect 27528 30200 27580 30252
rect 27896 30175 27948 30184
rect 27896 30141 27905 30175
rect 27905 30141 27939 30175
rect 27939 30141 27948 30175
rect 28908 30200 28960 30252
rect 27896 30132 27948 30141
rect 29092 30132 29144 30184
rect 28448 30064 28500 30116
rect 28540 30064 28592 30116
rect 29920 30243 29972 30252
rect 29920 30209 29929 30243
rect 29929 30209 29963 30243
rect 29963 30209 29972 30243
rect 29920 30200 29972 30209
rect 12900 29996 12952 30048
rect 20720 29996 20772 30048
rect 27528 29996 27580 30048
rect 5170 29894 5222 29946
rect 5234 29894 5286 29946
rect 5298 29894 5350 29946
rect 5362 29894 5414 29946
rect 5426 29894 5478 29946
rect 13611 29894 13663 29946
rect 13675 29894 13727 29946
rect 13739 29894 13791 29946
rect 13803 29894 13855 29946
rect 13867 29894 13919 29946
rect 22052 29894 22104 29946
rect 22116 29894 22168 29946
rect 22180 29894 22232 29946
rect 22244 29894 22296 29946
rect 22308 29894 22360 29946
rect 30493 29894 30545 29946
rect 30557 29894 30609 29946
rect 30621 29894 30673 29946
rect 30685 29894 30737 29946
rect 30749 29894 30801 29946
rect 10508 29792 10560 29844
rect 14832 29835 14884 29844
rect 14832 29801 14841 29835
rect 14841 29801 14875 29835
rect 14875 29801 14884 29835
rect 14832 29792 14884 29801
rect 26056 29792 26108 29844
rect 27436 29792 27488 29844
rect 29920 29792 29972 29844
rect 9956 29656 10008 29708
rect 12624 29656 12676 29708
rect 13084 29656 13136 29708
rect 10508 29588 10560 29640
rect 12900 29588 12952 29640
rect 10968 29520 11020 29572
rect 15016 29588 15068 29640
rect 19248 29588 19300 29640
rect 20536 29656 20588 29708
rect 21548 29699 21600 29708
rect 21548 29665 21557 29699
rect 21557 29665 21591 29699
rect 21591 29665 21600 29699
rect 21548 29656 21600 29665
rect 23296 29724 23348 29776
rect 27436 29656 27488 29708
rect 20168 29631 20220 29640
rect 20168 29597 20177 29631
rect 20177 29597 20211 29631
rect 20211 29597 20220 29631
rect 20168 29588 20220 29597
rect 20812 29588 20864 29640
rect 21272 29588 21324 29640
rect 21640 29588 21692 29640
rect 24768 29631 24820 29640
rect 24768 29597 24777 29631
rect 24777 29597 24811 29631
rect 24811 29597 24820 29631
rect 24768 29588 24820 29597
rect 27896 29724 27948 29776
rect 28080 29656 28132 29708
rect 27712 29631 27764 29640
rect 14280 29520 14332 29572
rect 15108 29563 15160 29572
rect 15108 29529 15117 29563
rect 15117 29529 15151 29563
rect 15151 29529 15160 29563
rect 15108 29520 15160 29529
rect 24584 29520 24636 29572
rect 27712 29597 27721 29631
rect 27721 29597 27755 29631
rect 27755 29597 27764 29631
rect 27712 29588 27764 29597
rect 28632 29656 28684 29708
rect 28264 29588 28316 29640
rect 25412 29520 25464 29572
rect 26056 29520 26108 29572
rect 28816 29588 28868 29640
rect 9312 29452 9364 29504
rect 10324 29495 10376 29504
rect 10324 29461 10333 29495
rect 10333 29461 10367 29495
rect 10367 29461 10376 29495
rect 10324 29452 10376 29461
rect 12808 29495 12860 29504
rect 12808 29461 12817 29495
rect 12817 29461 12851 29495
rect 12851 29461 12860 29495
rect 12808 29452 12860 29461
rect 19432 29452 19484 29504
rect 21456 29452 21508 29504
rect 29092 29452 29144 29504
rect 9390 29350 9442 29402
rect 9454 29350 9506 29402
rect 9518 29350 9570 29402
rect 9582 29350 9634 29402
rect 9646 29350 9698 29402
rect 17831 29350 17883 29402
rect 17895 29350 17947 29402
rect 17959 29350 18011 29402
rect 18023 29350 18075 29402
rect 18087 29350 18139 29402
rect 26272 29350 26324 29402
rect 26336 29350 26388 29402
rect 26400 29350 26452 29402
rect 26464 29350 26516 29402
rect 26528 29350 26580 29402
rect 34713 29350 34765 29402
rect 34777 29350 34829 29402
rect 34841 29350 34893 29402
rect 34905 29350 34957 29402
rect 34969 29350 35021 29402
rect 9312 29155 9364 29164
rect 9312 29121 9321 29155
rect 9321 29121 9355 29155
rect 9355 29121 9364 29155
rect 9312 29112 9364 29121
rect 12900 29248 12952 29300
rect 14556 29291 14608 29300
rect 14556 29257 14565 29291
rect 14565 29257 14599 29291
rect 14599 29257 14608 29291
rect 14556 29248 14608 29257
rect 14924 29248 14976 29300
rect 20260 29291 20312 29300
rect 11060 29112 11112 29164
rect 11796 29155 11848 29164
rect 11796 29121 11805 29155
rect 11805 29121 11839 29155
rect 11839 29121 11848 29155
rect 11796 29112 11848 29121
rect 15108 29180 15160 29232
rect 20260 29257 20269 29291
rect 20269 29257 20303 29291
rect 20303 29257 20312 29291
rect 20260 29248 20312 29257
rect 21732 29248 21784 29300
rect 12624 29155 12676 29164
rect 12624 29121 12633 29155
rect 12633 29121 12667 29155
rect 12667 29121 12676 29155
rect 12624 29112 12676 29121
rect 12808 29112 12860 29164
rect 13360 29112 13412 29164
rect 15568 29155 15620 29164
rect 15568 29121 15577 29155
rect 15577 29121 15611 29155
rect 15611 29121 15620 29155
rect 15568 29112 15620 29121
rect 15752 29155 15804 29164
rect 15752 29121 15761 29155
rect 15761 29121 15795 29155
rect 15795 29121 15804 29155
rect 15752 29112 15804 29121
rect 19340 29180 19392 29232
rect 19432 29155 19484 29164
rect 19432 29121 19441 29155
rect 19441 29121 19475 29155
rect 19475 29121 19484 29155
rect 19432 29112 19484 29121
rect 20444 29155 20496 29164
rect 20444 29121 20453 29155
rect 20453 29121 20487 29155
rect 20487 29121 20496 29155
rect 20444 29112 20496 29121
rect 20720 29155 20772 29164
rect 10324 29044 10376 29096
rect 15016 29044 15068 29096
rect 20168 29044 20220 29096
rect 20720 29121 20729 29155
rect 20729 29121 20763 29155
rect 20763 29121 20772 29155
rect 20720 29112 20772 29121
rect 20812 29155 20864 29164
rect 20812 29121 20821 29155
rect 20821 29121 20855 29155
rect 20855 29121 20864 29155
rect 21640 29180 21692 29232
rect 20812 29112 20864 29121
rect 22284 29155 22336 29164
rect 22284 29121 22293 29155
rect 22293 29121 22327 29155
rect 22327 29121 22336 29155
rect 22284 29112 22336 29121
rect 23480 29180 23532 29232
rect 24676 29180 24728 29232
rect 25320 29248 25372 29300
rect 27528 29291 27580 29300
rect 27528 29257 27537 29291
rect 27537 29257 27571 29291
rect 27571 29257 27580 29291
rect 27528 29248 27580 29257
rect 27620 29248 27672 29300
rect 28264 29291 28316 29300
rect 28264 29257 28289 29291
rect 28289 29257 28316 29291
rect 28264 29248 28316 29257
rect 28908 29248 28960 29300
rect 27988 29180 28040 29232
rect 28080 29223 28132 29232
rect 28080 29189 28089 29223
rect 28089 29189 28123 29223
rect 28123 29189 28132 29223
rect 28080 29180 28132 29189
rect 22744 29155 22796 29164
rect 22744 29121 22753 29155
rect 22753 29121 22787 29155
rect 22787 29121 22796 29155
rect 22744 29112 22796 29121
rect 23572 29112 23624 29164
rect 25780 29112 25832 29164
rect 27436 29155 27488 29164
rect 27436 29121 27445 29155
rect 27445 29121 27479 29155
rect 27479 29121 27488 29155
rect 27436 29112 27488 29121
rect 28908 29155 28960 29164
rect 21640 29044 21692 29096
rect 21456 28976 21508 29028
rect 23296 28976 23348 29028
rect 27896 28976 27948 29028
rect 28908 29121 28917 29155
rect 28917 29121 28951 29155
rect 28951 29121 28960 29155
rect 28908 29112 28960 29121
rect 29092 29155 29144 29164
rect 29092 29121 29101 29155
rect 29101 29121 29135 29155
rect 29135 29121 29144 29155
rect 29092 29112 29144 29121
rect 28632 29044 28684 29096
rect 30288 28976 30340 29028
rect 7748 28908 7800 28960
rect 9312 28908 9364 28960
rect 10416 28908 10468 28960
rect 27528 28908 27580 28960
rect 28816 28908 28868 28960
rect 5170 28806 5222 28858
rect 5234 28806 5286 28858
rect 5298 28806 5350 28858
rect 5362 28806 5414 28858
rect 5426 28806 5478 28858
rect 13611 28806 13663 28858
rect 13675 28806 13727 28858
rect 13739 28806 13791 28858
rect 13803 28806 13855 28858
rect 13867 28806 13919 28858
rect 22052 28806 22104 28858
rect 22116 28806 22168 28858
rect 22180 28806 22232 28858
rect 22244 28806 22296 28858
rect 22308 28806 22360 28858
rect 30493 28806 30545 28858
rect 30557 28806 30609 28858
rect 30621 28806 30673 28858
rect 30685 28806 30737 28858
rect 30749 28806 30801 28858
rect 13360 28704 13412 28756
rect 21088 28747 21140 28756
rect 11060 28636 11112 28688
rect 21088 28713 21097 28747
rect 21097 28713 21131 28747
rect 21131 28713 21140 28747
rect 21088 28704 21140 28713
rect 28816 28704 28868 28756
rect 11796 28568 11848 28620
rect 12532 28568 12584 28620
rect 13360 28611 13412 28620
rect 13360 28577 13369 28611
rect 13369 28577 13403 28611
rect 13403 28577 13412 28611
rect 13360 28568 13412 28577
rect 15016 28568 15068 28620
rect 15936 28568 15988 28620
rect 20812 28636 20864 28688
rect 21640 28636 21692 28688
rect 7748 28500 7800 28552
rect 9036 28500 9088 28552
rect 9312 28543 9364 28552
rect 9312 28509 9321 28543
rect 9321 28509 9355 28543
rect 9355 28509 9364 28543
rect 9312 28500 9364 28509
rect 10968 28500 11020 28552
rect 12808 28500 12860 28552
rect 12992 28500 13044 28552
rect 13268 28543 13320 28552
rect 13268 28509 13277 28543
rect 13277 28509 13311 28543
rect 13311 28509 13320 28543
rect 14556 28543 14608 28552
rect 13268 28500 13320 28509
rect 14556 28509 14565 28543
rect 14565 28509 14599 28543
rect 14599 28509 14608 28543
rect 14556 28500 14608 28509
rect 15108 28500 15160 28552
rect 15384 28543 15436 28552
rect 15384 28509 15393 28543
rect 15393 28509 15427 28543
rect 15427 28509 15436 28543
rect 15384 28500 15436 28509
rect 15476 28500 15528 28552
rect 19708 28543 19760 28552
rect 19708 28509 19717 28543
rect 19717 28509 19751 28543
rect 19751 28509 19760 28543
rect 19708 28500 19760 28509
rect 19892 28543 19944 28552
rect 19892 28509 19901 28543
rect 19901 28509 19935 28543
rect 19935 28509 19944 28543
rect 19892 28500 19944 28509
rect 21272 28568 21324 28620
rect 27160 28568 27212 28620
rect 27620 28568 27672 28620
rect 13360 28432 13412 28484
rect 15752 28432 15804 28484
rect 19248 28432 19300 28484
rect 22836 28543 22888 28552
rect 22836 28509 22845 28543
rect 22845 28509 22879 28543
rect 22879 28509 22888 28543
rect 22836 28500 22888 28509
rect 23296 28500 23348 28552
rect 23480 28500 23532 28552
rect 27896 28500 27948 28552
rect 29000 28543 29052 28552
rect 29000 28509 29009 28543
rect 29009 28509 29043 28543
rect 29043 28509 29052 28543
rect 29000 28500 29052 28509
rect 20720 28432 20772 28484
rect 21548 28432 21600 28484
rect 9220 28407 9272 28416
rect 9220 28373 9229 28407
rect 9229 28373 9263 28407
rect 9263 28373 9272 28407
rect 9220 28364 9272 28373
rect 12900 28407 12952 28416
rect 12900 28373 12909 28407
rect 12909 28373 12943 28407
rect 12943 28373 12952 28407
rect 12900 28364 12952 28373
rect 20536 28364 20588 28416
rect 22744 28364 22796 28416
rect 27252 28407 27304 28416
rect 27252 28373 27261 28407
rect 27261 28373 27295 28407
rect 27295 28373 27304 28407
rect 27252 28364 27304 28373
rect 9390 28262 9442 28314
rect 9454 28262 9506 28314
rect 9518 28262 9570 28314
rect 9582 28262 9634 28314
rect 9646 28262 9698 28314
rect 17831 28262 17883 28314
rect 17895 28262 17947 28314
rect 17959 28262 18011 28314
rect 18023 28262 18075 28314
rect 18087 28262 18139 28314
rect 26272 28262 26324 28314
rect 26336 28262 26388 28314
rect 26400 28262 26452 28314
rect 26464 28262 26516 28314
rect 26528 28262 26580 28314
rect 34713 28262 34765 28314
rect 34777 28262 34829 28314
rect 34841 28262 34893 28314
rect 34905 28262 34957 28314
rect 34969 28262 35021 28314
rect 7748 28067 7800 28076
rect 7748 28033 7757 28067
rect 7757 28033 7791 28067
rect 7791 28033 7800 28067
rect 7748 28024 7800 28033
rect 8760 28067 8812 28076
rect 8760 28033 8769 28067
rect 8769 28033 8803 28067
rect 8803 28033 8812 28067
rect 8760 28024 8812 28033
rect 9864 28160 9916 28212
rect 10968 28092 11020 28144
rect 12992 28160 13044 28212
rect 13360 28160 13412 28212
rect 15384 28203 15436 28212
rect 15384 28169 15393 28203
rect 15393 28169 15427 28203
rect 15427 28169 15436 28203
rect 15384 28160 15436 28169
rect 22376 28203 22428 28212
rect 22376 28169 22385 28203
rect 22385 28169 22419 28203
rect 22419 28169 22428 28203
rect 22376 28160 22428 28169
rect 9036 28067 9088 28076
rect 9036 28033 9045 28067
rect 9045 28033 9079 28067
rect 9079 28033 9088 28067
rect 9036 28024 9088 28033
rect 12532 28067 12584 28076
rect 12532 28033 12541 28067
rect 12541 28033 12575 28067
rect 12575 28033 12584 28067
rect 12532 28024 12584 28033
rect 15016 28092 15068 28144
rect 15568 28092 15620 28144
rect 16028 28092 16080 28144
rect 19892 28092 19944 28144
rect 13268 28024 13320 28076
rect 14004 28067 14056 28076
rect 14004 28033 14013 28067
rect 14013 28033 14047 28067
rect 14047 28033 14056 28067
rect 14004 28024 14056 28033
rect 14280 28024 14332 28076
rect 15476 28024 15528 28076
rect 19248 28067 19300 28076
rect 19248 28033 19257 28067
rect 19257 28033 19291 28067
rect 19291 28033 19300 28067
rect 19248 28024 19300 28033
rect 20720 28092 20772 28144
rect 22836 28135 22888 28144
rect 22836 28101 22845 28135
rect 22845 28101 22879 28135
rect 22879 28101 22888 28135
rect 22836 28092 22888 28101
rect 9312 27956 9364 28008
rect 12440 27999 12492 28008
rect 12440 27965 12449 27999
rect 12449 27965 12483 27999
rect 12483 27965 12492 27999
rect 12440 27956 12492 27965
rect 14556 27956 14608 28008
rect 19340 27956 19392 28008
rect 24676 28024 24728 28076
rect 25044 28067 25096 28076
rect 25044 28033 25053 28067
rect 25053 28033 25087 28067
rect 25087 28033 25096 28067
rect 25044 28024 25096 28033
rect 25228 28024 25280 28076
rect 27068 28024 27120 28076
rect 27712 28024 27764 28076
rect 29276 28024 29328 28076
rect 30288 28067 30340 28076
rect 30288 28033 30297 28067
rect 30297 28033 30331 28067
rect 30331 28033 30340 28067
rect 30288 28024 30340 28033
rect 32312 28024 32364 28076
rect 25136 27956 25188 28008
rect 25780 27999 25832 28008
rect 25780 27965 25789 27999
rect 25789 27965 25823 27999
rect 25823 27965 25832 27999
rect 25780 27956 25832 27965
rect 26240 27956 26292 28008
rect 12992 27888 13044 27940
rect 15384 27888 15436 27940
rect 23480 27888 23532 27940
rect 25872 27888 25924 27940
rect 9128 27820 9180 27872
rect 9312 27820 9364 27872
rect 9588 27820 9640 27872
rect 19708 27820 19760 27872
rect 26608 27820 26660 27872
rect 30012 27820 30064 27872
rect 5170 27718 5222 27770
rect 5234 27718 5286 27770
rect 5298 27718 5350 27770
rect 5362 27718 5414 27770
rect 5426 27718 5478 27770
rect 13611 27718 13663 27770
rect 13675 27718 13727 27770
rect 13739 27718 13791 27770
rect 13803 27718 13855 27770
rect 13867 27718 13919 27770
rect 22052 27718 22104 27770
rect 22116 27718 22168 27770
rect 22180 27718 22232 27770
rect 22244 27718 22296 27770
rect 22308 27718 22360 27770
rect 30493 27718 30545 27770
rect 30557 27718 30609 27770
rect 30621 27718 30673 27770
rect 30685 27718 30737 27770
rect 30749 27718 30801 27770
rect 16028 27548 16080 27600
rect 24584 27548 24636 27600
rect 27896 27591 27948 27600
rect 27896 27557 27905 27591
rect 27905 27557 27939 27591
rect 27939 27557 27948 27591
rect 27896 27548 27948 27557
rect 12532 27480 12584 27532
rect 13084 27480 13136 27532
rect 9128 27412 9180 27464
rect 9588 27412 9640 27464
rect 9772 27344 9824 27396
rect 8208 27276 8260 27328
rect 12348 27344 12400 27396
rect 13820 27412 13872 27464
rect 14004 27344 14056 27396
rect 15844 27412 15896 27464
rect 16028 27455 16080 27464
rect 16028 27421 16037 27455
rect 16037 27421 16071 27455
rect 16071 27421 16080 27455
rect 16028 27412 16080 27421
rect 18236 27455 18288 27464
rect 18236 27421 18245 27455
rect 18245 27421 18279 27455
rect 18279 27421 18288 27455
rect 18236 27412 18288 27421
rect 19248 27344 19300 27396
rect 20996 27344 21048 27396
rect 25872 27480 25924 27532
rect 23572 27412 23624 27464
rect 25688 27455 25740 27464
rect 25044 27344 25096 27396
rect 19800 27276 19852 27328
rect 25688 27421 25697 27455
rect 25697 27421 25731 27455
rect 25731 27421 25740 27455
rect 25688 27412 25740 27421
rect 25596 27344 25648 27396
rect 26148 27412 26200 27464
rect 27712 27455 27764 27464
rect 26240 27344 26292 27396
rect 27712 27421 27721 27455
rect 27721 27421 27755 27455
rect 27755 27421 27764 27455
rect 27712 27412 27764 27421
rect 27988 27412 28040 27464
rect 29000 27412 29052 27464
rect 29736 27455 29788 27464
rect 25780 27276 25832 27328
rect 26700 27276 26752 27328
rect 27068 27276 27120 27328
rect 29736 27421 29745 27455
rect 29745 27421 29779 27455
rect 29779 27421 29788 27455
rect 29736 27412 29788 27421
rect 29184 27344 29236 27396
rect 9390 27174 9442 27226
rect 9454 27174 9506 27226
rect 9518 27174 9570 27226
rect 9582 27174 9634 27226
rect 9646 27174 9698 27226
rect 17831 27174 17883 27226
rect 17895 27174 17947 27226
rect 17959 27174 18011 27226
rect 18023 27174 18075 27226
rect 18087 27174 18139 27226
rect 26272 27174 26324 27226
rect 26336 27174 26388 27226
rect 26400 27174 26452 27226
rect 26464 27174 26516 27226
rect 26528 27174 26580 27226
rect 34713 27174 34765 27226
rect 34777 27174 34829 27226
rect 34841 27174 34893 27226
rect 34905 27174 34957 27226
rect 34969 27174 35021 27226
rect 8760 27004 8812 27056
rect 8208 26979 8260 26988
rect 8208 26945 8217 26979
rect 8217 26945 8251 26979
rect 8251 26945 8260 26979
rect 8208 26936 8260 26945
rect 9220 26979 9272 26988
rect 9220 26945 9229 26979
rect 9229 26945 9263 26979
rect 9263 26945 9272 26979
rect 9220 26936 9272 26945
rect 12900 27072 12952 27124
rect 18236 27072 18288 27124
rect 20996 27072 21048 27124
rect 30288 27072 30340 27124
rect 13084 27004 13136 27056
rect 13820 27004 13872 27056
rect 14280 27004 14332 27056
rect 19800 27004 19852 27056
rect 12440 26936 12492 26988
rect 15660 26979 15712 26988
rect 15660 26945 15669 26979
rect 15669 26945 15703 26979
rect 15703 26945 15712 26979
rect 15660 26936 15712 26945
rect 15752 26979 15804 26988
rect 15752 26945 15761 26979
rect 15761 26945 15795 26979
rect 15795 26945 15804 26979
rect 15752 26936 15804 26945
rect 18328 26936 18380 26988
rect 20996 26979 21048 26988
rect 10692 26868 10744 26920
rect 12624 26868 12676 26920
rect 20536 26868 20588 26920
rect 20996 26945 21005 26979
rect 21005 26945 21039 26979
rect 21039 26945 21048 26979
rect 20996 26936 21048 26945
rect 24768 26936 24820 26988
rect 25136 26979 25188 26988
rect 25136 26945 25145 26979
rect 25145 26945 25179 26979
rect 25179 26945 25188 26979
rect 25136 26936 25188 26945
rect 25596 26979 25648 26988
rect 25596 26945 25605 26979
rect 25605 26945 25639 26979
rect 25639 26945 25648 26979
rect 25596 26936 25648 26945
rect 26148 27004 26200 27056
rect 25872 26979 25924 26988
rect 25872 26945 25881 26979
rect 25881 26945 25915 26979
rect 25915 26945 25924 26979
rect 25872 26936 25924 26945
rect 27252 26979 27304 26988
rect 27252 26945 27261 26979
rect 27261 26945 27295 26979
rect 27295 26945 27304 26979
rect 27252 26936 27304 26945
rect 27344 26979 27396 26988
rect 27344 26945 27353 26979
rect 27353 26945 27387 26979
rect 27387 26945 27396 26979
rect 30012 26979 30064 26988
rect 27344 26936 27396 26945
rect 30012 26945 30021 26979
rect 30021 26945 30055 26979
rect 30055 26945 30064 26979
rect 30012 26936 30064 26945
rect 22652 26911 22704 26920
rect 22652 26877 22661 26911
rect 22661 26877 22695 26911
rect 22695 26877 22704 26911
rect 22652 26868 22704 26877
rect 26148 26868 26200 26920
rect 27620 26868 27672 26920
rect 29736 26911 29788 26920
rect 29736 26877 29745 26911
rect 29745 26877 29779 26911
rect 29779 26877 29788 26911
rect 29736 26868 29788 26877
rect 29920 26868 29972 26920
rect 21548 26800 21600 26852
rect 9220 26732 9272 26784
rect 11152 26732 11204 26784
rect 22376 26732 22428 26784
rect 24584 26732 24636 26784
rect 27160 26732 27212 26784
rect 5170 26630 5222 26682
rect 5234 26630 5286 26682
rect 5298 26630 5350 26682
rect 5362 26630 5414 26682
rect 5426 26630 5478 26682
rect 13611 26630 13663 26682
rect 13675 26630 13727 26682
rect 13739 26630 13791 26682
rect 13803 26630 13855 26682
rect 13867 26630 13919 26682
rect 22052 26630 22104 26682
rect 22116 26630 22168 26682
rect 22180 26630 22232 26682
rect 22244 26630 22296 26682
rect 22308 26630 22360 26682
rect 30493 26630 30545 26682
rect 30557 26630 30609 26682
rect 30621 26630 30673 26682
rect 30685 26630 30737 26682
rect 30749 26630 30801 26682
rect 12440 26528 12492 26580
rect 12900 26528 12952 26580
rect 13360 26528 13412 26580
rect 25136 26528 25188 26580
rect 9312 26460 9364 26512
rect 25964 26528 26016 26580
rect 26608 26528 26660 26580
rect 26792 26528 26844 26580
rect 27068 26571 27120 26580
rect 27068 26537 27077 26571
rect 27077 26537 27111 26571
rect 27111 26537 27120 26571
rect 27068 26528 27120 26537
rect 29184 26571 29236 26580
rect 29184 26537 29193 26571
rect 29193 26537 29227 26571
rect 29227 26537 29236 26571
rect 29184 26528 29236 26537
rect 11152 26435 11204 26444
rect 11152 26401 11161 26435
rect 11161 26401 11195 26435
rect 11195 26401 11204 26435
rect 11152 26392 11204 26401
rect 27528 26460 27580 26512
rect 28632 26460 28684 26512
rect 12808 26392 12860 26444
rect 18236 26392 18288 26444
rect 12624 26367 12676 26376
rect 12624 26333 12633 26367
rect 12633 26333 12667 26367
rect 12667 26333 12676 26367
rect 12624 26324 12676 26333
rect 13084 26324 13136 26376
rect 9772 26256 9824 26308
rect 12532 26256 12584 26308
rect 13452 26299 13504 26308
rect 13452 26265 13463 26299
rect 13463 26265 13504 26299
rect 15844 26324 15896 26376
rect 17224 26324 17276 26376
rect 20996 26392 21048 26444
rect 21640 26392 21692 26444
rect 22744 26392 22796 26444
rect 21548 26324 21600 26376
rect 25044 26324 25096 26376
rect 25320 26324 25372 26376
rect 25504 26367 25556 26376
rect 25504 26333 25513 26367
rect 25513 26333 25547 26367
rect 25547 26333 25556 26367
rect 25504 26324 25556 26333
rect 25872 26367 25924 26376
rect 25872 26333 25881 26367
rect 25881 26333 25915 26367
rect 25915 26333 25924 26367
rect 25872 26324 25924 26333
rect 26516 26367 26568 26376
rect 26516 26333 26525 26367
rect 26525 26333 26559 26367
rect 26559 26333 26568 26367
rect 26516 26324 26568 26333
rect 13452 26256 13504 26265
rect 18420 26299 18472 26308
rect 18420 26265 18429 26299
rect 18429 26265 18463 26299
rect 18463 26265 18472 26299
rect 18420 26256 18472 26265
rect 19340 26256 19392 26308
rect 22560 26299 22612 26308
rect 22560 26265 22569 26299
rect 22569 26265 22603 26299
rect 22603 26265 22612 26299
rect 22560 26256 22612 26265
rect 22652 26256 22704 26308
rect 25136 26256 25188 26308
rect 26884 26367 26936 26376
rect 26884 26333 26893 26367
rect 26893 26333 26927 26367
rect 26927 26333 26936 26367
rect 26884 26324 26936 26333
rect 27160 26324 27212 26376
rect 28724 26367 28776 26376
rect 28724 26333 28733 26367
rect 28733 26333 28767 26367
rect 28767 26333 28776 26367
rect 28724 26324 28776 26333
rect 28908 26324 28960 26376
rect 27620 26256 27672 26308
rect 9312 26188 9364 26240
rect 15660 26188 15712 26240
rect 21180 26188 21232 26240
rect 26792 26188 26844 26240
rect 29092 26256 29144 26308
rect 29000 26188 29052 26240
rect 9390 26086 9442 26138
rect 9454 26086 9506 26138
rect 9518 26086 9570 26138
rect 9582 26086 9634 26138
rect 9646 26086 9698 26138
rect 17831 26086 17883 26138
rect 17895 26086 17947 26138
rect 17959 26086 18011 26138
rect 18023 26086 18075 26138
rect 18087 26086 18139 26138
rect 26272 26086 26324 26138
rect 26336 26086 26388 26138
rect 26400 26086 26452 26138
rect 26464 26086 26516 26138
rect 26528 26086 26580 26138
rect 34713 26086 34765 26138
rect 34777 26086 34829 26138
rect 34841 26086 34893 26138
rect 34905 26086 34957 26138
rect 34969 26086 35021 26138
rect 9772 25984 9824 26036
rect 12532 25984 12584 26036
rect 9312 25916 9364 25968
rect 12440 25959 12492 25968
rect 12440 25925 12449 25959
rect 12449 25925 12483 25959
rect 12483 25925 12492 25959
rect 12440 25916 12492 25925
rect 9772 25891 9824 25900
rect 9772 25857 9781 25891
rect 9781 25857 9815 25891
rect 9815 25857 9824 25891
rect 9772 25848 9824 25857
rect 10416 25891 10468 25900
rect 10416 25857 10425 25891
rect 10425 25857 10459 25891
rect 10459 25857 10468 25891
rect 10416 25848 10468 25857
rect 12256 25848 12308 25900
rect 12348 25891 12400 25900
rect 12348 25857 12357 25891
rect 12357 25857 12391 25891
rect 12391 25857 12400 25891
rect 14740 25984 14792 26036
rect 22652 25984 22704 26036
rect 23572 26027 23624 26036
rect 23572 25993 23581 26027
rect 23581 25993 23615 26027
rect 23615 25993 23624 26027
rect 23572 25984 23624 25993
rect 25688 25984 25740 26036
rect 27252 25984 27304 26036
rect 29920 26027 29972 26036
rect 29920 25993 29929 26027
rect 29929 25993 29963 26027
rect 29963 25993 29972 26027
rect 29920 25984 29972 25993
rect 13360 25959 13412 25968
rect 13360 25925 13369 25959
rect 13369 25925 13403 25959
rect 13403 25925 13412 25959
rect 13360 25916 13412 25925
rect 19248 25916 19300 25968
rect 20996 25916 21048 25968
rect 12348 25848 12400 25857
rect 9220 25780 9272 25832
rect 13452 25891 13504 25900
rect 13452 25857 13466 25891
rect 13466 25857 13500 25891
rect 13500 25857 13504 25891
rect 16948 25891 17000 25900
rect 13452 25848 13504 25857
rect 16948 25857 16957 25891
rect 16957 25857 16991 25891
rect 16991 25857 17000 25891
rect 16948 25848 17000 25857
rect 19616 25891 19668 25900
rect 19616 25857 19625 25891
rect 19625 25857 19659 25891
rect 19659 25857 19668 25891
rect 19616 25848 19668 25857
rect 25504 25916 25556 25968
rect 28632 25959 28684 25968
rect 28632 25925 28641 25959
rect 28641 25925 28675 25959
rect 28675 25925 28684 25959
rect 28632 25916 28684 25925
rect 21548 25848 21600 25900
rect 22376 25848 22428 25900
rect 24676 25891 24728 25900
rect 23664 25780 23716 25832
rect 24676 25857 24685 25891
rect 24685 25857 24719 25891
rect 24719 25857 24728 25891
rect 24676 25848 24728 25857
rect 25872 25848 25924 25900
rect 26516 25891 26568 25900
rect 26516 25857 26525 25891
rect 26525 25857 26559 25891
rect 26559 25857 26568 25891
rect 26516 25848 26568 25857
rect 27620 25891 27672 25900
rect 27620 25857 27629 25891
rect 27629 25857 27663 25891
rect 27663 25857 27672 25891
rect 27620 25848 27672 25857
rect 32312 25891 32364 25900
rect 32312 25857 32321 25891
rect 32321 25857 32355 25891
rect 32355 25857 32364 25891
rect 32312 25848 32364 25857
rect 32404 25891 32456 25900
rect 32404 25857 32413 25891
rect 32413 25857 32447 25891
rect 32447 25857 32456 25891
rect 32404 25848 32456 25857
rect 26056 25780 26108 25832
rect 26700 25780 26752 25832
rect 27068 25780 27120 25832
rect 10416 25712 10468 25764
rect 14464 25712 14516 25764
rect 21180 25712 21232 25764
rect 24860 25712 24912 25764
rect 26884 25712 26936 25764
rect 27528 25823 27580 25832
rect 27528 25789 27537 25823
rect 27537 25789 27571 25823
rect 27571 25789 27580 25823
rect 27528 25780 27580 25789
rect 32496 25780 32548 25832
rect 12716 25644 12768 25696
rect 13084 25687 13136 25696
rect 13084 25653 13093 25687
rect 13093 25653 13127 25687
rect 13127 25653 13136 25687
rect 13084 25644 13136 25653
rect 17224 25687 17276 25696
rect 17224 25653 17233 25687
rect 17233 25653 17267 25687
rect 17267 25653 17276 25687
rect 17224 25644 17276 25653
rect 18328 25687 18380 25696
rect 18328 25653 18337 25687
rect 18337 25653 18371 25687
rect 18371 25653 18380 25687
rect 18328 25644 18380 25653
rect 20904 25644 20956 25696
rect 32772 25687 32824 25696
rect 32772 25653 32781 25687
rect 32781 25653 32815 25687
rect 32815 25653 32824 25687
rect 32772 25644 32824 25653
rect 5170 25542 5222 25594
rect 5234 25542 5286 25594
rect 5298 25542 5350 25594
rect 5362 25542 5414 25594
rect 5426 25542 5478 25594
rect 13611 25542 13663 25594
rect 13675 25542 13727 25594
rect 13739 25542 13791 25594
rect 13803 25542 13855 25594
rect 13867 25542 13919 25594
rect 22052 25542 22104 25594
rect 22116 25542 22168 25594
rect 22180 25542 22232 25594
rect 22244 25542 22296 25594
rect 22308 25542 22360 25594
rect 30493 25542 30545 25594
rect 30557 25542 30609 25594
rect 30621 25542 30673 25594
rect 30685 25542 30737 25594
rect 30749 25542 30801 25594
rect 15660 25440 15712 25492
rect 19800 25483 19852 25492
rect 19800 25449 19809 25483
rect 19809 25449 19843 25483
rect 19843 25449 19852 25483
rect 19800 25440 19852 25449
rect 25964 25440 26016 25492
rect 26792 25440 26844 25492
rect 27620 25440 27672 25492
rect 3332 25304 3384 25356
rect 4160 25279 4212 25288
rect 4160 25245 4169 25279
rect 4169 25245 4203 25279
rect 4203 25245 4212 25279
rect 4160 25236 4212 25245
rect 6828 25236 6880 25288
rect 7472 25236 7524 25288
rect 12256 25279 12308 25288
rect 12256 25245 12265 25279
rect 12265 25245 12299 25279
rect 12299 25245 12308 25279
rect 12256 25236 12308 25245
rect 13084 25304 13136 25356
rect 16304 25415 16356 25424
rect 16304 25381 16313 25415
rect 16313 25381 16347 25415
rect 16347 25381 16356 25415
rect 16304 25372 16356 25381
rect 21180 25347 21232 25356
rect 12716 25279 12768 25288
rect 12716 25245 12725 25279
rect 12725 25245 12759 25279
rect 12759 25245 12768 25279
rect 12716 25236 12768 25245
rect 15292 25236 15344 25288
rect 15384 25236 15436 25288
rect 21180 25313 21189 25347
rect 21189 25313 21223 25347
rect 21223 25313 21232 25347
rect 21180 25304 21232 25313
rect 24676 25304 24728 25356
rect 26608 25347 26660 25356
rect 20904 25279 20956 25288
rect 20904 25245 20922 25279
rect 20922 25245 20956 25279
rect 20904 25236 20956 25245
rect 23480 25236 23532 25288
rect 24584 25279 24636 25288
rect 24584 25245 24593 25279
rect 24593 25245 24627 25279
rect 24627 25245 24636 25279
rect 24584 25236 24636 25245
rect 26608 25313 26617 25347
rect 26617 25313 26651 25347
rect 26651 25313 26660 25347
rect 26608 25304 26660 25313
rect 27252 25279 27304 25288
rect 27252 25245 27291 25279
rect 27291 25245 27304 25279
rect 27252 25236 27304 25245
rect 10232 25168 10284 25220
rect 15476 25168 15528 25220
rect 3976 25143 4028 25152
rect 3976 25109 3985 25143
rect 3985 25109 4019 25143
rect 4019 25109 4028 25143
rect 3976 25100 4028 25109
rect 5080 25100 5132 25152
rect 13452 25100 13504 25152
rect 15200 25143 15252 25152
rect 15200 25109 15209 25143
rect 15209 25109 15243 25143
rect 15243 25109 15252 25143
rect 15200 25100 15252 25109
rect 15384 25143 15436 25152
rect 15384 25109 15411 25143
rect 15411 25109 15436 25143
rect 15384 25100 15436 25109
rect 21088 25168 21140 25220
rect 26056 25168 26108 25220
rect 26516 25168 26568 25220
rect 28908 25236 28960 25288
rect 32404 25440 32456 25492
rect 30104 25279 30156 25288
rect 30104 25245 30113 25279
rect 30113 25245 30147 25279
rect 30147 25245 30156 25279
rect 30104 25236 30156 25245
rect 32772 25236 32824 25288
rect 16396 25100 16448 25152
rect 22560 25100 22612 25152
rect 27068 25143 27120 25152
rect 27068 25109 27077 25143
rect 27077 25109 27111 25143
rect 27111 25109 27120 25143
rect 27068 25100 27120 25109
rect 9390 24998 9442 25050
rect 9454 24998 9506 25050
rect 9518 24998 9570 25050
rect 9582 24998 9634 25050
rect 9646 24998 9698 25050
rect 17831 24998 17883 25050
rect 17895 24998 17947 25050
rect 17959 24998 18011 25050
rect 18023 24998 18075 25050
rect 18087 24998 18139 25050
rect 26272 24998 26324 25050
rect 26336 24998 26388 25050
rect 26400 24998 26452 25050
rect 26464 24998 26516 25050
rect 26528 24998 26580 25050
rect 34713 24998 34765 25050
rect 34777 24998 34829 25050
rect 34841 24998 34893 25050
rect 34905 24998 34957 25050
rect 34969 24998 35021 25050
rect 17224 24896 17276 24948
rect 23388 24896 23440 24948
rect 4712 24828 4764 24880
rect 3332 24760 3384 24812
rect 6828 24760 6880 24812
rect 7472 24760 7524 24812
rect 12808 24760 12860 24812
rect 3700 24735 3752 24744
rect 3700 24701 3709 24735
rect 3709 24701 3743 24735
rect 3743 24701 3752 24735
rect 3700 24692 3752 24701
rect 4068 24692 4120 24744
rect 4528 24692 4580 24744
rect 8484 24692 8536 24744
rect 15200 24803 15252 24812
rect 15200 24769 15209 24803
rect 15209 24769 15243 24803
rect 15243 24769 15252 24803
rect 15200 24760 15252 24769
rect 15384 24803 15436 24812
rect 15384 24769 15393 24803
rect 15393 24769 15427 24803
rect 15427 24769 15436 24803
rect 23664 24871 23716 24880
rect 15384 24760 15436 24769
rect 16304 24760 16356 24812
rect 18420 24760 18472 24812
rect 20444 24760 20496 24812
rect 17316 24692 17368 24744
rect 19340 24735 19392 24744
rect 19340 24701 19349 24735
rect 19349 24701 19383 24735
rect 19383 24701 19392 24735
rect 19340 24692 19392 24701
rect 20628 24692 20680 24744
rect 21180 24760 21232 24812
rect 15568 24624 15620 24676
rect 23664 24837 23673 24871
rect 23673 24837 23707 24871
rect 23707 24837 23716 24871
rect 23664 24828 23716 24837
rect 24860 24828 24912 24880
rect 25136 24803 25188 24812
rect 25136 24769 25145 24803
rect 25145 24769 25179 24803
rect 25179 24769 25188 24803
rect 25320 24803 25372 24812
rect 25136 24760 25188 24769
rect 25320 24769 25329 24803
rect 25329 24769 25363 24803
rect 25363 24769 25372 24803
rect 25320 24760 25372 24769
rect 27068 24828 27120 24880
rect 27160 24828 27212 24880
rect 28816 24871 28868 24880
rect 28816 24837 28825 24871
rect 28825 24837 28859 24871
rect 28859 24837 28868 24871
rect 28816 24828 28868 24837
rect 29092 24803 29144 24812
rect 29092 24769 29101 24803
rect 29101 24769 29135 24803
rect 29135 24769 29144 24803
rect 29092 24760 29144 24769
rect 30380 24803 30432 24812
rect 30380 24769 30414 24803
rect 30414 24769 30432 24803
rect 30380 24760 30432 24769
rect 27988 24692 28040 24744
rect 30104 24735 30156 24744
rect 30104 24701 30113 24735
rect 30113 24701 30147 24735
rect 30147 24701 30156 24735
rect 30104 24692 30156 24701
rect 3240 24556 3292 24608
rect 15200 24556 15252 24608
rect 16396 24556 16448 24608
rect 21272 24624 21324 24676
rect 20536 24556 20588 24608
rect 25964 24599 26016 24608
rect 25964 24565 25973 24599
rect 25973 24565 26007 24599
rect 26007 24565 26016 24599
rect 25964 24556 26016 24565
rect 26608 24556 26660 24608
rect 28908 24556 28960 24608
rect 31484 24599 31536 24608
rect 31484 24565 31493 24599
rect 31493 24565 31527 24599
rect 31527 24565 31536 24599
rect 31484 24556 31536 24565
rect 5170 24454 5222 24506
rect 5234 24454 5286 24506
rect 5298 24454 5350 24506
rect 5362 24454 5414 24506
rect 5426 24454 5478 24506
rect 13611 24454 13663 24506
rect 13675 24454 13727 24506
rect 13739 24454 13791 24506
rect 13803 24454 13855 24506
rect 13867 24454 13919 24506
rect 22052 24454 22104 24506
rect 22116 24454 22168 24506
rect 22180 24454 22232 24506
rect 22244 24454 22296 24506
rect 22308 24454 22360 24506
rect 30493 24454 30545 24506
rect 30557 24454 30609 24506
rect 30621 24454 30673 24506
rect 30685 24454 30737 24506
rect 30749 24454 30801 24506
rect 3332 24395 3384 24404
rect 3332 24361 3341 24395
rect 3341 24361 3375 24395
rect 3375 24361 3384 24395
rect 3332 24352 3384 24361
rect 3700 24352 3752 24404
rect 6828 24395 6880 24404
rect 6828 24361 6837 24395
rect 6837 24361 6871 24395
rect 6871 24361 6880 24395
rect 6828 24352 6880 24361
rect 14648 24352 14700 24404
rect 20536 24352 20588 24404
rect 3976 24259 4028 24268
rect 3976 24225 3985 24259
rect 3985 24225 4019 24259
rect 4019 24225 4028 24259
rect 3976 24216 4028 24225
rect 3240 24191 3292 24200
rect 2596 24123 2648 24132
rect 2596 24089 2605 24123
rect 2605 24089 2639 24123
rect 2639 24089 2648 24123
rect 2596 24080 2648 24089
rect 3240 24157 3249 24191
rect 3249 24157 3283 24191
rect 3283 24157 3292 24191
rect 3240 24148 3292 24157
rect 3792 24148 3844 24200
rect 9220 24284 9272 24336
rect 15752 24284 15804 24336
rect 15844 24284 15896 24336
rect 17960 24284 18012 24336
rect 20444 24284 20496 24336
rect 5172 24216 5224 24268
rect 13452 24216 13504 24268
rect 4436 24191 4488 24200
rect 4436 24157 4445 24191
rect 4445 24157 4479 24191
rect 4479 24157 4488 24191
rect 4436 24148 4488 24157
rect 4712 24148 4764 24200
rect 4160 24080 4212 24132
rect 4252 24080 4304 24132
rect 7196 24148 7248 24200
rect 7288 24080 7340 24132
rect 9312 24148 9364 24200
rect 11980 24191 12032 24200
rect 11980 24157 11989 24191
rect 11989 24157 12023 24191
rect 12023 24157 12032 24191
rect 11980 24148 12032 24157
rect 13084 24148 13136 24200
rect 8300 24080 8352 24132
rect 12256 24080 12308 24132
rect 14556 24191 14608 24200
rect 14556 24157 14565 24191
rect 14565 24157 14599 24191
rect 14599 24157 14608 24191
rect 14556 24148 14608 24157
rect 14832 24191 14884 24200
rect 14832 24157 14841 24191
rect 14841 24157 14875 24191
rect 14875 24157 14884 24191
rect 14832 24148 14884 24157
rect 15936 24191 15988 24200
rect 15660 24080 15712 24132
rect 4896 24012 4948 24064
rect 7564 24012 7616 24064
rect 12624 24012 12676 24064
rect 12900 24012 12952 24064
rect 15568 24055 15620 24064
rect 15568 24021 15577 24055
rect 15577 24021 15611 24055
rect 15611 24021 15620 24055
rect 15568 24012 15620 24021
rect 15936 24157 15945 24191
rect 15945 24157 15979 24191
rect 15979 24157 15988 24191
rect 15936 24148 15988 24157
rect 18052 24216 18104 24268
rect 18236 24216 18288 24268
rect 21180 24284 21232 24336
rect 23480 24284 23532 24336
rect 21088 24216 21140 24268
rect 17960 24148 18012 24200
rect 18696 24080 18748 24132
rect 17408 24012 17460 24064
rect 17592 24012 17644 24064
rect 20720 24191 20772 24200
rect 20720 24157 20729 24191
rect 20729 24157 20763 24191
rect 20763 24157 20772 24191
rect 20720 24148 20772 24157
rect 21272 24148 21324 24200
rect 23388 24191 23440 24200
rect 23388 24157 23397 24191
rect 23397 24157 23431 24191
rect 23431 24157 23440 24191
rect 23388 24148 23440 24157
rect 30380 24352 30432 24404
rect 23756 24148 23808 24200
rect 27528 24216 27580 24268
rect 28724 24216 28776 24268
rect 26700 24148 26752 24200
rect 30840 24148 30892 24200
rect 32312 24216 32364 24268
rect 21180 24012 21232 24064
rect 24492 24080 24544 24132
rect 29000 24080 29052 24132
rect 21732 24012 21784 24064
rect 23480 24012 23532 24064
rect 24676 24012 24728 24064
rect 25228 24055 25280 24064
rect 25228 24021 25237 24055
rect 25237 24021 25271 24055
rect 25271 24021 25280 24055
rect 25228 24012 25280 24021
rect 31484 24012 31536 24064
rect 9390 23910 9442 23962
rect 9454 23910 9506 23962
rect 9518 23910 9570 23962
rect 9582 23910 9634 23962
rect 9646 23910 9698 23962
rect 17831 23910 17883 23962
rect 17895 23910 17947 23962
rect 17959 23910 18011 23962
rect 18023 23910 18075 23962
rect 18087 23910 18139 23962
rect 26272 23910 26324 23962
rect 26336 23910 26388 23962
rect 26400 23910 26452 23962
rect 26464 23910 26516 23962
rect 26528 23910 26580 23962
rect 34713 23910 34765 23962
rect 34777 23910 34829 23962
rect 34841 23910 34893 23962
rect 34905 23910 34957 23962
rect 34969 23910 35021 23962
rect 2596 23808 2648 23860
rect 4344 23740 4396 23792
rect 4528 23740 4580 23792
rect 3424 23672 3476 23724
rect 8300 23808 8352 23860
rect 8576 23808 8628 23860
rect 9404 23808 9456 23860
rect 15384 23808 15436 23860
rect 20628 23808 20680 23860
rect 6736 23672 6788 23724
rect 8484 23740 8536 23792
rect 8944 23672 8996 23724
rect 9220 23715 9272 23724
rect 9220 23681 9229 23715
rect 9229 23681 9263 23715
rect 9263 23681 9272 23715
rect 9220 23672 9272 23681
rect 12900 23715 12952 23724
rect 3240 23536 3292 23588
rect 6644 23604 6696 23656
rect 7104 23647 7156 23656
rect 4068 23468 4120 23520
rect 7104 23613 7113 23647
rect 7113 23613 7147 23647
rect 7147 23613 7156 23647
rect 7104 23604 7156 23613
rect 7472 23604 7524 23656
rect 9404 23647 9456 23656
rect 9404 23613 9413 23647
rect 9413 23613 9447 23647
rect 9447 23613 9456 23647
rect 9404 23604 9456 23613
rect 7288 23468 7340 23520
rect 8300 23468 8352 23520
rect 12900 23681 12909 23715
rect 12909 23681 12943 23715
rect 12943 23681 12952 23715
rect 12900 23672 12952 23681
rect 12256 23647 12308 23656
rect 12256 23613 12265 23647
rect 12265 23613 12299 23647
rect 12299 23613 12308 23647
rect 12256 23604 12308 23613
rect 14648 23740 14700 23792
rect 15200 23740 15252 23792
rect 20904 23740 20956 23792
rect 21916 23740 21968 23792
rect 23480 23808 23532 23860
rect 29276 23808 29328 23860
rect 30104 23851 30156 23860
rect 30104 23817 30113 23851
rect 30113 23817 30147 23851
rect 30147 23817 30156 23851
rect 30104 23808 30156 23817
rect 23756 23740 23808 23792
rect 28632 23783 28684 23792
rect 28632 23749 28641 23783
rect 28641 23749 28675 23783
rect 28675 23749 28684 23783
rect 28632 23740 28684 23749
rect 13084 23672 13136 23724
rect 15568 23672 15620 23724
rect 15936 23672 15988 23724
rect 17408 23672 17460 23724
rect 20536 23715 20588 23724
rect 20536 23681 20545 23715
rect 20545 23681 20579 23715
rect 20579 23681 20588 23715
rect 20536 23672 20588 23681
rect 20720 23715 20772 23724
rect 20720 23681 20729 23715
rect 20729 23681 20763 23715
rect 20763 23681 20772 23715
rect 20720 23672 20772 23681
rect 13176 23647 13228 23656
rect 13176 23613 13185 23647
rect 13185 23613 13219 23647
rect 13219 23613 13228 23647
rect 13176 23604 13228 23613
rect 14740 23604 14792 23656
rect 15292 23647 15344 23656
rect 15292 23613 15301 23647
rect 15301 23613 15335 23647
rect 15335 23613 15344 23647
rect 15292 23604 15344 23613
rect 18420 23604 18472 23656
rect 20812 23647 20864 23656
rect 20812 23613 20821 23647
rect 20821 23613 20855 23647
rect 20855 23613 20864 23647
rect 20812 23604 20864 23613
rect 23664 23672 23716 23724
rect 27160 23604 27212 23656
rect 16580 23536 16632 23588
rect 19708 23536 19760 23588
rect 20076 23536 20128 23588
rect 28816 23536 28868 23588
rect 15292 23468 15344 23520
rect 24952 23468 25004 23520
rect 25964 23468 26016 23520
rect 5170 23366 5222 23418
rect 5234 23366 5286 23418
rect 5298 23366 5350 23418
rect 5362 23366 5414 23418
rect 5426 23366 5478 23418
rect 13611 23366 13663 23418
rect 13675 23366 13727 23418
rect 13739 23366 13791 23418
rect 13803 23366 13855 23418
rect 13867 23366 13919 23418
rect 22052 23366 22104 23418
rect 22116 23366 22168 23418
rect 22180 23366 22232 23418
rect 22244 23366 22296 23418
rect 22308 23366 22360 23418
rect 30493 23366 30545 23418
rect 30557 23366 30609 23418
rect 30621 23366 30673 23418
rect 30685 23366 30737 23418
rect 30749 23366 30801 23418
rect 4160 23264 4212 23316
rect 7104 23264 7156 23316
rect 7564 23264 7616 23316
rect 4436 23196 4488 23248
rect 6644 23196 6696 23248
rect 4252 23128 4304 23180
rect 4712 23171 4764 23180
rect 4712 23137 4721 23171
rect 4721 23137 4755 23171
rect 4755 23137 4764 23171
rect 4712 23128 4764 23137
rect 8576 23196 8628 23248
rect 8852 23128 8904 23180
rect 3424 23103 3476 23112
rect 3424 23069 3433 23103
rect 3433 23069 3467 23103
rect 3467 23069 3476 23103
rect 3424 23060 3476 23069
rect 5080 23060 5132 23112
rect 7104 23103 7156 23112
rect 7104 23069 7113 23103
rect 7113 23069 7147 23103
rect 7147 23069 7156 23103
rect 7104 23060 7156 23069
rect 7288 23103 7340 23112
rect 7288 23069 7297 23103
rect 7297 23069 7331 23103
rect 7331 23069 7340 23103
rect 7288 23060 7340 23069
rect 7564 23103 7616 23112
rect 7564 23069 7573 23103
rect 7573 23069 7607 23103
rect 7607 23069 7616 23103
rect 7564 23060 7616 23069
rect 8116 23103 8168 23112
rect 8116 23069 8125 23103
rect 8125 23069 8159 23103
rect 8159 23069 8168 23103
rect 8116 23060 8168 23069
rect 7012 22992 7064 23044
rect 8116 22924 8168 22976
rect 9404 23264 9456 23316
rect 9864 23264 9916 23316
rect 14004 23264 14056 23316
rect 18696 23307 18748 23316
rect 18696 23273 18705 23307
rect 18705 23273 18739 23307
rect 18739 23273 18748 23307
rect 18696 23264 18748 23273
rect 21916 23307 21968 23316
rect 21916 23273 21925 23307
rect 21925 23273 21959 23307
rect 21959 23273 21968 23307
rect 21916 23264 21968 23273
rect 19616 23196 19668 23248
rect 24676 23196 24728 23248
rect 15292 23171 15344 23180
rect 15292 23137 15301 23171
rect 15301 23137 15335 23171
rect 15335 23137 15344 23171
rect 15292 23128 15344 23137
rect 15384 23171 15436 23180
rect 15384 23137 15393 23171
rect 15393 23137 15427 23171
rect 15427 23137 15436 23171
rect 16580 23171 16632 23180
rect 15384 23128 15436 23137
rect 16580 23137 16589 23171
rect 16589 23137 16623 23171
rect 16623 23137 16632 23171
rect 16580 23128 16632 23137
rect 17316 23171 17368 23180
rect 17316 23137 17325 23171
rect 17325 23137 17359 23171
rect 17359 23137 17368 23171
rect 17316 23128 17368 23137
rect 25228 23171 25280 23180
rect 25228 23137 25237 23171
rect 25237 23137 25271 23171
rect 25271 23137 25280 23171
rect 25228 23128 25280 23137
rect 9312 23060 9364 23112
rect 12072 23103 12124 23112
rect 12072 23069 12081 23103
rect 12081 23069 12115 23103
rect 12115 23069 12124 23103
rect 12072 23060 12124 23069
rect 14740 23060 14792 23112
rect 15200 23103 15252 23112
rect 15200 23069 15209 23103
rect 15209 23069 15243 23103
rect 15243 23069 15252 23103
rect 15200 23060 15252 23069
rect 17592 23103 17644 23112
rect 17592 23069 17626 23103
rect 17626 23069 17644 23103
rect 9772 22992 9824 23044
rect 11888 22992 11940 23044
rect 12440 22992 12492 23044
rect 17592 23060 17644 23069
rect 19432 23103 19484 23112
rect 19432 23069 19441 23103
rect 19441 23069 19475 23103
rect 19475 23069 19484 23103
rect 19432 23060 19484 23069
rect 19708 23103 19760 23112
rect 19708 23069 19717 23103
rect 19717 23069 19751 23103
rect 19751 23069 19760 23103
rect 19708 23060 19760 23069
rect 20812 23060 20864 23112
rect 20996 23060 21048 23112
rect 27712 23128 27764 23180
rect 32680 23171 32732 23180
rect 32680 23137 32689 23171
rect 32689 23137 32723 23171
rect 32723 23137 32732 23171
rect 32680 23128 32732 23137
rect 33140 23171 33192 23180
rect 33140 23137 33149 23171
rect 33149 23137 33183 23171
rect 33183 23137 33192 23171
rect 33140 23128 33192 23137
rect 27528 23103 27580 23112
rect 27528 23069 27537 23103
rect 27537 23069 27571 23103
rect 27571 23069 27580 23103
rect 27528 23060 27580 23069
rect 27988 23103 28040 23112
rect 27988 23069 27997 23103
rect 27997 23069 28031 23103
rect 28031 23069 28040 23103
rect 27988 23060 28040 23069
rect 28264 23103 28316 23112
rect 28264 23069 28273 23103
rect 28273 23069 28307 23103
rect 28307 23069 28316 23103
rect 28264 23060 28316 23069
rect 31760 23103 31812 23112
rect 10140 22924 10192 22976
rect 10324 22967 10376 22976
rect 10324 22933 10333 22967
rect 10333 22933 10367 22967
rect 10367 22933 10376 22967
rect 10324 22924 10376 22933
rect 10416 22924 10468 22976
rect 12808 22924 12860 22976
rect 17500 22992 17552 23044
rect 25320 22992 25372 23044
rect 27620 22992 27672 23044
rect 31760 23069 31769 23103
rect 31769 23069 31803 23103
rect 31803 23069 31812 23103
rect 31760 23060 31812 23069
rect 32036 23103 32088 23112
rect 32036 23069 32045 23103
rect 32045 23069 32079 23103
rect 32079 23069 32088 23103
rect 32036 23060 32088 23069
rect 32404 23060 32456 23112
rect 33324 23060 33376 23112
rect 31300 22992 31352 23044
rect 14740 22924 14792 22976
rect 18512 22924 18564 22976
rect 20628 22924 20680 22976
rect 24860 22924 24912 22976
rect 25136 22967 25188 22976
rect 25136 22933 25145 22967
rect 25145 22933 25179 22967
rect 25179 22933 25188 22967
rect 25136 22924 25188 22933
rect 31116 22924 31168 22976
rect 33232 22924 33284 22976
rect 33508 22924 33560 22976
rect 9390 22822 9442 22874
rect 9454 22822 9506 22874
rect 9518 22822 9570 22874
rect 9582 22822 9634 22874
rect 9646 22822 9698 22874
rect 17831 22822 17883 22874
rect 17895 22822 17947 22874
rect 17959 22822 18011 22874
rect 18023 22822 18075 22874
rect 18087 22822 18139 22874
rect 26272 22822 26324 22874
rect 26336 22822 26388 22874
rect 26400 22822 26452 22874
rect 26464 22822 26516 22874
rect 26528 22822 26580 22874
rect 34713 22822 34765 22874
rect 34777 22822 34829 22874
rect 34841 22822 34893 22874
rect 34905 22822 34957 22874
rect 34969 22822 35021 22874
rect 4528 22720 4580 22772
rect 7564 22720 7616 22772
rect 3240 22652 3292 22704
rect 7104 22652 7156 22704
rect 8300 22695 8352 22704
rect 8300 22661 8309 22695
rect 8309 22661 8343 22695
rect 8343 22661 8352 22695
rect 8300 22652 8352 22661
rect 8484 22695 8536 22704
rect 8484 22661 8493 22695
rect 8493 22661 8527 22695
rect 8527 22661 8536 22695
rect 8484 22652 8536 22661
rect 4896 22627 4948 22636
rect 4896 22593 4905 22627
rect 4905 22593 4939 22627
rect 4939 22593 4948 22627
rect 4896 22584 4948 22593
rect 7472 22584 7524 22636
rect 8852 22584 8904 22636
rect 4988 22448 5040 22500
rect 12440 22720 12492 22772
rect 9772 22652 9824 22704
rect 9588 22584 9640 22636
rect 10416 22584 10468 22636
rect 11704 22627 11756 22636
rect 11704 22593 11713 22627
rect 11713 22593 11747 22627
rect 11747 22593 11756 22627
rect 11704 22584 11756 22593
rect 11796 22516 11848 22568
rect 12624 22584 12676 22636
rect 13268 22584 13320 22636
rect 31116 22720 31168 22772
rect 32036 22720 32088 22772
rect 15476 22652 15528 22704
rect 14740 22627 14792 22636
rect 12716 22516 12768 22568
rect 13084 22516 13136 22568
rect 14740 22593 14749 22627
rect 14749 22593 14783 22627
rect 14783 22593 14792 22627
rect 14740 22584 14792 22593
rect 15660 22627 15712 22636
rect 14096 22516 14148 22568
rect 14648 22516 14700 22568
rect 15660 22593 15669 22627
rect 15669 22593 15703 22627
rect 15703 22593 15712 22627
rect 15660 22584 15712 22593
rect 16396 22584 16448 22636
rect 17408 22627 17460 22636
rect 17408 22593 17417 22627
rect 17417 22593 17451 22627
rect 17451 22593 17460 22627
rect 17408 22584 17460 22593
rect 17500 22584 17552 22636
rect 18512 22652 18564 22704
rect 18696 22695 18748 22704
rect 18696 22661 18705 22695
rect 18705 22661 18739 22695
rect 18739 22661 18748 22695
rect 18696 22652 18748 22661
rect 25136 22652 25188 22704
rect 20076 22627 20128 22636
rect 20076 22593 20085 22627
rect 20085 22593 20119 22627
rect 20119 22593 20128 22627
rect 20076 22584 20128 22593
rect 11980 22448 12032 22500
rect 17960 22448 18012 22500
rect 20628 22584 20680 22636
rect 21180 22584 21232 22636
rect 21824 22584 21876 22636
rect 22192 22627 22244 22636
rect 22192 22593 22201 22627
rect 22201 22593 22235 22627
rect 22235 22593 22244 22627
rect 22192 22584 22244 22593
rect 27160 22584 27212 22636
rect 27988 22627 28040 22636
rect 27988 22593 27997 22627
rect 27997 22593 28031 22627
rect 28031 22593 28040 22627
rect 27988 22584 28040 22593
rect 28264 22584 28316 22636
rect 33140 22652 33192 22704
rect 33508 22695 33560 22704
rect 33508 22661 33517 22695
rect 33517 22661 33551 22695
rect 33551 22661 33560 22695
rect 33508 22652 33560 22661
rect 23848 22516 23900 22568
rect 26148 22516 26200 22568
rect 3608 22423 3660 22432
rect 3608 22389 3617 22423
rect 3617 22389 3651 22423
rect 3651 22389 3660 22423
rect 3608 22380 3660 22389
rect 3792 22423 3844 22432
rect 3792 22389 3801 22423
rect 3801 22389 3835 22423
rect 3835 22389 3844 22423
rect 3792 22380 3844 22389
rect 4344 22380 4396 22432
rect 4620 22380 4672 22432
rect 13176 22380 13228 22432
rect 18052 22423 18104 22432
rect 18052 22389 18061 22423
rect 18061 22389 18095 22423
rect 18095 22389 18104 22423
rect 18052 22380 18104 22389
rect 19892 22423 19944 22432
rect 19892 22389 19901 22423
rect 19901 22389 19935 22423
rect 19935 22389 19944 22423
rect 19892 22380 19944 22389
rect 23020 22380 23072 22432
rect 24584 22423 24636 22432
rect 24584 22389 24593 22423
rect 24593 22389 24627 22423
rect 24627 22389 24636 22423
rect 24584 22380 24636 22389
rect 26976 22380 27028 22432
rect 30380 22380 30432 22432
rect 31392 22584 31444 22636
rect 32680 22627 32732 22636
rect 32680 22593 32689 22627
rect 32689 22593 32723 22627
rect 32723 22593 32732 22627
rect 32680 22584 32732 22593
rect 33692 22627 33744 22636
rect 33692 22593 33701 22627
rect 33701 22593 33735 22627
rect 33735 22593 33744 22627
rect 33692 22584 33744 22593
rect 31300 22559 31352 22568
rect 31300 22525 31309 22559
rect 31309 22525 31343 22559
rect 31343 22525 31352 22559
rect 31300 22516 31352 22525
rect 32404 22516 32456 22568
rect 33324 22516 33376 22568
rect 31484 22448 31536 22500
rect 5170 22278 5222 22330
rect 5234 22278 5286 22330
rect 5298 22278 5350 22330
rect 5362 22278 5414 22330
rect 5426 22278 5478 22330
rect 13611 22278 13663 22330
rect 13675 22278 13727 22330
rect 13739 22278 13791 22330
rect 13803 22278 13855 22330
rect 13867 22278 13919 22330
rect 22052 22278 22104 22330
rect 22116 22278 22168 22330
rect 22180 22278 22232 22330
rect 22244 22278 22296 22330
rect 22308 22278 22360 22330
rect 30493 22278 30545 22330
rect 30557 22278 30609 22330
rect 30621 22278 30673 22330
rect 30685 22278 30737 22330
rect 30749 22278 30801 22330
rect 11704 22176 11756 22228
rect 16396 22176 16448 22228
rect 20076 22176 20128 22228
rect 20904 22176 20956 22228
rect 23020 22219 23072 22228
rect 23020 22185 23029 22219
rect 23029 22185 23063 22219
rect 23063 22185 23072 22219
rect 23020 22176 23072 22185
rect 6644 22108 6696 22160
rect 10324 22108 10376 22160
rect 12716 22108 12768 22160
rect 13084 22108 13136 22160
rect 13268 22108 13320 22160
rect 10784 22040 10836 22092
rect 7104 21972 7156 22024
rect 7472 21972 7524 22024
rect 9312 22015 9364 22024
rect 9312 21981 9321 22015
rect 9321 21981 9355 22015
rect 9355 21981 9364 22015
rect 9312 21972 9364 21981
rect 12072 22015 12124 22024
rect 12072 21981 12081 22015
rect 12081 21981 12115 22015
rect 12115 21981 12124 22015
rect 12072 21972 12124 21981
rect 11704 21904 11756 21956
rect 7196 21879 7248 21888
rect 7196 21845 7205 21879
rect 7205 21845 7239 21879
rect 7239 21845 7248 21879
rect 7196 21836 7248 21845
rect 8852 21836 8904 21888
rect 9036 21836 9088 21888
rect 10232 21836 10284 21888
rect 11060 21836 11112 21888
rect 18052 22040 18104 22092
rect 13176 21972 13228 22024
rect 17960 22015 18012 22024
rect 17960 21981 17969 22015
rect 17969 21981 18003 22015
rect 18003 21981 18012 22015
rect 17960 21972 18012 21981
rect 20444 22040 20496 22092
rect 18420 21972 18472 22024
rect 18788 21972 18840 22024
rect 22652 22108 22704 22160
rect 33692 22176 33744 22228
rect 24860 22083 24912 22092
rect 24860 22049 24869 22083
rect 24869 22049 24903 22083
rect 24903 22049 24912 22083
rect 24860 22040 24912 22049
rect 24952 22083 25004 22092
rect 24952 22049 24961 22083
rect 24961 22049 24995 22083
rect 24995 22049 25004 22083
rect 26976 22083 27028 22092
rect 24952 22040 25004 22049
rect 26976 22049 26985 22083
rect 26985 22049 27019 22083
rect 27019 22049 27028 22083
rect 26976 22040 27028 22049
rect 27252 22040 27304 22092
rect 29920 22040 29972 22092
rect 30380 22108 30432 22160
rect 33140 22083 33192 22092
rect 33140 22049 33149 22083
rect 33149 22049 33183 22083
rect 33183 22049 33192 22083
rect 33140 22040 33192 22049
rect 18236 21947 18288 21956
rect 18236 21913 18245 21947
rect 18245 21913 18279 21947
rect 18279 21913 18288 21947
rect 22836 21972 22888 22024
rect 24584 21972 24636 22024
rect 24768 22015 24820 22024
rect 24768 21981 24777 22015
rect 24777 21981 24811 22015
rect 24811 21981 24820 22015
rect 24768 21972 24820 21981
rect 25136 21972 25188 22024
rect 18236 21904 18288 21913
rect 18972 21836 19024 21888
rect 19800 21879 19852 21888
rect 19800 21845 19809 21879
rect 19809 21845 19843 21879
rect 19843 21845 19852 21879
rect 19800 21836 19852 21845
rect 21088 21904 21140 21956
rect 21548 21904 21600 21956
rect 27068 22015 27120 22024
rect 27068 21981 27077 22015
rect 27077 21981 27111 22015
rect 27111 21981 27120 22015
rect 27068 21972 27120 21981
rect 31024 22015 31076 22024
rect 27528 21904 27580 21956
rect 28448 21947 28500 21956
rect 28448 21913 28457 21947
rect 28457 21913 28491 21947
rect 28491 21913 28500 21947
rect 28448 21904 28500 21913
rect 31024 21981 31033 22015
rect 31033 21981 31067 22015
rect 31067 21981 31076 22015
rect 31392 22015 31444 22024
rect 31024 21972 31076 21981
rect 30380 21904 30432 21956
rect 31392 21981 31401 22015
rect 31401 21981 31435 22015
rect 31435 21981 31444 22015
rect 31392 21972 31444 21981
rect 31576 22015 31628 22024
rect 31576 21981 31585 22015
rect 31585 21981 31619 22015
rect 31619 21981 31628 22015
rect 31576 21972 31628 21981
rect 32404 22015 32456 22024
rect 32404 21981 32413 22015
rect 32413 21981 32447 22015
rect 32447 21981 32456 22015
rect 32404 21972 32456 21981
rect 32588 22015 32640 22024
rect 32588 21981 32597 22015
rect 32597 21981 32631 22015
rect 32631 21981 32640 22015
rect 32588 21972 32640 21981
rect 33324 22015 33376 22024
rect 33324 21981 33333 22015
rect 33333 21981 33367 22015
rect 33367 21981 33376 22015
rect 33324 21972 33376 21981
rect 21180 21836 21232 21888
rect 22284 21879 22336 21888
rect 22284 21845 22293 21879
rect 22293 21845 22327 21879
rect 22327 21845 22336 21879
rect 22284 21836 22336 21845
rect 25044 21836 25096 21888
rect 26884 21836 26936 21888
rect 26976 21836 27028 21888
rect 29736 21879 29788 21888
rect 29736 21845 29745 21879
rect 29745 21845 29779 21879
rect 29779 21845 29788 21879
rect 29736 21836 29788 21845
rect 9390 21734 9442 21786
rect 9454 21734 9506 21786
rect 9518 21734 9570 21786
rect 9582 21734 9634 21786
rect 9646 21734 9698 21786
rect 17831 21734 17883 21786
rect 17895 21734 17947 21786
rect 17959 21734 18011 21786
rect 18023 21734 18075 21786
rect 18087 21734 18139 21786
rect 26272 21734 26324 21786
rect 26336 21734 26388 21786
rect 26400 21734 26452 21786
rect 26464 21734 26516 21786
rect 26528 21734 26580 21786
rect 34713 21734 34765 21786
rect 34777 21734 34829 21786
rect 34841 21734 34893 21786
rect 34905 21734 34957 21786
rect 34969 21734 35021 21786
rect 18420 21632 18472 21684
rect 19432 21632 19484 21684
rect 11704 21607 11756 21616
rect 11704 21573 11713 21607
rect 11713 21573 11747 21607
rect 11747 21573 11756 21607
rect 11704 21564 11756 21573
rect 3608 21496 3660 21548
rect 7472 21496 7524 21548
rect 11796 21539 11848 21548
rect 11796 21505 11805 21539
rect 11805 21505 11839 21539
rect 11839 21505 11848 21539
rect 11796 21496 11848 21505
rect 11980 21539 12032 21548
rect 11980 21505 11989 21539
rect 11989 21505 12023 21539
rect 12023 21505 12032 21539
rect 11980 21496 12032 21505
rect 14004 21496 14056 21548
rect 15292 21539 15344 21548
rect 15292 21505 15301 21539
rect 15301 21505 15335 21539
rect 15335 21505 15344 21539
rect 15292 21496 15344 21505
rect 15752 21496 15804 21548
rect 17684 21496 17736 21548
rect 20536 21632 20588 21684
rect 26976 21632 27028 21684
rect 27160 21675 27212 21684
rect 27160 21641 27169 21675
rect 27169 21641 27203 21675
rect 27203 21641 27212 21675
rect 27160 21632 27212 21641
rect 27528 21632 27580 21684
rect 30380 21675 30432 21684
rect 30380 21641 30389 21675
rect 30389 21641 30423 21675
rect 30423 21641 30432 21675
rect 30380 21632 30432 21641
rect 31760 21632 31812 21684
rect 19892 21539 19944 21548
rect 19892 21505 19901 21539
rect 19901 21505 19935 21539
rect 19935 21505 19944 21539
rect 19892 21496 19944 21505
rect 26884 21564 26936 21616
rect 22284 21539 22336 21548
rect 3700 21428 3752 21480
rect 4436 21428 4488 21480
rect 18236 21428 18288 21480
rect 3056 21335 3108 21344
rect 3056 21301 3065 21335
rect 3065 21301 3099 21335
rect 3099 21301 3108 21335
rect 3608 21335 3660 21344
rect 3056 21292 3108 21301
rect 3608 21301 3617 21335
rect 3617 21301 3651 21335
rect 3651 21301 3660 21335
rect 3608 21292 3660 21301
rect 3700 21292 3752 21344
rect 4068 21360 4120 21412
rect 19248 21360 19300 21412
rect 22284 21505 22293 21539
rect 22293 21505 22327 21539
rect 22327 21505 22336 21539
rect 22284 21496 22336 21505
rect 27712 21496 27764 21548
rect 28448 21564 28500 21616
rect 22376 21471 22428 21480
rect 22376 21437 22385 21471
rect 22385 21437 22419 21471
rect 22419 21437 22428 21471
rect 22376 21428 22428 21437
rect 23204 21471 23256 21480
rect 23204 21437 23213 21471
rect 23213 21437 23247 21471
rect 23247 21437 23256 21471
rect 23204 21428 23256 21437
rect 23572 21428 23624 21480
rect 23940 21428 23992 21480
rect 27344 21428 27396 21480
rect 27620 21428 27672 21480
rect 29736 21496 29788 21548
rect 30472 21564 30524 21616
rect 31024 21564 31076 21616
rect 31392 21564 31444 21616
rect 31484 21539 31536 21548
rect 31484 21505 31493 21539
rect 31493 21505 31527 21539
rect 31527 21505 31536 21539
rect 31484 21496 31536 21505
rect 32588 21496 32640 21548
rect 15384 21292 15436 21344
rect 15844 21292 15896 21344
rect 15936 21292 15988 21344
rect 23848 21292 23900 21344
rect 27896 21292 27948 21344
rect 28448 21292 28500 21344
rect 5170 21190 5222 21242
rect 5234 21190 5286 21242
rect 5298 21190 5350 21242
rect 5362 21190 5414 21242
rect 5426 21190 5478 21242
rect 13611 21190 13663 21242
rect 13675 21190 13727 21242
rect 13739 21190 13791 21242
rect 13803 21190 13855 21242
rect 13867 21190 13919 21242
rect 22052 21190 22104 21242
rect 22116 21190 22168 21242
rect 22180 21190 22232 21242
rect 22244 21190 22296 21242
rect 22308 21190 22360 21242
rect 30493 21190 30545 21242
rect 30557 21190 30609 21242
rect 30621 21190 30673 21242
rect 30685 21190 30737 21242
rect 30749 21190 30801 21242
rect 13084 21088 13136 21140
rect 17316 21088 17368 21140
rect 18788 21131 18840 21140
rect 18788 21097 18797 21131
rect 18797 21097 18831 21131
rect 18831 21097 18840 21131
rect 18788 21088 18840 21097
rect 21272 21131 21324 21140
rect 21272 21097 21281 21131
rect 21281 21097 21315 21131
rect 21315 21097 21324 21131
rect 21272 21088 21324 21097
rect 23572 21131 23624 21140
rect 23572 21097 23581 21131
rect 23581 21097 23615 21131
rect 23615 21097 23624 21131
rect 23572 21088 23624 21097
rect 23756 21088 23808 21140
rect 30932 21088 30984 21140
rect 31484 21131 31536 21140
rect 31484 21097 31493 21131
rect 31493 21097 31527 21131
rect 31527 21097 31536 21131
rect 31484 21088 31536 21097
rect 32404 21131 32456 21140
rect 32404 21097 32413 21131
rect 32413 21097 32447 21131
rect 32447 21097 32456 21131
rect 32404 21088 32456 21097
rect 25872 21020 25924 21072
rect 25964 21020 26016 21072
rect 32496 21020 32548 21072
rect 7472 20952 7524 21004
rect 3240 20927 3292 20936
rect 3240 20893 3249 20927
rect 3249 20893 3283 20927
rect 3283 20893 3292 20927
rect 3240 20884 3292 20893
rect 4436 20884 4488 20936
rect 7288 20884 7340 20936
rect 7656 20927 7708 20936
rect 7656 20893 7665 20927
rect 7665 20893 7699 20927
rect 7699 20893 7708 20927
rect 7656 20884 7708 20893
rect 10140 20884 10192 20936
rect 10416 20927 10468 20936
rect 10416 20893 10425 20927
rect 10425 20893 10459 20927
rect 10459 20893 10468 20927
rect 10416 20884 10468 20893
rect 10784 20884 10836 20936
rect 13452 20884 13504 20936
rect 14464 20927 14516 20936
rect 14464 20893 14473 20927
rect 14473 20893 14507 20927
rect 14507 20893 14516 20927
rect 14464 20884 14516 20893
rect 18328 20884 18380 20936
rect 11888 20816 11940 20868
rect 15936 20816 15988 20868
rect 20076 20952 20128 21004
rect 21456 20952 21508 21004
rect 19248 20884 19300 20936
rect 28448 20952 28500 21004
rect 22560 20927 22612 20936
rect 22560 20893 22569 20927
rect 22569 20893 22603 20927
rect 22603 20893 22612 20927
rect 22560 20884 22612 20893
rect 23756 20927 23808 20936
rect 3148 20748 3200 20800
rect 7380 20791 7432 20800
rect 7380 20757 7389 20791
rect 7389 20757 7423 20791
rect 7423 20757 7432 20791
rect 7380 20748 7432 20757
rect 10232 20791 10284 20800
rect 10232 20757 10241 20791
rect 10241 20757 10275 20791
rect 10275 20757 10284 20791
rect 10232 20748 10284 20757
rect 14280 20791 14332 20800
rect 14280 20757 14289 20791
rect 14289 20757 14323 20791
rect 14323 20757 14332 20791
rect 14280 20748 14332 20757
rect 15844 20748 15896 20800
rect 21180 20816 21232 20868
rect 23756 20893 23765 20927
rect 23765 20893 23799 20927
rect 23799 20893 23808 20927
rect 23756 20884 23808 20893
rect 23940 20927 23992 20936
rect 23940 20893 23949 20927
rect 23949 20893 23983 20927
rect 23983 20893 23992 20927
rect 23940 20884 23992 20893
rect 23388 20748 23440 20800
rect 23940 20748 23992 20800
rect 24676 20884 24728 20936
rect 24124 20816 24176 20868
rect 25504 20884 25556 20936
rect 28724 20884 28776 20936
rect 32220 20927 32272 20936
rect 27344 20816 27396 20868
rect 29092 20816 29144 20868
rect 32220 20893 32229 20927
rect 32229 20893 32263 20927
rect 32263 20893 32272 20927
rect 32220 20884 32272 20893
rect 32312 20884 32364 20936
rect 32956 20927 33008 20936
rect 32956 20893 32965 20927
rect 32965 20893 32999 20927
rect 32999 20893 33008 20927
rect 32956 20884 33008 20893
rect 32772 20816 32824 20868
rect 33048 20816 33100 20868
rect 24952 20791 25004 20800
rect 24952 20757 24961 20791
rect 24961 20757 24995 20791
rect 24995 20757 25004 20791
rect 24952 20748 25004 20757
rect 32220 20748 32272 20800
rect 32404 20748 32456 20800
rect 9390 20646 9442 20698
rect 9454 20646 9506 20698
rect 9518 20646 9570 20698
rect 9582 20646 9634 20698
rect 9646 20646 9698 20698
rect 17831 20646 17883 20698
rect 17895 20646 17947 20698
rect 17959 20646 18011 20698
rect 18023 20646 18075 20698
rect 18087 20646 18139 20698
rect 26272 20646 26324 20698
rect 26336 20646 26388 20698
rect 26400 20646 26452 20698
rect 26464 20646 26516 20698
rect 26528 20646 26580 20698
rect 34713 20646 34765 20698
rect 34777 20646 34829 20698
rect 34841 20646 34893 20698
rect 34905 20646 34957 20698
rect 34969 20646 35021 20698
rect 8300 20544 8352 20596
rect 20996 20587 21048 20596
rect 3608 20519 3660 20528
rect 3608 20485 3617 20519
rect 3617 20485 3651 20519
rect 3651 20485 3660 20519
rect 3608 20476 3660 20485
rect 7748 20476 7800 20528
rect 20996 20553 21005 20587
rect 21005 20553 21039 20587
rect 21039 20553 21048 20587
rect 20996 20544 21048 20553
rect 21640 20544 21692 20596
rect 22284 20544 22336 20596
rect 24676 20544 24728 20596
rect 25964 20544 26016 20596
rect 31576 20587 31628 20596
rect 31576 20553 31585 20587
rect 31585 20553 31619 20587
rect 31619 20553 31628 20587
rect 31576 20544 31628 20553
rect 32588 20587 32640 20596
rect 32588 20553 32597 20587
rect 32597 20553 32631 20587
rect 32631 20553 32640 20587
rect 32588 20544 32640 20553
rect 3148 20451 3200 20460
rect 3148 20417 3157 20451
rect 3157 20417 3191 20451
rect 3191 20417 3200 20451
rect 3148 20408 3200 20417
rect 3976 20408 4028 20460
rect 3056 20340 3108 20392
rect 3424 20340 3476 20392
rect 4068 20383 4120 20392
rect 4068 20349 4077 20383
rect 4077 20349 4111 20383
rect 4111 20349 4120 20383
rect 4068 20340 4120 20349
rect 4344 20383 4396 20392
rect 4344 20349 4353 20383
rect 4353 20349 4387 20383
rect 4387 20349 4396 20383
rect 4344 20340 4396 20349
rect 1860 20272 1912 20324
rect 7288 20408 7340 20460
rect 8024 20408 8076 20460
rect 8484 20451 8536 20460
rect 8484 20417 8493 20451
rect 8493 20417 8527 20451
rect 8527 20417 8536 20451
rect 8484 20408 8536 20417
rect 10232 20408 10284 20460
rect 11060 20451 11112 20460
rect 11060 20417 11069 20451
rect 11069 20417 11103 20451
rect 11103 20417 11112 20451
rect 11060 20408 11112 20417
rect 14280 20476 14332 20528
rect 16212 20476 16264 20528
rect 19708 20476 19760 20528
rect 20720 20519 20772 20528
rect 20720 20485 20729 20519
rect 20729 20485 20763 20519
rect 20763 20485 20772 20519
rect 20720 20476 20772 20485
rect 22376 20476 22428 20528
rect 15108 20451 15160 20460
rect 8944 20340 8996 20392
rect 10416 20383 10468 20392
rect 10416 20349 10425 20383
rect 10425 20349 10459 20383
rect 10459 20349 10468 20383
rect 10416 20340 10468 20349
rect 5080 20272 5132 20324
rect 6920 20272 6972 20324
rect 7840 20272 7892 20324
rect 13728 20340 13780 20392
rect 13176 20272 13228 20324
rect 2780 20204 2832 20256
rect 12900 20204 12952 20256
rect 15108 20417 15117 20451
rect 15117 20417 15151 20451
rect 15151 20417 15160 20451
rect 15108 20408 15160 20417
rect 15384 20408 15436 20460
rect 15752 20408 15804 20460
rect 20352 20408 20404 20460
rect 14096 20272 14148 20324
rect 16948 20340 17000 20392
rect 17224 20340 17276 20392
rect 17316 20340 17368 20392
rect 20536 20408 20588 20460
rect 20996 20408 21048 20460
rect 27988 20451 28040 20460
rect 27988 20417 27997 20451
rect 27997 20417 28031 20451
rect 28031 20417 28040 20451
rect 27988 20408 28040 20417
rect 27896 20383 27948 20392
rect 27896 20349 27905 20383
rect 27905 20349 27939 20383
rect 27939 20349 27948 20383
rect 27896 20340 27948 20349
rect 32588 20408 32640 20460
rect 32772 20451 32824 20460
rect 32772 20417 32781 20451
rect 32781 20417 32815 20451
rect 32815 20417 32824 20451
rect 32772 20408 32824 20417
rect 33048 20451 33100 20460
rect 33048 20417 33057 20451
rect 33057 20417 33091 20451
rect 33091 20417 33100 20451
rect 33048 20408 33100 20417
rect 31944 20340 31996 20392
rect 14832 20272 14884 20324
rect 17408 20204 17460 20256
rect 18696 20247 18748 20256
rect 18696 20213 18705 20247
rect 18705 20213 18739 20247
rect 18739 20213 18748 20247
rect 18696 20204 18748 20213
rect 20812 20272 20864 20324
rect 32312 20272 32364 20324
rect 32956 20315 33008 20324
rect 32956 20281 32965 20315
rect 32965 20281 32999 20315
rect 32999 20281 33008 20315
rect 32956 20272 33008 20281
rect 28080 20204 28132 20256
rect 5170 20102 5222 20154
rect 5234 20102 5286 20154
rect 5298 20102 5350 20154
rect 5362 20102 5414 20154
rect 5426 20102 5478 20154
rect 13611 20102 13663 20154
rect 13675 20102 13727 20154
rect 13739 20102 13791 20154
rect 13803 20102 13855 20154
rect 13867 20102 13919 20154
rect 22052 20102 22104 20154
rect 22116 20102 22168 20154
rect 22180 20102 22232 20154
rect 22244 20102 22296 20154
rect 22308 20102 22360 20154
rect 30493 20102 30545 20154
rect 30557 20102 30609 20154
rect 30621 20102 30673 20154
rect 30685 20102 30737 20154
rect 30749 20102 30801 20154
rect 3976 20043 4028 20052
rect 3976 20009 3985 20043
rect 3985 20009 4019 20043
rect 4019 20009 4028 20043
rect 3976 20000 4028 20009
rect 4712 20000 4764 20052
rect 5080 20043 5132 20052
rect 5080 20009 5089 20043
rect 5089 20009 5123 20043
rect 5123 20009 5132 20043
rect 5080 20000 5132 20009
rect 3792 19932 3844 19984
rect 4344 19864 4396 19916
rect 1860 19839 1912 19848
rect 1860 19805 1869 19839
rect 1869 19805 1903 19839
rect 1903 19805 1912 19839
rect 1860 19796 1912 19805
rect 3240 19728 3292 19780
rect 3976 19728 4028 19780
rect 3332 19660 3384 19712
rect 4160 19839 4212 19848
rect 4160 19805 4169 19839
rect 4169 19805 4203 19839
rect 4203 19805 4212 19839
rect 4160 19796 4212 19805
rect 4252 19771 4304 19780
rect 4252 19737 4261 19771
rect 4261 19737 4295 19771
rect 4295 19737 4304 19771
rect 4252 19728 4304 19737
rect 4436 19660 4488 19712
rect 4620 19839 4672 19848
rect 4620 19805 4629 19839
rect 4629 19805 4663 19839
rect 4663 19805 4672 19839
rect 4620 19796 4672 19805
rect 6644 19932 6696 19984
rect 7104 19975 7156 19984
rect 7104 19941 7113 19975
rect 7113 19941 7147 19975
rect 7147 19941 7156 19975
rect 7104 19932 7156 19941
rect 7656 20000 7708 20052
rect 15292 20000 15344 20052
rect 24768 20000 24820 20052
rect 7748 19975 7800 19984
rect 7748 19941 7757 19975
rect 7757 19941 7791 19975
rect 7791 19941 7800 19975
rect 7748 19932 7800 19941
rect 5448 19839 5500 19848
rect 5448 19805 5457 19839
rect 5457 19805 5491 19839
rect 5491 19805 5500 19839
rect 5448 19796 5500 19805
rect 6552 19728 6604 19780
rect 7380 19796 7432 19848
rect 8024 19839 8076 19848
rect 8024 19805 8033 19839
rect 8033 19805 8067 19839
rect 8067 19805 8076 19839
rect 8024 19796 8076 19805
rect 8484 19796 8536 19848
rect 11888 19907 11940 19916
rect 9956 19796 10008 19848
rect 10416 19839 10468 19848
rect 10416 19805 10425 19839
rect 10425 19805 10459 19839
rect 10459 19805 10468 19839
rect 10416 19796 10468 19805
rect 11888 19873 11897 19907
rect 11897 19873 11931 19907
rect 11931 19873 11940 19907
rect 11888 19864 11940 19873
rect 15108 19864 15160 19916
rect 10876 19839 10928 19848
rect 10876 19805 10885 19839
rect 10885 19805 10919 19839
rect 10919 19805 10928 19839
rect 10876 19796 10928 19805
rect 12716 19796 12768 19848
rect 13176 19796 13228 19848
rect 13452 19796 13504 19848
rect 14464 19839 14516 19848
rect 14464 19805 14473 19839
rect 14473 19805 14507 19839
rect 14507 19805 14516 19839
rect 14464 19796 14516 19805
rect 17040 19864 17092 19916
rect 20996 19932 21048 19984
rect 32312 19975 32364 19984
rect 32312 19941 32321 19975
rect 32321 19941 32355 19975
rect 32355 19941 32364 19975
rect 32312 19932 32364 19941
rect 19340 19864 19392 19916
rect 7288 19728 7340 19780
rect 8944 19728 8996 19780
rect 9772 19728 9824 19780
rect 10232 19728 10284 19780
rect 12440 19728 12492 19780
rect 15752 19796 15804 19848
rect 15844 19796 15896 19848
rect 17132 19796 17184 19848
rect 18236 19796 18288 19848
rect 19432 19839 19484 19848
rect 19432 19805 19441 19839
rect 19441 19805 19475 19839
rect 19475 19805 19484 19839
rect 19432 19796 19484 19805
rect 19524 19839 19576 19848
rect 19524 19805 19534 19839
rect 19534 19805 19568 19839
rect 19568 19805 19576 19839
rect 19800 19839 19852 19848
rect 19524 19796 19576 19805
rect 19800 19805 19809 19839
rect 19809 19805 19843 19839
rect 19843 19805 19852 19839
rect 19800 19796 19852 19805
rect 20536 19864 20588 19916
rect 23204 19864 23256 19916
rect 28816 19839 28868 19848
rect 16764 19771 16816 19780
rect 16764 19737 16773 19771
rect 16773 19737 16807 19771
rect 16807 19737 16816 19771
rect 16764 19728 16816 19737
rect 17684 19728 17736 19780
rect 19708 19771 19760 19780
rect 19708 19737 19717 19771
rect 19717 19737 19751 19771
rect 19751 19737 19760 19771
rect 19708 19728 19760 19737
rect 20812 19771 20864 19780
rect 20812 19737 20821 19771
rect 20821 19737 20855 19771
rect 20855 19737 20864 19771
rect 20812 19728 20864 19737
rect 28816 19805 28825 19839
rect 28825 19805 28859 19839
rect 28859 19805 28868 19839
rect 28816 19796 28868 19805
rect 28908 19796 28960 19848
rect 31760 19796 31812 19848
rect 31944 19839 31996 19848
rect 31944 19805 31953 19839
rect 31953 19805 31987 19839
rect 31987 19805 31996 19839
rect 31944 19796 31996 19805
rect 32220 19839 32272 19848
rect 32220 19805 32229 19839
rect 32229 19805 32263 19839
rect 32263 19805 32272 19839
rect 32220 19796 32272 19805
rect 32404 19839 32456 19848
rect 32404 19805 32413 19839
rect 32413 19805 32447 19839
rect 32447 19805 32456 19839
rect 32404 19796 32456 19805
rect 32588 19839 32640 19848
rect 32588 19805 32597 19839
rect 32597 19805 32631 19839
rect 32631 19805 32640 19839
rect 32588 19796 32640 19805
rect 28724 19728 28776 19780
rect 7472 19660 7524 19712
rect 11520 19703 11572 19712
rect 11520 19669 11529 19703
rect 11529 19669 11563 19703
rect 11563 19669 11572 19703
rect 11520 19660 11572 19669
rect 15292 19660 15344 19712
rect 17316 19660 17368 19712
rect 19432 19660 19484 19712
rect 20260 19660 20312 19712
rect 28172 19660 28224 19712
rect 9390 19558 9442 19610
rect 9454 19558 9506 19610
rect 9518 19558 9570 19610
rect 9582 19558 9634 19610
rect 9646 19558 9698 19610
rect 17831 19558 17883 19610
rect 17895 19558 17947 19610
rect 17959 19558 18011 19610
rect 18023 19558 18075 19610
rect 18087 19558 18139 19610
rect 26272 19558 26324 19610
rect 26336 19558 26388 19610
rect 26400 19558 26452 19610
rect 26464 19558 26516 19610
rect 26528 19558 26580 19610
rect 34713 19558 34765 19610
rect 34777 19558 34829 19610
rect 34841 19558 34893 19610
rect 34905 19558 34957 19610
rect 34969 19558 35021 19610
rect 4068 19456 4120 19508
rect 4896 19456 4948 19508
rect 6920 19456 6972 19508
rect 19524 19456 19576 19508
rect 20720 19456 20772 19508
rect 2780 19363 2832 19372
rect 2780 19329 2789 19363
rect 2789 19329 2823 19363
rect 2823 19329 2832 19363
rect 2780 19320 2832 19329
rect 3516 19320 3568 19372
rect 3884 19320 3936 19372
rect 4712 19388 4764 19440
rect 16764 19388 16816 19440
rect 23020 19456 23072 19508
rect 32220 19456 32272 19508
rect 33048 19456 33100 19508
rect 4804 19363 4856 19372
rect 4804 19329 4813 19363
rect 4813 19329 4847 19363
rect 4847 19329 4856 19363
rect 4804 19320 4856 19329
rect 4896 19363 4948 19372
rect 4896 19329 4905 19363
rect 4905 19329 4939 19363
rect 4939 19329 4948 19363
rect 4896 19320 4948 19329
rect 7656 19320 7708 19372
rect 8944 19320 8996 19372
rect 9772 19320 9824 19372
rect 10324 19320 10376 19372
rect 12440 19363 12492 19372
rect 12440 19329 12449 19363
rect 12449 19329 12483 19363
rect 12483 19329 12492 19363
rect 12440 19320 12492 19329
rect 13268 19320 13320 19372
rect 24952 19388 25004 19440
rect 17132 19320 17184 19372
rect 18696 19320 18748 19372
rect 11060 19252 11112 19304
rect 11520 19252 11572 19304
rect 14740 19252 14792 19304
rect 20996 19320 21048 19372
rect 22376 19320 22428 19372
rect 23204 19320 23256 19372
rect 27344 19320 27396 19372
rect 27436 19363 27488 19372
rect 27436 19329 27445 19363
rect 27445 19329 27479 19363
rect 27479 19329 27488 19363
rect 27436 19320 27488 19329
rect 29092 19363 29144 19372
rect 23388 19295 23440 19304
rect 23388 19261 23397 19295
rect 23397 19261 23431 19295
rect 23431 19261 23440 19295
rect 23388 19252 23440 19261
rect 28724 19295 28776 19304
rect 28724 19261 28733 19295
rect 28733 19261 28767 19295
rect 28767 19261 28776 19295
rect 28724 19252 28776 19261
rect 29092 19329 29101 19363
rect 29101 19329 29135 19363
rect 29135 19329 29144 19363
rect 29092 19320 29144 19329
rect 29736 19363 29788 19372
rect 29736 19329 29745 19363
rect 29745 19329 29779 19363
rect 29779 19329 29788 19363
rect 29736 19320 29788 19329
rect 31208 19363 31260 19372
rect 31208 19329 31217 19363
rect 31217 19329 31251 19363
rect 31251 19329 31260 19363
rect 31208 19320 31260 19329
rect 31944 19388 31996 19440
rect 32404 19388 32456 19440
rect 32588 19363 32640 19372
rect 32588 19329 32597 19363
rect 32597 19329 32631 19363
rect 32631 19329 32640 19363
rect 32588 19320 32640 19329
rect 4620 19227 4672 19236
rect 4620 19193 4629 19227
rect 4629 19193 4663 19227
rect 4663 19193 4672 19227
rect 4620 19184 4672 19193
rect 4252 19116 4304 19168
rect 5448 19116 5500 19168
rect 9772 19184 9824 19236
rect 31760 19252 31812 19304
rect 32680 19252 32732 19304
rect 8208 19116 8260 19168
rect 9128 19159 9180 19168
rect 9128 19125 9137 19159
rect 9137 19125 9171 19159
rect 9171 19125 9180 19159
rect 9128 19116 9180 19125
rect 10232 19159 10284 19168
rect 10232 19125 10241 19159
rect 10241 19125 10275 19159
rect 10275 19125 10284 19159
rect 10232 19116 10284 19125
rect 10692 19159 10744 19168
rect 10692 19125 10701 19159
rect 10701 19125 10735 19159
rect 10735 19125 10744 19159
rect 10692 19116 10744 19125
rect 26424 19116 26476 19168
rect 5170 19014 5222 19066
rect 5234 19014 5286 19066
rect 5298 19014 5350 19066
rect 5362 19014 5414 19066
rect 5426 19014 5478 19066
rect 13611 19014 13663 19066
rect 13675 19014 13727 19066
rect 13739 19014 13791 19066
rect 13803 19014 13855 19066
rect 13867 19014 13919 19066
rect 22052 19014 22104 19066
rect 22116 19014 22168 19066
rect 22180 19014 22232 19066
rect 22244 19014 22296 19066
rect 22308 19014 22360 19066
rect 30493 19014 30545 19066
rect 30557 19014 30609 19066
rect 30621 19014 30673 19066
rect 30685 19014 30737 19066
rect 30749 19014 30801 19066
rect 7656 18955 7708 18964
rect 7656 18921 7665 18955
rect 7665 18921 7699 18955
rect 7699 18921 7708 18955
rect 7656 18912 7708 18921
rect 17316 18912 17368 18964
rect 17408 18912 17460 18964
rect 25872 18955 25924 18964
rect 25872 18921 25881 18955
rect 25881 18921 25915 18955
rect 25915 18921 25924 18955
rect 25872 18912 25924 18921
rect 28264 18955 28316 18964
rect 28264 18921 28273 18955
rect 28273 18921 28307 18955
rect 28307 18921 28316 18955
rect 28264 18912 28316 18921
rect 33324 18912 33376 18964
rect 2964 18844 3016 18896
rect 7104 18776 7156 18828
rect 8484 18844 8536 18896
rect 9128 18776 9180 18828
rect 27804 18844 27856 18896
rect 3332 18751 3384 18760
rect 3332 18717 3341 18751
rect 3341 18717 3375 18751
rect 3375 18717 3384 18751
rect 3332 18708 3384 18717
rect 3424 18751 3476 18760
rect 3424 18717 3433 18751
rect 3433 18717 3467 18751
rect 3467 18717 3476 18751
rect 3424 18708 3476 18717
rect 10232 18708 10284 18760
rect 3240 18640 3292 18692
rect 7196 18640 7248 18692
rect 8208 18640 8260 18692
rect 10692 18708 10744 18760
rect 12440 18708 12492 18760
rect 14740 18708 14792 18760
rect 15292 18708 15344 18760
rect 21732 18708 21784 18760
rect 24492 18708 24544 18760
rect 26424 18776 26476 18828
rect 28724 18819 28776 18828
rect 28724 18785 28733 18819
rect 28733 18785 28767 18819
rect 28767 18785 28776 18819
rect 28724 18776 28776 18785
rect 28908 18819 28960 18828
rect 28908 18785 28917 18819
rect 28917 18785 28951 18819
rect 28951 18785 28960 18819
rect 28908 18776 28960 18785
rect 29092 18776 29144 18828
rect 25228 18708 25280 18760
rect 25504 18708 25556 18760
rect 26240 18751 26292 18760
rect 26240 18717 26249 18751
rect 26249 18717 26283 18751
rect 26283 18717 26292 18751
rect 26240 18708 26292 18717
rect 27344 18751 27396 18760
rect 16212 18640 16264 18692
rect 17316 18640 17368 18692
rect 19524 18640 19576 18692
rect 20904 18640 20956 18692
rect 25688 18640 25740 18692
rect 27344 18717 27353 18751
rect 27353 18717 27387 18751
rect 27387 18717 27396 18751
rect 27344 18708 27396 18717
rect 27436 18708 27488 18760
rect 27620 18708 27672 18760
rect 28816 18708 28868 18760
rect 29828 18751 29880 18760
rect 29828 18717 29837 18751
rect 29837 18717 29871 18751
rect 29871 18717 29880 18751
rect 32496 18776 32548 18828
rect 32588 18776 32640 18828
rect 29828 18708 29880 18717
rect 29460 18640 29512 18692
rect 32864 18708 32916 18760
rect 32404 18640 32456 18692
rect 19340 18572 19392 18624
rect 20352 18572 20404 18624
rect 23480 18572 23532 18624
rect 24216 18572 24268 18624
rect 24584 18615 24636 18624
rect 24584 18581 24593 18615
rect 24593 18581 24627 18615
rect 24627 18581 24636 18615
rect 24584 18572 24636 18581
rect 25136 18572 25188 18624
rect 26240 18572 26292 18624
rect 27068 18572 27120 18624
rect 9390 18470 9442 18522
rect 9454 18470 9506 18522
rect 9518 18470 9570 18522
rect 9582 18470 9634 18522
rect 9646 18470 9698 18522
rect 17831 18470 17883 18522
rect 17895 18470 17947 18522
rect 17959 18470 18011 18522
rect 18023 18470 18075 18522
rect 18087 18470 18139 18522
rect 26272 18470 26324 18522
rect 26336 18470 26388 18522
rect 26400 18470 26452 18522
rect 26464 18470 26516 18522
rect 26528 18470 26580 18522
rect 34713 18470 34765 18522
rect 34777 18470 34829 18522
rect 34841 18470 34893 18522
rect 34905 18470 34957 18522
rect 34969 18470 35021 18522
rect 8944 18368 8996 18420
rect 17684 18368 17736 18420
rect 19800 18368 19852 18420
rect 21088 18368 21140 18420
rect 7196 18300 7248 18352
rect 11980 18300 12032 18352
rect 14740 18343 14792 18352
rect 6644 18232 6696 18284
rect 8208 18275 8260 18284
rect 8208 18241 8217 18275
rect 8217 18241 8251 18275
rect 8251 18241 8260 18275
rect 8208 18232 8260 18241
rect 11060 18232 11112 18284
rect 11796 18232 11848 18284
rect 12348 18275 12400 18284
rect 12348 18241 12357 18275
rect 12357 18241 12391 18275
rect 12391 18241 12400 18275
rect 12348 18232 12400 18241
rect 14740 18309 14749 18343
rect 14749 18309 14783 18343
rect 14783 18309 14792 18343
rect 14740 18300 14792 18309
rect 15292 18300 15344 18352
rect 12992 18275 13044 18284
rect 12992 18241 13001 18275
rect 13001 18241 13035 18275
rect 13035 18241 13044 18275
rect 12992 18232 13044 18241
rect 16672 18300 16724 18352
rect 17316 18343 17368 18352
rect 17316 18309 17325 18343
rect 17325 18309 17359 18343
rect 17359 18309 17368 18343
rect 17316 18300 17368 18309
rect 18972 18343 19024 18352
rect 18972 18309 19006 18343
rect 19006 18309 19024 18343
rect 18972 18300 19024 18309
rect 24492 18368 24544 18420
rect 25688 18411 25740 18420
rect 25688 18377 25697 18411
rect 25697 18377 25731 18411
rect 25731 18377 25740 18411
rect 25688 18368 25740 18377
rect 27620 18368 27672 18420
rect 32864 18368 32916 18420
rect 18696 18275 18748 18284
rect 6736 18207 6788 18216
rect 6736 18173 6745 18207
rect 6745 18173 6779 18207
rect 6779 18173 6788 18207
rect 6736 18164 6788 18173
rect 6920 18207 6972 18216
rect 6920 18173 6929 18207
rect 6929 18173 6963 18207
rect 6963 18173 6972 18207
rect 6920 18164 6972 18173
rect 12164 18207 12216 18216
rect 12164 18173 12173 18207
rect 12173 18173 12207 18207
rect 12207 18173 12216 18207
rect 12164 18164 12216 18173
rect 7288 18139 7340 18148
rect 7288 18105 7297 18139
rect 7297 18105 7331 18139
rect 7331 18105 7340 18139
rect 7288 18096 7340 18105
rect 18696 18241 18705 18275
rect 18705 18241 18739 18275
rect 18739 18241 18748 18275
rect 18696 18232 18748 18241
rect 24216 18300 24268 18352
rect 29092 18300 29144 18352
rect 20904 18232 20956 18284
rect 23480 18275 23532 18284
rect 23480 18241 23489 18275
rect 23489 18241 23523 18275
rect 23523 18241 23532 18275
rect 23480 18232 23532 18241
rect 25320 18275 25372 18284
rect 25320 18241 25329 18275
rect 25329 18241 25363 18275
rect 25363 18241 25372 18275
rect 25320 18232 25372 18241
rect 28172 18275 28224 18284
rect 28172 18241 28181 18275
rect 28181 18241 28215 18275
rect 28215 18241 28224 18275
rect 28172 18232 28224 18241
rect 28540 18232 28592 18284
rect 28816 18232 28868 18284
rect 29184 18275 29236 18284
rect 29184 18241 29193 18275
rect 29193 18241 29227 18275
rect 29227 18241 29236 18275
rect 29184 18232 29236 18241
rect 29276 18275 29328 18284
rect 29276 18241 29285 18275
rect 29285 18241 29319 18275
rect 29319 18241 29328 18275
rect 32496 18275 32548 18284
rect 29276 18232 29328 18241
rect 32496 18241 32505 18275
rect 32505 18241 32539 18275
rect 32539 18241 32548 18275
rect 32496 18232 32548 18241
rect 23112 18164 23164 18216
rect 25412 18207 25464 18216
rect 25412 18173 25421 18207
rect 25421 18173 25455 18207
rect 25455 18173 25464 18207
rect 25412 18164 25464 18173
rect 27344 18164 27396 18216
rect 29460 18164 29512 18216
rect 32312 18207 32364 18216
rect 32312 18173 32321 18207
rect 32321 18173 32355 18207
rect 32355 18173 32364 18207
rect 32312 18164 32364 18173
rect 32864 18207 32916 18216
rect 32864 18173 32873 18207
rect 32873 18173 32907 18207
rect 32907 18173 32916 18207
rect 32864 18164 32916 18173
rect 34336 18207 34388 18216
rect 34336 18173 34345 18207
rect 34345 18173 34379 18207
rect 34379 18173 34388 18207
rect 34336 18164 34388 18173
rect 17316 18096 17368 18148
rect 10232 18071 10284 18080
rect 10232 18037 10241 18071
rect 10241 18037 10275 18071
rect 10275 18037 10284 18071
rect 10232 18028 10284 18037
rect 15844 18071 15896 18080
rect 15844 18037 15853 18071
rect 15853 18037 15887 18071
rect 15887 18037 15896 18071
rect 15844 18028 15896 18037
rect 16948 18071 17000 18080
rect 16948 18037 16957 18071
rect 16957 18037 16991 18071
rect 16991 18037 17000 18071
rect 16948 18028 17000 18037
rect 17408 18028 17460 18080
rect 20536 18071 20588 18080
rect 20536 18037 20545 18071
rect 20545 18037 20579 18071
rect 20579 18037 20588 18071
rect 20536 18028 20588 18037
rect 24952 18028 25004 18080
rect 5170 17926 5222 17978
rect 5234 17926 5286 17978
rect 5298 17926 5350 17978
rect 5362 17926 5414 17978
rect 5426 17926 5478 17978
rect 13611 17926 13663 17978
rect 13675 17926 13727 17978
rect 13739 17926 13791 17978
rect 13803 17926 13855 17978
rect 13867 17926 13919 17978
rect 22052 17926 22104 17978
rect 22116 17926 22168 17978
rect 22180 17926 22232 17978
rect 22244 17926 22296 17978
rect 22308 17926 22360 17978
rect 30493 17926 30545 17978
rect 30557 17926 30609 17978
rect 30621 17926 30673 17978
rect 30685 17926 30737 17978
rect 30749 17926 30801 17978
rect 6736 17824 6788 17876
rect 27988 17867 28040 17876
rect 27988 17833 27997 17867
rect 27997 17833 28031 17867
rect 28031 17833 28040 17867
rect 27988 17824 28040 17833
rect 29276 17824 29328 17876
rect 3516 17756 3568 17808
rect 11336 17688 11388 17740
rect 12072 17688 12124 17740
rect 27620 17731 27672 17740
rect 3240 17663 3292 17672
rect 3240 17629 3249 17663
rect 3249 17629 3283 17663
rect 3283 17629 3292 17663
rect 3240 17620 3292 17629
rect 6368 17663 6420 17672
rect 6368 17629 6377 17663
rect 6377 17629 6411 17663
rect 6411 17629 6420 17663
rect 6368 17620 6420 17629
rect 6552 17663 6604 17672
rect 6552 17629 6561 17663
rect 6561 17629 6595 17663
rect 6595 17629 6604 17663
rect 6552 17620 6604 17629
rect 27620 17697 27629 17731
rect 27629 17697 27663 17731
rect 27663 17697 27672 17731
rect 27620 17688 27672 17697
rect 29460 17756 29512 17808
rect 13544 17620 13596 17672
rect 16948 17663 17000 17672
rect 16948 17629 16957 17663
rect 16957 17629 16991 17663
rect 16991 17629 17000 17663
rect 16948 17620 17000 17629
rect 18696 17620 18748 17672
rect 20536 17620 20588 17672
rect 25228 17663 25280 17672
rect 25228 17629 25237 17663
rect 25237 17629 25271 17663
rect 25271 17629 25280 17663
rect 25228 17620 25280 17629
rect 25688 17620 25740 17672
rect 28540 17663 28592 17672
rect 2688 17552 2740 17604
rect 12164 17552 12216 17604
rect 12900 17552 12952 17604
rect 3056 17527 3108 17536
rect 3056 17493 3065 17527
rect 3065 17493 3099 17527
rect 3099 17493 3108 17527
rect 3056 17484 3108 17493
rect 3148 17527 3200 17536
rect 3148 17493 3157 17527
rect 3157 17493 3191 17527
rect 3191 17493 3200 17527
rect 3148 17484 3200 17493
rect 10968 17484 11020 17536
rect 12992 17484 13044 17536
rect 24492 17552 24544 17604
rect 28540 17629 28549 17663
rect 28549 17629 28583 17663
rect 28583 17629 28592 17663
rect 28540 17620 28592 17629
rect 29276 17620 29328 17672
rect 30932 17663 30984 17672
rect 30932 17629 30941 17663
rect 30941 17629 30975 17663
rect 30975 17629 30984 17663
rect 32312 17756 32364 17808
rect 30932 17620 30984 17629
rect 32588 17663 32640 17672
rect 32588 17629 32597 17663
rect 32597 17629 32631 17663
rect 32631 17629 32640 17663
rect 32588 17620 32640 17629
rect 33416 17663 33468 17672
rect 33416 17629 33425 17663
rect 33425 17629 33459 17663
rect 33459 17629 33468 17663
rect 33416 17620 33468 17629
rect 26148 17552 26200 17604
rect 27804 17552 27856 17604
rect 29184 17552 29236 17604
rect 29828 17552 29880 17604
rect 31116 17595 31168 17604
rect 31116 17561 31125 17595
rect 31125 17561 31159 17595
rect 31159 17561 31168 17595
rect 31116 17552 31168 17561
rect 21088 17484 21140 17536
rect 9390 17382 9442 17434
rect 9454 17382 9506 17434
rect 9518 17382 9570 17434
rect 9582 17382 9634 17434
rect 9646 17382 9698 17434
rect 17831 17382 17883 17434
rect 17895 17382 17947 17434
rect 17959 17382 18011 17434
rect 18023 17382 18075 17434
rect 18087 17382 18139 17434
rect 26272 17382 26324 17434
rect 26336 17382 26388 17434
rect 26400 17382 26452 17434
rect 26464 17382 26516 17434
rect 26528 17382 26580 17434
rect 34713 17382 34765 17434
rect 34777 17382 34829 17434
rect 34841 17382 34893 17434
rect 34905 17382 34957 17434
rect 34969 17382 35021 17434
rect 6920 17280 6972 17332
rect 2964 17255 3016 17264
rect 2964 17221 2973 17255
rect 2973 17221 3007 17255
rect 3007 17221 3016 17255
rect 2964 17212 3016 17221
rect 4252 17144 4304 17196
rect 6736 17187 6788 17196
rect 6736 17153 6745 17187
rect 6745 17153 6779 17187
rect 6779 17153 6788 17187
rect 6736 17144 6788 17153
rect 6828 17144 6880 17196
rect 7472 17144 7524 17196
rect 7748 17144 7800 17196
rect 8852 17212 8904 17264
rect 10324 17280 10376 17332
rect 14464 17280 14516 17332
rect 25136 17280 25188 17332
rect 25688 17323 25740 17332
rect 25688 17289 25697 17323
rect 25697 17289 25731 17323
rect 25731 17289 25740 17323
rect 25688 17280 25740 17289
rect 29828 17323 29880 17332
rect 29828 17289 29837 17323
rect 29837 17289 29871 17323
rect 29871 17289 29880 17323
rect 29828 17280 29880 17289
rect 30012 17280 30064 17332
rect 30932 17323 30984 17332
rect 30932 17289 30941 17323
rect 30941 17289 30975 17323
rect 30975 17289 30984 17323
rect 30932 17280 30984 17289
rect 12256 17212 12308 17264
rect 13360 17212 13412 17264
rect 9864 17187 9916 17196
rect 9864 17153 9873 17187
rect 9873 17153 9907 17187
rect 9907 17153 9916 17187
rect 9864 17144 9916 17153
rect 13544 17187 13596 17196
rect 13544 17153 13553 17187
rect 13553 17153 13587 17187
rect 13587 17153 13596 17187
rect 16212 17187 16264 17196
rect 13544 17144 13596 17153
rect 16212 17153 16221 17187
rect 16221 17153 16255 17187
rect 16255 17153 16264 17187
rect 16212 17144 16264 17153
rect 19432 17144 19484 17196
rect 20720 17144 20772 17196
rect 21732 17212 21784 17264
rect 24584 17212 24636 17264
rect 23756 17144 23808 17196
rect 25964 17212 26016 17264
rect 31668 17280 31720 17332
rect 32864 17280 32916 17332
rect 33416 17280 33468 17332
rect 25044 17187 25096 17196
rect 25044 17153 25053 17187
rect 25053 17153 25087 17187
rect 25087 17153 25096 17187
rect 25044 17144 25096 17153
rect 2688 17119 2740 17128
rect 2688 17085 2697 17119
rect 2697 17085 2731 17119
rect 2731 17085 2740 17119
rect 2688 17076 2740 17085
rect 6644 17119 6696 17128
rect 6644 17085 6653 17119
rect 6653 17085 6687 17119
rect 6687 17085 6696 17119
rect 6644 17076 6696 17085
rect 9772 17119 9824 17128
rect 9772 17085 9781 17119
rect 9781 17085 9815 17119
rect 9815 17085 9824 17119
rect 9772 17076 9824 17085
rect 16304 17076 16356 17128
rect 18696 17076 18748 17128
rect 22560 17076 22612 17128
rect 23112 17119 23164 17128
rect 23112 17085 23121 17119
rect 23121 17085 23155 17119
rect 23155 17085 23164 17119
rect 23112 17076 23164 17085
rect 25504 17187 25556 17196
rect 25504 17153 25518 17187
rect 25518 17153 25552 17187
rect 25552 17153 25556 17187
rect 25504 17144 25556 17153
rect 30288 17076 30340 17128
rect 31300 17144 31352 17196
rect 8208 16983 8260 16992
rect 8208 16949 8217 16983
rect 8217 16949 8251 16983
rect 8251 16949 8260 16983
rect 8208 16940 8260 16949
rect 8300 16940 8352 16992
rect 10048 16983 10100 16992
rect 10048 16949 10057 16983
rect 10057 16949 10091 16983
rect 10091 16949 10100 16983
rect 10048 16940 10100 16949
rect 11152 16940 11204 16992
rect 19800 16940 19852 16992
rect 22376 16940 22428 16992
rect 23296 16940 23348 16992
rect 30012 17008 30064 17060
rect 32588 17144 32640 17196
rect 32588 16940 32640 16992
rect 5170 16838 5222 16890
rect 5234 16838 5286 16890
rect 5298 16838 5350 16890
rect 5362 16838 5414 16890
rect 5426 16838 5478 16890
rect 13611 16838 13663 16890
rect 13675 16838 13727 16890
rect 13739 16838 13791 16890
rect 13803 16838 13855 16890
rect 13867 16838 13919 16890
rect 22052 16838 22104 16890
rect 22116 16838 22168 16890
rect 22180 16838 22232 16890
rect 22244 16838 22296 16890
rect 22308 16838 22360 16890
rect 30493 16838 30545 16890
rect 30557 16838 30609 16890
rect 30621 16838 30673 16890
rect 30685 16838 30737 16890
rect 30749 16838 30801 16890
rect 2688 16736 2740 16788
rect 3240 16779 3292 16788
rect 3240 16745 3249 16779
rect 3249 16745 3283 16779
rect 3283 16745 3292 16779
rect 3240 16736 3292 16745
rect 4252 16779 4304 16788
rect 4252 16745 4261 16779
rect 4261 16745 4295 16779
rect 4295 16745 4304 16779
rect 4252 16736 4304 16745
rect 6276 16736 6328 16788
rect 6920 16736 6972 16788
rect 7196 16711 7248 16720
rect 7196 16677 7205 16711
rect 7205 16677 7239 16711
rect 7239 16677 7248 16711
rect 7196 16668 7248 16677
rect 8208 16736 8260 16788
rect 12256 16779 12308 16788
rect 12256 16745 12265 16779
rect 12265 16745 12299 16779
rect 12299 16745 12308 16779
rect 12256 16736 12308 16745
rect 19432 16779 19484 16788
rect 19432 16745 19441 16779
rect 19441 16745 19475 16779
rect 19475 16745 19484 16779
rect 19432 16736 19484 16745
rect 10968 16668 11020 16720
rect 15200 16668 15252 16720
rect 16304 16668 16356 16720
rect 22376 16736 22428 16788
rect 25780 16736 25832 16788
rect 31116 16736 31168 16788
rect 31668 16736 31720 16788
rect 6552 16600 6604 16652
rect 4068 16575 4120 16584
rect 4068 16541 4077 16575
rect 4077 16541 4111 16575
rect 4111 16541 4120 16575
rect 4068 16532 4120 16541
rect 4344 16575 4396 16584
rect 4344 16541 4353 16575
rect 4353 16541 4387 16575
rect 4387 16541 4396 16575
rect 4344 16532 4396 16541
rect 6460 16532 6512 16584
rect 11980 16600 12032 16652
rect 9956 16532 10008 16584
rect 10048 16575 10100 16584
rect 10048 16541 10057 16575
rect 10057 16541 10091 16575
rect 10091 16541 10100 16575
rect 14740 16600 14792 16652
rect 19984 16600 20036 16652
rect 10048 16532 10100 16541
rect 12440 16575 12492 16584
rect 12440 16541 12449 16575
rect 12449 16541 12483 16575
rect 12483 16541 12492 16575
rect 12440 16532 12492 16541
rect 3056 16464 3108 16516
rect 6552 16464 6604 16516
rect 11152 16464 11204 16516
rect 15292 16464 15344 16516
rect 15844 16532 15896 16584
rect 17224 16575 17276 16584
rect 17224 16541 17233 16575
rect 17233 16541 17267 16575
rect 17267 16541 17276 16575
rect 17224 16532 17276 16541
rect 19800 16575 19852 16584
rect 16120 16464 16172 16516
rect 16304 16464 16356 16516
rect 17316 16464 17368 16516
rect 19800 16541 19809 16575
rect 19809 16541 19843 16575
rect 19843 16541 19852 16575
rect 19800 16532 19852 16541
rect 19892 16575 19944 16584
rect 19892 16541 19901 16575
rect 19901 16541 19935 16575
rect 19935 16541 19944 16575
rect 24584 16575 24636 16584
rect 19892 16532 19944 16541
rect 24584 16541 24593 16575
rect 24593 16541 24627 16575
rect 24627 16541 24636 16575
rect 24584 16532 24636 16541
rect 24676 16532 24728 16584
rect 29092 16532 29144 16584
rect 30012 16575 30064 16584
rect 30012 16541 30021 16575
rect 30021 16541 30055 16575
rect 30055 16541 30064 16575
rect 30012 16532 30064 16541
rect 30104 16532 30156 16584
rect 32220 16600 32272 16652
rect 32496 16600 32548 16652
rect 20720 16464 20772 16516
rect 20996 16507 21048 16516
rect 20996 16473 21030 16507
rect 21030 16473 21048 16507
rect 20996 16464 21048 16473
rect 25872 16464 25924 16516
rect 26148 16464 26200 16516
rect 29736 16507 29788 16516
rect 29736 16473 29745 16507
rect 29745 16473 29779 16507
rect 29779 16473 29788 16507
rect 29736 16464 29788 16473
rect 30380 16464 30432 16516
rect 31300 16464 31352 16516
rect 6368 16396 6420 16448
rect 10416 16396 10468 16448
rect 14464 16439 14516 16448
rect 14464 16405 14473 16439
rect 14473 16405 14507 16439
rect 14507 16405 14516 16439
rect 14464 16396 14516 16405
rect 16672 16439 16724 16448
rect 16672 16405 16681 16439
rect 16681 16405 16715 16439
rect 16715 16405 16724 16439
rect 16672 16396 16724 16405
rect 17500 16396 17552 16448
rect 19892 16396 19944 16448
rect 20904 16396 20956 16448
rect 26056 16396 26108 16448
rect 30104 16439 30156 16448
rect 30104 16405 30113 16439
rect 30113 16405 30147 16439
rect 30147 16405 30156 16439
rect 30288 16439 30340 16448
rect 30104 16396 30156 16405
rect 30288 16405 30297 16439
rect 30297 16405 30331 16439
rect 30331 16405 30340 16439
rect 30288 16396 30340 16405
rect 32404 16575 32456 16584
rect 32404 16541 32413 16575
rect 32413 16541 32447 16575
rect 32447 16541 32456 16575
rect 32404 16532 32456 16541
rect 9390 16294 9442 16346
rect 9454 16294 9506 16346
rect 9518 16294 9570 16346
rect 9582 16294 9634 16346
rect 9646 16294 9698 16346
rect 17831 16294 17883 16346
rect 17895 16294 17947 16346
rect 17959 16294 18011 16346
rect 18023 16294 18075 16346
rect 18087 16294 18139 16346
rect 26272 16294 26324 16346
rect 26336 16294 26388 16346
rect 26400 16294 26452 16346
rect 26464 16294 26516 16346
rect 26528 16294 26580 16346
rect 34713 16294 34765 16346
rect 34777 16294 34829 16346
rect 34841 16294 34893 16346
rect 34905 16294 34957 16346
rect 34969 16294 35021 16346
rect 6736 16235 6788 16244
rect 6736 16201 6745 16235
rect 6745 16201 6779 16235
rect 6779 16201 6788 16235
rect 6736 16192 6788 16201
rect 12348 16192 12400 16244
rect 13268 16192 13320 16244
rect 18696 16235 18748 16244
rect 5724 16167 5776 16176
rect 5724 16133 5733 16167
rect 5733 16133 5767 16167
rect 5767 16133 5776 16167
rect 5724 16124 5776 16133
rect 6828 16124 6880 16176
rect 11336 16124 11388 16176
rect 13452 16124 13504 16176
rect 15200 16167 15252 16176
rect 15200 16133 15234 16167
rect 15234 16133 15252 16167
rect 15200 16124 15252 16133
rect 6552 16099 6604 16108
rect 6552 16065 6561 16099
rect 6561 16065 6595 16099
rect 6595 16065 6604 16099
rect 6552 16056 6604 16065
rect 6920 16056 6972 16108
rect 7380 16099 7432 16108
rect 7380 16065 7389 16099
rect 7389 16065 7423 16099
rect 7423 16065 7432 16099
rect 7380 16056 7432 16065
rect 7472 16056 7524 16108
rect 10416 16099 10468 16108
rect 10416 16065 10425 16099
rect 10425 16065 10459 16099
rect 10459 16065 10468 16099
rect 10416 16056 10468 16065
rect 10968 16099 11020 16108
rect 10968 16065 10977 16099
rect 10977 16065 11011 16099
rect 11011 16065 11020 16099
rect 10968 16056 11020 16065
rect 11152 16099 11204 16108
rect 11152 16065 11161 16099
rect 11161 16065 11195 16099
rect 11195 16065 11204 16099
rect 11152 16056 11204 16065
rect 7196 15988 7248 16040
rect 5540 15920 5592 15972
rect 6460 15920 6512 15972
rect 14280 16099 14332 16108
rect 14280 16065 14289 16099
rect 14289 16065 14323 16099
rect 14323 16065 14332 16099
rect 14280 16056 14332 16065
rect 16304 16056 16356 16108
rect 17408 16099 17460 16108
rect 17408 16065 17417 16099
rect 17417 16065 17451 16099
rect 17451 16065 17460 16099
rect 17408 16056 17460 16065
rect 17592 16099 17644 16108
rect 17592 16065 17601 16099
rect 17601 16065 17635 16099
rect 17635 16065 17644 16099
rect 17592 16056 17644 16065
rect 18696 16201 18705 16235
rect 18705 16201 18739 16235
rect 18739 16201 18748 16235
rect 18696 16192 18748 16201
rect 22652 16235 22704 16244
rect 19340 16124 19392 16176
rect 20352 16124 20404 16176
rect 20168 16056 20220 16108
rect 20444 16099 20496 16108
rect 20444 16065 20453 16099
rect 20453 16065 20487 16099
rect 20487 16065 20496 16099
rect 20444 16056 20496 16065
rect 14740 15988 14792 16040
rect 19800 15988 19852 16040
rect 21088 16124 21140 16176
rect 22652 16201 22661 16235
rect 22661 16201 22695 16235
rect 22695 16201 22704 16235
rect 22652 16192 22704 16201
rect 25872 16192 25924 16244
rect 21640 16056 21692 16108
rect 22008 16099 22060 16108
rect 22008 16065 22017 16099
rect 22017 16065 22051 16099
rect 22051 16065 22060 16099
rect 22008 16056 22060 16065
rect 26056 16124 26108 16176
rect 32496 16192 32548 16244
rect 33048 16192 33100 16244
rect 20628 15920 20680 15972
rect 22376 16099 22428 16108
rect 22376 16065 22385 16099
rect 22385 16065 22419 16099
rect 22419 16065 22428 16099
rect 22376 16056 22428 16065
rect 22652 16056 22704 16108
rect 25136 16099 25188 16108
rect 25136 16065 25145 16099
rect 25145 16065 25179 16099
rect 25179 16065 25188 16099
rect 25136 16056 25188 16065
rect 25780 16056 25832 16108
rect 30380 16124 30432 16176
rect 28448 16099 28500 16108
rect 24492 15988 24544 16040
rect 28448 16065 28457 16099
rect 28457 16065 28491 16099
rect 28491 16065 28500 16099
rect 28448 16056 28500 16065
rect 29092 16056 29144 16108
rect 27712 15988 27764 16040
rect 27804 15988 27856 16040
rect 28356 16031 28408 16040
rect 28356 15997 28365 16031
rect 28365 15997 28399 16031
rect 28399 15997 28408 16031
rect 29736 16056 29788 16108
rect 33876 16056 33928 16108
rect 28356 15988 28408 15997
rect 7748 15895 7800 15904
rect 7748 15861 7757 15895
rect 7757 15861 7791 15895
rect 7791 15861 7800 15895
rect 7748 15852 7800 15861
rect 14464 15852 14516 15904
rect 20076 15852 20128 15904
rect 22008 15852 22060 15904
rect 24584 15852 24636 15904
rect 25228 15852 25280 15904
rect 30104 15988 30156 16040
rect 32312 16031 32364 16040
rect 32312 15997 32321 16031
rect 32321 15997 32355 16031
rect 32355 15997 32364 16031
rect 32312 15988 32364 15997
rect 5170 15750 5222 15802
rect 5234 15750 5286 15802
rect 5298 15750 5350 15802
rect 5362 15750 5414 15802
rect 5426 15750 5478 15802
rect 13611 15750 13663 15802
rect 13675 15750 13727 15802
rect 13739 15750 13791 15802
rect 13803 15750 13855 15802
rect 13867 15750 13919 15802
rect 22052 15750 22104 15802
rect 22116 15750 22168 15802
rect 22180 15750 22232 15802
rect 22244 15750 22296 15802
rect 22308 15750 22360 15802
rect 30493 15750 30545 15802
rect 30557 15750 30609 15802
rect 30621 15750 30673 15802
rect 30685 15750 30737 15802
rect 30749 15750 30801 15802
rect 4804 15648 4856 15700
rect 7748 15648 7800 15700
rect 19248 15648 19300 15700
rect 19892 15691 19944 15700
rect 19892 15657 19901 15691
rect 19901 15657 19935 15691
rect 19935 15657 19944 15691
rect 19892 15648 19944 15657
rect 25136 15648 25188 15700
rect 26056 15648 26108 15700
rect 28356 15648 28408 15700
rect 31760 15648 31812 15700
rect 32312 15648 32364 15700
rect 33876 15691 33928 15700
rect 33876 15657 33885 15691
rect 33885 15657 33919 15691
rect 33919 15657 33928 15691
rect 33876 15648 33928 15657
rect 18236 15580 18288 15632
rect 22376 15580 22428 15632
rect 32680 15580 32732 15632
rect 4344 15512 4396 15564
rect 6552 15512 6604 15564
rect 13268 15512 13320 15564
rect 4068 15444 4120 15496
rect 6092 15487 6144 15496
rect 6092 15453 6101 15487
rect 6101 15453 6135 15487
rect 6135 15453 6144 15487
rect 6092 15444 6144 15453
rect 6276 15487 6328 15496
rect 6276 15453 6285 15487
rect 6285 15453 6319 15487
rect 6319 15453 6328 15487
rect 6276 15444 6328 15453
rect 6736 15487 6788 15496
rect 6736 15453 6745 15487
rect 6745 15453 6779 15487
rect 6779 15453 6788 15487
rect 6736 15444 6788 15453
rect 9772 15444 9824 15496
rect 16580 15512 16632 15564
rect 17408 15512 17460 15564
rect 17500 15512 17552 15564
rect 21180 15512 21232 15564
rect 22560 15555 22612 15564
rect 22560 15521 22569 15555
rect 22569 15521 22603 15555
rect 22603 15521 22612 15555
rect 22560 15512 22612 15521
rect 29552 15512 29604 15564
rect 2964 15419 3016 15428
rect 2964 15385 2973 15419
rect 2973 15385 3007 15419
rect 3007 15385 3016 15419
rect 2964 15376 3016 15385
rect 5540 15376 5592 15428
rect 4436 15308 4488 15360
rect 7380 15376 7432 15428
rect 16304 15444 16356 15496
rect 18328 15444 18380 15496
rect 20812 15487 20864 15496
rect 20812 15453 20821 15487
rect 20821 15453 20855 15487
rect 20855 15453 20864 15487
rect 20812 15444 20864 15453
rect 23020 15444 23072 15496
rect 23388 15487 23440 15496
rect 23388 15453 23397 15487
rect 23397 15453 23431 15487
rect 23431 15453 23440 15487
rect 23388 15444 23440 15453
rect 24492 15444 24544 15496
rect 30288 15444 30340 15496
rect 33416 15487 33468 15496
rect 33416 15453 33425 15487
rect 33425 15453 33459 15487
rect 33459 15453 33468 15487
rect 33416 15444 33468 15453
rect 15292 15376 15344 15428
rect 17132 15376 17184 15428
rect 17408 15376 17460 15428
rect 17592 15376 17644 15428
rect 20168 15419 20220 15428
rect 20168 15385 20177 15419
rect 20177 15385 20211 15419
rect 20211 15385 20220 15419
rect 20168 15376 20220 15385
rect 20536 15376 20588 15428
rect 24676 15376 24728 15428
rect 25228 15419 25280 15428
rect 25228 15385 25237 15419
rect 25237 15385 25271 15419
rect 25271 15385 25280 15419
rect 25228 15376 25280 15385
rect 25780 15376 25832 15428
rect 29000 15376 29052 15428
rect 33600 15376 33652 15428
rect 6828 15351 6880 15360
rect 6828 15317 6837 15351
rect 6837 15317 6871 15351
rect 6871 15317 6880 15351
rect 6828 15308 6880 15317
rect 16396 15351 16448 15360
rect 16396 15317 16405 15351
rect 16405 15317 16439 15351
rect 16439 15317 16448 15351
rect 16396 15308 16448 15317
rect 17316 15308 17368 15360
rect 17500 15308 17552 15360
rect 20996 15308 21048 15360
rect 22928 15308 22980 15360
rect 23480 15308 23532 15360
rect 25964 15308 26016 15360
rect 33048 15308 33100 15360
rect 9390 15206 9442 15258
rect 9454 15206 9506 15258
rect 9518 15206 9570 15258
rect 9582 15206 9634 15258
rect 9646 15206 9698 15258
rect 17831 15206 17883 15258
rect 17895 15206 17947 15258
rect 17959 15206 18011 15258
rect 18023 15206 18075 15258
rect 18087 15206 18139 15258
rect 26272 15206 26324 15258
rect 26336 15206 26388 15258
rect 26400 15206 26452 15258
rect 26464 15206 26516 15258
rect 26528 15206 26580 15258
rect 34713 15206 34765 15258
rect 34777 15206 34829 15258
rect 34841 15206 34893 15258
rect 34905 15206 34957 15258
rect 34969 15206 35021 15258
rect 5724 15104 5776 15156
rect 18420 15104 18472 15156
rect 2964 15036 3016 15088
rect 6276 15036 6328 15088
rect 11796 15036 11848 15088
rect 16948 15036 17000 15088
rect 17868 15036 17920 15088
rect 21824 15104 21876 15156
rect 22928 15147 22980 15156
rect 22928 15113 22937 15147
rect 22937 15113 22971 15147
rect 22971 15113 22980 15147
rect 22928 15104 22980 15113
rect 23296 15147 23348 15156
rect 23296 15113 23305 15147
rect 23305 15113 23339 15147
rect 23339 15113 23348 15147
rect 23296 15104 23348 15113
rect 23388 15104 23440 15156
rect 25136 15104 25188 15156
rect 29552 15104 29604 15156
rect 33600 15147 33652 15156
rect 33600 15113 33609 15147
rect 33609 15113 33643 15147
rect 33643 15113 33652 15147
rect 33600 15104 33652 15113
rect 19984 15079 20036 15088
rect 1676 14943 1728 14952
rect 1676 14909 1685 14943
rect 1685 14909 1719 14943
rect 1719 14909 1728 14943
rect 1676 14900 1728 14909
rect 2688 14900 2740 14952
rect 3240 14832 3292 14884
rect 4528 14968 4580 15020
rect 9036 15011 9088 15020
rect 9036 14977 9045 15011
rect 9045 14977 9079 15011
rect 9079 14977 9088 15011
rect 9036 14968 9088 14977
rect 9956 14968 10008 15020
rect 10692 15011 10744 15020
rect 8944 14943 8996 14952
rect 8944 14909 8953 14943
rect 8953 14909 8987 14943
rect 8987 14909 8996 14943
rect 8944 14900 8996 14909
rect 9864 14900 9916 14952
rect 10324 14900 10376 14952
rect 10692 14977 10701 15011
rect 10701 14977 10735 15011
rect 10735 14977 10744 15011
rect 10692 14968 10744 14977
rect 12164 14968 12216 15020
rect 16212 14968 16264 15020
rect 16672 14968 16724 15020
rect 19984 15045 19993 15079
rect 19993 15045 20027 15079
rect 20027 15045 20036 15079
rect 19984 15036 20036 15045
rect 18236 15011 18288 15020
rect 12072 14900 12124 14952
rect 18236 14977 18245 15011
rect 18245 14977 18279 15011
rect 18279 14977 18288 15011
rect 18236 14968 18288 14977
rect 18512 14968 18564 15020
rect 19800 14968 19852 15020
rect 17224 14900 17276 14952
rect 19892 14900 19944 14952
rect 13452 14832 13504 14884
rect 15108 14832 15160 14884
rect 22192 15011 22244 15020
rect 22192 14977 22201 15011
rect 22201 14977 22235 15011
rect 22235 14977 22244 15011
rect 22192 14968 22244 14977
rect 22376 15011 22428 15020
rect 22376 14977 22385 15011
rect 22385 14977 22419 15011
rect 22419 14977 22428 15011
rect 22376 14968 22428 14977
rect 22468 15011 22520 15020
rect 22468 14977 22477 15011
rect 22477 14977 22511 15011
rect 22511 14977 22520 15011
rect 22468 14968 22520 14977
rect 23020 14968 23072 15020
rect 26148 15036 26200 15088
rect 25044 15011 25096 15020
rect 25044 14977 25062 15011
rect 25062 14977 25096 15011
rect 25044 14968 25096 14977
rect 30012 14968 30064 15020
rect 20720 14943 20772 14952
rect 20720 14909 20729 14943
rect 20729 14909 20763 14943
rect 20763 14909 20772 14943
rect 20720 14900 20772 14909
rect 21916 14900 21968 14952
rect 26424 14900 26476 14952
rect 29644 14832 29696 14884
rect 2964 14764 3016 14816
rect 6092 14764 6144 14816
rect 9956 14764 10008 14816
rect 10692 14764 10744 14816
rect 19892 14764 19944 14816
rect 23664 14764 23716 14816
rect 5170 14662 5222 14714
rect 5234 14662 5286 14714
rect 5298 14662 5350 14714
rect 5362 14662 5414 14714
rect 5426 14662 5478 14714
rect 13611 14662 13663 14714
rect 13675 14662 13727 14714
rect 13739 14662 13791 14714
rect 13803 14662 13855 14714
rect 13867 14662 13919 14714
rect 22052 14662 22104 14714
rect 22116 14662 22168 14714
rect 22180 14662 22232 14714
rect 22244 14662 22296 14714
rect 22308 14662 22360 14714
rect 30493 14662 30545 14714
rect 30557 14662 30609 14714
rect 30621 14662 30673 14714
rect 30685 14662 30737 14714
rect 30749 14662 30801 14714
rect 6828 14560 6880 14612
rect 1400 14424 1452 14476
rect 6276 14492 6328 14544
rect 7380 14560 7432 14612
rect 14372 14603 14424 14612
rect 14372 14569 14381 14603
rect 14381 14569 14415 14603
rect 14415 14569 14424 14603
rect 14372 14560 14424 14569
rect 8668 14492 8720 14544
rect 9220 14535 9272 14544
rect 9220 14501 9229 14535
rect 9229 14501 9263 14535
rect 9263 14501 9272 14535
rect 9220 14492 9272 14501
rect 2688 14399 2740 14408
rect 2688 14365 2697 14399
rect 2697 14365 2731 14399
rect 2731 14365 2740 14399
rect 2688 14356 2740 14365
rect 3056 14356 3108 14408
rect 6276 14356 6328 14408
rect 3148 14288 3200 14340
rect 5724 14288 5776 14340
rect 6460 14288 6512 14340
rect 7932 14331 7984 14340
rect 7932 14297 7941 14331
rect 7941 14297 7975 14331
rect 7975 14297 7984 14331
rect 9588 14356 9640 14408
rect 7932 14288 7984 14297
rect 6920 14220 6972 14272
rect 7196 14263 7248 14272
rect 7196 14229 7221 14263
rect 7221 14229 7248 14263
rect 7196 14220 7248 14229
rect 7748 14220 7800 14272
rect 7840 14220 7892 14272
rect 8300 14288 8352 14340
rect 10232 14356 10284 14408
rect 11980 14356 12032 14408
rect 18512 14467 18564 14476
rect 18512 14433 18521 14467
rect 18521 14433 18555 14467
rect 18555 14433 18564 14467
rect 18512 14424 18564 14433
rect 19984 14560 20036 14612
rect 21732 14560 21784 14612
rect 23664 14560 23716 14612
rect 9956 14288 10008 14340
rect 11704 14288 11756 14340
rect 12440 14288 12492 14340
rect 13084 14331 13136 14340
rect 13084 14297 13093 14331
rect 13093 14297 13127 14331
rect 13127 14297 13136 14331
rect 13084 14288 13136 14297
rect 17408 14356 17460 14408
rect 17868 14356 17920 14408
rect 21640 14399 21692 14408
rect 21640 14365 21649 14399
rect 21649 14365 21683 14399
rect 21683 14365 21692 14399
rect 21640 14356 21692 14365
rect 21732 14399 21784 14408
rect 21732 14365 21741 14399
rect 21741 14365 21775 14399
rect 21775 14365 21784 14399
rect 22100 14492 22152 14544
rect 25228 14560 25280 14612
rect 25964 14603 26016 14612
rect 25964 14569 25973 14603
rect 25973 14569 26007 14603
rect 26007 14569 26016 14603
rect 25964 14560 26016 14569
rect 26700 14560 26752 14612
rect 21732 14356 21784 14365
rect 22376 14356 22428 14408
rect 19892 14331 19944 14340
rect 9864 14220 9916 14272
rect 19892 14297 19926 14331
rect 19926 14297 19944 14331
rect 19892 14288 19944 14297
rect 20628 14288 20680 14340
rect 21824 14331 21876 14340
rect 20812 14220 20864 14272
rect 21824 14297 21833 14331
rect 21833 14297 21867 14331
rect 21867 14297 21876 14331
rect 23756 14424 23808 14476
rect 24584 14467 24636 14476
rect 24584 14433 24593 14467
rect 24593 14433 24627 14467
rect 24627 14433 24636 14467
rect 24584 14424 24636 14433
rect 23480 14356 23532 14408
rect 26424 14399 26476 14408
rect 26424 14365 26433 14399
rect 26433 14365 26467 14399
rect 26467 14365 26476 14399
rect 26424 14356 26476 14365
rect 26976 14356 27028 14408
rect 27712 14356 27764 14408
rect 28632 14356 28684 14408
rect 32496 14560 32548 14612
rect 31760 14424 31812 14476
rect 32312 14424 32364 14476
rect 30104 14356 30156 14408
rect 32128 14399 32180 14408
rect 32128 14365 32137 14399
rect 32137 14365 32171 14399
rect 32171 14365 32180 14399
rect 32128 14356 32180 14365
rect 23572 14331 23624 14340
rect 21824 14288 21876 14297
rect 23572 14297 23581 14331
rect 23581 14297 23615 14331
rect 23615 14297 23624 14331
rect 23572 14288 23624 14297
rect 26700 14331 26752 14340
rect 26700 14297 26734 14331
rect 26734 14297 26752 14331
rect 26700 14288 26752 14297
rect 27620 14288 27672 14340
rect 29092 14288 29144 14340
rect 29736 14331 29788 14340
rect 29736 14297 29745 14331
rect 29745 14297 29779 14331
rect 29779 14297 29788 14331
rect 29736 14288 29788 14297
rect 24032 14220 24084 14272
rect 27712 14220 27764 14272
rect 29000 14220 29052 14272
rect 29920 14220 29972 14272
rect 31300 14220 31352 14272
rect 33048 14220 33100 14272
rect 9390 14118 9442 14170
rect 9454 14118 9506 14170
rect 9518 14118 9570 14170
rect 9582 14118 9634 14170
rect 9646 14118 9698 14170
rect 17831 14118 17883 14170
rect 17895 14118 17947 14170
rect 17959 14118 18011 14170
rect 18023 14118 18075 14170
rect 18087 14118 18139 14170
rect 26272 14118 26324 14170
rect 26336 14118 26388 14170
rect 26400 14118 26452 14170
rect 26464 14118 26516 14170
rect 26528 14118 26580 14170
rect 34713 14118 34765 14170
rect 34777 14118 34829 14170
rect 34841 14118 34893 14170
rect 34905 14118 34957 14170
rect 34969 14118 35021 14170
rect 1676 14016 1728 14068
rect 3148 14016 3200 14068
rect 4436 13991 4488 14000
rect 4436 13957 4445 13991
rect 4445 13957 4479 13991
rect 4479 13957 4488 13991
rect 4436 13948 4488 13957
rect 3056 13880 3108 13932
rect 5540 13880 5592 13932
rect 7932 14016 7984 14068
rect 8300 14059 8352 14068
rect 8300 14025 8309 14059
rect 8309 14025 8343 14059
rect 8343 14025 8352 14059
rect 8300 14016 8352 14025
rect 6460 13948 6512 14000
rect 7196 13948 7248 14000
rect 7472 13948 7524 14000
rect 9312 13948 9364 14000
rect 9864 13948 9916 14000
rect 11060 14016 11112 14068
rect 11796 14016 11848 14068
rect 8392 13880 8444 13932
rect 11980 13948 12032 14000
rect 22376 14016 22428 14068
rect 23664 14016 23716 14068
rect 25044 14059 25096 14068
rect 25044 14025 25053 14059
rect 25053 14025 25087 14059
rect 25087 14025 25096 14059
rect 25044 14016 25096 14025
rect 27804 14016 27856 14068
rect 30012 14016 30064 14068
rect 30104 14059 30156 14068
rect 30104 14025 30113 14059
rect 30113 14025 30147 14059
rect 30147 14025 30156 14059
rect 30104 14016 30156 14025
rect 32588 14016 32640 14068
rect 13084 13948 13136 14000
rect 16672 13948 16724 14000
rect 4160 13855 4212 13864
rect 4160 13821 4169 13855
rect 4169 13821 4203 13855
rect 4203 13821 4212 13855
rect 4160 13812 4212 13821
rect 4068 13744 4120 13796
rect 5080 13812 5132 13864
rect 11704 13880 11756 13932
rect 14004 13880 14056 13932
rect 14556 13880 14608 13932
rect 15200 13923 15252 13932
rect 15200 13889 15209 13923
rect 15209 13889 15243 13923
rect 15243 13889 15252 13923
rect 15200 13880 15252 13889
rect 15568 13923 15620 13932
rect 15568 13889 15577 13923
rect 15577 13889 15611 13923
rect 15611 13889 15620 13923
rect 15568 13880 15620 13889
rect 17592 13948 17644 14000
rect 19524 13948 19576 14000
rect 19616 13991 19668 14000
rect 19616 13957 19625 13991
rect 19625 13957 19659 13991
rect 19659 13957 19668 13991
rect 19616 13948 19668 13957
rect 21824 13948 21876 14000
rect 27620 13991 27672 14000
rect 27620 13957 27629 13991
rect 27629 13957 27663 13991
rect 27663 13957 27672 13991
rect 28724 13991 28776 14000
rect 27620 13948 27672 13957
rect 28724 13957 28733 13991
rect 28733 13957 28767 13991
rect 28767 13957 28776 13991
rect 28724 13948 28776 13957
rect 17316 13923 17368 13932
rect 17316 13889 17325 13923
rect 17325 13889 17359 13923
rect 17359 13889 17368 13923
rect 17316 13880 17368 13889
rect 20536 13923 20588 13932
rect 20536 13889 20545 13923
rect 20545 13889 20579 13923
rect 20579 13889 20588 13923
rect 20536 13880 20588 13889
rect 21640 13880 21692 13932
rect 24032 13880 24084 13932
rect 24492 13880 24544 13932
rect 11796 13855 11848 13864
rect 11796 13821 11805 13855
rect 11805 13821 11839 13855
rect 11839 13821 11848 13855
rect 11796 13812 11848 13821
rect 17684 13812 17736 13864
rect 16212 13744 16264 13796
rect 6828 13676 6880 13728
rect 10140 13719 10192 13728
rect 10140 13685 10149 13719
rect 10149 13685 10183 13719
rect 10183 13685 10192 13719
rect 10140 13676 10192 13685
rect 19524 13676 19576 13728
rect 20720 13744 20772 13796
rect 24676 13744 24728 13796
rect 25044 13880 25096 13932
rect 26700 13812 26752 13864
rect 27804 13880 27856 13932
rect 29644 13923 29696 13932
rect 29644 13889 29653 13923
rect 29653 13889 29687 13923
rect 29687 13889 29696 13923
rect 29644 13880 29696 13889
rect 29736 13923 29788 13932
rect 29736 13889 29745 13923
rect 29745 13889 29779 13923
rect 29779 13889 29788 13923
rect 29736 13880 29788 13889
rect 29920 13923 29972 13932
rect 29920 13889 29929 13923
rect 29929 13889 29963 13923
rect 29963 13889 29972 13923
rect 29920 13880 29972 13889
rect 30288 13812 30340 13864
rect 19800 13719 19852 13728
rect 19800 13685 19809 13719
rect 19809 13685 19843 13719
rect 19843 13685 19852 13719
rect 19800 13676 19852 13685
rect 28540 13676 28592 13728
rect 29460 13676 29512 13728
rect 32312 13855 32364 13864
rect 32312 13821 32321 13855
rect 32321 13821 32355 13855
rect 32355 13821 32364 13855
rect 32312 13812 32364 13821
rect 33416 13676 33468 13728
rect 5170 13574 5222 13626
rect 5234 13574 5286 13626
rect 5298 13574 5350 13626
rect 5362 13574 5414 13626
rect 5426 13574 5478 13626
rect 13611 13574 13663 13626
rect 13675 13574 13727 13626
rect 13739 13574 13791 13626
rect 13803 13574 13855 13626
rect 13867 13574 13919 13626
rect 22052 13574 22104 13626
rect 22116 13574 22168 13626
rect 22180 13574 22232 13626
rect 22244 13574 22296 13626
rect 22308 13574 22360 13626
rect 30493 13574 30545 13626
rect 30557 13574 30609 13626
rect 30621 13574 30673 13626
rect 30685 13574 30737 13626
rect 30749 13574 30801 13626
rect 4160 13472 4212 13524
rect 5540 13472 5592 13524
rect 12808 13472 12860 13524
rect 13268 13472 13320 13524
rect 14280 13472 14332 13524
rect 17316 13472 17368 13524
rect 26976 13472 27028 13524
rect 32312 13472 32364 13524
rect 2964 13311 3016 13320
rect 2964 13277 2973 13311
rect 2973 13277 3007 13311
rect 3007 13277 3016 13311
rect 2964 13268 3016 13277
rect 2412 13175 2464 13184
rect 2412 13141 2421 13175
rect 2421 13141 2455 13175
rect 2455 13141 2464 13175
rect 2412 13132 2464 13141
rect 3884 13268 3936 13320
rect 4344 13336 4396 13388
rect 5080 13268 5132 13320
rect 7748 13336 7800 13388
rect 9128 13379 9180 13388
rect 9128 13345 9137 13379
rect 9137 13345 9171 13379
rect 9171 13345 9180 13379
rect 11796 13379 11848 13388
rect 9128 13336 9180 13345
rect 11796 13345 11805 13379
rect 11805 13345 11839 13379
rect 11839 13345 11848 13379
rect 11796 13336 11848 13345
rect 12072 13379 12124 13388
rect 12072 13345 12081 13379
rect 12081 13345 12115 13379
rect 12115 13345 12124 13379
rect 12072 13336 12124 13345
rect 12808 13336 12860 13388
rect 15568 13336 15620 13388
rect 8300 13311 8352 13320
rect 8300 13277 8309 13311
rect 8309 13277 8343 13311
rect 8343 13277 8352 13311
rect 8300 13268 8352 13277
rect 3424 13200 3476 13252
rect 14004 13268 14056 13320
rect 8484 13200 8536 13252
rect 8668 13200 8720 13252
rect 10140 13200 10192 13252
rect 14372 13200 14424 13252
rect 14556 13200 14608 13252
rect 15752 13268 15804 13320
rect 18328 13404 18380 13456
rect 21640 13336 21692 13388
rect 18328 13311 18380 13320
rect 18328 13277 18337 13311
rect 18337 13277 18371 13311
rect 18371 13277 18380 13311
rect 18328 13268 18380 13277
rect 19800 13268 19852 13320
rect 26056 13311 26108 13320
rect 26056 13277 26065 13311
rect 26065 13277 26099 13311
rect 26099 13277 26108 13311
rect 26056 13268 26108 13277
rect 33600 13268 33652 13320
rect 4436 13132 4488 13184
rect 7380 13132 7432 13184
rect 9036 13132 9088 13184
rect 12808 13132 12860 13184
rect 13084 13132 13136 13184
rect 15200 13132 15252 13184
rect 18236 13132 18288 13184
rect 9390 13030 9442 13082
rect 9454 13030 9506 13082
rect 9518 13030 9570 13082
rect 9582 13030 9634 13082
rect 9646 13030 9698 13082
rect 17831 13030 17883 13082
rect 17895 13030 17947 13082
rect 17959 13030 18011 13082
rect 18023 13030 18075 13082
rect 18087 13030 18139 13082
rect 26272 13030 26324 13082
rect 26336 13030 26388 13082
rect 26400 13030 26452 13082
rect 26464 13030 26516 13082
rect 26528 13030 26580 13082
rect 34713 13030 34765 13082
rect 34777 13030 34829 13082
rect 34841 13030 34893 13082
rect 34905 13030 34957 13082
rect 34969 13030 35021 13082
rect 4344 12928 4396 12980
rect 4436 12971 4488 12980
rect 4436 12937 4445 12971
rect 4445 12937 4479 12971
rect 4479 12937 4488 12971
rect 20444 12971 20496 12980
rect 4436 12928 4488 12937
rect 20444 12937 20453 12971
rect 20453 12937 20487 12971
rect 20487 12937 20496 12971
rect 20444 12928 20496 12937
rect 2412 12903 2464 12912
rect 2412 12869 2421 12903
rect 2421 12869 2455 12903
rect 2455 12869 2464 12903
rect 2412 12860 2464 12869
rect 3148 12860 3200 12912
rect 8484 12860 8536 12912
rect 9220 12860 9272 12912
rect 12992 12903 13044 12912
rect 12992 12869 13001 12903
rect 13001 12869 13035 12903
rect 13035 12869 13044 12903
rect 12992 12860 13044 12869
rect 14740 12903 14792 12912
rect 14740 12869 14749 12903
rect 14749 12869 14783 12903
rect 14783 12869 14792 12903
rect 14740 12860 14792 12869
rect 3056 12724 3108 12776
rect 3976 12792 4028 12844
rect 4528 12835 4580 12844
rect 4528 12801 4537 12835
rect 4537 12801 4571 12835
rect 4571 12801 4580 12835
rect 4528 12792 4580 12801
rect 15108 12792 15160 12844
rect 16948 12835 17000 12844
rect 3884 12767 3936 12776
rect 3884 12733 3893 12767
rect 3893 12733 3927 12767
rect 3927 12733 3936 12767
rect 3884 12724 3936 12733
rect 9128 12724 9180 12776
rect 14556 12724 14608 12776
rect 16948 12801 16957 12835
rect 16957 12801 16991 12835
rect 16991 12801 17000 12835
rect 16948 12792 17000 12801
rect 17408 12792 17460 12844
rect 22652 12860 22704 12912
rect 18328 12792 18380 12844
rect 16580 12724 16632 12776
rect 19616 12724 19668 12776
rect 20720 12835 20772 12844
rect 20720 12801 20729 12835
rect 20729 12801 20763 12835
rect 20763 12801 20772 12835
rect 20904 12835 20956 12844
rect 20720 12792 20772 12801
rect 20904 12801 20913 12835
rect 20913 12801 20947 12835
rect 20947 12801 20956 12835
rect 20904 12792 20956 12801
rect 20996 12835 21048 12844
rect 20996 12801 21005 12835
rect 21005 12801 21039 12835
rect 21039 12801 21048 12835
rect 20996 12792 21048 12801
rect 26608 12792 26660 12844
rect 27712 12928 27764 12980
rect 28356 12928 28408 12980
rect 32128 12928 32180 12980
rect 33048 12928 33100 12980
rect 27804 12860 27856 12912
rect 28448 12860 28500 12912
rect 24032 12724 24084 12776
rect 25504 12724 25556 12776
rect 17408 12656 17460 12708
rect 20536 12656 20588 12708
rect 29000 12724 29052 12776
rect 29644 12792 29696 12844
rect 32496 12835 32548 12844
rect 32496 12801 32505 12835
rect 32505 12801 32539 12835
rect 32539 12801 32548 12835
rect 32496 12792 32548 12801
rect 33416 12792 33468 12844
rect 30196 12724 30248 12776
rect 27896 12656 27948 12708
rect 30380 12656 30432 12708
rect 7472 12588 7524 12640
rect 14556 12588 14608 12640
rect 17500 12588 17552 12640
rect 21364 12588 21416 12640
rect 21456 12588 21508 12640
rect 25044 12588 25096 12640
rect 28356 12631 28408 12640
rect 28356 12597 28365 12631
rect 28365 12597 28399 12631
rect 28399 12597 28408 12631
rect 28356 12588 28408 12597
rect 5170 12486 5222 12538
rect 5234 12486 5286 12538
rect 5298 12486 5350 12538
rect 5362 12486 5414 12538
rect 5426 12486 5478 12538
rect 13611 12486 13663 12538
rect 13675 12486 13727 12538
rect 13739 12486 13791 12538
rect 13803 12486 13855 12538
rect 13867 12486 13919 12538
rect 22052 12486 22104 12538
rect 22116 12486 22168 12538
rect 22180 12486 22232 12538
rect 22244 12486 22296 12538
rect 22308 12486 22360 12538
rect 30493 12486 30545 12538
rect 30557 12486 30609 12538
rect 30621 12486 30673 12538
rect 30685 12486 30737 12538
rect 30749 12486 30801 12538
rect 3148 12427 3200 12436
rect 3148 12393 3157 12427
rect 3157 12393 3191 12427
rect 3191 12393 3200 12427
rect 3148 12384 3200 12393
rect 14004 12384 14056 12436
rect 15108 12384 15160 12436
rect 4344 12248 4396 12300
rect 16948 12316 17000 12368
rect 20904 12316 20956 12368
rect 3424 12180 3476 12232
rect 14556 12223 14608 12232
rect 14556 12189 14565 12223
rect 14565 12189 14599 12223
rect 14599 12189 14608 12223
rect 14556 12180 14608 12189
rect 15108 12180 15160 12232
rect 15752 12180 15804 12232
rect 16304 12180 16356 12232
rect 17592 12223 17644 12232
rect 17592 12189 17601 12223
rect 17601 12189 17635 12223
rect 17635 12189 17644 12223
rect 17592 12180 17644 12189
rect 18328 12248 18380 12300
rect 22560 12291 22612 12300
rect 22560 12257 22569 12291
rect 22569 12257 22603 12291
rect 22603 12257 22612 12291
rect 22560 12248 22612 12257
rect 21364 12180 21416 12232
rect 28632 12248 28684 12300
rect 28080 12223 28132 12232
rect 28080 12189 28084 12223
rect 28084 12189 28118 12223
rect 28118 12189 28132 12223
rect 19156 12112 19208 12164
rect 20812 12155 20864 12164
rect 20812 12121 20821 12155
rect 20821 12121 20855 12155
rect 20855 12121 20864 12155
rect 20812 12112 20864 12121
rect 23664 12112 23716 12164
rect 24492 12112 24544 12164
rect 28080 12180 28132 12189
rect 28448 12223 28500 12232
rect 28448 12189 28456 12223
rect 28456 12189 28490 12223
rect 28490 12189 28500 12223
rect 28448 12180 28500 12189
rect 28540 12223 28592 12232
rect 28540 12189 28549 12223
rect 28549 12189 28583 12223
rect 28583 12189 28592 12223
rect 28540 12180 28592 12189
rect 17132 12044 17184 12096
rect 17316 12044 17368 12096
rect 24584 12087 24636 12096
rect 24584 12053 24593 12087
rect 24593 12053 24627 12087
rect 24627 12053 24636 12087
rect 24584 12044 24636 12053
rect 24952 12087 25004 12096
rect 24952 12053 24961 12087
rect 24961 12053 24995 12087
rect 24995 12053 25004 12087
rect 24952 12044 25004 12053
rect 28632 12112 28684 12164
rect 31300 12044 31352 12096
rect 9390 11942 9442 11994
rect 9454 11942 9506 11994
rect 9518 11942 9570 11994
rect 9582 11942 9634 11994
rect 9646 11942 9698 11994
rect 17831 11942 17883 11994
rect 17895 11942 17947 11994
rect 17959 11942 18011 11994
rect 18023 11942 18075 11994
rect 18087 11942 18139 11994
rect 26272 11942 26324 11994
rect 26336 11942 26388 11994
rect 26400 11942 26452 11994
rect 26464 11942 26516 11994
rect 26528 11942 26580 11994
rect 34713 11942 34765 11994
rect 34777 11942 34829 11994
rect 34841 11942 34893 11994
rect 34905 11942 34957 11994
rect 34969 11942 35021 11994
rect 15752 11815 15804 11824
rect 15752 11781 15761 11815
rect 15761 11781 15795 11815
rect 15795 11781 15804 11815
rect 15752 11772 15804 11781
rect 15200 11704 15252 11756
rect 16304 11704 16356 11756
rect 16580 11704 16632 11756
rect 18420 11772 18472 11824
rect 20536 11840 20588 11892
rect 20720 11840 20772 11892
rect 22468 11840 22520 11892
rect 28172 11840 28224 11892
rect 28448 11840 28500 11892
rect 31300 11883 31352 11892
rect 31300 11849 31309 11883
rect 31309 11849 31343 11883
rect 31343 11849 31352 11883
rect 31300 11840 31352 11849
rect 32680 11883 32732 11892
rect 32680 11849 32689 11883
rect 32689 11849 32723 11883
rect 32723 11849 32732 11883
rect 32680 11840 32732 11849
rect 33692 11840 33744 11892
rect 19708 11747 19760 11756
rect 16856 11636 16908 11688
rect 19708 11713 19717 11747
rect 19717 11713 19751 11747
rect 19751 11713 19760 11747
rect 19708 11704 19760 11713
rect 20444 11704 20496 11756
rect 22560 11772 22612 11824
rect 22744 11772 22796 11824
rect 21548 11636 21600 11688
rect 24584 11704 24636 11756
rect 25320 11704 25372 11756
rect 28356 11772 28408 11824
rect 30380 11772 30432 11824
rect 28632 11704 28684 11756
rect 30196 11704 30248 11756
rect 23848 11679 23900 11688
rect 23848 11645 23857 11679
rect 23857 11645 23891 11679
rect 23891 11645 23900 11679
rect 23848 11636 23900 11645
rect 27344 11679 27396 11688
rect 27344 11645 27353 11679
rect 27353 11645 27387 11679
rect 27387 11645 27396 11679
rect 27344 11636 27396 11645
rect 31852 11704 31904 11756
rect 32496 11747 32548 11756
rect 32496 11713 32505 11747
rect 32505 11713 32539 11747
rect 32539 11713 32548 11747
rect 32496 11704 32548 11713
rect 33416 11636 33468 11688
rect 22652 11500 22704 11552
rect 22928 11500 22980 11552
rect 23480 11500 23532 11552
rect 24952 11500 25004 11552
rect 26056 11543 26108 11552
rect 26056 11509 26065 11543
rect 26065 11509 26099 11543
rect 26099 11509 26108 11543
rect 26056 11500 26108 11509
rect 29368 11500 29420 11552
rect 31668 11543 31720 11552
rect 31668 11509 31677 11543
rect 31677 11509 31711 11543
rect 31711 11509 31720 11543
rect 31668 11500 31720 11509
rect 32404 11500 32456 11552
rect 5170 11398 5222 11450
rect 5234 11398 5286 11450
rect 5298 11398 5350 11450
rect 5362 11398 5414 11450
rect 5426 11398 5478 11450
rect 13611 11398 13663 11450
rect 13675 11398 13727 11450
rect 13739 11398 13791 11450
rect 13803 11398 13855 11450
rect 13867 11398 13919 11450
rect 22052 11398 22104 11450
rect 22116 11398 22168 11450
rect 22180 11398 22232 11450
rect 22244 11398 22296 11450
rect 22308 11398 22360 11450
rect 30493 11398 30545 11450
rect 30557 11398 30609 11450
rect 30621 11398 30673 11450
rect 30685 11398 30737 11450
rect 30749 11398 30801 11450
rect 4528 11296 4580 11348
rect 17316 11296 17368 11348
rect 21088 11296 21140 11348
rect 21548 11339 21600 11348
rect 21548 11305 21557 11339
rect 21557 11305 21591 11339
rect 21591 11305 21600 11339
rect 21548 11296 21600 11305
rect 15936 11228 15988 11280
rect 22468 11296 22520 11348
rect 22836 11339 22888 11348
rect 22836 11305 22845 11339
rect 22845 11305 22879 11339
rect 22879 11305 22888 11339
rect 22836 11296 22888 11305
rect 2964 11160 3016 11212
rect 3332 11160 3384 11212
rect 3240 11135 3292 11144
rect 3240 11101 3249 11135
rect 3249 11101 3283 11135
rect 3283 11101 3292 11135
rect 3240 11092 3292 11101
rect 12164 11160 12216 11212
rect 17684 11160 17736 11212
rect 2504 11024 2556 11076
rect 3976 11067 4028 11076
rect 3976 11033 3985 11067
rect 3985 11033 4019 11067
rect 4019 11033 4028 11067
rect 3976 11024 4028 11033
rect 6092 11092 6144 11144
rect 10416 11092 10468 11144
rect 11060 11092 11112 11144
rect 12532 11092 12584 11144
rect 12900 11092 12952 11144
rect 13084 11135 13136 11144
rect 13084 11101 13093 11135
rect 13093 11101 13127 11135
rect 13127 11101 13136 11135
rect 13084 11092 13136 11101
rect 16856 11135 16908 11144
rect 16856 11101 16865 11135
rect 16865 11101 16899 11135
rect 16899 11101 16908 11135
rect 16856 11092 16908 11101
rect 16948 11092 17000 11144
rect 17592 11135 17644 11144
rect 17592 11101 17601 11135
rect 17601 11101 17635 11135
rect 17635 11101 17644 11135
rect 17592 11092 17644 11101
rect 19984 11135 20036 11144
rect 5632 11024 5684 11076
rect 9220 11024 9272 11076
rect 3148 10956 3200 11008
rect 4344 10999 4396 11008
rect 4344 10965 4353 10999
rect 4353 10965 4387 10999
rect 4387 10965 4396 10999
rect 4344 10956 4396 10965
rect 6920 10999 6972 11008
rect 6920 10965 6929 10999
rect 6929 10965 6963 10999
rect 6963 10965 6972 10999
rect 6920 10956 6972 10965
rect 7104 10956 7156 11008
rect 8852 10956 8904 11008
rect 8944 10956 8996 11008
rect 9956 10956 10008 11008
rect 12440 11024 12492 11076
rect 12624 11067 12676 11076
rect 12624 11033 12633 11067
rect 12633 11033 12667 11067
rect 12667 11033 12676 11067
rect 12624 11024 12676 11033
rect 13452 11067 13504 11076
rect 13452 11033 13461 11067
rect 13461 11033 13495 11067
rect 13495 11033 13504 11067
rect 13452 11024 13504 11033
rect 16764 11067 16816 11076
rect 16764 11033 16773 11067
rect 16773 11033 16807 11067
rect 16807 11033 16816 11067
rect 16764 11024 16816 11033
rect 19984 11101 19993 11135
rect 19993 11101 20027 11135
rect 20027 11101 20036 11135
rect 19984 11092 20036 11101
rect 20076 11135 20128 11144
rect 20076 11101 20086 11135
rect 20086 11101 20120 11135
rect 20120 11101 20128 11135
rect 20076 11092 20128 11101
rect 19892 11024 19944 11076
rect 20536 11092 20588 11144
rect 21088 11135 21140 11144
rect 21088 11101 21097 11135
rect 21097 11101 21131 11135
rect 21131 11101 21140 11135
rect 21088 11092 21140 11101
rect 21364 11135 21416 11144
rect 21364 11101 21373 11135
rect 21373 11101 21407 11135
rect 21407 11101 21416 11135
rect 21364 11092 21416 11101
rect 22192 11135 22244 11144
rect 22192 11101 22201 11135
rect 22201 11101 22235 11135
rect 22235 11101 22244 11135
rect 22192 11092 22244 11101
rect 22284 11135 22336 11144
rect 22284 11101 22294 11135
rect 22294 11101 22328 11135
rect 22328 11101 22336 11135
rect 22284 11092 22336 11101
rect 22652 11092 22704 11144
rect 25320 11296 25372 11348
rect 31300 11296 31352 11348
rect 23572 11135 23624 11144
rect 23572 11101 23581 11135
rect 23581 11101 23615 11135
rect 23615 11101 23624 11135
rect 23940 11160 23992 11212
rect 24676 11160 24728 11212
rect 23572 11092 23624 11101
rect 12716 10956 12768 11008
rect 20996 10956 21048 11008
rect 21180 11067 21232 11076
rect 21180 11033 21189 11067
rect 21189 11033 21223 11067
rect 21223 11033 21232 11067
rect 21180 11024 21232 11033
rect 23480 11024 23532 11076
rect 25872 11092 25924 11144
rect 26056 11135 26108 11144
rect 26056 11101 26065 11135
rect 26065 11101 26099 11135
rect 26099 11101 26108 11135
rect 26056 11092 26108 11101
rect 26608 11092 26660 11144
rect 26792 11092 26844 11144
rect 29552 11092 29604 11144
rect 30196 11135 30248 11144
rect 24860 11024 24912 11076
rect 28080 11024 28132 11076
rect 29460 11024 29512 11076
rect 30196 11101 30205 11135
rect 30205 11101 30239 11135
rect 30239 11101 30248 11135
rect 30196 11092 30248 11101
rect 32312 11092 32364 11144
rect 30840 11024 30892 11076
rect 31668 11024 31720 11076
rect 26608 10956 26660 11008
rect 29736 10999 29788 11008
rect 29736 10965 29745 10999
rect 29745 10965 29779 10999
rect 29779 10965 29788 10999
rect 29736 10956 29788 10965
rect 30104 10999 30156 11008
rect 30104 10965 30113 10999
rect 30113 10965 30147 10999
rect 30147 10965 30156 10999
rect 30104 10956 30156 10965
rect 9390 10854 9442 10906
rect 9454 10854 9506 10906
rect 9518 10854 9570 10906
rect 9582 10854 9634 10906
rect 9646 10854 9698 10906
rect 17831 10854 17883 10906
rect 17895 10854 17947 10906
rect 17959 10854 18011 10906
rect 18023 10854 18075 10906
rect 18087 10854 18139 10906
rect 26272 10854 26324 10906
rect 26336 10854 26388 10906
rect 26400 10854 26452 10906
rect 26464 10854 26516 10906
rect 26528 10854 26580 10906
rect 34713 10854 34765 10906
rect 34777 10854 34829 10906
rect 34841 10854 34893 10906
rect 34905 10854 34957 10906
rect 34969 10854 35021 10906
rect 4344 10752 4396 10804
rect 6644 10752 6696 10804
rect 6736 10727 6788 10736
rect 2688 10616 2740 10668
rect 3148 10659 3200 10668
rect 3148 10625 3157 10659
rect 3157 10625 3191 10659
rect 3191 10625 3200 10659
rect 3148 10616 3200 10625
rect 6736 10693 6745 10727
rect 6745 10693 6779 10727
rect 6779 10693 6788 10727
rect 6736 10684 6788 10693
rect 6920 10684 6972 10736
rect 7472 10727 7524 10736
rect 7472 10693 7481 10727
rect 7481 10693 7515 10727
rect 7515 10693 7524 10727
rect 7472 10684 7524 10693
rect 8208 10752 8260 10804
rect 8484 10752 8536 10804
rect 8944 10752 8996 10804
rect 4252 10616 4304 10668
rect 7104 10659 7156 10668
rect 7104 10625 7113 10659
rect 7113 10625 7147 10659
rect 7147 10625 7156 10659
rect 7104 10616 7156 10625
rect 2964 10548 3016 10600
rect 3424 10591 3476 10600
rect 2136 10480 2188 10532
rect 3424 10557 3433 10591
rect 3433 10557 3467 10591
rect 3467 10557 3476 10591
rect 3424 10548 3476 10557
rect 6644 10548 6696 10600
rect 9220 10684 9272 10736
rect 9772 10752 9824 10804
rect 9956 10752 10008 10804
rect 19708 10795 19760 10804
rect 19708 10761 19717 10795
rect 19717 10761 19751 10795
rect 19751 10761 19760 10795
rect 19708 10752 19760 10761
rect 20444 10795 20496 10804
rect 20444 10761 20453 10795
rect 20453 10761 20487 10795
rect 20487 10761 20496 10795
rect 20444 10752 20496 10761
rect 20720 10752 20772 10804
rect 22192 10752 22244 10804
rect 11888 10684 11940 10736
rect 12348 10684 12400 10736
rect 12532 10727 12584 10736
rect 12532 10693 12541 10727
rect 12541 10693 12575 10727
rect 12575 10693 12584 10727
rect 12532 10684 12584 10693
rect 12900 10727 12952 10736
rect 12900 10693 12909 10727
rect 12909 10693 12943 10727
rect 12943 10693 12952 10727
rect 12900 10684 12952 10693
rect 14004 10684 14056 10736
rect 18236 10727 18288 10736
rect 18236 10693 18245 10727
rect 18245 10693 18279 10727
rect 18279 10693 18288 10727
rect 18236 10684 18288 10693
rect 19892 10684 19944 10736
rect 23572 10752 23624 10804
rect 25872 10752 25924 10804
rect 29000 10752 29052 10804
rect 30104 10752 30156 10804
rect 33692 10795 33744 10804
rect 33692 10761 33701 10795
rect 33701 10761 33735 10795
rect 33735 10761 33744 10795
rect 33692 10752 33744 10761
rect 9036 10659 9088 10668
rect 9036 10625 9045 10659
rect 9045 10625 9079 10659
rect 9079 10625 9088 10659
rect 9036 10616 9088 10625
rect 12440 10616 12492 10668
rect 19340 10616 19392 10668
rect 11152 10548 11204 10600
rect 12164 10548 12216 10600
rect 22376 10616 22428 10668
rect 23756 10684 23808 10736
rect 24860 10727 24912 10736
rect 24860 10693 24894 10727
rect 24894 10693 24912 10727
rect 24860 10684 24912 10693
rect 28080 10684 28132 10736
rect 29460 10684 29512 10736
rect 22928 10659 22980 10668
rect 22928 10625 22937 10659
rect 22937 10625 22971 10659
rect 22971 10625 22980 10659
rect 22928 10616 22980 10625
rect 29736 10616 29788 10668
rect 32404 10616 32456 10668
rect 8668 10480 8720 10532
rect 23480 10548 23532 10600
rect 24584 10591 24636 10600
rect 24584 10557 24593 10591
rect 24593 10557 24627 10591
rect 24627 10557 24636 10591
rect 24584 10548 24636 10557
rect 27344 10591 27396 10600
rect 27344 10557 27353 10591
rect 27353 10557 27387 10591
rect 27387 10557 27396 10591
rect 27344 10548 27396 10557
rect 32312 10591 32364 10600
rect 32312 10557 32321 10591
rect 32321 10557 32355 10591
rect 32355 10557 32364 10591
rect 32312 10548 32364 10557
rect 22652 10480 22704 10532
rect 2872 10412 2924 10464
rect 4068 10412 4120 10464
rect 5540 10412 5592 10464
rect 7932 10412 7984 10464
rect 10048 10455 10100 10464
rect 10048 10421 10057 10455
rect 10057 10421 10091 10455
rect 10091 10421 10100 10455
rect 10048 10412 10100 10421
rect 14372 10412 14424 10464
rect 29368 10412 29420 10464
rect 31024 10412 31076 10464
rect 5170 10310 5222 10362
rect 5234 10310 5286 10362
rect 5298 10310 5350 10362
rect 5362 10310 5414 10362
rect 5426 10310 5478 10362
rect 13611 10310 13663 10362
rect 13675 10310 13727 10362
rect 13739 10310 13791 10362
rect 13803 10310 13855 10362
rect 13867 10310 13919 10362
rect 22052 10310 22104 10362
rect 22116 10310 22168 10362
rect 22180 10310 22232 10362
rect 22244 10310 22296 10362
rect 22308 10310 22360 10362
rect 30493 10310 30545 10362
rect 30557 10310 30609 10362
rect 30621 10310 30673 10362
rect 30685 10310 30737 10362
rect 30749 10310 30801 10362
rect 2688 10251 2740 10260
rect 2688 10217 2697 10251
rect 2697 10217 2731 10251
rect 2731 10217 2740 10251
rect 2688 10208 2740 10217
rect 3056 10208 3108 10260
rect 4160 10251 4212 10260
rect 4160 10217 4169 10251
rect 4169 10217 4203 10251
rect 4203 10217 4212 10251
rect 4160 10208 4212 10217
rect 2872 10115 2924 10124
rect 1768 10047 1820 10056
rect 1768 10013 1777 10047
rect 1777 10013 1811 10047
rect 1811 10013 1820 10047
rect 1768 10004 1820 10013
rect 2872 10081 2881 10115
rect 2881 10081 2915 10115
rect 2915 10081 2924 10115
rect 2872 10072 2924 10081
rect 3240 10115 3292 10124
rect 3240 10081 3249 10115
rect 3249 10081 3283 10115
rect 3283 10081 3292 10115
rect 3240 10072 3292 10081
rect 3332 10115 3384 10124
rect 3332 10081 3341 10115
rect 3341 10081 3375 10115
rect 3375 10081 3384 10115
rect 5540 10208 5592 10260
rect 6736 10251 6788 10260
rect 6736 10217 6745 10251
rect 6745 10217 6779 10251
rect 6779 10217 6788 10251
rect 6736 10208 6788 10217
rect 9036 10208 9088 10260
rect 12624 10251 12676 10260
rect 12624 10217 12633 10251
rect 12633 10217 12667 10251
rect 12667 10217 12676 10251
rect 12624 10208 12676 10217
rect 23848 10208 23900 10260
rect 24584 10208 24636 10260
rect 25412 10208 25464 10260
rect 27344 10251 27396 10260
rect 27344 10217 27353 10251
rect 27353 10217 27387 10251
rect 27387 10217 27396 10251
rect 27344 10208 27396 10217
rect 28264 10251 28316 10260
rect 28264 10217 28273 10251
rect 28273 10217 28307 10251
rect 28307 10217 28316 10251
rect 28264 10208 28316 10217
rect 32312 10208 32364 10260
rect 8668 10140 8720 10192
rect 11152 10140 11204 10192
rect 3332 10072 3384 10081
rect 10416 10072 10468 10124
rect 4344 10004 4396 10056
rect 6092 10004 6144 10056
rect 7472 10047 7524 10056
rect 7472 10013 7506 10047
rect 7506 10013 7524 10047
rect 2136 9868 2188 9920
rect 5632 9979 5684 9988
rect 5632 9945 5666 9979
rect 5666 9945 5684 9979
rect 2964 9868 3016 9920
rect 3056 9911 3108 9920
rect 3056 9877 3065 9911
rect 3065 9877 3099 9911
rect 3099 9877 3108 9911
rect 5632 9936 5684 9945
rect 7472 10004 7524 10013
rect 24768 10004 24820 10056
rect 25320 10047 25372 10056
rect 25320 10013 25329 10047
rect 25329 10013 25363 10047
rect 25363 10013 25372 10047
rect 25320 10004 25372 10013
rect 11796 9936 11848 9988
rect 12072 9936 12124 9988
rect 25228 9979 25280 9988
rect 25228 9945 25237 9979
rect 25237 9945 25271 9979
rect 25271 9945 25280 9979
rect 25228 9936 25280 9945
rect 25872 9936 25924 9988
rect 26608 10004 26660 10056
rect 28632 10047 28684 10056
rect 3056 9868 3108 9877
rect 4252 9868 4304 9920
rect 7840 9868 7892 9920
rect 13360 9868 13412 9920
rect 27896 9936 27948 9988
rect 28264 9936 28316 9988
rect 28632 10013 28641 10047
rect 28641 10013 28675 10047
rect 28675 10013 28684 10047
rect 28632 10004 28684 10013
rect 29000 10072 29052 10124
rect 28908 10047 28960 10056
rect 28908 10013 28917 10047
rect 28917 10013 28951 10047
rect 28951 10013 28960 10047
rect 28908 10004 28960 10013
rect 29460 10004 29512 10056
rect 30288 10047 30340 10056
rect 30288 10013 30297 10047
rect 30297 10013 30331 10047
rect 30331 10013 30340 10047
rect 30288 10004 30340 10013
rect 33416 10047 33468 10056
rect 33416 10013 33425 10047
rect 33425 10013 33459 10047
rect 33459 10013 33468 10047
rect 33416 10004 33468 10013
rect 33600 10004 33652 10056
rect 28540 9979 28592 9988
rect 28540 9945 28549 9979
rect 28549 9945 28583 9979
rect 28583 9945 28592 9979
rect 28540 9936 28592 9945
rect 32312 9868 32364 9920
rect 33692 9868 33744 9920
rect 33876 9911 33928 9920
rect 33876 9877 33885 9911
rect 33885 9877 33919 9911
rect 33919 9877 33928 9911
rect 33876 9868 33928 9877
rect 9390 9766 9442 9818
rect 9454 9766 9506 9818
rect 9518 9766 9570 9818
rect 9582 9766 9634 9818
rect 9646 9766 9698 9818
rect 17831 9766 17883 9818
rect 17895 9766 17947 9818
rect 17959 9766 18011 9818
rect 18023 9766 18075 9818
rect 18087 9766 18139 9818
rect 26272 9766 26324 9818
rect 26336 9766 26388 9818
rect 26400 9766 26452 9818
rect 26464 9766 26516 9818
rect 26528 9766 26580 9818
rect 34713 9766 34765 9818
rect 34777 9766 34829 9818
rect 34841 9766 34893 9818
rect 34905 9766 34957 9818
rect 34969 9766 35021 9818
rect 1768 9664 1820 9716
rect 4160 9707 4212 9716
rect 4160 9673 4169 9707
rect 4169 9673 4203 9707
rect 4203 9673 4212 9707
rect 4160 9664 4212 9673
rect 4252 9664 4304 9716
rect 8484 9707 8536 9716
rect 8484 9673 8493 9707
rect 8493 9673 8527 9707
rect 8527 9673 8536 9707
rect 8484 9664 8536 9673
rect 10048 9664 10100 9716
rect 17040 9664 17092 9716
rect 2136 9571 2188 9580
rect 2136 9537 2145 9571
rect 2145 9537 2179 9571
rect 2179 9537 2188 9571
rect 2136 9528 2188 9537
rect 7472 9596 7524 9648
rect 16396 9596 16448 9648
rect 28908 9664 28960 9716
rect 31392 9707 31444 9716
rect 4068 9571 4120 9580
rect 3148 9460 3200 9512
rect 4068 9537 4077 9571
rect 4077 9537 4111 9571
rect 4111 9537 4120 9571
rect 4068 9528 4120 9537
rect 4712 9571 4764 9580
rect 4712 9537 4721 9571
rect 4721 9537 4755 9571
rect 4755 9537 4764 9571
rect 4712 9528 4764 9537
rect 5540 9528 5592 9580
rect 6828 9528 6880 9580
rect 11796 9528 11848 9580
rect 17132 9528 17184 9580
rect 17316 9571 17368 9580
rect 17316 9537 17325 9571
rect 17325 9537 17359 9571
rect 17359 9537 17368 9571
rect 17316 9528 17368 9537
rect 17592 9528 17644 9580
rect 18420 9571 18472 9580
rect 10784 9460 10836 9512
rect 16764 9460 16816 9512
rect 18420 9537 18429 9571
rect 18429 9537 18463 9571
rect 18463 9537 18472 9571
rect 18420 9528 18472 9537
rect 19064 9528 19116 9580
rect 12716 9392 12768 9444
rect 2872 9367 2924 9376
rect 2872 9333 2881 9367
rect 2881 9333 2915 9367
rect 2915 9333 2924 9367
rect 2872 9324 2924 9333
rect 15292 9324 15344 9376
rect 19156 9460 19208 9512
rect 19708 9571 19760 9580
rect 19708 9537 19717 9571
rect 19717 9537 19751 9571
rect 19751 9537 19760 9571
rect 19708 9528 19760 9537
rect 19892 9528 19944 9580
rect 20628 9571 20680 9580
rect 20628 9537 20637 9571
rect 20637 9537 20671 9571
rect 20671 9537 20680 9571
rect 20628 9528 20680 9537
rect 21272 9596 21324 9648
rect 23572 9596 23624 9648
rect 24768 9596 24820 9648
rect 31392 9673 31401 9707
rect 31401 9673 31435 9707
rect 31435 9673 31444 9707
rect 31392 9664 31444 9673
rect 21456 9528 21508 9580
rect 22468 9571 22520 9580
rect 22468 9537 22477 9571
rect 22477 9537 22511 9571
rect 22511 9537 22520 9571
rect 22468 9528 22520 9537
rect 25964 9528 26016 9580
rect 31024 9596 31076 9648
rect 27988 9528 28040 9580
rect 30104 9528 30156 9580
rect 31576 9571 31628 9580
rect 31576 9537 31585 9571
rect 31585 9537 31619 9571
rect 31619 9537 31628 9571
rect 31576 9528 31628 9537
rect 18788 9435 18840 9444
rect 18788 9401 18797 9435
rect 18797 9401 18831 9435
rect 18831 9401 18840 9435
rect 18788 9392 18840 9401
rect 18880 9392 18932 9444
rect 23940 9460 23992 9512
rect 19984 9435 20036 9444
rect 19984 9401 19993 9435
rect 19993 9401 20027 9435
rect 20027 9401 20036 9435
rect 19984 9392 20036 9401
rect 20720 9392 20772 9444
rect 25044 9392 25096 9444
rect 30196 9392 30248 9444
rect 33600 9460 33652 9512
rect 20168 9324 20220 9376
rect 30840 9324 30892 9376
rect 31576 9324 31628 9376
rect 31760 9367 31812 9376
rect 31760 9333 31769 9367
rect 31769 9333 31803 9367
rect 31803 9333 31812 9367
rect 31760 9324 31812 9333
rect 33692 9324 33744 9376
rect 5170 9222 5222 9274
rect 5234 9222 5286 9274
rect 5298 9222 5350 9274
rect 5362 9222 5414 9274
rect 5426 9222 5478 9274
rect 13611 9222 13663 9274
rect 13675 9222 13727 9274
rect 13739 9222 13791 9274
rect 13803 9222 13855 9274
rect 13867 9222 13919 9274
rect 22052 9222 22104 9274
rect 22116 9222 22168 9274
rect 22180 9222 22232 9274
rect 22244 9222 22296 9274
rect 22308 9222 22360 9274
rect 30493 9222 30545 9274
rect 30557 9222 30609 9274
rect 30621 9222 30673 9274
rect 30685 9222 30737 9274
rect 30749 9222 30801 9274
rect 2964 9163 3016 9172
rect 2964 9129 2973 9163
rect 2973 9129 3007 9163
rect 3007 9129 3016 9163
rect 2964 9120 3016 9129
rect 12532 9120 12584 9172
rect 16396 9163 16448 9172
rect 16396 9129 16405 9163
rect 16405 9129 16439 9163
rect 16439 9129 16448 9163
rect 16396 9120 16448 9129
rect 18788 9120 18840 9172
rect 20260 9120 20312 9172
rect 21272 9163 21324 9172
rect 21272 9129 21281 9163
rect 21281 9129 21315 9163
rect 21315 9129 21324 9163
rect 21272 9120 21324 9129
rect 22836 9120 22888 9172
rect 26700 9120 26752 9172
rect 32312 9163 32364 9172
rect 32312 9129 32321 9163
rect 32321 9129 32355 9163
rect 32355 9129 32364 9163
rect 32312 9120 32364 9129
rect 21088 9052 21140 9104
rect 4712 8984 4764 9036
rect 6828 8984 6880 9036
rect 10784 9027 10836 9036
rect 10784 8993 10793 9027
rect 10793 8993 10827 9027
rect 10827 8993 10836 9027
rect 10784 8984 10836 8993
rect 4344 8916 4396 8968
rect 11060 8959 11112 8968
rect 11060 8925 11094 8959
rect 11094 8925 11112 8959
rect 11060 8916 11112 8925
rect 15108 8916 15160 8968
rect 15292 8959 15344 8968
rect 15292 8925 15326 8959
rect 15326 8925 15344 8959
rect 15292 8916 15344 8925
rect 16856 8959 16908 8968
rect 16856 8925 16865 8959
rect 16865 8925 16899 8959
rect 16899 8925 16908 8959
rect 16856 8916 16908 8925
rect 19524 8916 19576 8968
rect 19892 8959 19944 8968
rect 19892 8925 19901 8959
rect 19901 8925 19935 8959
rect 19935 8925 19944 8959
rect 19892 8916 19944 8925
rect 20168 8959 20220 8968
rect 20168 8925 20202 8959
rect 20202 8925 20220 8959
rect 20168 8916 20220 8925
rect 22652 8959 22704 8968
rect 22652 8925 22661 8959
rect 22661 8925 22695 8959
rect 22695 8925 22704 8959
rect 22652 8916 22704 8925
rect 22836 8959 22888 8968
rect 22836 8925 22845 8959
rect 22845 8925 22879 8959
rect 22879 8925 22888 8959
rect 22836 8916 22888 8925
rect 23388 9052 23440 9104
rect 26792 9052 26844 9104
rect 30196 9052 30248 9104
rect 23664 8916 23716 8968
rect 24584 8959 24636 8968
rect 24584 8925 24593 8959
rect 24593 8925 24627 8959
rect 24627 8925 24636 8959
rect 24584 8916 24636 8925
rect 2872 8848 2924 8900
rect 3056 8848 3108 8900
rect 3424 8848 3476 8900
rect 17224 8848 17276 8900
rect 19708 8848 19760 8900
rect 28908 8916 28960 8968
rect 30196 8959 30248 8968
rect 4344 8823 4396 8832
rect 4344 8789 4353 8823
rect 4353 8789 4387 8823
rect 4387 8789 4396 8823
rect 4344 8780 4396 8789
rect 18788 8780 18840 8832
rect 21916 8780 21968 8832
rect 28172 8848 28224 8900
rect 30196 8925 30205 8959
rect 30205 8925 30239 8959
rect 30239 8925 30248 8959
rect 30196 8916 30248 8925
rect 32312 8916 32364 8968
rect 30288 8848 30340 8900
rect 33876 8848 33928 8900
rect 23664 8780 23716 8832
rect 25044 8823 25096 8832
rect 25044 8789 25053 8823
rect 25053 8789 25087 8823
rect 25087 8789 25096 8823
rect 25044 8780 25096 8789
rect 29184 8823 29236 8832
rect 29184 8789 29193 8823
rect 29193 8789 29227 8823
rect 29227 8789 29236 8823
rect 29184 8780 29236 8789
rect 29736 8823 29788 8832
rect 29736 8789 29745 8823
rect 29745 8789 29779 8823
rect 29779 8789 29788 8823
rect 29736 8780 29788 8789
rect 9390 8678 9442 8730
rect 9454 8678 9506 8730
rect 9518 8678 9570 8730
rect 9582 8678 9634 8730
rect 9646 8678 9698 8730
rect 17831 8678 17883 8730
rect 17895 8678 17947 8730
rect 17959 8678 18011 8730
rect 18023 8678 18075 8730
rect 18087 8678 18139 8730
rect 26272 8678 26324 8730
rect 26336 8678 26388 8730
rect 26400 8678 26452 8730
rect 26464 8678 26516 8730
rect 26528 8678 26580 8730
rect 34713 8678 34765 8730
rect 34777 8678 34829 8730
rect 34841 8678 34893 8730
rect 34905 8678 34957 8730
rect 34969 8678 35021 8730
rect 16212 8576 16264 8628
rect 9312 8508 9364 8560
rect 16396 8508 16448 8560
rect 9864 8304 9916 8356
rect 16856 8440 16908 8492
rect 17684 8619 17736 8628
rect 17684 8585 17693 8619
rect 17693 8585 17727 8619
rect 17727 8585 17736 8619
rect 17684 8576 17736 8585
rect 19064 8576 19116 8628
rect 19156 8576 19208 8628
rect 18880 8508 18932 8560
rect 17592 8372 17644 8424
rect 16304 8304 16356 8356
rect 17132 8236 17184 8288
rect 18696 8440 18748 8492
rect 18788 8440 18840 8492
rect 19892 8372 19944 8424
rect 20536 8372 20588 8424
rect 23388 8576 23440 8628
rect 23664 8619 23716 8628
rect 23664 8585 23673 8619
rect 23673 8585 23707 8619
rect 23707 8585 23716 8619
rect 23664 8576 23716 8585
rect 23940 8576 23992 8628
rect 22744 8551 22796 8560
rect 22744 8517 22753 8551
rect 22753 8517 22787 8551
rect 22787 8517 22796 8551
rect 22744 8508 22796 8517
rect 23572 8508 23624 8560
rect 25044 8508 25096 8560
rect 25228 8576 25280 8628
rect 25872 8619 25924 8628
rect 25872 8585 25881 8619
rect 25881 8585 25915 8619
rect 25915 8585 25924 8619
rect 25872 8576 25924 8585
rect 28908 8576 28960 8628
rect 21456 8440 21508 8492
rect 24952 8440 25004 8492
rect 26056 8440 26108 8492
rect 29092 8508 29144 8560
rect 30288 8576 30340 8628
rect 30932 8576 30984 8628
rect 31392 8576 31444 8628
rect 29736 8440 29788 8492
rect 30196 8440 30248 8492
rect 31760 8508 31812 8560
rect 20904 8372 20956 8424
rect 25044 8415 25096 8424
rect 25044 8381 25053 8415
rect 25053 8381 25087 8415
rect 25087 8381 25096 8415
rect 25044 8372 25096 8381
rect 31852 8440 31904 8492
rect 32312 8483 32364 8492
rect 32312 8449 32321 8483
rect 32321 8449 32355 8483
rect 32355 8449 32364 8483
rect 32312 8440 32364 8449
rect 24032 8304 24084 8356
rect 19340 8236 19392 8288
rect 29368 8236 29420 8288
rect 5170 8134 5222 8186
rect 5234 8134 5286 8186
rect 5298 8134 5350 8186
rect 5362 8134 5414 8186
rect 5426 8134 5478 8186
rect 13611 8134 13663 8186
rect 13675 8134 13727 8186
rect 13739 8134 13791 8186
rect 13803 8134 13855 8186
rect 13867 8134 13919 8186
rect 22052 8134 22104 8186
rect 22116 8134 22168 8186
rect 22180 8134 22232 8186
rect 22244 8134 22296 8186
rect 22308 8134 22360 8186
rect 30493 8134 30545 8186
rect 30557 8134 30609 8186
rect 30621 8134 30673 8186
rect 30685 8134 30737 8186
rect 30749 8134 30801 8186
rect 15660 8032 15712 8084
rect 18696 8032 18748 8084
rect 29368 8032 29420 8084
rect 32312 8032 32364 8084
rect 19340 7964 19392 8016
rect 4068 7828 4120 7880
rect 20628 7896 20680 7948
rect 25136 7896 25188 7948
rect 9864 7871 9916 7880
rect 9864 7837 9873 7871
rect 9873 7837 9907 7871
rect 9907 7837 9916 7871
rect 9864 7828 9916 7837
rect 7380 7803 7432 7812
rect 7380 7769 7389 7803
rect 7389 7769 7423 7803
rect 7423 7769 7432 7803
rect 7380 7760 7432 7769
rect 8208 7760 8260 7812
rect 24032 7828 24084 7880
rect 33692 7871 33744 7880
rect 33692 7837 33701 7871
rect 33701 7837 33735 7871
rect 33735 7837 33744 7871
rect 33692 7828 33744 7837
rect 10232 7803 10284 7812
rect 10232 7769 10241 7803
rect 10241 7769 10275 7803
rect 10275 7769 10284 7803
rect 10232 7760 10284 7769
rect 15568 7760 15620 7812
rect 17316 7760 17368 7812
rect 17500 7735 17552 7744
rect 17500 7701 17509 7735
rect 17509 7701 17543 7735
rect 17543 7701 17552 7735
rect 17500 7692 17552 7701
rect 19156 7692 19208 7744
rect 20812 7760 20864 7812
rect 28080 7803 28132 7812
rect 28080 7769 28089 7803
rect 28089 7769 28123 7803
rect 28123 7769 28132 7803
rect 28080 7760 28132 7769
rect 28448 7760 28500 7812
rect 23388 7692 23440 7744
rect 28264 7735 28316 7744
rect 28264 7701 28273 7735
rect 28273 7701 28307 7735
rect 28307 7701 28316 7735
rect 28264 7692 28316 7701
rect 30380 7692 30432 7744
rect 9390 7590 9442 7642
rect 9454 7590 9506 7642
rect 9518 7590 9570 7642
rect 9582 7590 9634 7642
rect 9646 7590 9698 7642
rect 17831 7590 17883 7642
rect 17895 7590 17947 7642
rect 17959 7590 18011 7642
rect 18023 7590 18075 7642
rect 18087 7590 18139 7642
rect 26272 7590 26324 7642
rect 26336 7590 26388 7642
rect 26400 7590 26452 7642
rect 26464 7590 26516 7642
rect 26528 7590 26580 7642
rect 34713 7590 34765 7642
rect 34777 7590 34829 7642
rect 34841 7590 34893 7642
rect 34905 7590 34957 7642
rect 34969 7590 35021 7642
rect 10692 7531 10744 7540
rect 10692 7497 10701 7531
rect 10701 7497 10735 7531
rect 10735 7497 10744 7531
rect 10692 7488 10744 7497
rect 15568 7531 15620 7540
rect 15568 7497 15577 7531
rect 15577 7497 15611 7531
rect 15611 7497 15620 7531
rect 15568 7488 15620 7497
rect 16764 7488 16816 7540
rect 17500 7488 17552 7540
rect 18788 7488 18840 7540
rect 19524 7531 19576 7540
rect 19524 7497 19533 7531
rect 19533 7497 19567 7531
rect 19567 7497 19576 7531
rect 19524 7488 19576 7497
rect 20720 7488 20772 7540
rect 20904 7488 20956 7540
rect 25964 7531 26016 7540
rect 25964 7497 25973 7531
rect 25973 7497 26007 7531
rect 26007 7497 26016 7531
rect 25964 7488 26016 7497
rect 29092 7531 29144 7540
rect 29092 7497 29101 7531
rect 29101 7497 29135 7531
rect 29135 7497 29144 7531
rect 29092 7488 29144 7497
rect 5632 7420 5684 7472
rect 7380 7420 7432 7472
rect 10232 7420 10284 7472
rect 17316 7420 17368 7472
rect 2504 7395 2556 7404
rect 2504 7361 2513 7395
rect 2513 7361 2547 7395
rect 2547 7361 2556 7395
rect 2504 7352 2556 7361
rect 8392 7352 8444 7404
rect 8944 7395 8996 7404
rect 8944 7361 8953 7395
rect 8953 7361 8987 7395
rect 8987 7361 8996 7395
rect 8944 7352 8996 7361
rect 17500 7395 17552 7404
rect 17500 7361 17509 7395
rect 17509 7361 17543 7395
rect 17543 7361 17552 7395
rect 17500 7352 17552 7361
rect 17868 7352 17920 7404
rect 19340 7352 19392 7404
rect 20628 7395 20680 7404
rect 20628 7361 20637 7395
rect 20637 7361 20671 7395
rect 20671 7361 20680 7395
rect 20628 7352 20680 7361
rect 22284 7420 22336 7472
rect 23388 7463 23440 7472
rect 23388 7429 23397 7463
rect 23397 7429 23431 7463
rect 23431 7429 23440 7463
rect 23388 7420 23440 7429
rect 25044 7463 25096 7472
rect 25044 7429 25053 7463
rect 25053 7429 25087 7463
rect 25087 7429 25096 7463
rect 25044 7420 25096 7429
rect 11060 7284 11112 7336
rect 11152 7284 11204 7336
rect 11888 7327 11940 7336
rect 11888 7293 11897 7327
rect 11897 7293 11931 7327
rect 11931 7293 11940 7327
rect 11888 7284 11940 7293
rect 13084 7284 13136 7336
rect 17224 7284 17276 7336
rect 25136 7352 25188 7404
rect 26056 7395 26108 7404
rect 26056 7361 26065 7395
rect 26065 7361 26099 7395
rect 26099 7361 26108 7395
rect 26056 7352 26108 7361
rect 30380 7395 30432 7404
rect 30380 7361 30389 7395
rect 30389 7361 30423 7395
rect 30423 7361 30432 7395
rect 30380 7352 30432 7361
rect 23756 7284 23808 7336
rect 24032 7284 24084 7336
rect 24584 7284 24636 7336
rect 2596 7191 2648 7200
rect 2596 7157 2605 7191
rect 2605 7157 2639 7191
rect 2639 7157 2648 7191
rect 2596 7148 2648 7157
rect 8300 7191 8352 7200
rect 8300 7157 8309 7191
rect 8309 7157 8343 7191
rect 8343 7157 8352 7191
rect 8300 7148 8352 7157
rect 12532 7191 12584 7200
rect 12532 7157 12541 7191
rect 12541 7157 12575 7191
rect 12575 7157 12584 7191
rect 12532 7148 12584 7157
rect 15108 7148 15160 7200
rect 15660 7148 15712 7200
rect 20444 7191 20496 7200
rect 20444 7157 20453 7191
rect 20453 7157 20487 7191
rect 20487 7157 20496 7191
rect 20444 7148 20496 7157
rect 20720 7148 20772 7200
rect 25596 7191 25648 7200
rect 25596 7157 25605 7191
rect 25605 7157 25639 7191
rect 25639 7157 25648 7191
rect 25596 7148 25648 7157
rect 5170 7046 5222 7098
rect 5234 7046 5286 7098
rect 5298 7046 5350 7098
rect 5362 7046 5414 7098
rect 5426 7046 5478 7098
rect 13611 7046 13663 7098
rect 13675 7046 13727 7098
rect 13739 7046 13791 7098
rect 13803 7046 13855 7098
rect 13867 7046 13919 7098
rect 22052 7046 22104 7098
rect 22116 7046 22168 7098
rect 22180 7046 22232 7098
rect 22244 7046 22296 7098
rect 22308 7046 22360 7098
rect 30493 7046 30545 7098
rect 30557 7046 30609 7098
rect 30621 7046 30673 7098
rect 30685 7046 30737 7098
rect 30749 7046 30801 7098
rect 2504 6944 2556 6996
rect 2596 6944 2648 6996
rect 13084 6987 13136 6996
rect 13084 6953 13093 6987
rect 13093 6953 13127 6987
rect 13127 6953 13136 6987
rect 13084 6944 13136 6953
rect 20812 6987 20864 6996
rect 20812 6953 20821 6987
rect 20821 6953 20855 6987
rect 20855 6953 20864 6987
rect 20812 6944 20864 6953
rect 4344 6808 4396 6860
rect 5080 6808 5132 6860
rect 3424 6783 3476 6792
rect 3424 6749 3433 6783
rect 3433 6749 3467 6783
rect 3467 6749 3476 6783
rect 3424 6740 3476 6749
rect 4068 6740 4120 6792
rect 5724 6783 5776 6792
rect 5724 6749 5758 6783
rect 5758 6749 5776 6783
rect 5724 6740 5776 6749
rect 17224 6876 17276 6928
rect 17868 6876 17920 6928
rect 2688 6672 2740 6724
rect 6920 6604 6972 6656
rect 8300 6808 8352 6860
rect 10324 6808 10376 6860
rect 15108 6808 15160 6860
rect 10416 6740 10468 6792
rect 10692 6672 10744 6724
rect 11152 6740 11204 6792
rect 11704 6783 11756 6792
rect 11704 6749 11713 6783
rect 11713 6749 11747 6783
rect 11747 6749 11756 6783
rect 11704 6740 11756 6749
rect 11060 6672 11112 6724
rect 12808 6672 12860 6724
rect 15660 6740 15712 6792
rect 16304 6740 16356 6792
rect 16396 6740 16448 6792
rect 19340 6808 19392 6860
rect 20536 6808 20588 6860
rect 17868 6783 17920 6792
rect 17868 6749 17877 6783
rect 17877 6749 17911 6783
rect 17911 6749 17920 6783
rect 17868 6740 17920 6749
rect 19524 6740 19576 6792
rect 20444 6740 20496 6792
rect 21916 6740 21968 6792
rect 23756 6783 23808 6792
rect 23756 6749 23765 6783
rect 23765 6749 23799 6783
rect 23799 6749 23808 6783
rect 23756 6740 23808 6749
rect 24032 6783 24084 6792
rect 24032 6749 24041 6783
rect 24041 6749 24075 6783
rect 24075 6749 24084 6783
rect 24032 6740 24084 6749
rect 28908 6783 28960 6792
rect 28908 6749 28926 6783
rect 28926 6749 28960 6783
rect 28908 6740 28960 6749
rect 29092 6740 29144 6792
rect 29828 6740 29880 6792
rect 17224 6672 17276 6724
rect 17500 6672 17552 6724
rect 23480 6672 23532 6724
rect 24952 6672 25004 6724
rect 25044 6672 25096 6724
rect 29276 6672 29328 6724
rect 13636 6647 13688 6656
rect 13636 6613 13645 6647
rect 13645 6613 13679 6647
rect 13679 6613 13688 6647
rect 13636 6604 13688 6613
rect 17684 6604 17736 6656
rect 22836 6604 22888 6656
rect 23572 6647 23624 6656
rect 23572 6613 23581 6647
rect 23581 6613 23615 6647
rect 23615 6613 23624 6647
rect 23572 6604 23624 6613
rect 25872 6604 25924 6656
rect 27804 6647 27856 6656
rect 27804 6613 27813 6647
rect 27813 6613 27847 6647
rect 27847 6613 27856 6647
rect 27804 6604 27856 6613
rect 28540 6604 28592 6656
rect 9390 6502 9442 6554
rect 9454 6502 9506 6554
rect 9518 6502 9570 6554
rect 9582 6502 9634 6554
rect 9646 6502 9698 6554
rect 17831 6502 17883 6554
rect 17895 6502 17947 6554
rect 17959 6502 18011 6554
rect 18023 6502 18075 6554
rect 18087 6502 18139 6554
rect 26272 6502 26324 6554
rect 26336 6502 26388 6554
rect 26400 6502 26452 6554
rect 26464 6502 26516 6554
rect 26528 6502 26580 6554
rect 34713 6502 34765 6554
rect 34777 6502 34829 6554
rect 34841 6502 34893 6554
rect 34905 6502 34957 6554
rect 34969 6502 35021 6554
rect 2504 6400 2556 6452
rect 6920 6443 6972 6452
rect 2688 6332 2740 6384
rect 6920 6409 6929 6443
rect 6929 6409 6963 6443
rect 6963 6409 6972 6443
rect 6920 6400 6972 6409
rect 12532 6400 12584 6452
rect 20904 6443 20956 6452
rect 20904 6409 20913 6443
rect 20913 6409 20947 6443
rect 20947 6409 20956 6443
rect 20904 6400 20956 6409
rect 27804 6400 27856 6452
rect 30932 6400 30984 6452
rect 7012 6332 7064 6384
rect 13636 6332 13688 6384
rect 20720 6332 20772 6384
rect 23572 6332 23624 6384
rect 29184 6332 29236 6384
rect 2964 6307 3016 6316
rect 2964 6273 2973 6307
rect 2973 6273 3007 6307
rect 3007 6273 3016 6307
rect 2964 6264 3016 6273
rect 3424 6264 3476 6316
rect 5724 6196 5776 6248
rect 12348 6196 12400 6248
rect 19524 6239 19576 6248
rect 19524 6205 19533 6239
rect 19533 6205 19567 6239
rect 19567 6205 19576 6239
rect 19524 6196 19576 6205
rect 29828 6239 29880 6248
rect 18420 6128 18472 6180
rect 23480 6128 23532 6180
rect 3976 6060 4028 6112
rect 20168 6060 20220 6112
rect 24676 6060 24728 6112
rect 29828 6205 29837 6239
rect 29837 6205 29871 6239
rect 29871 6205 29880 6239
rect 29828 6196 29880 6205
rect 28172 6128 28224 6180
rect 5170 5958 5222 6010
rect 5234 5958 5286 6010
rect 5298 5958 5350 6010
rect 5362 5958 5414 6010
rect 5426 5958 5478 6010
rect 13611 5958 13663 6010
rect 13675 5958 13727 6010
rect 13739 5958 13791 6010
rect 13803 5958 13855 6010
rect 13867 5958 13919 6010
rect 22052 5958 22104 6010
rect 22116 5958 22168 6010
rect 22180 5958 22232 6010
rect 22244 5958 22296 6010
rect 22308 5958 22360 6010
rect 30493 5958 30545 6010
rect 30557 5958 30609 6010
rect 30621 5958 30673 6010
rect 30685 5958 30737 6010
rect 30749 5958 30801 6010
rect 25964 5899 26016 5908
rect 25964 5865 25973 5899
rect 25973 5865 26007 5899
rect 26007 5865 26016 5899
rect 25964 5856 26016 5865
rect 29276 5856 29328 5908
rect 3976 5763 4028 5772
rect 3976 5729 3985 5763
rect 3985 5729 4019 5763
rect 4019 5729 4028 5763
rect 3976 5720 4028 5729
rect 5540 5720 5592 5772
rect 5724 5763 5776 5772
rect 5724 5729 5733 5763
rect 5733 5729 5767 5763
rect 5767 5729 5776 5763
rect 5724 5720 5776 5729
rect 11888 5720 11940 5772
rect 12348 5652 12400 5704
rect 12716 5695 12768 5704
rect 12716 5661 12725 5695
rect 12725 5661 12759 5695
rect 12759 5661 12768 5695
rect 12716 5652 12768 5661
rect 24676 5652 24728 5704
rect 25596 5652 25648 5704
rect 29000 5788 29052 5840
rect 30840 5652 30892 5704
rect 4712 5584 4764 5636
rect 28540 5584 28592 5636
rect 14280 5516 14332 5568
rect 9390 5414 9442 5466
rect 9454 5414 9506 5466
rect 9518 5414 9570 5466
rect 9582 5414 9634 5466
rect 9646 5414 9698 5466
rect 17831 5414 17883 5466
rect 17895 5414 17947 5466
rect 17959 5414 18011 5466
rect 18023 5414 18075 5466
rect 18087 5414 18139 5466
rect 26272 5414 26324 5466
rect 26336 5414 26388 5466
rect 26400 5414 26452 5466
rect 26464 5414 26516 5466
rect 26528 5414 26580 5466
rect 34713 5414 34765 5466
rect 34777 5414 34829 5466
rect 34841 5414 34893 5466
rect 34905 5414 34957 5466
rect 34969 5414 35021 5466
rect 5540 5312 5592 5364
rect 4712 5244 4764 5296
rect 10232 5312 10284 5364
rect 10416 5355 10468 5364
rect 10416 5321 10425 5355
rect 10425 5321 10459 5355
rect 10459 5321 10468 5355
rect 10416 5312 10468 5321
rect 12716 5312 12768 5364
rect 19524 5355 19576 5364
rect 19524 5321 19533 5355
rect 19533 5321 19567 5355
rect 19567 5321 19576 5355
rect 19524 5312 19576 5321
rect 24676 5355 24728 5364
rect 24676 5321 24685 5355
rect 24685 5321 24719 5355
rect 24719 5321 24728 5355
rect 24676 5312 24728 5321
rect 6644 5244 6696 5296
rect 4068 5219 4120 5228
rect 4068 5185 4077 5219
rect 4077 5185 4111 5219
rect 4111 5185 4120 5219
rect 4068 5176 4120 5185
rect 5724 5219 5776 5228
rect 2964 5108 3016 5160
rect 5724 5185 5733 5219
rect 5733 5185 5767 5219
rect 5767 5185 5776 5219
rect 5724 5176 5776 5185
rect 8208 5108 8260 5160
rect 9220 5244 9272 5296
rect 18696 5244 18748 5296
rect 23388 5287 23440 5296
rect 23388 5253 23397 5287
rect 23397 5253 23431 5287
rect 23431 5253 23440 5287
rect 23388 5244 23440 5253
rect 26056 5244 26108 5296
rect 10876 5176 10928 5228
rect 11796 5176 11848 5228
rect 15200 5219 15252 5228
rect 15200 5185 15209 5219
rect 15209 5185 15243 5219
rect 15243 5185 15252 5219
rect 15200 5176 15252 5185
rect 26240 5176 26292 5228
rect 9312 5108 9364 5160
rect 11704 5151 11756 5160
rect 7196 5040 7248 5092
rect 11704 5117 11713 5151
rect 11713 5117 11747 5151
rect 11747 5117 11756 5151
rect 11704 5108 11756 5117
rect 14832 4972 14884 5024
rect 14924 4972 14976 5024
rect 25596 5015 25648 5024
rect 25596 4981 25605 5015
rect 25605 4981 25639 5015
rect 25639 4981 25648 5015
rect 25596 4972 25648 4981
rect 5170 4870 5222 4922
rect 5234 4870 5286 4922
rect 5298 4870 5350 4922
rect 5362 4870 5414 4922
rect 5426 4870 5478 4922
rect 13611 4870 13663 4922
rect 13675 4870 13727 4922
rect 13739 4870 13791 4922
rect 13803 4870 13855 4922
rect 13867 4870 13919 4922
rect 22052 4870 22104 4922
rect 22116 4870 22168 4922
rect 22180 4870 22232 4922
rect 22244 4870 22296 4922
rect 22308 4870 22360 4922
rect 30493 4870 30545 4922
rect 30557 4870 30609 4922
rect 30621 4870 30673 4922
rect 30685 4870 30737 4922
rect 30749 4870 30801 4922
rect 10876 4811 10928 4820
rect 10876 4777 10885 4811
rect 10885 4777 10919 4811
rect 10919 4777 10928 4811
rect 10876 4768 10928 4777
rect 11888 4768 11940 4820
rect 13268 4768 13320 4820
rect 5080 4632 5132 4684
rect 7196 4675 7248 4684
rect 7196 4641 7205 4675
rect 7205 4641 7239 4675
rect 7239 4641 7248 4675
rect 7196 4632 7248 4641
rect 8944 4632 8996 4684
rect 7472 4607 7524 4616
rect 7472 4573 7506 4607
rect 7506 4573 7524 4607
rect 7472 4564 7524 4573
rect 20720 4700 20772 4752
rect 14188 4632 14240 4684
rect 12348 4564 12400 4616
rect 14280 4607 14332 4616
rect 14280 4573 14289 4607
rect 14289 4573 14323 4607
rect 14323 4573 14332 4607
rect 14280 4564 14332 4573
rect 20444 4675 20496 4684
rect 20444 4641 20453 4675
rect 20453 4641 20487 4675
rect 20487 4641 20496 4675
rect 20444 4632 20496 4641
rect 26240 4768 26292 4820
rect 26608 4768 26660 4820
rect 24952 4743 25004 4752
rect 24952 4709 24961 4743
rect 24961 4709 24995 4743
rect 24995 4709 25004 4743
rect 24952 4700 25004 4709
rect 15936 4607 15988 4616
rect 15936 4573 15945 4607
rect 15945 4573 15979 4607
rect 15979 4573 15988 4607
rect 15936 4564 15988 4573
rect 17316 4564 17368 4616
rect 18420 4607 18472 4616
rect 18420 4573 18429 4607
rect 18429 4573 18463 4607
rect 18463 4573 18472 4607
rect 18420 4564 18472 4573
rect 20168 4607 20220 4616
rect 20168 4573 20177 4607
rect 20177 4573 20211 4607
rect 20211 4573 20220 4607
rect 20168 4564 20220 4573
rect 20904 4564 20956 4616
rect 25872 4607 25924 4616
rect 25872 4573 25881 4607
rect 25881 4573 25915 4607
rect 25915 4573 25924 4607
rect 25872 4564 25924 4573
rect 8576 4471 8628 4480
rect 8576 4437 8585 4471
rect 8585 4437 8619 4471
rect 8619 4437 8628 4471
rect 8576 4428 8628 4437
rect 10416 4496 10468 4548
rect 26148 4539 26200 4548
rect 26148 4505 26182 4539
rect 26182 4505 26200 4539
rect 26148 4496 26200 4505
rect 11796 4428 11848 4480
rect 15568 4471 15620 4480
rect 15568 4437 15577 4471
rect 15577 4437 15611 4471
rect 15611 4437 15620 4471
rect 15568 4428 15620 4437
rect 16304 4428 16356 4480
rect 17500 4471 17552 4480
rect 17500 4437 17509 4471
rect 17509 4437 17543 4471
rect 17543 4437 17552 4471
rect 17500 4428 17552 4437
rect 18236 4428 18288 4480
rect 19064 4428 19116 4480
rect 19800 4471 19852 4480
rect 19800 4437 19809 4471
rect 19809 4437 19843 4471
rect 19843 4437 19852 4471
rect 19800 4428 19852 4437
rect 20812 4428 20864 4480
rect 21548 4471 21600 4480
rect 21548 4437 21557 4471
rect 21557 4437 21591 4471
rect 21591 4437 21600 4471
rect 21548 4428 21600 4437
rect 22100 4428 22152 4480
rect 25044 4471 25096 4480
rect 25044 4437 25053 4471
rect 25053 4437 25087 4471
rect 25087 4437 25096 4471
rect 25044 4428 25096 4437
rect 27252 4471 27304 4480
rect 27252 4437 27261 4471
rect 27261 4437 27295 4471
rect 27295 4437 27304 4471
rect 27252 4428 27304 4437
rect 9390 4326 9442 4378
rect 9454 4326 9506 4378
rect 9518 4326 9570 4378
rect 9582 4326 9634 4378
rect 9646 4326 9698 4378
rect 17831 4326 17883 4378
rect 17895 4326 17947 4378
rect 17959 4326 18011 4378
rect 18023 4326 18075 4378
rect 18087 4326 18139 4378
rect 26272 4326 26324 4378
rect 26336 4326 26388 4378
rect 26400 4326 26452 4378
rect 26464 4326 26516 4378
rect 26528 4326 26580 4378
rect 34713 4326 34765 4378
rect 34777 4326 34829 4378
rect 34841 4326 34893 4378
rect 34905 4326 34957 4378
rect 34969 4326 35021 4378
rect 7472 4224 7524 4276
rect 8576 4224 8628 4276
rect 13360 4267 13412 4276
rect 13360 4233 13369 4267
rect 13369 4233 13403 4267
rect 13403 4233 13412 4267
rect 13360 4224 13412 4233
rect 14832 4224 14884 4276
rect 22468 4224 22520 4276
rect 26148 4267 26200 4276
rect 26148 4233 26157 4267
rect 26157 4233 26191 4267
rect 26191 4233 26200 4267
rect 26148 4224 26200 4233
rect 7932 4156 7984 4208
rect 9220 4156 9272 4208
rect 15568 4156 15620 4208
rect 8944 4088 8996 4140
rect 10416 4131 10468 4140
rect 10416 4097 10425 4131
rect 10425 4097 10459 4131
rect 10459 4097 10468 4131
rect 10416 4088 10468 4097
rect 10508 4131 10560 4140
rect 10508 4097 10517 4131
rect 10517 4097 10551 4131
rect 10551 4097 10560 4131
rect 10784 4131 10836 4140
rect 10508 4088 10560 4097
rect 10784 4097 10793 4131
rect 10793 4097 10827 4131
rect 10827 4097 10836 4131
rect 10784 4088 10836 4097
rect 14004 4088 14056 4140
rect 14924 4131 14976 4140
rect 14924 4097 14933 4131
rect 14933 4097 14967 4131
rect 14967 4097 14976 4131
rect 14924 4088 14976 4097
rect 17316 4088 17368 4140
rect 17500 4088 17552 4140
rect 17960 4131 18012 4140
rect 17960 4097 17994 4131
rect 17994 4097 18012 4131
rect 17960 4088 18012 4097
rect 25596 4156 25648 4208
rect 20904 4088 20956 4140
rect 21180 4131 21232 4140
rect 21180 4097 21198 4131
rect 21198 4097 21232 4131
rect 21180 4088 21232 4097
rect 21548 4088 21600 4140
rect 22100 4088 22152 4140
rect 22284 4131 22336 4140
rect 22284 4097 22318 4131
rect 22318 4097 22336 4131
rect 22284 4088 22336 4097
rect 25872 4088 25924 4140
rect 28264 4131 28316 4140
rect 28264 4097 28282 4131
rect 28282 4097 28316 4131
rect 28264 4088 28316 4097
rect 28448 4088 28500 4140
rect 11888 4020 11940 4072
rect 14188 4020 14240 4072
rect 26608 4063 26660 4072
rect 26608 4029 26617 4063
rect 26617 4029 26651 4063
rect 26651 4029 26660 4063
rect 26608 4020 26660 4029
rect 9312 3952 9364 4004
rect 26240 3995 26292 4004
rect 26240 3961 26249 3995
rect 26249 3961 26283 3995
rect 26283 3961 26292 3995
rect 26240 3952 26292 3961
rect 12992 3927 13044 3936
rect 12992 3893 13001 3927
rect 13001 3893 13035 3927
rect 13035 3893 13044 3927
rect 12992 3884 13044 3893
rect 16304 3927 16356 3936
rect 16304 3893 16313 3927
rect 16313 3893 16347 3927
rect 16347 3893 16356 3927
rect 16304 3884 16356 3893
rect 16672 3884 16724 3936
rect 19064 3927 19116 3936
rect 19064 3893 19073 3927
rect 19073 3893 19107 3927
rect 19107 3893 19116 3927
rect 19064 3884 19116 3893
rect 21088 3884 21140 3936
rect 23388 3927 23440 3936
rect 23388 3893 23397 3927
rect 23397 3893 23431 3927
rect 23431 3893 23440 3927
rect 23388 3884 23440 3893
rect 24952 3884 25004 3936
rect 27620 3884 27672 3936
rect 5170 3782 5222 3834
rect 5234 3782 5286 3834
rect 5298 3782 5350 3834
rect 5362 3782 5414 3834
rect 5426 3782 5478 3834
rect 13611 3782 13663 3834
rect 13675 3782 13727 3834
rect 13739 3782 13791 3834
rect 13803 3782 13855 3834
rect 13867 3782 13919 3834
rect 22052 3782 22104 3834
rect 22116 3782 22168 3834
rect 22180 3782 22232 3834
rect 22244 3782 22296 3834
rect 22308 3782 22360 3834
rect 30493 3782 30545 3834
rect 30557 3782 30609 3834
rect 30621 3782 30673 3834
rect 30685 3782 30737 3834
rect 30749 3782 30801 3834
rect 7932 3723 7984 3732
rect 7932 3689 7941 3723
rect 7941 3689 7975 3723
rect 7975 3689 7984 3723
rect 7932 3680 7984 3689
rect 14004 3680 14056 3732
rect 20812 3680 20864 3732
rect 22376 3680 22428 3732
rect 26792 3723 26844 3732
rect 26792 3689 26801 3723
rect 26801 3689 26835 3723
rect 26835 3689 26844 3723
rect 26792 3680 26844 3689
rect 9864 3544 9916 3596
rect 10784 3544 10836 3596
rect 16672 3587 16724 3596
rect 16672 3553 16681 3587
rect 16681 3553 16715 3587
rect 16715 3553 16724 3587
rect 16672 3544 16724 3553
rect 8208 3476 8260 3528
rect 10508 3476 10560 3528
rect 12348 3519 12400 3528
rect 12348 3485 12357 3519
rect 12357 3485 12391 3519
rect 12391 3485 12400 3519
rect 12348 3476 12400 3485
rect 12992 3476 13044 3528
rect 15660 3519 15712 3528
rect 15660 3485 15669 3519
rect 15669 3485 15703 3519
rect 15703 3485 15712 3519
rect 15660 3476 15712 3485
rect 16764 3476 16816 3528
rect 19524 3519 19576 3528
rect 14740 3408 14792 3460
rect 16948 3451 17000 3460
rect 16948 3417 16982 3451
rect 16982 3417 17000 3451
rect 19524 3485 19533 3519
rect 19533 3485 19567 3519
rect 19567 3485 19576 3519
rect 19524 3476 19576 3485
rect 19800 3519 19852 3528
rect 19800 3485 19834 3519
rect 19834 3485 19852 3519
rect 19800 3476 19852 3485
rect 20904 3476 20956 3528
rect 22744 3587 22796 3596
rect 22744 3553 22753 3587
rect 22753 3553 22787 3587
rect 22787 3553 22796 3587
rect 22744 3544 22796 3553
rect 22468 3519 22520 3528
rect 22468 3485 22477 3519
rect 22477 3485 22511 3519
rect 22511 3485 22520 3519
rect 25596 3612 25648 3664
rect 28264 3680 28316 3732
rect 26240 3544 26292 3596
rect 27252 3612 27304 3664
rect 27896 3655 27948 3664
rect 27896 3621 27905 3655
rect 27905 3621 27939 3655
rect 27939 3621 27948 3655
rect 27896 3612 27948 3621
rect 22468 3476 22520 3485
rect 25872 3476 25924 3528
rect 26056 3476 26108 3528
rect 27620 3544 27672 3596
rect 28356 3544 28408 3596
rect 16948 3408 17000 3417
rect 14280 3383 14332 3392
rect 14280 3349 14289 3383
rect 14289 3349 14323 3383
rect 14323 3349 14332 3383
rect 14280 3340 14332 3349
rect 18236 3340 18288 3392
rect 23388 3408 23440 3460
rect 25044 3408 25096 3460
rect 25964 3383 26016 3392
rect 25964 3349 25973 3383
rect 25973 3349 26007 3383
rect 26007 3349 26016 3383
rect 25964 3340 26016 3349
rect 26240 3340 26292 3392
rect 26608 3340 26660 3392
rect 9390 3238 9442 3290
rect 9454 3238 9506 3290
rect 9518 3238 9570 3290
rect 9582 3238 9634 3290
rect 9646 3238 9698 3290
rect 17831 3238 17883 3290
rect 17895 3238 17947 3290
rect 17959 3238 18011 3290
rect 18023 3238 18075 3290
rect 18087 3238 18139 3290
rect 26272 3238 26324 3290
rect 26336 3238 26388 3290
rect 26400 3238 26452 3290
rect 26464 3238 26516 3290
rect 26528 3238 26580 3290
rect 34713 3238 34765 3290
rect 34777 3238 34829 3290
rect 34841 3238 34893 3290
rect 34905 3238 34957 3290
rect 34969 3238 35021 3290
rect 12348 3136 12400 3188
rect 14372 3179 14424 3188
rect 14372 3145 14381 3179
rect 14381 3145 14415 3179
rect 14415 3145 14424 3179
rect 14372 3136 14424 3145
rect 14740 3179 14792 3188
rect 14740 3145 14749 3179
rect 14749 3145 14783 3179
rect 14783 3145 14792 3179
rect 14740 3136 14792 3145
rect 15660 3136 15712 3188
rect 16948 3179 17000 3188
rect 16948 3145 16957 3179
rect 16957 3145 16991 3179
rect 16991 3145 17000 3179
rect 16948 3136 17000 3145
rect 17040 3136 17092 3188
rect 18236 3136 18288 3188
rect 19524 3136 19576 3188
rect 20904 3136 20956 3188
rect 21088 3179 21140 3188
rect 21088 3145 21097 3179
rect 21097 3145 21131 3179
rect 21131 3145 21140 3179
rect 21088 3136 21140 3145
rect 29828 3136 29880 3188
rect 30380 3111 30432 3120
rect 10784 3000 10836 3052
rect 15200 3043 15252 3052
rect 15200 3009 15209 3043
rect 15209 3009 15243 3043
rect 15243 3009 15252 3043
rect 15200 3000 15252 3009
rect 30380 3077 30389 3111
rect 30389 3077 30423 3111
rect 30423 3077 30432 3111
rect 30380 3068 30432 3077
rect 20720 3000 20772 3052
rect 14188 2975 14240 2984
rect 14188 2941 14197 2975
rect 14197 2941 14231 2975
rect 14231 2941 14240 2975
rect 14188 2932 14240 2941
rect 14280 2975 14332 2984
rect 14280 2941 14289 2975
rect 14289 2941 14323 2975
rect 14323 2941 14332 2975
rect 14280 2932 14332 2941
rect 15476 2932 15528 2984
rect 20444 2932 20496 2984
rect 22744 3000 22796 3052
rect 26792 3000 26844 3052
rect 25964 2932 26016 2984
rect 26240 2932 26292 2984
rect 21180 2864 21232 2916
rect 24952 2864 25004 2916
rect 25596 2907 25648 2916
rect 25596 2873 25605 2907
rect 25605 2873 25639 2907
rect 25639 2873 25648 2907
rect 25596 2864 25648 2873
rect 26056 2864 26108 2916
rect 5170 2694 5222 2746
rect 5234 2694 5286 2746
rect 5298 2694 5350 2746
rect 5362 2694 5414 2746
rect 5426 2694 5478 2746
rect 13611 2694 13663 2746
rect 13675 2694 13727 2746
rect 13739 2694 13791 2746
rect 13803 2694 13855 2746
rect 13867 2694 13919 2746
rect 22052 2694 22104 2746
rect 22116 2694 22168 2746
rect 22180 2694 22232 2746
rect 22244 2694 22296 2746
rect 22308 2694 22360 2746
rect 30493 2694 30545 2746
rect 30557 2694 30609 2746
rect 30621 2694 30673 2746
rect 30685 2694 30737 2746
rect 30749 2694 30801 2746
rect 1216 2320 1268 2372
rect 2504 2320 2556 2372
rect 3792 2320 3844 2372
rect 15936 2592 15988 2644
rect 10048 2524 10100 2576
rect 5080 2320 5132 2372
rect 6368 2388 6420 2440
rect 7656 2388 7708 2440
rect 8944 2388 8996 2440
rect 10232 2388 10284 2440
rect 11520 2388 11572 2440
rect 12808 2388 12860 2440
rect 14004 2388 14056 2440
rect 15476 2431 15528 2440
rect 15476 2397 15485 2431
rect 15485 2397 15519 2431
rect 15519 2397 15528 2431
rect 15476 2388 15528 2397
rect 16304 2388 16356 2440
rect 18236 2456 18288 2508
rect 20904 2456 20956 2508
rect 19064 2388 19116 2440
rect 21088 2388 21140 2440
rect 23388 2388 23440 2440
rect 25596 2388 25648 2440
rect 26240 2431 26292 2440
rect 26240 2397 26249 2431
rect 26249 2397 26283 2431
rect 26283 2397 26292 2431
rect 26240 2388 26292 2397
rect 27896 2388 27948 2440
rect 28356 2431 28408 2440
rect 28356 2397 28365 2431
rect 28365 2397 28399 2431
rect 28399 2397 28408 2431
rect 28356 2388 28408 2397
rect 29552 2388 29604 2440
rect 30840 2388 30892 2440
rect 32128 2388 32180 2440
rect 33416 2388 33468 2440
rect 7840 2320 7892 2372
rect 14096 2320 14148 2372
rect 15384 2320 15436 2372
rect 16672 2320 16724 2372
rect 18236 2320 18288 2372
rect 19248 2320 19300 2372
rect 20536 2320 20588 2372
rect 21824 2320 21876 2372
rect 23112 2320 23164 2372
rect 24400 2320 24452 2372
rect 25688 2320 25740 2372
rect 26976 2320 27028 2372
rect 28264 2320 28316 2372
rect 14372 2252 14424 2304
rect 34612 2252 34664 2304
rect 9390 2150 9442 2202
rect 9454 2150 9506 2202
rect 9518 2150 9570 2202
rect 9582 2150 9634 2202
rect 9646 2150 9698 2202
rect 17831 2150 17883 2202
rect 17895 2150 17947 2202
rect 17959 2150 18011 2202
rect 18023 2150 18075 2202
rect 18087 2150 18139 2202
rect 26272 2150 26324 2202
rect 26336 2150 26388 2202
rect 26400 2150 26452 2202
rect 26464 2150 26516 2202
rect 26528 2150 26580 2202
rect 34713 2150 34765 2202
rect 34777 2150 34829 2202
rect 34841 2150 34893 2202
rect 34905 2150 34957 2202
rect 34969 2150 35021 2202
<< metal2 >>
rect 1766 35306 1822 36000
rect 1412 35278 1822 35306
rect 1412 14482 1440 35278
rect 1766 35200 1822 35278
rect 4710 35306 4766 36000
rect 7654 35306 7710 36000
rect 4710 35278 4936 35306
rect 4710 35200 4766 35278
rect 4908 33590 4936 35278
rect 7654 35278 7880 35306
rect 7654 35200 7710 35278
rect 7852 33590 7880 35278
rect 10598 35200 10654 36000
rect 13542 35306 13598 36000
rect 13542 35278 13768 35306
rect 13542 35200 13598 35278
rect 9390 33756 9698 33765
rect 9390 33754 9396 33756
rect 9452 33754 9476 33756
rect 9532 33754 9556 33756
rect 9612 33754 9636 33756
rect 9692 33754 9698 33756
rect 9452 33702 9454 33754
rect 9634 33702 9636 33754
rect 9390 33700 9396 33702
rect 9452 33700 9476 33702
rect 9532 33700 9556 33702
rect 9612 33700 9636 33702
rect 9692 33700 9698 33702
rect 9390 33691 9698 33700
rect 10612 33590 10640 35200
rect 4896 33584 4948 33590
rect 4896 33526 4948 33532
rect 7840 33584 7892 33590
rect 7840 33526 7892 33532
rect 10600 33584 10652 33590
rect 13740 33572 13768 35278
rect 16486 35200 16542 36000
rect 19430 35200 19486 36000
rect 22374 35306 22430 36000
rect 25318 35306 25374 36000
rect 22374 35278 22692 35306
rect 22374 35200 22430 35278
rect 13820 33584 13872 33590
rect 13740 33544 13820 33572
rect 10600 33526 10652 33532
rect 16500 33572 16528 35200
rect 17831 33756 18139 33765
rect 17831 33754 17837 33756
rect 17893 33754 17917 33756
rect 17973 33754 17997 33756
rect 18053 33754 18077 33756
rect 18133 33754 18139 33756
rect 17893 33702 17895 33754
rect 18075 33702 18077 33754
rect 17831 33700 17837 33702
rect 17893 33700 17917 33702
rect 17973 33700 17997 33702
rect 18053 33700 18077 33702
rect 18133 33700 18139 33702
rect 17831 33691 18139 33700
rect 19444 33590 19472 35200
rect 22664 33590 22692 35278
rect 25318 35278 25636 35306
rect 25318 35200 25374 35278
rect 25608 33590 25636 35278
rect 28262 35200 28318 36000
rect 31206 35306 31262 36000
rect 34150 35306 34206 36000
rect 31206 35278 31524 35306
rect 31206 35200 31262 35278
rect 26272 33756 26580 33765
rect 26272 33754 26278 33756
rect 26334 33754 26358 33756
rect 26414 33754 26438 33756
rect 26494 33754 26518 33756
rect 26574 33754 26580 33756
rect 26334 33702 26336 33754
rect 26516 33702 26518 33754
rect 26272 33700 26278 33702
rect 26334 33700 26358 33702
rect 26414 33700 26438 33702
rect 26494 33700 26518 33702
rect 26574 33700 26580 33702
rect 26272 33691 26580 33700
rect 28276 33590 28304 35200
rect 31496 33590 31524 35278
rect 34150 35278 34284 35306
rect 34150 35200 34206 35278
rect 34256 33590 34284 35278
rect 34713 33756 35021 33765
rect 34713 33754 34719 33756
rect 34775 33754 34799 33756
rect 34855 33754 34879 33756
rect 34935 33754 34959 33756
rect 35015 33754 35021 33756
rect 34775 33702 34777 33754
rect 34957 33702 34959 33754
rect 34713 33700 34719 33702
rect 34775 33700 34799 33702
rect 34855 33700 34879 33702
rect 34935 33700 34959 33702
rect 35015 33700 35021 33702
rect 34713 33691 35021 33700
rect 16580 33584 16632 33590
rect 16500 33544 16580 33572
rect 13820 33526 13872 33532
rect 16580 33526 16632 33532
rect 19432 33584 19484 33590
rect 19432 33526 19484 33532
rect 22652 33584 22704 33590
rect 22652 33526 22704 33532
rect 25596 33584 25648 33590
rect 25596 33526 25648 33532
rect 28264 33584 28316 33590
rect 28264 33526 28316 33532
rect 31484 33584 31536 33590
rect 31484 33526 31536 33532
rect 34244 33584 34296 33590
rect 34244 33526 34296 33532
rect 8024 33380 8076 33386
rect 8024 33322 8076 33328
rect 12256 33380 12308 33386
rect 12256 33322 12308 33328
rect 14280 33380 14332 33386
rect 14280 33322 14332 33328
rect 16856 33380 16908 33386
rect 16856 33322 16908 33328
rect 19524 33380 19576 33386
rect 19524 33322 19576 33328
rect 22468 33380 22520 33386
rect 22468 33322 22520 33328
rect 25412 33380 25464 33386
rect 25412 33322 25464 33328
rect 28356 33380 28408 33386
rect 28356 33322 28408 33328
rect 31300 33380 31352 33386
rect 31300 33322 31352 33328
rect 33416 33380 33468 33386
rect 33416 33322 33468 33328
rect 4988 33312 5040 33318
rect 4988 33254 5040 33260
rect 3332 25356 3384 25362
rect 3332 25298 3384 25304
rect 3344 24818 3372 25298
rect 4160 25288 4212 25294
rect 4160 25230 4212 25236
rect 3976 25152 4028 25158
rect 3976 25094 4028 25100
rect 3332 24812 3384 24818
rect 3332 24754 3384 24760
rect 3240 24608 3292 24614
rect 3240 24550 3292 24556
rect 3252 24206 3280 24550
rect 3344 24410 3372 24754
rect 3700 24744 3752 24750
rect 3700 24686 3752 24692
rect 3712 24410 3740 24686
rect 3332 24404 3384 24410
rect 3332 24346 3384 24352
rect 3700 24404 3752 24410
rect 3700 24346 3752 24352
rect 3988 24274 4016 25094
rect 4068 24744 4120 24750
rect 4068 24686 4120 24692
rect 3976 24268 4028 24274
rect 3976 24210 4028 24216
rect 3240 24200 3292 24206
rect 3240 24142 3292 24148
rect 3792 24200 3844 24206
rect 3792 24142 3844 24148
rect 2596 24132 2648 24138
rect 2596 24074 2648 24080
rect 2608 23866 2636 24074
rect 2596 23860 2648 23866
rect 2596 23802 2648 23808
rect 3252 23594 3280 24142
rect 3424 23724 3476 23730
rect 3424 23666 3476 23672
rect 3240 23588 3292 23594
rect 3240 23530 3292 23536
rect 3252 22710 3280 23530
rect 3436 23118 3464 23666
rect 3424 23112 3476 23118
rect 3424 23054 3476 23060
rect 3240 22704 3292 22710
rect 3240 22646 3292 22652
rect 3804 22438 3832 24142
rect 4080 23526 4108 24686
rect 4172 24138 4200 25230
rect 4712 24880 4764 24886
rect 4712 24822 4764 24828
rect 4528 24744 4580 24750
rect 4528 24686 4580 24692
rect 4436 24200 4488 24206
rect 4436 24142 4488 24148
rect 4160 24132 4212 24138
rect 4160 24074 4212 24080
rect 4252 24132 4304 24138
rect 4252 24074 4304 24080
rect 4068 23520 4120 23526
rect 4068 23462 4120 23468
rect 3608 22432 3660 22438
rect 3608 22374 3660 22380
rect 3792 22432 3844 22438
rect 3792 22374 3844 22380
rect 3620 21554 3648 22374
rect 3608 21548 3660 21554
rect 3608 21490 3660 21496
rect 3700 21480 3752 21486
rect 3700 21422 3752 21428
rect 3712 21350 3740 21422
rect 3056 21344 3108 21350
rect 3056 21286 3108 21292
rect 3608 21344 3660 21350
rect 3608 21286 3660 21292
rect 3700 21344 3752 21350
rect 3700 21286 3752 21292
rect 3068 20398 3096 21286
rect 3240 20936 3292 20942
rect 3240 20878 3292 20884
rect 3148 20800 3200 20806
rect 3148 20742 3200 20748
rect 3160 20466 3188 20742
rect 3148 20460 3200 20466
rect 3148 20402 3200 20408
rect 3056 20392 3108 20398
rect 3056 20334 3108 20340
rect 1860 20324 1912 20330
rect 1860 20266 1912 20272
rect 1872 19854 1900 20266
rect 2780 20256 2832 20262
rect 2780 20198 2832 20204
rect 1860 19848 1912 19854
rect 1860 19790 1912 19796
rect 2792 19378 2820 20198
rect 3252 19786 3280 20878
rect 3620 20534 3648 21286
rect 3608 20528 3660 20534
rect 3608 20470 3660 20476
rect 3424 20392 3476 20398
rect 3424 20334 3476 20340
rect 3240 19780 3292 19786
rect 3240 19722 3292 19728
rect 3332 19712 3384 19718
rect 3332 19654 3384 19660
rect 2780 19372 2832 19378
rect 2780 19314 2832 19320
rect 2964 18896 3016 18902
rect 2964 18838 3016 18844
rect 2688 17604 2740 17610
rect 2688 17546 2740 17552
rect 2700 17134 2728 17546
rect 2976 17270 3004 18838
rect 3344 18766 3372 19654
rect 3436 18766 3464 20334
rect 3804 19990 3832 22374
rect 4080 22094 4108 23462
rect 4172 23322 4200 24074
rect 4160 23316 4212 23322
rect 4160 23258 4212 23264
rect 4264 23186 4292 24074
rect 4344 23792 4396 23798
rect 4344 23734 4396 23740
rect 4252 23180 4304 23186
rect 4252 23122 4304 23128
rect 4356 22438 4384 23734
rect 4448 23254 4476 24142
rect 4540 23798 4568 24686
rect 4724 24206 4752 24822
rect 4712 24200 4764 24206
rect 4712 24142 4764 24148
rect 4528 23792 4580 23798
rect 4528 23734 4580 23740
rect 4436 23248 4488 23254
rect 4436 23190 4488 23196
rect 4344 22432 4396 22438
rect 4344 22374 4396 22380
rect 3896 22066 4108 22094
rect 3792 19984 3844 19990
rect 3792 19926 3844 19932
rect 3896 19378 3924 22066
rect 4448 21486 4476 23190
rect 4540 22778 4568 23734
rect 4724 23186 4752 24142
rect 4896 24064 4948 24070
rect 4896 24006 4948 24012
rect 4712 23180 4764 23186
rect 4712 23122 4764 23128
rect 4528 22772 4580 22778
rect 4528 22714 4580 22720
rect 4908 22642 4936 24006
rect 4896 22636 4948 22642
rect 4896 22578 4948 22584
rect 5000 22506 5028 33254
rect 5170 33212 5478 33221
rect 5170 33210 5176 33212
rect 5232 33210 5256 33212
rect 5312 33210 5336 33212
rect 5392 33210 5416 33212
rect 5472 33210 5478 33212
rect 5232 33158 5234 33210
rect 5414 33158 5416 33210
rect 5170 33156 5176 33158
rect 5232 33156 5256 33158
rect 5312 33156 5336 33158
rect 5392 33156 5416 33158
rect 5472 33156 5478 33158
rect 5170 33147 5478 33156
rect 5170 32124 5478 32133
rect 5170 32122 5176 32124
rect 5232 32122 5256 32124
rect 5312 32122 5336 32124
rect 5392 32122 5416 32124
rect 5472 32122 5478 32124
rect 5232 32070 5234 32122
rect 5414 32070 5416 32122
rect 5170 32068 5176 32070
rect 5232 32068 5256 32070
rect 5312 32068 5336 32070
rect 5392 32068 5416 32070
rect 5472 32068 5478 32070
rect 5170 32059 5478 32068
rect 8036 31686 8064 33322
rect 10508 32904 10560 32910
rect 10508 32846 10560 32852
rect 10140 32768 10192 32774
rect 10140 32710 10192 32716
rect 9390 32668 9698 32677
rect 9390 32666 9396 32668
rect 9452 32666 9476 32668
rect 9532 32666 9556 32668
rect 9612 32666 9636 32668
rect 9692 32666 9698 32668
rect 9452 32614 9454 32666
rect 9634 32614 9636 32666
rect 9390 32612 9396 32614
rect 9452 32612 9476 32614
rect 9532 32612 9556 32614
rect 9612 32612 9636 32614
rect 9692 32612 9698 32614
rect 9390 32603 9698 32612
rect 8576 32292 8628 32298
rect 8576 32234 8628 32240
rect 8588 31958 8616 32234
rect 10048 32224 10100 32230
rect 10048 32166 10100 32172
rect 8576 31952 8628 31958
rect 8576 31894 8628 31900
rect 8760 31952 8812 31958
rect 8760 31894 8812 31900
rect 8024 31680 8076 31686
rect 8024 31622 8076 31628
rect 5170 31036 5478 31045
rect 5170 31034 5176 31036
rect 5232 31034 5256 31036
rect 5312 31034 5336 31036
rect 5392 31034 5416 31036
rect 5472 31034 5478 31036
rect 5232 30982 5234 31034
rect 5414 30982 5416 31034
rect 5170 30980 5176 30982
rect 5232 30980 5256 30982
rect 5312 30980 5336 30982
rect 5392 30980 5416 30982
rect 5472 30980 5478 30982
rect 5170 30971 5478 30980
rect 5170 29948 5478 29957
rect 5170 29946 5176 29948
rect 5232 29946 5256 29948
rect 5312 29946 5336 29948
rect 5392 29946 5416 29948
rect 5472 29946 5478 29948
rect 5232 29894 5234 29946
rect 5414 29894 5416 29946
rect 5170 29892 5176 29894
rect 5232 29892 5256 29894
rect 5312 29892 5336 29894
rect 5392 29892 5416 29894
rect 5472 29892 5478 29894
rect 5170 29883 5478 29892
rect 7748 28960 7800 28966
rect 7748 28902 7800 28908
rect 5170 28860 5478 28869
rect 5170 28858 5176 28860
rect 5232 28858 5256 28860
rect 5312 28858 5336 28860
rect 5392 28858 5416 28860
rect 5472 28858 5478 28860
rect 5232 28806 5234 28858
rect 5414 28806 5416 28858
rect 5170 28804 5176 28806
rect 5232 28804 5256 28806
rect 5312 28804 5336 28806
rect 5392 28804 5416 28806
rect 5472 28804 5478 28806
rect 5170 28795 5478 28804
rect 7760 28558 7788 28902
rect 7748 28552 7800 28558
rect 7748 28494 7800 28500
rect 7760 28082 7788 28494
rect 8772 28082 8800 31894
rect 9864 31884 9916 31890
rect 9864 31826 9916 31832
rect 9390 31580 9698 31589
rect 9390 31578 9396 31580
rect 9452 31578 9476 31580
rect 9532 31578 9556 31580
rect 9612 31578 9636 31580
rect 9692 31578 9698 31580
rect 9452 31526 9454 31578
rect 9634 31526 9636 31578
rect 9390 31524 9396 31526
rect 9452 31524 9476 31526
rect 9532 31524 9556 31526
rect 9612 31524 9636 31526
rect 9692 31524 9698 31526
rect 9390 31515 9698 31524
rect 9876 31482 9904 31826
rect 10060 31754 10088 32166
rect 10152 31822 10180 32710
rect 10520 32434 10548 32846
rect 12268 32570 12296 33322
rect 13611 33212 13919 33221
rect 13611 33210 13617 33212
rect 13673 33210 13697 33212
rect 13753 33210 13777 33212
rect 13833 33210 13857 33212
rect 13913 33210 13919 33212
rect 13673 33158 13675 33210
rect 13855 33158 13857 33210
rect 13611 33156 13617 33158
rect 13673 33156 13697 33158
rect 13753 33156 13777 33158
rect 13833 33156 13857 33158
rect 13913 33156 13919 33158
rect 13611 33147 13919 33156
rect 13268 32768 13320 32774
rect 13268 32710 13320 32716
rect 12256 32564 12308 32570
rect 12256 32506 12308 32512
rect 13280 32502 13308 32710
rect 14292 32570 14320 33322
rect 16868 32978 16896 33322
rect 16856 32972 16908 32978
rect 16856 32914 16908 32920
rect 16212 32836 16264 32842
rect 16212 32778 16264 32784
rect 16764 32836 16816 32842
rect 16764 32778 16816 32784
rect 14280 32564 14332 32570
rect 14280 32506 14332 32512
rect 10692 32496 10744 32502
rect 10692 32438 10744 32444
rect 13268 32496 13320 32502
rect 13268 32438 13320 32444
rect 10508 32428 10560 32434
rect 10508 32370 10560 32376
rect 10520 32026 10548 32370
rect 10600 32224 10652 32230
rect 10600 32166 10652 32172
rect 10508 32020 10560 32026
rect 10508 31962 10560 31968
rect 10140 31816 10192 31822
rect 10140 31758 10192 31764
rect 10048 31748 10100 31754
rect 10048 31690 10100 31696
rect 9864 31476 9916 31482
rect 9864 31418 9916 31424
rect 10060 31414 10088 31690
rect 10048 31408 10100 31414
rect 10048 31350 10100 31356
rect 9864 31340 9916 31346
rect 9864 31282 9916 31288
rect 10232 31340 10284 31346
rect 10232 31282 10284 31288
rect 9404 31272 9456 31278
rect 9404 31214 9456 31220
rect 9416 30938 9444 31214
rect 9404 30932 9456 30938
rect 9404 30874 9456 30880
rect 9390 30492 9698 30501
rect 9390 30490 9396 30492
rect 9452 30490 9476 30492
rect 9532 30490 9556 30492
rect 9612 30490 9636 30492
rect 9692 30490 9698 30492
rect 9452 30438 9454 30490
rect 9634 30438 9636 30490
rect 9390 30436 9396 30438
rect 9452 30436 9476 30438
rect 9532 30436 9556 30438
rect 9612 30436 9636 30438
rect 9692 30436 9698 30438
rect 9390 30427 9698 30436
rect 9312 29504 9364 29510
rect 9312 29446 9364 29452
rect 9324 29170 9352 29446
rect 9390 29404 9698 29413
rect 9390 29402 9396 29404
rect 9452 29402 9476 29404
rect 9532 29402 9556 29404
rect 9612 29402 9636 29404
rect 9692 29402 9698 29404
rect 9452 29350 9454 29402
rect 9634 29350 9636 29402
rect 9390 29348 9396 29350
rect 9452 29348 9476 29350
rect 9532 29348 9556 29350
rect 9612 29348 9636 29350
rect 9692 29348 9698 29350
rect 9390 29339 9698 29348
rect 9312 29164 9364 29170
rect 9312 29106 9364 29112
rect 9312 28960 9364 28966
rect 9312 28902 9364 28908
rect 9324 28558 9352 28902
rect 9036 28552 9088 28558
rect 9036 28494 9088 28500
rect 9312 28552 9364 28558
rect 9312 28494 9364 28500
rect 9048 28082 9076 28494
rect 9220 28416 9272 28422
rect 9220 28358 9272 28364
rect 7748 28076 7800 28082
rect 7748 28018 7800 28024
rect 8760 28076 8812 28082
rect 8760 28018 8812 28024
rect 9036 28076 9088 28082
rect 9036 28018 9088 28024
rect 5170 27772 5478 27781
rect 5170 27770 5176 27772
rect 5232 27770 5256 27772
rect 5312 27770 5336 27772
rect 5392 27770 5416 27772
rect 5472 27770 5478 27772
rect 5232 27718 5234 27770
rect 5414 27718 5416 27770
rect 5170 27716 5176 27718
rect 5232 27716 5256 27718
rect 5312 27716 5336 27718
rect 5392 27716 5416 27718
rect 5472 27716 5478 27718
rect 5170 27707 5478 27716
rect 8208 27328 8260 27334
rect 8208 27270 8260 27276
rect 8220 26994 8248 27270
rect 8772 27062 8800 28018
rect 9128 27872 9180 27878
rect 9128 27814 9180 27820
rect 9140 27470 9168 27814
rect 9128 27464 9180 27470
rect 9128 27406 9180 27412
rect 8760 27056 8812 27062
rect 8760 26998 8812 27004
rect 9232 26994 9260 28358
rect 9324 28014 9352 28494
rect 9390 28316 9698 28325
rect 9390 28314 9396 28316
rect 9452 28314 9476 28316
rect 9532 28314 9556 28316
rect 9612 28314 9636 28316
rect 9692 28314 9698 28316
rect 9452 28262 9454 28314
rect 9634 28262 9636 28314
rect 9390 28260 9396 28262
rect 9452 28260 9476 28262
rect 9532 28260 9556 28262
rect 9612 28260 9636 28262
rect 9692 28260 9698 28262
rect 9390 28251 9698 28260
rect 9876 28218 9904 31282
rect 10048 31272 10100 31278
rect 10048 31214 10100 31220
rect 10060 30938 10088 31214
rect 10244 30938 10272 31282
rect 10416 31272 10468 31278
rect 10416 31214 10468 31220
rect 10048 30932 10100 30938
rect 10048 30874 10100 30880
rect 10232 30932 10284 30938
rect 10232 30874 10284 30880
rect 9956 30728 10008 30734
rect 9956 30670 10008 30676
rect 9968 29714 9996 30670
rect 10428 30666 10456 31214
rect 10520 30802 10548 31962
rect 10612 31414 10640 32166
rect 10600 31408 10652 31414
rect 10600 31350 10652 31356
rect 10704 31142 10732 32438
rect 12348 32360 12400 32366
rect 14004 32360 14056 32366
rect 12348 32302 12400 32308
rect 11980 32224 12032 32230
rect 11980 32166 12032 32172
rect 11704 31952 11756 31958
rect 11704 31894 11756 31900
rect 10968 31204 11020 31210
rect 10968 31146 11020 31152
rect 10692 31136 10744 31142
rect 10692 31078 10744 31084
rect 10508 30796 10560 30802
rect 10508 30738 10560 30744
rect 10704 30734 10732 31078
rect 10692 30728 10744 30734
rect 10692 30670 10744 30676
rect 10416 30660 10468 30666
rect 10416 30602 10468 30608
rect 10508 30660 10560 30666
rect 10508 30602 10560 30608
rect 9956 29708 10008 29714
rect 9956 29650 10008 29656
rect 10324 29504 10376 29510
rect 10324 29446 10376 29452
rect 10336 29102 10364 29446
rect 10324 29096 10376 29102
rect 10324 29038 10376 29044
rect 10428 28966 10456 30602
rect 10520 29850 10548 30602
rect 10508 29844 10560 29850
rect 10508 29786 10560 29792
rect 10520 29646 10548 29786
rect 10508 29640 10560 29646
rect 10508 29582 10560 29588
rect 10416 28960 10468 28966
rect 10416 28902 10468 28908
rect 9864 28212 9916 28218
rect 9864 28154 9916 28160
rect 9312 28008 9364 28014
rect 9312 27950 9364 27956
rect 9312 27872 9364 27878
rect 9312 27814 9364 27820
rect 9588 27872 9640 27878
rect 9588 27814 9640 27820
rect 8208 26988 8260 26994
rect 8208 26930 8260 26936
rect 9220 26988 9272 26994
rect 9220 26930 9272 26936
rect 9220 26784 9272 26790
rect 9220 26726 9272 26732
rect 5170 26684 5478 26693
rect 5170 26682 5176 26684
rect 5232 26682 5256 26684
rect 5312 26682 5336 26684
rect 5392 26682 5416 26684
rect 5472 26682 5478 26684
rect 5232 26630 5234 26682
rect 5414 26630 5416 26682
rect 5170 26628 5176 26630
rect 5232 26628 5256 26630
rect 5312 26628 5336 26630
rect 5392 26628 5416 26630
rect 5472 26628 5478 26630
rect 5170 26619 5478 26628
rect 9232 25838 9260 26726
rect 9324 26518 9352 27814
rect 9600 27470 9628 27814
rect 9588 27464 9640 27470
rect 9588 27406 9640 27412
rect 9772 27396 9824 27402
rect 9772 27338 9824 27344
rect 9390 27228 9698 27237
rect 9390 27226 9396 27228
rect 9452 27226 9476 27228
rect 9532 27226 9556 27228
rect 9612 27226 9636 27228
rect 9692 27226 9698 27228
rect 9452 27174 9454 27226
rect 9634 27174 9636 27226
rect 9390 27172 9396 27174
rect 9452 27172 9476 27174
rect 9532 27172 9556 27174
rect 9612 27172 9636 27174
rect 9692 27172 9698 27174
rect 9390 27163 9698 27172
rect 9312 26512 9364 26518
rect 9312 26454 9364 26460
rect 9784 26314 9812 27338
rect 10704 26926 10732 30670
rect 10980 29578 11008 31146
rect 10968 29572 11020 29578
rect 10968 29514 11020 29520
rect 10980 28558 11008 29514
rect 11060 29164 11112 29170
rect 11060 29106 11112 29112
rect 11072 28694 11100 29106
rect 11060 28688 11112 28694
rect 11060 28630 11112 28636
rect 10968 28552 11020 28558
rect 10968 28494 11020 28500
rect 10980 28150 11008 28494
rect 10968 28144 11020 28150
rect 10968 28086 11020 28092
rect 10692 26920 10744 26926
rect 10692 26862 10744 26868
rect 11152 26784 11204 26790
rect 11152 26726 11204 26732
rect 11164 26450 11192 26726
rect 11152 26444 11204 26450
rect 11152 26386 11204 26392
rect 9772 26308 9824 26314
rect 9772 26250 9824 26256
rect 9312 26240 9364 26246
rect 9312 26182 9364 26188
rect 9324 25974 9352 26182
rect 9390 26140 9698 26149
rect 9390 26138 9396 26140
rect 9452 26138 9476 26140
rect 9532 26138 9556 26140
rect 9612 26138 9636 26140
rect 9692 26138 9698 26140
rect 9452 26086 9454 26138
rect 9634 26086 9636 26138
rect 9390 26084 9396 26086
rect 9452 26084 9476 26086
rect 9532 26084 9556 26086
rect 9612 26084 9636 26086
rect 9692 26084 9698 26086
rect 9390 26075 9698 26084
rect 9772 26036 9824 26042
rect 9772 25978 9824 25984
rect 9312 25968 9364 25974
rect 9312 25910 9364 25916
rect 9784 25906 9812 25978
rect 9772 25900 9824 25906
rect 9772 25842 9824 25848
rect 10416 25900 10468 25906
rect 10416 25842 10468 25848
rect 9220 25832 9272 25838
rect 9220 25774 9272 25780
rect 10428 25770 10456 25842
rect 10416 25764 10468 25770
rect 10416 25706 10468 25712
rect 5170 25596 5478 25605
rect 5170 25594 5176 25596
rect 5232 25594 5256 25596
rect 5312 25594 5336 25596
rect 5392 25594 5416 25596
rect 5472 25594 5478 25596
rect 5232 25542 5234 25594
rect 5414 25542 5416 25594
rect 5170 25540 5176 25542
rect 5232 25540 5256 25542
rect 5312 25540 5336 25542
rect 5392 25540 5416 25542
rect 5472 25540 5478 25542
rect 5170 25531 5478 25540
rect 6828 25288 6880 25294
rect 6828 25230 6880 25236
rect 7472 25288 7524 25294
rect 7472 25230 7524 25236
rect 5080 25152 5132 25158
rect 5080 25094 5132 25100
rect 5092 24290 5120 25094
rect 6840 24818 6868 25230
rect 7484 24818 7512 25230
rect 10232 25220 10284 25226
rect 10232 25162 10284 25168
rect 9390 25052 9698 25061
rect 9390 25050 9396 25052
rect 9452 25050 9476 25052
rect 9532 25050 9556 25052
rect 9612 25050 9636 25052
rect 9692 25050 9698 25052
rect 9452 24998 9454 25050
rect 9634 24998 9636 25050
rect 9390 24996 9396 24998
rect 9452 24996 9476 24998
rect 9532 24996 9556 24998
rect 9612 24996 9636 24998
rect 9692 24996 9698 24998
rect 9390 24987 9698 24996
rect 6828 24812 6880 24818
rect 6828 24754 6880 24760
rect 7472 24812 7524 24818
rect 7472 24754 7524 24760
rect 5170 24508 5478 24517
rect 5170 24506 5176 24508
rect 5232 24506 5256 24508
rect 5312 24506 5336 24508
rect 5392 24506 5416 24508
rect 5472 24506 5478 24508
rect 5232 24454 5234 24506
rect 5414 24454 5416 24506
rect 5170 24452 5176 24454
rect 5232 24452 5256 24454
rect 5312 24452 5336 24454
rect 5392 24452 5416 24454
rect 5472 24452 5478 24454
rect 5170 24443 5478 24452
rect 6840 24410 6868 24754
rect 6828 24404 6880 24410
rect 6828 24346 6880 24352
rect 5092 24274 5212 24290
rect 5092 24268 5224 24274
rect 5092 24262 5172 24268
rect 5092 23118 5120 24262
rect 5172 24210 5224 24216
rect 7196 24200 7248 24206
rect 7196 24142 7248 24148
rect 6748 23730 7052 23746
rect 6736 23724 7052 23730
rect 6788 23718 7052 23724
rect 6736 23666 6788 23672
rect 6644 23656 6696 23662
rect 6644 23598 6696 23604
rect 5170 23420 5478 23429
rect 5170 23418 5176 23420
rect 5232 23418 5256 23420
rect 5312 23418 5336 23420
rect 5392 23418 5416 23420
rect 5472 23418 5478 23420
rect 5232 23366 5234 23418
rect 5414 23366 5416 23418
rect 5170 23364 5176 23366
rect 5232 23364 5256 23366
rect 5312 23364 5336 23366
rect 5392 23364 5416 23366
rect 5472 23364 5478 23366
rect 5170 23355 5478 23364
rect 6656 23254 6684 23598
rect 6644 23248 6696 23254
rect 6644 23190 6696 23196
rect 5080 23112 5132 23118
rect 5080 23054 5132 23060
rect 4988 22500 5040 22506
rect 4988 22442 5040 22448
rect 4620 22432 4672 22438
rect 4620 22374 4672 22380
rect 4436 21480 4488 21486
rect 4436 21422 4488 21428
rect 4068 21412 4120 21418
rect 4068 21354 4120 21360
rect 3976 20460 4028 20466
rect 3976 20402 4028 20408
rect 3988 20058 4016 20402
rect 4080 20398 4108 21354
rect 4632 21026 4660 22374
rect 5170 22332 5478 22341
rect 5170 22330 5176 22332
rect 5232 22330 5256 22332
rect 5312 22330 5336 22332
rect 5392 22330 5416 22332
rect 5472 22330 5478 22332
rect 5232 22278 5234 22330
rect 5414 22278 5416 22330
rect 5170 22276 5176 22278
rect 5232 22276 5256 22278
rect 5312 22276 5336 22278
rect 5392 22276 5416 22278
rect 5472 22276 5478 22278
rect 5170 22267 5478 22276
rect 6656 22166 6684 23190
rect 7024 23050 7052 23718
rect 7104 23656 7156 23662
rect 7104 23598 7156 23604
rect 7116 23322 7144 23598
rect 7104 23316 7156 23322
rect 7104 23258 7156 23264
rect 7104 23112 7156 23118
rect 7104 23054 7156 23060
rect 7012 23044 7064 23050
rect 7012 22986 7064 22992
rect 7024 22522 7052 22986
rect 7116 22710 7144 23054
rect 7104 22704 7156 22710
rect 7104 22646 7156 22652
rect 7024 22494 7144 22522
rect 6644 22160 6696 22166
rect 6644 22102 6696 22108
rect 5170 21244 5478 21253
rect 5170 21242 5176 21244
rect 5232 21242 5256 21244
rect 5312 21242 5336 21244
rect 5392 21242 5416 21244
rect 5472 21242 5478 21244
rect 5232 21190 5234 21242
rect 5414 21190 5416 21242
rect 5170 21188 5176 21190
rect 5232 21188 5256 21190
rect 5312 21188 5336 21190
rect 5392 21188 5416 21190
rect 5472 21188 5478 21190
rect 5170 21179 5478 21188
rect 4448 20998 4660 21026
rect 4448 20942 4476 20998
rect 4436 20936 4488 20942
rect 4436 20878 4488 20884
rect 4068 20392 4120 20398
rect 4068 20334 4120 20340
rect 4344 20392 4396 20398
rect 4344 20334 4396 20340
rect 3976 20052 4028 20058
rect 3976 19994 4028 20000
rect 4356 19922 4384 20334
rect 4344 19916 4396 19922
rect 4344 19858 4396 19864
rect 4160 19848 4212 19854
rect 4080 19808 4160 19836
rect 3976 19780 4028 19786
rect 4080 19768 4108 19808
rect 4160 19790 4212 19796
rect 4028 19740 4108 19768
rect 3976 19722 4028 19728
rect 4080 19514 4108 19740
rect 4252 19780 4304 19786
rect 4252 19722 4304 19728
rect 4068 19508 4120 19514
rect 4068 19450 4120 19456
rect 3516 19372 3568 19378
rect 3516 19314 3568 19320
rect 3884 19372 3936 19378
rect 3884 19314 3936 19320
rect 3332 18760 3384 18766
rect 3332 18702 3384 18708
rect 3424 18760 3476 18766
rect 3424 18702 3476 18708
rect 3240 18692 3292 18698
rect 3240 18634 3292 18640
rect 3252 17678 3280 18634
rect 3528 17814 3556 19314
rect 4264 19174 4292 19722
rect 4448 19718 4476 20878
rect 5080 20324 5132 20330
rect 5080 20266 5132 20272
rect 5092 20058 5120 20266
rect 5170 20156 5478 20165
rect 5170 20154 5176 20156
rect 5232 20154 5256 20156
rect 5312 20154 5336 20156
rect 5392 20154 5416 20156
rect 5472 20154 5478 20156
rect 5232 20102 5234 20154
rect 5414 20102 5416 20154
rect 5170 20100 5176 20102
rect 5232 20100 5256 20102
rect 5312 20100 5336 20102
rect 5392 20100 5416 20102
rect 5472 20100 5478 20102
rect 5170 20091 5478 20100
rect 6656 20074 6684 22102
rect 7116 22030 7144 22494
rect 7104 22024 7156 22030
rect 7104 21966 7156 21972
rect 7208 21894 7236 24142
rect 7288 24132 7340 24138
rect 7288 24074 7340 24080
rect 7300 23526 7328 24074
rect 7484 23662 7512 24754
rect 8484 24744 8536 24750
rect 8484 24686 8536 24692
rect 8300 24132 8352 24138
rect 8300 24074 8352 24080
rect 7564 24064 7616 24070
rect 7564 24006 7616 24012
rect 7472 23656 7524 23662
rect 7472 23598 7524 23604
rect 7288 23520 7340 23526
rect 7288 23462 7340 23468
rect 7300 23118 7328 23462
rect 7288 23112 7340 23118
rect 7288 23054 7340 23060
rect 7484 22642 7512 23598
rect 7576 23322 7604 24006
rect 8312 23866 8340 24074
rect 8300 23860 8352 23866
rect 8300 23802 8352 23808
rect 8496 23798 8524 24686
rect 9220 24336 9272 24342
rect 9220 24278 9272 24284
rect 8576 23860 8628 23866
rect 8576 23802 8628 23808
rect 8484 23792 8536 23798
rect 8484 23734 8536 23740
rect 8300 23520 8352 23526
rect 8300 23462 8352 23468
rect 7564 23316 7616 23322
rect 7564 23258 7616 23264
rect 7564 23112 7616 23118
rect 7564 23054 7616 23060
rect 8116 23112 8168 23118
rect 8116 23054 8168 23060
rect 7576 22778 7604 23054
rect 8128 22982 8156 23054
rect 8116 22976 8168 22982
rect 8116 22918 8168 22924
rect 7564 22772 7616 22778
rect 7564 22714 7616 22720
rect 8312 22710 8340 23462
rect 8496 22710 8524 23734
rect 8588 23254 8616 23802
rect 9232 23730 9260 24278
rect 9312 24200 9364 24206
rect 9312 24142 9364 24148
rect 8944 23724 8996 23730
rect 8944 23666 8996 23672
rect 9220 23724 9272 23730
rect 9220 23666 9272 23672
rect 8576 23248 8628 23254
rect 8576 23190 8628 23196
rect 8852 23180 8904 23186
rect 8852 23122 8904 23128
rect 8300 22704 8352 22710
rect 8300 22646 8352 22652
rect 8484 22704 8536 22710
rect 8484 22646 8536 22652
rect 7472 22636 7524 22642
rect 7472 22578 7524 22584
rect 7472 22024 7524 22030
rect 7472 21966 7524 21972
rect 7196 21888 7248 21894
rect 7196 21830 7248 21836
rect 6920 20324 6972 20330
rect 6920 20266 6972 20272
rect 4712 20052 4764 20058
rect 4712 19994 4764 20000
rect 5080 20052 5132 20058
rect 5080 19994 5132 20000
rect 6564 20046 6684 20074
rect 4620 19848 4672 19854
rect 4620 19790 4672 19796
rect 4436 19712 4488 19718
rect 4436 19654 4488 19660
rect 4252 19168 4304 19174
rect 4252 19110 4304 19116
rect 4448 19122 4476 19654
rect 4632 19242 4660 19790
rect 4724 19446 4752 19994
rect 5448 19848 5500 19854
rect 5448 19790 5500 19796
rect 4896 19508 4948 19514
rect 4896 19450 4948 19456
rect 4712 19440 4764 19446
rect 4712 19382 4764 19388
rect 4908 19378 4936 19450
rect 4804 19372 4856 19378
rect 4804 19314 4856 19320
rect 4896 19372 4948 19378
rect 4896 19314 4948 19320
rect 4620 19236 4672 19242
rect 4620 19178 4672 19184
rect 4816 19122 4844 19314
rect 5460 19174 5488 19790
rect 6564 19786 6592 20046
rect 6644 19984 6696 19990
rect 6644 19926 6696 19932
rect 6552 19780 6604 19786
rect 6552 19722 6604 19728
rect 4448 19094 4844 19122
rect 5448 19168 5500 19174
rect 5448 19110 5500 19116
rect 3516 17808 3568 17814
rect 3516 17750 3568 17756
rect 3240 17672 3292 17678
rect 3240 17614 3292 17620
rect 3056 17536 3108 17542
rect 3056 17478 3108 17484
rect 3148 17536 3200 17542
rect 3148 17478 3200 17484
rect 2964 17264 3016 17270
rect 2964 17206 3016 17212
rect 2688 17128 2740 17134
rect 2688 17070 2740 17076
rect 2700 16794 2728 17070
rect 2688 16788 2740 16794
rect 2688 16730 2740 16736
rect 3068 16522 3096 17478
rect 3160 16776 3188 17478
rect 4252 17196 4304 17202
rect 4252 17138 4304 17144
rect 4264 16794 4292 17138
rect 3240 16788 3292 16794
rect 3160 16748 3240 16776
rect 3240 16730 3292 16736
rect 4252 16788 4304 16794
rect 4252 16730 4304 16736
rect 3056 16516 3108 16522
rect 3056 16458 3108 16464
rect 2964 15428 3016 15434
rect 2964 15370 3016 15376
rect 2976 15094 3004 15370
rect 2964 15088 3016 15094
rect 2964 15030 3016 15036
rect 1676 14952 1728 14958
rect 1676 14894 1728 14900
rect 2688 14952 2740 14958
rect 2688 14894 2740 14900
rect 1400 14476 1452 14482
rect 1400 14418 1452 14424
rect 1688 14074 1716 14894
rect 2700 14414 2728 14894
rect 2964 14816 3016 14822
rect 2964 14758 3016 14764
rect 2688 14408 2740 14414
rect 2688 14350 2740 14356
rect 1676 14068 1728 14074
rect 1676 14010 1728 14016
rect 2976 13326 3004 14758
rect 3068 14414 3096 16458
rect 3252 14890 3280 16730
rect 4068 16584 4120 16590
rect 4068 16526 4120 16532
rect 4344 16584 4396 16590
rect 4344 16526 4396 16532
rect 4080 15502 4108 16526
rect 4356 15570 4384 16526
rect 4816 15706 4844 19094
rect 5170 19068 5478 19077
rect 5170 19066 5176 19068
rect 5232 19066 5256 19068
rect 5312 19066 5336 19068
rect 5392 19066 5416 19068
rect 5472 19066 5478 19068
rect 5232 19014 5234 19066
rect 5414 19014 5416 19066
rect 5170 19012 5176 19014
rect 5232 19012 5256 19014
rect 5312 19012 5336 19014
rect 5392 19012 5416 19014
rect 5472 19012 5478 19014
rect 5170 19003 5478 19012
rect 5170 17980 5478 17989
rect 5170 17978 5176 17980
rect 5232 17978 5256 17980
rect 5312 17978 5336 17980
rect 5392 17978 5416 17980
rect 5472 17978 5478 17980
rect 5232 17926 5234 17978
rect 5414 17926 5416 17978
rect 5170 17924 5176 17926
rect 5232 17924 5256 17926
rect 5312 17924 5336 17926
rect 5392 17924 5416 17926
rect 5472 17924 5478 17926
rect 5170 17915 5478 17924
rect 6564 17678 6592 19722
rect 6656 18290 6684 19926
rect 6932 19514 6960 20266
rect 7104 19984 7156 19990
rect 7104 19926 7156 19932
rect 6920 19508 6972 19514
rect 6920 19450 6972 19456
rect 7116 18834 7144 19926
rect 7104 18828 7156 18834
rect 7104 18770 7156 18776
rect 7208 18698 7236 21830
rect 7484 21554 7512 21966
rect 7472 21548 7524 21554
rect 7472 21490 7524 21496
rect 7484 21010 7512 21490
rect 7472 21004 7524 21010
rect 7472 20946 7524 20952
rect 7288 20936 7340 20942
rect 7288 20878 7340 20884
rect 7300 20466 7328 20878
rect 7380 20800 7432 20806
rect 7380 20742 7432 20748
rect 7288 20460 7340 20466
rect 7288 20402 7340 20408
rect 7300 19786 7328 20402
rect 7392 19854 7420 20742
rect 7380 19848 7432 19854
rect 7380 19790 7432 19796
rect 7288 19780 7340 19786
rect 7288 19722 7340 19728
rect 7196 18692 7248 18698
rect 7196 18634 7248 18640
rect 7196 18352 7248 18358
rect 7196 18294 7248 18300
rect 6644 18284 6696 18290
rect 6644 18226 6696 18232
rect 6368 17672 6420 17678
rect 6368 17614 6420 17620
rect 6552 17672 6604 17678
rect 6552 17614 6604 17620
rect 5170 16892 5478 16901
rect 5170 16890 5176 16892
rect 5232 16890 5256 16892
rect 5312 16890 5336 16892
rect 5392 16890 5416 16892
rect 5472 16890 5478 16892
rect 5232 16838 5234 16890
rect 5414 16838 5416 16890
rect 5170 16836 5176 16838
rect 5232 16836 5256 16838
rect 5312 16836 5336 16838
rect 5392 16836 5416 16838
rect 5472 16836 5478 16838
rect 5170 16827 5478 16836
rect 6276 16788 6328 16794
rect 6276 16730 6328 16736
rect 5724 16176 5776 16182
rect 5724 16118 5776 16124
rect 5540 15972 5592 15978
rect 5540 15914 5592 15920
rect 5170 15804 5478 15813
rect 5170 15802 5176 15804
rect 5232 15802 5256 15804
rect 5312 15802 5336 15804
rect 5392 15802 5416 15804
rect 5472 15802 5478 15804
rect 5232 15750 5234 15802
rect 5414 15750 5416 15802
rect 5170 15748 5176 15750
rect 5232 15748 5256 15750
rect 5312 15748 5336 15750
rect 5392 15748 5416 15750
rect 5472 15748 5478 15750
rect 5170 15739 5478 15748
rect 4804 15700 4856 15706
rect 4804 15642 4856 15648
rect 4344 15564 4396 15570
rect 4344 15506 4396 15512
rect 4068 15496 4120 15502
rect 4068 15438 4120 15444
rect 3240 14884 3292 14890
rect 3240 14826 3292 14832
rect 3056 14408 3108 14414
rect 3056 14350 3108 14356
rect 3068 13938 3096 14350
rect 3148 14340 3200 14346
rect 3148 14282 3200 14288
rect 3160 14074 3188 14282
rect 3148 14068 3200 14074
rect 3148 14010 3200 14016
rect 3160 13954 3188 14010
rect 3056 13932 3108 13938
rect 3160 13926 3280 13954
rect 3056 13874 3108 13880
rect 2964 13320 3016 13326
rect 2964 13262 3016 13268
rect 2412 13184 2464 13190
rect 2412 13126 2464 13132
rect 2424 12918 2452 13126
rect 2412 12912 2464 12918
rect 2412 12854 2464 12860
rect 2976 11218 3004 13262
rect 3068 12782 3096 13874
rect 3148 12912 3200 12918
rect 3148 12854 3200 12860
rect 3056 12776 3108 12782
rect 3056 12718 3108 12724
rect 3160 12442 3188 12854
rect 3148 12436 3200 12442
rect 3148 12378 3200 12384
rect 2964 11212 3016 11218
rect 2964 11154 3016 11160
rect 3252 11150 3280 13926
rect 4080 13802 4108 15438
rect 4160 13864 4212 13870
rect 4160 13806 4212 13812
rect 4068 13796 4120 13802
rect 4068 13738 4120 13744
rect 4172 13530 4200 13806
rect 4160 13524 4212 13530
rect 4160 13466 4212 13472
rect 4356 13394 4384 15506
rect 5552 15434 5580 15914
rect 5540 15428 5592 15434
rect 5540 15370 5592 15376
rect 4436 15360 4488 15366
rect 4436 15302 4488 15308
rect 4448 14006 4476 15302
rect 5736 15162 5764 16118
rect 6288 15502 6316 16730
rect 6380 16454 6408 17614
rect 6564 17218 6592 17614
rect 6472 17190 6592 17218
rect 6472 16590 6500 17190
rect 6656 17134 6684 18226
rect 6736 18216 6788 18222
rect 6736 18158 6788 18164
rect 6920 18216 6972 18222
rect 6920 18158 6972 18164
rect 6748 17882 6776 18158
rect 6736 17876 6788 17882
rect 6736 17818 6788 17824
rect 6932 17338 6960 18158
rect 6920 17332 6972 17338
rect 6920 17274 6972 17280
rect 6736 17196 6788 17202
rect 6736 17138 6788 17144
rect 6828 17196 6880 17202
rect 6828 17138 6880 17144
rect 6644 17128 6696 17134
rect 6564 17088 6644 17116
rect 6564 16658 6592 17088
rect 6644 17070 6696 17076
rect 6552 16652 6604 16658
rect 6552 16594 6604 16600
rect 6460 16584 6512 16590
rect 6460 16526 6512 16532
rect 6368 16448 6420 16454
rect 6368 16390 6420 16396
rect 6472 15978 6500 16526
rect 6552 16516 6604 16522
rect 6552 16458 6604 16464
rect 6564 16114 6592 16458
rect 6748 16250 6776 17138
rect 6736 16244 6788 16250
rect 6736 16186 6788 16192
rect 6552 16108 6604 16114
rect 6552 16050 6604 16056
rect 6460 15972 6512 15978
rect 6460 15914 6512 15920
rect 6564 15570 6592 16050
rect 6552 15564 6604 15570
rect 6552 15506 6604 15512
rect 6748 15502 6776 16186
rect 6840 16182 6868 17138
rect 6920 16788 6972 16794
rect 6920 16730 6972 16736
rect 6828 16176 6880 16182
rect 6828 16118 6880 16124
rect 6932 16114 6960 16730
rect 7208 16726 7236 18294
rect 7300 18154 7328 19722
rect 7484 19718 7512 20946
rect 7656 20936 7708 20942
rect 7656 20878 7708 20884
rect 7668 20058 7696 20878
rect 8312 20602 8340 22646
rect 8864 22642 8892 23122
rect 8852 22636 8904 22642
rect 8852 22578 8904 22584
rect 8864 21894 8892 22578
rect 8852 21888 8904 21894
rect 8852 21830 8904 21836
rect 8300 20596 8352 20602
rect 8300 20538 8352 20544
rect 7748 20528 7800 20534
rect 8956 20482 8984 23666
rect 9324 23118 9352 24142
rect 9390 23964 9698 23973
rect 9390 23962 9396 23964
rect 9452 23962 9476 23964
rect 9532 23962 9556 23964
rect 9612 23962 9636 23964
rect 9692 23962 9698 23964
rect 9452 23910 9454 23962
rect 9634 23910 9636 23962
rect 9390 23908 9396 23910
rect 9452 23908 9476 23910
rect 9532 23908 9556 23910
rect 9612 23908 9636 23910
rect 9692 23908 9698 23910
rect 9390 23899 9698 23908
rect 9404 23860 9456 23866
rect 9404 23802 9456 23808
rect 9416 23662 9444 23802
rect 9404 23656 9456 23662
rect 9404 23598 9456 23604
rect 9416 23322 9444 23598
rect 9404 23316 9456 23322
rect 9404 23258 9456 23264
rect 9864 23316 9916 23322
rect 9864 23258 9916 23264
rect 9312 23112 9364 23118
rect 9312 23054 9364 23060
rect 9324 22658 9352 23054
rect 9772 23044 9824 23050
rect 9772 22986 9824 22992
rect 9390 22876 9698 22885
rect 9390 22874 9396 22876
rect 9452 22874 9476 22876
rect 9532 22874 9556 22876
rect 9612 22874 9636 22876
rect 9692 22874 9698 22876
rect 9452 22822 9454 22874
rect 9634 22822 9636 22874
rect 9390 22820 9396 22822
rect 9452 22820 9476 22822
rect 9532 22820 9556 22822
rect 9612 22820 9636 22822
rect 9692 22820 9698 22822
rect 9390 22811 9698 22820
rect 9784 22710 9812 22986
rect 9772 22704 9824 22710
rect 9324 22642 9628 22658
rect 9772 22646 9824 22652
rect 9324 22636 9640 22642
rect 9324 22630 9588 22636
rect 9324 22030 9352 22630
rect 9588 22578 9640 22584
rect 9312 22024 9364 22030
rect 9312 21966 9364 21972
rect 9036 21888 9088 21894
rect 9036 21830 9088 21836
rect 7748 20470 7800 20476
rect 7656 20052 7708 20058
rect 7656 19994 7708 20000
rect 7760 19990 7788 20470
rect 8024 20460 8076 20466
rect 8024 20402 8076 20408
rect 8484 20460 8536 20466
rect 8484 20402 8536 20408
rect 8864 20454 8984 20482
rect 7840 20324 7892 20330
rect 7840 20266 7892 20272
rect 7748 19984 7800 19990
rect 7748 19926 7800 19932
rect 7472 19712 7524 19718
rect 7472 19654 7524 19660
rect 7288 18148 7340 18154
rect 7288 18090 7340 18096
rect 7484 17202 7512 19654
rect 7656 19372 7708 19378
rect 7656 19314 7708 19320
rect 7668 18970 7696 19314
rect 7656 18964 7708 18970
rect 7656 18906 7708 18912
rect 7472 17196 7524 17202
rect 7472 17138 7524 17144
rect 7748 17196 7800 17202
rect 7748 17138 7800 17144
rect 7196 16720 7248 16726
rect 7196 16662 7248 16668
rect 6920 16108 6972 16114
rect 6920 16050 6972 16056
rect 7208 16046 7236 16662
rect 7380 16108 7432 16114
rect 7380 16050 7432 16056
rect 7472 16108 7524 16114
rect 7472 16050 7524 16056
rect 7196 16040 7248 16046
rect 7196 15982 7248 15988
rect 6092 15496 6144 15502
rect 6092 15438 6144 15444
rect 6276 15496 6328 15502
rect 6276 15438 6328 15444
rect 6736 15496 6788 15502
rect 6736 15438 6788 15444
rect 5724 15156 5776 15162
rect 5724 15098 5776 15104
rect 4528 15020 4580 15026
rect 4528 14962 4580 14968
rect 4436 14000 4488 14006
rect 4436 13942 4488 13948
rect 4344 13388 4396 13394
rect 4344 13330 4396 13336
rect 3884 13320 3936 13326
rect 3884 13262 3936 13268
rect 3424 13252 3476 13258
rect 3424 13194 3476 13200
rect 3436 12238 3464 13194
rect 3896 12782 3924 13262
rect 4356 12986 4384 13330
rect 4436 13184 4488 13190
rect 4436 13126 4488 13132
rect 4448 12986 4476 13126
rect 4344 12980 4396 12986
rect 4344 12922 4396 12928
rect 4436 12980 4488 12986
rect 4436 12922 4488 12928
rect 3976 12844 4028 12850
rect 3976 12786 4028 12792
rect 3884 12776 3936 12782
rect 3884 12718 3936 12724
rect 3424 12232 3476 12238
rect 3424 12174 3476 12180
rect 3332 11212 3384 11218
rect 3332 11154 3384 11160
rect 3240 11144 3292 11150
rect 3240 11086 3292 11092
rect 2504 11076 2556 11082
rect 2504 11018 2556 11024
rect 2136 10532 2188 10538
rect 2136 10474 2188 10480
rect 1768 10056 1820 10062
rect 1768 9998 1820 10004
rect 1780 9722 1808 9998
rect 2148 9926 2176 10474
rect 2136 9920 2188 9926
rect 2136 9862 2188 9868
rect 1768 9716 1820 9722
rect 1768 9658 1820 9664
rect 2148 9586 2176 9862
rect 2136 9580 2188 9586
rect 2136 9522 2188 9528
rect 2516 7410 2544 11018
rect 3148 11008 3200 11014
rect 3148 10950 3200 10956
rect 3160 10674 3188 10950
rect 2688 10668 2740 10674
rect 2688 10610 2740 10616
rect 3148 10668 3200 10674
rect 3148 10610 3200 10616
rect 2700 10266 2728 10610
rect 2964 10600 3016 10606
rect 2964 10542 3016 10548
rect 2872 10464 2924 10470
rect 2872 10406 2924 10412
rect 2688 10260 2740 10266
rect 2688 10202 2740 10208
rect 2884 10130 2912 10406
rect 2872 10124 2924 10130
rect 2872 10066 2924 10072
rect 2976 9926 3004 10542
rect 3056 10260 3108 10266
rect 3056 10202 3108 10208
rect 3068 9926 3096 10202
rect 2964 9920 3016 9926
rect 2964 9862 3016 9868
rect 3056 9920 3108 9926
rect 3056 9862 3108 9868
rect 2872 9376 2924 9382
rect 2872 9318 2924 9324
rect 2884 8906 2912 9318
rect 2976 9178 3004 9862
rect 3160 9518 3188 10610
rect 3252 10130 3280 11086
rect 3344 10130 3372 11154
rect 3436 10606 3464 12174
rect 3988 11082 4016 12786
rect 4356 12306 4384 12922
rect 4540 12850 4568 14962
rect 5170 14716 5478 14725
rect 5170 14714 5176 14716
rect 5232 14714 5256 14716
rect 5312 14714 5336 14716
rect 5392 14714 5416 14716
rect 5472 14714 5478 14716
rect 5232 14662 5234 14714
rect 5414 14662 5416 14714
rect 5170 14660 5176 14662
rect 5232 14660 5256 14662
rect 5312 14660 5336 14662
rect 5392 14660 5416 14662
rect 5472 14660 5478 14662
rect 5170 14651 5478 14660
rect 5736 14346 5764 15098
rect 6104 14822 6132 15438
rect 6288 15094 6316 15438
rect 7392 15434 7420 16050
rect 7380 15428 7432 15434
rect 7380 15370 7432 15376
rect 6828 15360 6880 15366
rect 6828 15302 6880 15308
rect 6276 15088 6328 15094
rect 6276 15030 6328 15036
rect 6092 14816 6144 14822
rect 6092 14758 6144 14764
rect 6840 14618 6868 15302
rect 7392 14618 7420 15370
rect 6828 14612 6880 14618
rect 6828 14554 6880 14560
rect 7380 14612 7432 14618
rect 7380 14554 7432 14560
rect 6276 14544 6328 14550
rect 6276 14486 6328 14492
rect 6288 14414 6316 14486
rect 6276 14408 6328 14414
rect 6276 14350 6328 14356
rect 5724 14340 5776 14346
rect 5724 14282 5776 14288
rect 6460 14340 6512 14346
rect 6460 14282 6512 14288
rect 6472 14006 6500 14282
rect 6460 14000 6512 14006
rect 6460 13942 6512 13948
rect 5540 13932 5592 13938
rect 5540 13874 5592 13880
rect 5080 13864 5132 13870
rect 5080 13806 5132 13812
rect 5092 13326 5120 13806
rect 5170 13628 5478 13637
rect 5170 13626 5176 13628
rect 5232 13626 5256 13628
rect 5312 13626 5336 13628
rect 5392 13626 5416 13628
rect 5472 13626 5478 13628
rect 5232 13574 5234 13626
rect 5414 13574 5416 13626
rect 5170 13572 5176 13574
rect 5232 13572 5256 13574
rect 5312 13572 5336 13574
rect 5392 13572 5416 13574
rect 5472 13572 5478 13574
rect 5170 13563 5478 13572
rect 5552 13530 5580 13874
rect 6840 13734 6868 14554
rect 6920 14272 6972 14278
rect 6920 14214 6972 14220
rect 7196 14272 7248 14278
rect 7196 14214 7248 14220
rect 6828 13728 6880 13734
rect 6828 13670 6880 13676
rect 5540 13524 5592 13530
rect 5540 13466 5592 13472
rect 5080 13320 5132 13326
rect 5080 13262 5132 13268
rect 4528 12844 4580 12850
rect 4528 12786 4580 12792
rect 4344 12300 4396 12306
rect 4344 12242 4396 12248
rect 4540 11354 4568 12786
rect 5170 12540 5478 12549
rect 5170 12538 5176 12540
rect 5232 12538 5256 12540
rect 5312 12538 5336 12540
rect 5392 12538 5416 12540
rect 5472 12538 5478 12540
rect 5232 12486 5234 12538
rect 5414 12486 5416 12538
rect 5170 12484 5176 12486
rect 5232 12484 5256 12486
rect 5312 12484 5336 12486
rect 5392 12484 5416 12486
rect 5472 12484 5478 12486
rect 5170 12475 5478 12484
rect 6932 12434 6960 14214
rect 7208 14006 7236 14214
rect 7484 14006 7512 16050
rect 7760 15910 7788 17138
rect 7748 15904 7800 15910
rect 7748 15846 7800 15852
rect 7760 15706 7788 15846
rect 7748 15700 7800 15706
rect 7748 15642 7800 15648
rect 7852 14278 7880 20266
rect 8036 19854 8064 20402
rect 8496 19854 8524 20402
rect 8024 19848 8076 19854
rect 8024 19790 8076 19796
rect 8484 19848 8536 19854
rect 8484 19790 8536 19796
rect 8208 19168 8260 19174
rect 8208 19110 8260 19116
rect 8220 18698 8248 19110
rect 8496 18902 8524 19790
rect 8484 18896 8536 18902
rect 8484 18838 8536 18844
rect 8208 18692 8260 18698
rect 8208 18634 8260 18640
rect 8220 18290 8248 18634
rect 8208 18284 8260 18290
rect 8208 18226 8260 18232
rect 8220 17082 8248 18226
rect 8864 17270 8892 20454
rect 8944 20392 8996 20398
rect 8944 20334 8996 20340
rect 8956 19786 8984 20334
rect 8944 19780 8996 19786
rect 8944 19722 8996 19728
rect 8956 19378 8984 19722
rect 8944 19372 8996 19378
rect 8944 19314 8996 19320
rect 8956 18426 8984 19314
rect 8944 18420 8996 18426
rect 8944 18362 8996 18368
rect 8852 17264 8904 17270
rect 8852 17206 8904 17212
rect 8220 17054 8340 17082
rect 8312 16998 8340 17054
rect 8208 16992 8260 16998
rect 8208 16934 8260 16940
rect 8300 16992 8352 16998
rect 8300 16934 8352 16940
rect 8220 16794 8248 16934
rect 8208 16788 8260 16794
rect 8208 16730 8260 16736
rect 8312 16674 8340 16934
rect 8220 16646 8340 16674
rect 7932 14340 7984 14346
rect 7932 14282 7984 14288
rect 7748 14272 7800 14278
rect 7748 14214 7800 14220
rect 7840 14272 7892 14278
rect 7840 14214 7892 14220
rect 7196 14000 7248 14006
rect 7196 13942 7248 13948
rect 7472 14000 7524 14006
rect 7472 13942 7524 13948
rect 7760 13394 7788 14214
rect 7944 14074 7972 14282
rect 8220 14226 8248 16646
rect 9048 15026 9076 21830
rect 9390 21788 9698 21797
rect 9390 21786 9396 21788
rect 9452 21786 9476 21788
rect 9532 21786 9556 21788
rect 9612 21786 9636 21788
rect 9692 21786 9698 21788
rect 9452 21734 9454 21786
rect 9634 21734 9636 21786
rect 9390 21732 9396 21734
rect 9452 21732 9476 21734
rect 9532 21732 9556 21734
rect 9612 21732 9636 21734
rect 9692 21732 9698 21734
rect 9390 21723 9698 21732
rect 9390 20700 9698 20709
rect 9390 20698 9396 20700
rect 9452 20698 9476 20700
rect 9532 20698 9556 20700
rect 9612 20698 9636 20700
rect 9692 20698 9698 20700
rect 9452 20646 9454 20698
rect 9634 20646 9636 20698
rect 9390 20644 9396 20646
rect 9452 20644 9476 20646
rect 9532 20644 9556 20646
rect 9612 20644 9636 20646
rect 9692 20644 9698 20646
rect 9390 20635 9698 20644
rect 9772 19780 9824 19786
rect 9772 19722 9824 19728
rect 9390 19612 9698 19621
rect 9390 19610 9396 19612
rect 9452 19610 9476 19612
rect 9532 19610 9556 19612
rect 9612 19610 9636 19612
rect 9692 19610 9698 19612
rect 9452 19558 9454 19610
rect 9634 19558 9636 19610
rect 9390 19556 9396 19558
rect 9452 19556 9476 19558
rect 9532 19556 9556 19558
rect 9612 19556 9636 19558
rect 9692 19556 9698 19558
rect 9390 19547 9698 19556
rect 9784 19378 9812 19722
rect 9772 19372 9824 19378
rect 9772 19314 9824 19320
rect 9772 19236 9824 19242
rect 9772 19178 9824 19184
rect 9128 19168 9180 19174
rect 9128 19110 9180 19116
rect 9140 18834 9168 19110
rect 9128 18828 9180 18834
rect 9128 18770 9180 18776
rect 9390 18524 9698 18533
rect 9390 18522 9396 18524
rect 9452 18522 9476 18524
rect 9532 18522 9556 18524
rect 9612 18522 9636 18524
rect 9692 18522 9698 18524
rect 9452 18470 9454 18522
rect 9634 18470 9636 18522
rect 9390 18468 9396 18470
rect 9452 18468 9476 18470
rect 9532 18468 9556 18470
rect 9612 18468 9636 18470
rect 9692 18468 9698 18470
rect 9390 18459 9698 18468
rect 9390 17436 9698 17445
rect 9390 17434 9396 17436
rect 9452 17434 9476 17436
rect 9532 17434 9556 17436
rect 9612 17434 9636 17436
rect 9692 17434 9698 17436
rect 9452 17382 9454 17434
rect 9634 17382 9636 17434
rect 9390 17380 9396 17382
rect 9452 17380 9476 17382
rect 9532 17380 9556 17382
rect 9612 17380 9636 17382
rect 9692 17380 9698 17382
rect 9390 17371 9698 17380
rect 9784 17134 9812 19178
rect 9876 17202 9904 23258
rect 10140 22976 10192 22982
rect 10140 22918 10192 22924
rect 10152 20942 10180 22918
rect 10244 21894 10272 25162
rect 10324 22976 10376 22982
rect 10324 22918 10376 22924
rect 10416 22976 10468 22982
rect 10416 22918 10468 22924
rect 10336 22166 10364 22918
rect 10428 22642 10456 22918
rect 11716 22642 11744 31894
rect 11796 29164 11848 29170
rect 11796 29106 11848 29112
rect 11808 28626 11836 29106
rect 11796 28620 11848 28626
rect 11796 28562 11848 28568
rect 11992 24206 12020 32166
rect 12360 31822 12388 32302
rect 13464 32298 13676 32314
rect 14004 32302 14056 32308
rect 13452 32292 13688 32298
rect 13504 32286 13636 32292
rect 13452 32234 13504 32240
rect 13636 32234 13688 32240
rect 13176 32224 13228 32230
rect 13176 32166 13228 32172
rect 12348 31816 12400 31822
rect 12348 31758 12400 31764
rect 13084 31340 13136 31346
rect 13084 31282 13136 31288
rect 12900 30048 12952 30054
rect 12900 29990 12952 29996
rect 12624 29708 12676 29714
rect 12624 29650 12676 29656
rect 12636 29170 12664 29650
rect 12912 29646 12940 29990
rect 13096 29714 13124 31282
rect 13084 29708 13136 29714
rect 13084 29650 13136 29656
rect 12900 29640 12952 29646
rect 12900 29582 12952 29588
rect 12808 29504 12860 29510
rect 12808 29446 12860 29452
rect 12820 29170 12848 29446
rect 12912 29306 12940 29582
rect 12900 29300 12952 29306
rect 12900 29242 12952 29248
rect 12624 29164 12676 29170
rect 12624 29106 12676 29112
rect 12808 29164 12860 29170
rect 12808 29106 12860 29112
rect 12532 28620 12584 28626
rect 12532 28562 12584 28568
rect 12544 28082 12572 28562
rect 12820 28558 12848 29106
rect 12808 28552 12860 28558
rect 12808 28494 12860 28500
rect 12992 28552 13044 28558
rect 12992 28494 13044 28500
rect 12900 28416 12952 28422
rect 12900 28358 12952 28364
rect 12532 28076 12584 28082
rect 12532 28018 12584 28024
rect 12440 28008 12492 28014
rect 12440 27950 12492 27956
rect 12348 27396 12400 27402
rect 12348 27338 12400 27344
rect 12360 25906 12388 27338
rect 12452 26994 12480 27950
rect 12544 27538 12572 28018
rect 12532 27532 12584 27538
rect 12532 27474 12584 27480
rect 12912 27130 12940 28358
rect 13004 28218 13032 28494
rect 12992 28212 13044 28218
rect 12992 28154 13044 28160
rect 13004 27946 13032 28154
rect 12992 27940 13044 27946
rect 12992 27882 13044 27888
rect 13096 27538 13124 29650
rect 13084 27532 13136 27538
rect 13084 27474 13136 27480
rect 12900 27124 12952 27130
rect 12900 27066 12952 27072
rect 12440 26988 12492 26994
rect 12440 26930 12492 26936
rect 12452 26738 12480 26930
rect 12624 26920 12676 26926
rect 12624 26862 12676 26868
rect 12452 26710 12572 26738
rect 12440 26580 12492 26586
rect 12440 26522 12492 26528
rect 12452 25974 12480 26522
rect 12544 26314 12572 26710
rect 12636 26382 12664 26862
rect 12912 26586 12940 27066
rect 13096 27062 13124 27474
rect 13084 27056 13136 27062
rect 13084 26998 13136 27004
rect 12900 26580 12952 26586
rect 12900 26522 12952 26528
rect 12808 26444 12860 26450
rect 12808 26386 12860 26392
rect 12624 26376 12676 26382
rect 12624 26318 12676 26324
rect 12532 26308 12584 26314
rect 12532 26250 12584 26256
rect 12544 26042 12572 26250
rect 12532 26036 12584 26042
rect 12532 25978 12584 25984
rect 12440 25968 12492 25974
rect 12440 25910 12492 25916
rect 12256 25900 12308 25906
rect 12256 25842 12308 25848
rect 12348 25900 12400 25906
rect 12348 25842 12400 25848
rect 12268 25294 12296 25842
rect 12716 25696 12768 25702
rect 12716 25638 12768 25644
rect 12728 25294 12756 25638
rect 12256 25288 12308 25294
rect 12256 25230 12308 25236
rect 12716 25288 12768 25294
rect 12716 25230 12768 25236
rect 12820 24818 12848 26386
rect 13096 26382 13124 26998
rect 13084 26376 13136 26382
rect 13084 26318 13136 26324
rect 13084 25696 13136 25702
rect 13084 25638 13136 25644
rect 13096 25362 13124 25638
rect 13084 25356 13136 25362
rect 13084 25298 13136 25304
rect 12808 24812 12860 24818
rect 12808 24754 12860 24760
rect 11980 24200 12032 24206
rect 11980 24142 12032 24148
rect 13084 24200 13136 24206
rect 13084 24142 13136 24148
rect 11992 23066 12020 24142
rect 12256 24132 12308 24138
rect 12256 24074 12308 24080
rect 12268 23662 12296 24074
rect 12624 24064 12676 24070
rect 12624 24006 12676 24012
rect 12900 24064 12952 24070
rect 12900 24006 12952 24012
rect 12256 23656 12308 23662
rect 12256 23598 12308 23604
rect 11900 23050 12020 23066
rect 12072 23112 12124 23118
rect 12072 23054 12124 23060
rect 11888 23044 12020 23050
rect 11940 23038 12020 23044
rect 11888 22986 11940 22992
rect 10416 22636 10468 22642
rect 10416 22578 10468 22584
rect 11704 22636 11756 22642
rect 11704 22578 11756 22584
rect 11716 22234 11744 22578
rect 11796 22568 11848 22574
rect 11796 22510 11848 22516
rect 11704 22228 11756 22234
rect 11704 22170 11756 22176
rect 10324 22160 10376 22166
rect 10324 22102 10376 22108
rect 10232 21888 10284 21894
rect 10232 21830 10284 21836
rect 10140 20936 10192 20942
rect 10140 20878 10192 20884
rect 10232 20800 10284 20806
rect 10232 20742 10284 20748
rect 10244 20466 10272 20742
rect 10232 20460 10284 20466
rect 10232 20402 10284 20408
rect 9956 19848 10008 19854
rect 9956 19790 10008 19796
rect 9864 17196 9916 17202
rect 9864 17138 9916 17144
rect 9772 17128 9824 17134
rect 9772 17070 9824 17076
rect 9390 16348 9698 16357
rect 9390 16346 9396 16348
rect 9452 16346 9476 16348
rect 9532 16346 9556 16348
rect 9612 16346 9636 16348
rect 9692 16346 9698 16348
rect 9452 16294 9454 16346
rect 9634 16294 9636 16346
rect 9390 16292 9396 16294
rect 9452 16292 9476 16294
rect 9532 16292 9556 16294
rect 9612 16292 9636 16294
rect 9692 16292 9698 16294
rect 9390 16283 9698 16292
rect 9784 15502 9812 17070
rect 9772 15496 9824 15502
rect 9772 15438 9824 15444
rect 9390 15260 9698 15269
rect 9390 15258 9396 15260
rect 9452 15258 9476 15260
rect 9532 15258 9556 15260
rect 9612 15258 9636 15260
rect 9692 15258 9698 15260
rect 9452 15206 9454 15258
rect 9634 15206 9636 15258
rect 9390 15204 9396 15206
rect 9452 15204 9476 15206
rect 9532 15204 9556 15206
rect 9612 15204 9636 15206
rect 9692 15204 9698 15206
rect 9390 15195 9698 15204
rect 9036 15020 9088 15026
rect 9036 14962 9088 14968
rect 8944 14952 8996 14958
rect 8944 14894 8996 14900
rect 8668 14544 8720 14550
rect 8668 14486 8720 14492
rect 8300 14340 8352 14346
rect 8300 14282 8352 14288
rect 8312 14226 8340 14282
rect 8220 14198 8340 14226
rect 7932 14068 7984 14074
rect 7932 14010 7984 14016
rect 7748 13388 7800 13394
rect 7748 13330 7800 13336
rect 7380 13184 7432 13190
rect 7380 13126 7432 13132
rect 6932 12406 7052 12434
rect 5170 11452 5478 11461
rect 5170 11450 5176 11452
rect 5232 11450 5256 11452
rect 5312 11450 5336 11452
rect 5392 11450 5416 11452
rect 5472 11450 5478 11452
rect 5232 11398 5234 11450
rect 5414 11398 5416 11450
rect 5170 11396 5176 11398
rect 5232 11396 5256 11398
rect 5312 11396 5336 11398
rect 5392 11396 5416 11398
rect 5472 11396 5478 11398
rect 5170 11387 5478 11396
rect 4528 11348 4580 11354
rect 4528 11290 4580 11296
rect 6092 11144 6144 11150
rect 6092 11086 6144 11092
rect 3976 11076 4028 11082
rect 3976 11018 4028 11024
rect 5632 11076 5684 11082
rect 5632 11018 5684 11024
rect 4344 11008 4396 11014
rect 4344 10950 4396 10956
rect 4356 10810 4384 10950
rect 4344 10804 4396 10810
rect 4344 10746 4396 10752
rect 4252 10668 4304 10674
rect 4252 10610 4304 10616
rect 3424 10600 3476 10606
rect 3424 10542 3476 10548
rect 3240 10124 3292 10130
rect 3240 10066 3292 10072
rect 3332 10124 3384 10130
rect 3332 10066 3384 10072
rect 3148 9512 3200 9518
rect 3148 9454 3200 9460
rect 2964 9172 3016 9178
rect 2964 9114 3016 9120
rect 3436 8906 3464 10542
rect 4068 10464 4120 10470
rect 4068 10406 4120 10412
rect 4080 9586 4108 10406
rect 4160 10260 4212 10266
rect 4160 10202 4212 10208
rect 4172 9722 4200 10202
rect 4264 9926 4292 10610
rect 4356 10062 4384 10746
rect 5540 10464 5592 10470
rect 5540 10406 5592 10412
rect 5170 10364 5478 10373
rect 5170 10362 5176 10364
rect 5232 10362 5256 10364
rect 5312 10362 5336 10364
rect 5392 10362 5416 10364
rect 5472 10362 5478 10364
rect 5232 10310 5234 10362
rect 5414 10310 5416 10362
rect 5170 10308 5176 10310
rect 5232 10308 5256 10310
rect 5312 10308 5336 10310
rect 5392 10308 5416 10310
rect 5472 10308 5478 10310
rect 5170 10299 5478 10308
rect 5552 10266 5580 10406
rect 5540 10260 5592 10266
rect 5540 10202 5592 10208
rect 4344 10056 4396 10062
rect 4344 9998 4396 10004
rect 4252 9920 4304 9926
rect 4252 9862 4304 9868
rect 4264 9722 4292 9862
rect 4160 9716 4212 9722
rect 4160 9658 4212 9664
rect 4252 9716 4304 9722
rect 4252 9658 4304 9664
rect 4068 9580 4120 9586
rect 4068 9522 4120 9528
rect 4356 8974 4384 9998
rect 5552 9586 5580 10202
rect 5644 9994 5672 11018
rect 6104 10062 6132 11086
rect 6920 11008 6972 11014
rect 6920 10950 6972 10956
rect 6644 10804 6696 10810
rect 6644 10746 6696 10752
rect 6656 10606 6684 10746
rect 6932 10742 6960 10950
rect 6736 10736 6788 10742
rect 6736 10678 6788 10684
rect 6920 10736 6972 10742
rect 6920 10678 6972 10684
rect 6644 10600 6696 10606
rect 6644 10542 6696 10548
rect 6092 10056 6144 10062
rect 6092 9998 6144 10004
rect 5632 9988 5684 9994
rect 5632 9930 5684 9936
rect 4712 9580 4764 9586
rect 4712 9522 4764 9528
rect 5540 9580 5592 9586
rect 5540 9522 5592 9528
rect 4724 9042 4752 9522
rect 5170 9276 5478 9285
rect 5170 9274 5176 9276
rect 5232 9274 5256 9276
rect 5312 9274 5336 9276
rect 5392 9274 5416 9276
rect 5472 9274 5478 9276
rect 5232 9222 5234 9274
rect 5414 9222 5416 9274
rect 5170 9220 5176 9222
rect 5232 9220 5256 9222
rect 5312 9220 5336 9222
rect 5392 9220 5416 9222
rect 5472 9220 5478 9222
rect 5170 9211 5478 9220
rect 4712 9036 4764 9042
rect 4712 8978 4764 8984
rect 4344 8968 4396 8974
rect 4344 8910 4396 8916
rect 2872 8900 2924 8906
rect 2872 8842 2924 8848
rect 3056 8900 3108 8906
rect 3056 8842 3108 8848
rect 3424 8900 3476 8906
rect 3424 8842 3476 8848
rect 3068 8786 3096 8842
rect 2976 8758 3096 8786
rect 4344 8832 4396 8838
rect 4344 8774 4396 8780
rect 2504 7404 2556 7410
rect 2504 7346 2556 7352
rect 2516 7002 2544 7346
rect 2596 7200 2648 7206
rect 2596 7142 2648 7148
rect 2608 7002 2636 7142
rect 2504 6996 2556 7002
rect 2504 6938 2556 6944
rect 2596 6996 2648 7002
rect 2596 6938 2648 6944
rect 2516 6458 2544 6938
rect 2688 6724 2740 6730
rect 2688 6666 2740 6672
rect 2504 6452 2556 6458
rect 2504 6394 2556 6400
rect 2700 6390 2728 6666
rect 2688 6384 2740 6390
rect 2688 6326 2740 6332
rect 2976 6322 3004 8758
rect 4068 7880 4120 7886
rect 4068 7822 4120 7828
rect 4080 6798 4108 7822
rect 4356 6866 4384 8774
rect 5170 8188 5478 8197
rect 5170 8186 5176 8188
rect 5232 8186 5256 8188
rect 5312 8186 5336 8188
rect 5392 8186 5416 8188
rect 5472 8186 5478 8188
rect 5232 8134 5234 8186
rect 5414 8134 5416 8186
rect 5170 8132 5176 8134
rect 5232 8132 5256 8134
rect 5312 8132 5336 8134
rect 5392 8132 5416 8134
rect 5472 8132 5478 8134
rect 5170 8123 5478 8132
rect 5644 7478 5672 9930
rect 5632 7472 5684 7478
rect 5632 7414 5684 7420
rect 5170 7100 5478 7109
rect 5170 7098 5176 7100
rect 5232 7098 5256 7100
rect 5312 7098 5336 7100
rect 5392 7098 5416 7100
rect 5472 7098 5478 7100
rect 5232 7046 5234 7098
rect 5414 7046 5416 7098
rect 5170 7044 5176 7046
rect 5232 7044 5256 7046
rect 5312 7044 5336 7046
rect 5392 7044 5416 7046
rect 5472 7044 5478 7046
rect 5170 7035 5478 7044
rect 5644 6882 5672 7414
rect 4344 6860 4396 6866
rect 4344 6802 4396 6808
rect 5080 6860 5132 6866
rect 5644 6854 5764 6882
rect 5080 6802 5132 6808
rect 3424 6792 3476 6798
rect 3424 6734 3476 6740
rect 4068 6792 4120 6798
rect 4068 6734 4120 6740
rect 3436 6322 3464 6734
rect 2964 6316 3016 6322
rect 2964 6258 3016 6264
rect 3424 6316 3476 6322
rect 3424 6258 3476 6264
rect 2976 5166 3004 6258
rect 3976 6112 4028 6118
rect 3976 6054 4028 6060
rect 3988 5778 4016 6054
rect 3976 5772 4028 5778
rect 3976 5714 4028 5720
rect 4080 5234 4108 6734
rect 4712 5636 4764 5642
rect 4712 5578 4764 5584
rect 4724 5302 4752 5578
rect 4712 5296 4764 5302
rect 4712 5238 4764 5244
rect 4068 5228 4120 5234
rect 4068 5170 4120 5176
rect 2964 5160 3016 5166
rect 2964 5102 3016 5108
rect 5092 4690 5120 6802
rect 5736 6798 5764 6854
rect 5724 6792 5776 6798
rect 5724 6734 5776 6740
rect 5724 6248 5776 6254
rect 5724 6190 5776 6196
rect 5170 6012 5478 6021
rect 5170 6010 5176 6012
rect 5232 6010 5256 6012
rect 5312 6010 5336 6012
rect 5392 6010 5416 6012
rect 5472 6010 5478 6012
rect 5232 5958 5234 6010
rect 5414 5958 5416 6010
rect 5170 5956 5176 5958
rect 5232 5956 5256 5958
rect 5312 5956 5336 5958
rect 5392 5956 5416 5958
rect 5472 5956 5478 5958
rect 5170 5947 5478 5956
rect 5736 5778 5764 6190
rect 5540 5772 5592 5778
rect 5540 5714 5592 5720
rect 5724 5772 5776 5778
rect 5724 5714 5776 5720
rect 5552 5370 5580 5714
rect 5540 5364 5592 5370
rect 5540 5306 5592 5312
rect 5736 5234 5764 5714
rect 6656 5302 6684 10542
rect 6748 10266 6776 10678
rect 6736 10260 6788 10266
rect 6736 10202 6788 10208
rect 6828 9580 6880 9586
rect 6828 9522 6880 9528
rect 6840 9042 6868 9522
rect 6828 9036 6880 9042
rect 6828 8978 6880 8984
rect 6920 6656 6972 6662
rect 6920 6598 6972 6604
rect 6932 6458 6960 6598
rect 6920 6452 6972 6458
rect 6920 6394 6972 6400
rect 7024 6390 7052 12406
rect 7104 11008 7156 11014
rect 7104 10950 7156 10956
rect 7116 10674 7144 10950
rect 7104 10668 7156 10674
rect 7104 10610 7156 10616
rect 7392 10146 7420 13126
rect 7472 12640 7524 12646
rect 7472 12582 7524 12588
rect 7484 10742 7512 12582
rect 8220 10810 8248 14198
rect 8300 14068 8352 14074
rect 8300 14010 8352 14016
rect 8312 13326 8340 14010
rect 8392 13932 8444 13938
rect 8392 13874 8444 13880
rect 8300 13320 8352 13326
rect 8300 13262 8352 13268
rect 8208 10804 8260 10810
rect 8208 10746 8260 10752
rect 7472 10736 7524 10742
rect 7472 10678 7524 10684
rect 7932 10464 7984 10470
rect 7932 10406 7984 10412
rect 7944 10146 7972 10406
rect 7392 10118 7512 10146
rect 7484 10062 7512 10118
rect 7852 10118 7972 10146
rect 7472 10056 7524 10062
rect 7472 9998 7524 10004
rect 7484 9654 7512 9998
rect 7852 9926 7880 10118
rect 7840 9920 7892 9926
rect 7840 9862 7892 9868
rect 7472 9648 7524 9654
rect 7472 9590 7524 9596
rect 7380 7812 7432 7818
rect 7380 7754 7432 7760
rect 7392 7478 7420 7754
rect 7380 7472 7432 7478
rect 7380 7414 7432 7420
rect 7012 6384 7064 6390
rect 7012 6326 7064 6332
rect 6644 5296 6696 5302
rect 6644 5238 6696 5244
rect 5724 5228 5776 5234
rect 5724 5170 5776 5176
rect 7196 5092 7248 5098
rect 7196 5034 7248 5040
rect 5170 4924 5478 4933
rect 5170 4922 5176 4924
rect 5232 4922 5256 4924
rect 5312 4922 5336 4924
rect 5392 4922 5416 4924
rect 5472 4922 5478 4924
rect 5232 4870 5234 4922
rect 5414 4870 5416 4922
rect 5170 4868 5176 4870
rect 5232 4868 5256 4870
rect 5312 4868 5336 4870
rect 5392 4868 5416 4870
rect 5472 4868 5478 4870
rect 5170 4859 5478 4868
rect 7208 4690 7236 5034
rect 5080 4684 5132 4690
rect 5080 4626 5132 4632
rect 7196 4684 7248 4690
rect 7196 4626 7248 4632
rect 7484 4622 7512 9590
rect 7472 4616 7524 4622
rect 7472 4558 7524 4564
rect 7484 4282 7512 4558
rect 7472 4276 7524 4282
rect 7472 4218 7524 4224
rect 5170 3836 5478 3845
rect 5170 3834 5176 3836
rect 5232 3834 5256 3836
rect 5312 3834 5336 3836
rect 5392 3834 5416 3836
rect 5472 3834 5478 3836
rect 5232 3782 5234 3834
rect 5414 3782 5416 3834
rect 5170 3780 5176 3782
rect 5232 3780 5256 3782
rect 5312 3780 5336 3782
rect 5392 3780 5416 3782
rect 5472 3780 5478 3782
rect 5170 3771 5478 3780
rect 5170 2748 5478 2757
rect 5170 2746 5176 2748
rect 5232 2746 5256 2748
rect 5312 2746 5336 2748
rect 5392 2746 5416 2748
rect 5472 2746 5478 2748
rect 5232 2694 5234 2746
rect 5414 2694 5416 2746
rect 5170 2692 5176 2694
rect 5232 2692 5256 2694
rect 5312 2692 5336 2694
rect 5392 2692 5416 2694
rect 5472 2692 5478 2694
rect 5170 2683 5478 2692
rect 6368 2440 6420 2446
rect 6368 2382 6420 2388
rect 7656 2440 7708 2446
rect 7656 2382 7708 2388
rect 1216 2372 1268 2378
rect 1216 2314 1268 2320
rect 2504 2372 2556 2378
rect 2504 2314 2556 2320
rect 3792 2372 3844 2378
rect 3792 2314 3844 2320
rect 5080 2372 5132 2378
rect 5080 2314 5132 2320
rect 1228 800 1256 2314
rect 2516 800 2544 2314
rect 3804 800 3832 2314
rect 5092 800 5120 2314
rect 6380 800 6408 2382
rect 7668 800 7696 2382
rect 7852 2378 7880 9862
rect 8208 7812 8260 7818
rect 8208 7754 8260 7760
rect 8220 5166 8248 7754
rect 8404 7410 8432 13874
rect 8680 13258 8708 14486
rect 8484 13252 8536 13258
rect 8484 13194 8536 13200
rect 8668 13252 8720 13258
rect 8668 13194 8720 13200
rect 8496 12918 8524 13194
rect 8484 12912 8536 12918
rect 8484 12854 8536 12860
rect 8956 11014 8984 14894
rect 9220 14544 9272 14550
rect 9220 14486 9272 14492
rect 9128 13388 9180 13394
rect 9128 13330 9180 13336
rect 9036 13184 9088 13190
rect 9036 13126 9088 13132
rect 9048 12434 9076 13126
rect 9140 12782 9168 13330
rect 9232 12918 9260 14486
rect 9588 14408 9640 14414
rect 9784 14396 9812 15438
rect 9876 14958 9904 17138
rect 9968 16590 9996 19790
rect 10244 19786 10272 20402
rect 10232 19780 10284 19786
rect 10232 19722 10284 19728
rect 10336 19378 10364 22102
rect 10784 22092 10836 22098
rect 10784 22034 10836 22040
rect 10796 20942 10824 22034
rect 11704 21956 11756 21962
rect 11704 21898 11756 21904
rect 11060 21888 11112 21894
rect 11060 21830 11112 21836
rect 10416 20936 10468 20942
rect 10416 20878 10468 20884
rect 10784 20936 10836 20942
rect 10784 20878 10836 20884
rect 10428 20398 10456 20878
rect 10416 20392 10468 20398
rect 10416 20334 10468 20340
rect 10428 19854 10456 20334
rect 10416 19848 10468 19854
rect 10796 19836 10824 20878
rect 11072 20466 11100 21830
rect 11716 21622 11744 21898
rect 11704 21616 11756 21622
rect 11704 21558 11756 21564
rect 11808 21554 11836 22510
rect 11980 22500 12032 22506
rect 11980 22442 12032 22448
rect 11992 21554 12020 22442
rect 12084 22030 12112 23054
rect 12072 22024 12124 22030
rect 12072 21966 12124 21972
rect 11796 21548 11848 21554
rect 11796 21490 11848 21496
rect 11980 21548 12032 21554
rect 11980 21490 12032 21496
rect 11060 20460 11112 20466
rect 11060 20402 11112 20408
rect 10876 19848 10928 19854
rect 10796 19808 10876 19836
rect 10416 19790 10468 19796
rect 10876 19790 10928 19796
rect 11520 19712 11572 19718
rect 11520 19654 11572 19660
rect 10324 19372 10376 19378
rect 10324 19314 10376 19320
rect 11532 19310 11560 19654
rect 11060 19304 11112 19310
rect 11060 19246 11112 19252
rect 11520 19304 11572 19310
rect 11520 19246 11572 19252
rect 10232 19168 10284 19174
rect 10232 19110 10284 19116
rect 10692 19168 10744 19174
rect 10692 19110 10744 19116
rect 10244 18766 10272 19110
rect 10704 18766 10732 19110
rect 10232 18760 10284 18766
rect 10232 18702 10284 18708
rect 10692 18760 10744 18766
rect 10692 18702 10744 18708
rect 11072 18290 11100 19246
rect 11808 18290 11836 21490
rect 11888 20868 11940 20874
rect 11888 20810 11940 20816
rect 11900 19922 11928 20810
rect 11888 19916 11940 19922
rect 11888 19858 11940 19864
rect 11992 18358 12020 21490
rect 11980 18352 12032 18358
rect 11980 18294 12032 18300
rect 11060 18284 11112 18290
rect 11060 18226 11112 18232
rect 11796 18284 11848 18290
rect 11796 18226 11848 18232
rect 10232 18080 10284 18086
rect 10232 18022 10284 18028
rect 10048 16992 10100 16998
rect 10048 16934 10100 16940
rect 10060 16590 10088 16934
rect 9956 16584 10008 16590
rect 9956 16526 10008 16532
rect 10048 16584 10100 16590
rect 10048 16526 10100 16532
rect 9956 15020 10008 15026
rect 9956 14962 10008 14968
rect 9864 14952 9916 14958
rect 9864 14894 9916 14900
rect 9968 14822 9996 14962
rect 9956 14816 10008 14822
rect 9956 14758 10008 14764
rect 9640 14368 9812 14396
rect 9588 14350 9640 14356
rect 9390 14172 9698 14181
rect 9390 14170 9396 14172
rect 9452 14170 9476 14172
rect 9532 14170 9556 14172
rect 9612 14170 9636 14172
rect 9692 14170 9698 14172
rect 9452 14118 9454 14170
rect 9634 14118 9636 14170
rect 9390 14116 9396 14118
rect 9452 14116 9476 14118
rect 9532 14116 9556 14118
rect 9612 14116 9636 14118
rect 9692 14116 9698 14118
rect 9390 14107 9698 14116
rect 9312 14000 9364 14006
rect 9312 13942 9364 13948
rect 9220 12912 9272 12918
rect 9220 12854 9272 12860
rect 9128 12776 9180 12782
rect 9128 12718 9180 12724
rect 9048 12406 9168 12434
rect 8852 11008 8904 11014
rect 8852 10950 8904 10956
rect 8944 11008 8996 11014
rect 8944 10950 8996 10956
rect 8864 10826 8892 10950
rect 8864 10810 8984 10826
rect 8484 10804 8536 10810
rect 8864 10804 8996 10810
rect 8864 10798 8944 10804
rect 8484 10746 8536 10752
rect 8944 10746 8996 10752
rect 8496 9722 8524 10746
rect 9140 10724 9168 12406
rect 9232 11082 9260 12854
rect 9220 11076 9272 11082
rect 9220 11018 9272 11024
rect 9220 10736 9272 10742
rect 9140 10696 9220 10724
rect 9220 10678 9272 10684
rect 9036 10668 9088 10674
rect 9036 10610 9088 10616
rect 8668 10532 8720 10538
rect 8668 10474 8720 10480
rect 8680 10198 8708 10474
rect 9048 10266 9076 10610
rect 9036 10260 9088 10266
rect 9036 10202 9088 10208
rect 8668 10192 8720 10198
rect 8668 10134 8720 10140
rect 8484 9716 8536 9722
rect 8484 9658 8536 9664
rect 9324 8566 9352 13942
rect 9390 13084 9698 13093
rect 9390 13082 9396 13084
rect 9452 13082 9476 13084
rect 9532 13082 9556 13084
rect 9612 13082 9636 13084
rect 9692 13082 9698 13084
rect 9452 13030 9454 13082
rect 9634 13030 9636 13082
rect 9390 13028 9396 13030
rect 9452 13028 9476 13030
rect 9532 13028 9556 13030
rect 9612 13028 9636 13030
rect 9692 13028 9698 13030
rect 9390 13019 9698 13028
rect 9390 11996 9698 12005
rect 9390 11994 9396 11996
rect 9452 11994 9476 11996
rect 9532 11994 9556 11996
rect 9612 11994 9636 11996
rect 9692 11994 9698 11996
rect 9452 11942 9454 11994
rect 9634 11942 9636 11994
rect 9390 11940 9396 11942
rect 9452 11940 9476 11942
rect 9532 11940 9556 11942
rect 9612 11940 9636 11942
rect 9692 11940 9698 11942
rect 9390 11931 9698 11940
rect 9390 10908 9698 10917
rect 9390 10906 9396 10908
rect 9452 10906 9476 10908
rect 9532 10906 9556 10908
rect 9612 10906 9636 10908
rect 9692 10906 9698 10908
rect 9452 10854 9454 10906
rect 9634 10854 9636 10906
rect 9390 10852 9396 10854
rect 9452 10852 9476 10854
rect 9532 10852 9556 10854
rect 9612 10852 9636 10854
rect 9692 10852 9698 10854
rect 9390 10843 9698 10852
rect 9784 10810 9812 14368
rect 9968 14346 9996 14758
rect 10244 14414 10272 18022
rect 11336 17740 11388 17746
rect 11336 17682 11388 17688
rect 10968 17536 11020 17542
rect 10968 17478 11020 17484
rect 10324 17332 10376 17338
rect 10324 17274 10376 17280
rect 10336 14958 10364 17274
rect 10980 16726 11008 17478
rect 11152 16992 11204 16998
rect 11152 16934 11204 16940
rect 10968 16720 11020 16726
rect 10968 16662 11020 16668
rect 10416 16448 10468 16454
rect 10416 16390 10468 16396
rect 10428 16114 10456 16390
rect 10980 16114 11008 16662
rect 11164 16522 11192 16934
rect 11152 16516 11204 16522
rect 11152 16458 11204 16464
rect 11164 16114 11192 16458
rect 11348 16182 11376 17682
rect 11992 16658 12020 18294
rect 12084 17746 12112 21966
rect 12164 18216 12216 18222
rect 12164 18158 12216 18164
rect 12072 17740 12124 17746
rect 12072 17682 12124 17688
rect 12176 17610 12204 18158
rect 12164 17604 12216 17610
rect 12164 17546 12216 17552
rect 12268 17490 12296 23598
rect 12440 23044 12492 23050
rect 12440 22986 12492 22992
rect 12452 22778 12480 22986
rect 12440 22772 12492 22778
rect 12440 22714 12492 22720
rect 12636 22642 12664 24006
rect 12912 23730 12940 24006
rect 13096 23730 13124 24142
rect 12900 23724 12952 23730
rect 12900 23666 12952 23672
rect 13084 23724 13136 23730
rect 13084 23666 13136 23672
rect 12808 22976 12860 22982
rect 12808 22918 12860 22924
rect 12624 22636 12676 22642
rect 12624 22578 12676 22584
rect 12716 22568 12768 22574
rect 12716 22510 12768 22516
rect 12728 22166 12756 22510
rect 12716 22160 12768 22166
rect 12716 22102 12768 22108
rect 12728 19854 12756 22102
rect 12716 19848 12768 19854
rect 12716 19790 12768 19796
rect 12440 19780 12492 19786
rect 12440 19722 12492 19728
rect 12452 19378 12480 19722
rect 12440 19372 12492 19378
rect 12440 19314 12492 19320
rect 12452 18766 12480 19314
rect 12440 18760 12492 18766
rect 12440 18702 12492 18708
rect 12348 18284 12400 18290
rect 12348 18226 12400 18232
rect 12176 17462 12296 17490
rect 11980 16652 12032 16658
rect 11980 16594 12032 16600
rect 11336 16176 11388 16182
rect 11336 16118 11388 16124
rect 10416 16108 10468 16114
rect 10416 16050 10468 16056
rect 10968 16108 11020 16114
rect 10968 16050 11020 16056
rect 11152 16108 11204 16114
rect 11152 16050 11204 16056
rect 11796 15088 11848 15094
rect 11796 15030 11848 15036
rect 10692 15020 10744 15026
rect 10692 14962 10744 14968
rect 10324 14952 10376 14958
rect 10324 14894 10376 14900
rect 10704 14822 10732 14962
rect 10692 14816 10744 14822
rect 10692 14758 10744 14764
rect 10232 14408 10284 14414
rect 10232 14350 10284 14356
rect 9956 14340 10008 14346
rect 9956 14282 10008 14288
rect 11704 14340 11756 14346
rect 11704 14282 11756 14288
rect 9864 14272 9916 14278
rect 9864 14214 9916 14220
rect 9876 14006 9904 14214
rect 9864 14000 9916 14006
rect 9864 13942 9916 13948
rect 9968 12434 9996 14282
rect 11060 14068 11112 14074
rect 11060 14010 11112 14016
rect 10140 13728 10192 13734
rect 10140 13670 10192 13676
rect 10152 13258 10180 13670
rect 10140 13252 10192 13258
rect 10140 13194 10192 13200
rect 9968 12406 10364 12434
rect 9956 11008 10008 11014
rect 9956 10950 10008 10956
rect 9968 10810 9996 10950
rect 9772 10804 9824 10810
rect 9772 10746 9824 10752
rect 9956 10804 10008 10810
rect 9956 10746 10008 10752
rect 10048 10464 10100 10470
rect 10048 10406 10100 10412
rect 9390 9820 9698 9829
rect 9390 9818 9396 9820
rect 9452 9818 9476 9820
rect 9532 9818 9556 9820
rect 9612 9818 9636 9820
rect 9692 9818 9698 9820
rect 9452 9766 9454 9818
rect 9634 9766 9636 9818
rect 9390 9764 9396 9766
rect 9452 9764 9476 9766
rect 9532 9764 9556 9766
rect 9612 9764 9636 9766
rect 9692 9764 9698 9766
rect 9390 9755 9698 9764
rect 10060 9722 10088 10406
rect 10048 9716 10100 9722
rect 10048 9658 10100 9664
rect 9390 8732 9698 8741
rect 9390 8730 9396 8732
rect 9452 8730 9476 8732
rect 9532 8730 9556 8732
rect 9612 8730 9636 8732
rect 9692 8730 9698 8732
rect 9452 8678 9454 8730
rect 9634 8678 9636 8730
rect 9390 8676 9396 8678
rect 9452 8676 9476 8678
rect 9532 8676 9556 8678
rect 9612 8676 9636 8678
rect 9692 8676 9698 8678
rect 9390 8667 9698 8676
rect 9312 8560 9364 8566
rect 9312 8502 9364 8508
rect 9864 8356 9916 8362
rect 9864 8298 9916 8304
rect 9876 7886 9904 8298
rect 9864 7880 9916 7886
rect 9864 7822 9916 7828
rect 9390 7644 9698 7653
rect 9390 7642 9396 7644
rect 9452 7642 9476 7644
rect 9532 7642 9556 7644
rect 9612 7642 9636 7644
rect 9692 7642 9698 7644
rect 9452 7590 9454 7642
rect 9634 7590 9636 7642
rect 9390 7588 9396 7590
rect 9452 7588 9476 7590
rect 9532 7588 9556 7590
rect 9612 7588 9636 7590
rect 9692 7588 9698 7590
rect 9390 7579 9698 7588
rect 8392 7404 8444 7410
rect 8392 7346 8444 7352
rect 8944 7404 8996 7410
rect 8944 7346 8996 7352
rect 8300 7200 8352 7206
rect 8300 7142 8352 7148
rect 8312 6866 8340 7142
rect 8300 6860 8352 6866
rect 8300 6802 8352 6808
rect 8208 5160 8260 5166
rect 8208 5102 8260 5108
rect 7932 4208 7984 4214
rect 7932 4150 7984 4156
rect 7944 3738 7972 4150
rect 7932 3732 7984 3738
rect 7932 3674 7984 3680
rect 8220 3534 8248 5102
rect 8956 4690 8984 7346
rect 9390 6556 9698 6565
rect 9390 6554 9396 6556
rect 9452 6554 9476 6556
rect 9532 6554 9556 6556
rect 9612 6554 9636 6556
rect 9692 6554 9698 6556
rect 9452 6502 9454 6554
rect 9634 6502 9636 6554
rect 9390 6500 9396 6502
rect 9452 6500 9476 6502
rect 9532 6500 9556 6502
rect 9612 6500 9636 6502
rect 9692 6500 9698 6502
rect 9390 6491 9698 6500
rect 9390 5468 9698 5477
rect 9390 5466 9396 5468
rect 9452 5466 9476 5468
rect 9532 5466 9556 5468
rect 9612 5466 9636 5468
rect 9692 5466 9698 5468
rect 9452 5414 9454 5466
rect 9634 5414 9636 5466
rect 9390 5412 9396 5414
rect 9452 5412 9476 5414
rect 9532 5412 9556 5414
rect 9612 5412 9636 5414
rect 9692 5412 9698 5414
rect 9390 5403 9698 5412
rect 9220 5296 9272 5302
rect 9220 5238 9272 5244
rect 8944 4684 8996 4690
rect 8944 4626 8996 4632
rect 8576 4480 8628 4486
rect 8576 4422 8628 4428
rect 8588 4282 8616 4422
rect 8576 4276 8628 4282
rect 8576 4218 8628 4224
rect 8956 4146 8984 4626
rect 9232 4214 9260 5238
rect 9312 5160 9364 5166
rect 9312 5102 9364 5108
rect 9220 4208 9272 4214
rect 9220 4150 9272 4156
rect 8944 4140 8996 4146
rect 8944 4082 8996 4088
rect 9324 4010 9352 5102
rect 9390 4380 9698 4389
rect 9390 4378 9396 4380
rect 9452 4378 9476 4380
rect 9532 4378 9556 4380
rect 9612 4378 9636 4380
rect 9692 4378 9698 4380
rect 9452 4326 9454 4378
rect 9634 4326 9636 4378
rect 9390 4324 9396 4326
rect 9452 4324 9476 4326
rect 9532 4324 9556 4326
rect 9612 4324 9636 4326
rect 9692 4324 9698 4326
rect 9390 4315 9698 4324
rect 9312 4004 9364 4010
rect 9312 3946 9364 3952
rect 9876 3602 9904 7822
rect 9864 3596 9916 3602
rect 9864 3538 9916 3544
rect 8208 3528 8260 3534
rect 8208 3470 8260 3476
rect 9390 3292 9698 3301
rect 9390 3290 9396 3292
rect 9452 3290 9476 3292
rect 9532 3290 9556 3292
rect 9612 3290 9636 3292
rect 9692 3290 9698 3292
rect 9452 3238 9454 3290
rect 9634 3238 9636 3290
rect 9390 3236 9396 3238
rect 9452 3236 9476 3238
rect 9532 3236 9556 3238
rect 9612 3236 9636 3238
rect 9692 3236 9698 3238
rect 9390 3227 9698 3236
rect 10060 2582 10088 9658
rect 10232 7812 10284 7818
rect 10232 7754 10284 7760
rect 10244 7478 10272 7754
rect 10232 7472 10284 7478
rect 10232 7414 10284 7420
rect 10336 6866 10364 12406
rect 11072 11150 11100 14010
rect 11716 13938 11744 14282
rect 11808 14074 11836 15030
rect 11992 14414 12020 16594
rect 12176 15026 12204 17462
rect 12256 17264 12308 17270
rect 12256 17206 12308 17212
rect 12268 16794 12296 17206
rect 12256 16788 12308 16794
rect 12256 16730 12308 16736
rect 12360 16572 12388 18226
rect 12440 16584 12492 16590
rect 12360 16544 12440 16572
rect 12440 16526 12492 16532
rect 12348 16244 12400 16250
rect 12348 16186 12400 16192
rect 12164 15020 12216 15026
rect 12164 14962 12216 14968
rect 12072 14952 12124 14958
rect 12072 14894 12124 14900
rect 11980 14408 12032 14414
rect 11980 14350 12032 14356
rect 11796 14068 11848 14074
rect 11796 14010 11848 14016
rect 11992 14006 12020 14350
rect 11980 14000 12032 14006
rect 11980 13942 12032 13948
rect 11704 13932 11756 13938
rect 11704 13874 11756 13880
rect 11796 13864 11848 13870
rect 11796 13806 11848 13812
rect 11808 13394 11836 13806
rect 12084 13394 12112 14894
rect 11796 13388 11848 13394
rect 11796 13330 11848 13336
rect 12072 13388 12124 13394
rect 12072 13330 12124 13336
rect 10416 11144 10468 11150
rect 10416 11086 10468 11092
rect 11060 11144 11112 11150
rect 11060 11086 11112 11092
rect 10428 10130 10456 11086
rect 10416 10124 10468 10130
rect 10416 10066 10468 10072
rect 10784 9512 10836 9518
rect 10784 9454 10836 9460
rect 10796 9042 10824 9454
rect 10784 9036 10836 9042
rect 10784 8978 10836 8984
rect 11072 8974 11100 11086
rect 11888 10736 11940 10742
rect 11888 10678 11940 10684
rect 11152 10600 11204 10606
rect 11152 10542 11204 10548
rect 11164 10198 11192 10542
rect 11152 10192 11204 10198
rect 11152 10134 11204 10140
rect 11796 9988 11848 9994
rect 11796 9930 11848 9936
rect 11808 9586 11836 9930
rect 11796 9580 11848 9586
rect 11796 9522 11848 9528
rect 11060 8968 11112 8974
rect 11060 8910 11112 8916
rect 10692 7540 10744 7546
rect 10692 7482 10744 7488
rect 10324 6860 10376 6866
rect 10324 6802 10376 6808
rect 10232 5364 10284 5370
rect 10336 5352 10364 6802
rect 10416 6792 10468 6798
rect 10416 6734 10468 6740
rect 10428 5370 10456 6734
rect 10704 6730 10732 7482
rect 11072 7342 11100 8910
rect 11060 7336 11112 7342
rect 11060 7278 11112 7284
rect 11152 7336 11204 7342
rect 11152 7278 11204 7284
rect 11072 6730 11100 7278
rect 11164 6798 11192 7278
rect 11152 6792 11204 6798
rect 11152 6734 11204 6740
rect 11704 6792 11756 6798
rect 11704 6734 11756 6740
rect 10692 6724 10744 6730
rect 10692 6666 10744 6672
rect 11060 6724 11112 6730
rect 11060 6666 11112 6672
rect 10284 5324 10364 5352
rect 10416 5364 10468 5370
rect 10232 5306 10284 5312
rect 10416 5306 10468 5312
rect 10876 5228 10928 5234
rect 10876 5170 10928 5176
rect 10888 4826 10916 5170
rect 11716 5166 11744 6734
rect 11808 5234 11836 9522
rect 11900 7342 11928 10678
rect 12084 9994 12112 13330
rect 12360 11370 12388 16186
rect 12452 14346 12480 16526
rect 12440 14340 12492 14346
rect 12440 14282 12492 14288
rect 12728 12434 12756 19790
rect 12820 13530 12848 22918
rect 13096 22574 13124 23666
rect 13188 23662 13216 32166
rect 13611 32124 13919 32133
rect 13611 32122 13617 32124
rect 13673 32122 13697 32124
rect 13753 32122 13777 32124
rect 13833 32122 13857 32124
rect 13913 32122 13919 32124
rect 13673 32070 13675 32122
rect 13855 32070 13857 32122
rect 13611 32068 13617 32070
rect 13673 32068 13697 32070
rect 13753 32068 13777 32070
rect 13833 32068 13857 32070
rect 13913 32068 13919 32070
rect 13611 32059 13919 32068
rect 14016 31958 14044 32302
rect 16120 32020 16172 32026
rect 16120 31962 16172 31968
rect 14004 31952 14056 31958
rect 14004 31894 14056 31900
rect 14004 31816 14056 31822
rect 14004 31758 14056 31764
rect 14280 31816 14332 31822
rect 14280 31758 14332 31764
rect 14648 31816 14700 31822
rect 14648 31758 14700 31764
rect 13268 31272 13320 31278
rect 13268 31214 13320 31220
rect 13280 30938 13308 31214
rect 13611 31036 13919 31045
rect 13611 31034 13617 31036
rect 13673 31034 13697 31036
rect 13753 31034 13777 31036
rect 13833 31034 13857 31036
rect 13913 31034 13919 31036
rect 13673 30982 13675 31034
rect 13855 30982 13857 31034
rect 13611 30980 13617 30982
rect 13673 30980 13697 30982
rect 13753 30980 13777 30982
rect 13833 30980 13857 30982
rect 13913 30980 13919 30982
rect 13611 30971 13919 30980
rect 13268 30932 13320 30938
rect 13268 30874 13320 30880
rect 14016 30598 14044 31758
rect 14292 31482 14320 31758
rect 14280 31476 14332 31482
rect 14280 31418 14332 31424
rect 14096 31340 14148 31346
rect 14096 31282 14148 31288
rect 14108 30734 14136 31282
rect 14660 31278 14688 31758
rect 16132 31754 16160 31962
rect 15568 31748 15620 31754
rect 15568 31690 15620 31696
rect 16120 31748 16172 31754
rect 16120 31690 16172 31696
rect 15580 31414 15608 31690
rect 15752 31680 15804 31686
rect 15752 31622 15804 31628
rect 15568 31408 15620 31414
rect 15568 31350 15620 31356
rect 14832 31340 14884 31346
rect 14832 31282 14884 31288
rect 15476 31340 15528 31346
rect 15476 31282 15528 31288
rect 14648 31272 14700 31278
rect 14648 31214 14700 31220
rect 14280 31136 14332 31142
rect 14280 31078 14332 31084
rect 14096 30728 14148 30734
rect 14096 30670 14148 30676
rect 14004 30592 14056 30598
rect 14004 30534 14056 30540
rect 14292 30258 14320 31078
rect 14556 30728 14608 30734
rect 14556 30670 14608 30676
rect 14280 30252 14332 30258
rect 14280 30194 14332 30200
rect 13611 29948 13919 29957
rect 13611 29946 13617 29948
rect 13673 29946 13697 29948
rect 13753 29946 13777 29948
rect 13833 29946 13857 29948
rect 13913 29946 13919 29948
rect 13673 29894 13675 29946
rect 13855 29894 13857 29946
rect 13611 29892 13617 29894
rect 13673 29892 13697 29894
rect 13753 29892 13777 29894
rect 13833 29892 13857 29894
rect 13913 29892 13919 29894
rect 13611 29883 13919 29892
rect 14280 29572 14332 29578
rect 14280 29514 14332 29520
rect 13360 29164 13412 29170
rect 13360 29106 13412 29112
rect 13372 28762 13400 29106
rect 13611 28860 13919 28869
rect 13611 28858 13617 28860
rect 13673 28858 13697 28860
rect 13753 28858 13777 28860
rect 13833 28858 13857 28860
rect 13913 28858 13919 28860
rect 13673 28806 13675 28858
rect 13855 28806 13857 28858
rect 13611 28804 13617 28806
rect 13673 28804 13697 28806
rect 13753 28804 13777 28806
rect 13833 28804 13857 28806
rect 13913 28804 13919 28806
rect 13611 28795 13919 28804
rect 13360 28756 13412 28762
rect 13360 28698 13412 28704
rect 13372 28626 13400 28698
rect 13360 28620 13412 28626
rect 13360 28562 13412 28568
rect 13268 28552 13320 28558
rect 13268 28494 13320 28500
rect 13280 28082 13308 28494
rect 13372 28490 13400 28562
rect 13360 28484 13412 28490
rect 13360 28426 13412 28432
rect 13372 28218 13400 28426
rect 13360 28212 13412 28218
rect 13360 28154 13412 28160
rect 14292 28082 14320 29514
rect 14568 29306 14596 30670
rect 14556 29300 14608 29306
rect 14556 29242 14608 29248
rect 14660 29186 14688 31214
rect 14844 30870 14872 31282
rect 14832 30864 14884 30870
rect 14832 30806 14884 30812
rect 14844 29850 14872 30806
rect 15488 30734 15516 31282
rect 15764 31278 15792 31622
rect 16132 31482 16160 31690
rect 16120 31476 16172 31482
rect 16120 31418 16172 31424
rect 15752 31272 15804 31278
rect 15752 31214 15804 31220
rect 15764 30802 15792 31214
rect 15752 30796 15804 30802
rect 15752 30738 15804 30744
rect 14924 30728 14976 30734
rect 14924 30670 14976 30676
rect 15476 30728 15528 30734
rect 15476 30670 15528 30676
rect 14936 30258 14964 30670
rect 14924 30252 14976 30258
rect 14924 30194 14976 30200
rect 14832 29844 14884 29850
rect 14832 29786 14884 29792
rect 14936 29306 14964 30194
rect 15016 29640 15068 29646
rect 15016 29582 15068 29588
rect 14924 29300 14976 29306
rect 14924 29242 14976 29248
rect 14568 29158 14688 29186
rect 14568 28558 14596 29158
rect 15028 29102 15056 29582
rect 15108 29572 15160 29578
rect 15108 29514 15160 29520
rect 15120 29238 15148 29514
rect 15108 29232 15160 29238
rect 15108 29174 15160 29180
rect 15016 29096 15068 29102
rect 15016 29038 15068 29044
rect 15028 28626 15056 29038
rect 15016 28620 15068 28626
rect 15016 28562 15068 28568
rect 14556 28552 14608 28558
rect 14556 28494 14608 28500
rect 13268 28076 13320 28082
rect 13268 28018 13320 28024
rect 14004 28076 14056 28082
rect 14004 28018 14056 28024
rect 14280 28076 14332 28082
rect 14280 28018 14332 28024
rect 13611 27772 13919 27781
rect 13611 27770 13617 27772
rect 13673 27770 13697 27772
rect 13753 27770 13777 27772
rect 13833 27770 13857 27772
rect 13913 27770 13919 27772
rect 13673 27718 13675 27770
rect 13855 27718 13857 27770
rect 13611 27716 13617 27718
rect 13673 27716 13697 27718
rect 13753 27716 13777 27718
rect 13833 27716 13857 27718
rect 13913 27716 13919 27718
rect 13611 27707 13919 27716
rect 13820 27464 13872 27470
rect 13820 27406 13872 27412
rect 13832 27062 13860 27406
rect 14016 27402 14044 28018
rect 14004 27396 14056 27402
rect 14004 27338 14056 27344
rect 14292 27062 14320 28018
rect 14568 28014 14596 28494
rect 15028 28150 15056 28562
rect 15120 28558 15148 29174
rect 15568 29164 15620 29170
rect 15568 29106 15620 29112
rect 15752 29164 15804 29170
rect 15752 29106 15804 29112
rect 15108 28552 15160 28558
rect 15108 28494 15160 28500
rect 15384 28552 15436 28558
rect 15384 28494 15436 28500
rect 15476 28552 15528 28558
rect 15476 28494 15528 28500
rect 15396 28218 15424 28494
rect 15384 28212 15436 28218
rect 15384 28154 15436 28160
rect 15016 28144 15068 28150
rect 15016 28086 15068 28092
rect 15488 28082 15516 28494
rect 15580 28150 15608 29106
rect 15764 28490 15792 29106
rect 15936 28620 15988 28626
rect 15936 28562 15988 28568
rect 15752 28484 15804 28490
rect 15752 28426 15804 28432
rect 15568 28144 15620 28150
rect 15568 28086 15620 28092
rect 15476 28076 15528 28082
rect 15476 28018 15528 28024
rect 14556 28008 14608 28014
rect 14556 27950 14608 27956
rect 13820 27056 13872 27062
rect 13820 26998 13872 27004
rect 14280 27056 14332 27062
rect 14280 26998 14332 27004
rect 13611 26684 13919 26693
rect 13611 26682 13617 26684
rect 13673 26682 13697 26684
rect 13753 26682 13777 26684
rect 13833 26682 13857 26684
rect 13913 26682 13919 26684
rect 13673 26630 13675 26682
rect 13855 26630 13857 26682
rect 13611 26628 13617 26630
rect 13673 26628 13697 26630
rect 13753 26628 13777 26630
rect 13833 26628 13857 26630
rect 13913 26628 13919 26630
rect 13611 26619 13919 26628
rect 13360 26580 13412 26586
rect 13360 26522 13412 26528
rect 13372 25974 13400 26522
rect 13452 26308 13504 26314
rect 13452 26250 13504 26256
rect 13360 25968 13412 25974
rect 13360 25910 13412 25916
rect 13464 25906 13492 26250
rect 13452 25900 13504 25906
rect 13452 25842 13504 25848
rect 14464 25764 14516 25770
rect 14464 25706 14516 25712
rect 13611 25596 13919 25605
rect 13611 25594 13617 25596
rect 13673 25594 13697 25596
rect 13753 25594 13777 25596
rect 13833 25594 13857 25596
rect 13913 25594 13919 25596
rect 13673 25542 13675 25594
rect 13855 25542 13857 25594
rect 13611 25540 13617 25542
rect 13673 25540 13697 25542
rect 13753 25540 13777 25542
rect 13833 25540 13857 25542
rect 13913 25540 13919 25542
rect 13611 25531 13919 25540
rect 13452 25152 13504 25158
rect 13452 25094 13504 25100
rect 13464 24274 13492 25094
rect 13611 24508 13919 24517
rect 13611 24506 13617 24508
rect 13673 24506 13697 24508
rect 13753 24506 13777 24508
rect 13833 24506 13857 24508
rect 13913 24506 13919 24508
rect 13673 24454 13675 24506
rect 13855 24454 13857 24506
rect 13611 24452 13617 24454
rect 13673 24452 13697 24454
rect 13753 24452 13777 24454
rect 13833 24452 13857 24454
rect 13913 24452 13919 24454
rect 13611 24443 13919 24452
rect 13452 24268 13504 24274
rect 13452 24210 13504 24216
rect 13176 23656 13228 23662
rect 13228 23616 13400 23644
rect 13176 23598 13228 23604
rect 13268 22636 13320 22642
rect 13268 22578 13320 22584
rect 13084 22568 13136 22574
rect 13084 22510 13136 22516
rect 13176 22432 13228 22438
rect 13176 22374 13228 22380
rect 13084 22160 13136 22166
rect 13084 22102 13136 22108
rect 13096 21146 13124 22102
rect 13188 22030 13216 22374
rect 13280 22166 13308 22578
rect 13268 22160 13320 22166
rect 13268 22102 13320 22108
rect 13176 22024 13228 22030
rect 13176 21966 13228 21972
rect 13084 21140 13136 21146
rect 13084 21082 13136 21088
rect 13176 20324 13228 20330
rect 13176 20266 13228 20272
rect 12900 20256 12952 20262
rect 12900 20198 12952 20204
rect 12912 17610 12940 20198
rect 13188 19854 13216 20266
rect 13176 19848 13228 19854
rect 13176 19790 13228 19796
rect 13268 19372 13320 19378
rect 13268 19314 13320 19320
rect 12992 18284 13044 18290
rect 12992 18226 13044 18232
rect 12900 17604 12952 17610
rect 12900 17546 12952 17552
rect 13004 17542 13032 18226
rect 12992 17536 13044 17542
rect 12992 17478 13044 17484
rect 12808 13524 12860 13530
rect 12808 13466 12860 13472
rect 12808 13388 12860 13394
rect 12808 13330 12860 13336
rect 12820 13190 12848 13330
rect 12808 13184 12860 13190
rect 12808 13126 12860 13132
rect 13004 12918 13032 17478
rect 13280 16250 13308 19314
rect 13372 17270 13400 23616
rect 13611 23420 13919 23429
rect 13611 23418 13617 23420
rect 13673 23418 13697 23420
rect 13753 23418 13777 23420
rect 13833 23418 13857 23420
rect 13913 23418 13919 23420
rect 13673 23366 13675 23418
rect 13855 23366 13857 23418
rect 13611 23364 13617 23366
rect 13673 23364 13697 23366
rect 13753 23364 13777 23366
rect 13833 23364 13857 23366
rect 13913 23364 13919 23366
rect 13611 23355 13919 23364
rect 14004 23316 14056 23322
rect 14004 23258 14056 23264
rect 13611 22332 13919 22341
rect 13611 22330 13617 22332
rect 13673 22330 13697 22332
rect 13753 22330 13777 22332
rect 13833 22330 13857 22332
rect 13913 22330 13919 22332
rect 13673 22278 13675 22330
rect 13855 22278 13857 22330
rect 13611 22276 13617 22278
rect 13673 22276 13697 22278
rect 13753 22276 13777 22278
rect 13833 22276 13857 22278
rect 13913 22276 13919 22278
rect 13611 22267 13919 22276
rect 14016 21554 14044 23258
rect 14096 22568 14148 22574
rect 14096 22510 14148 22516
rect 14004 21548 14056 21554
rect 14004 21490 14056 21496
rect 13611 21244 13919 21253
rect 13611 21242 13617 21244
rect 13673 21242 13697 21244
rect 13753 21242 13777 21244
rect 13833 21242 13857 21244
rect 13913 21242 13919 21244
rect 13673 21190 13675 21242
rect 13855 21190 13857 21242
rect 13611 21188 13617 21190
rect 13673 21188 13697 21190
rect 13753 21188 13777 21190
rect 13833 21188 13857 21190
rect 13913 21188 13919 21190
rect 13611 21179 13919 21188
rect 13452 20936 13504 20942
rect 13452 20878 13504 20884
rect 13464 19854 13492 20878
rect 13728 20392 13780 20398
rect 14108 20346 14136 22510
rect 14476 20942 14504 25706
rect 14568 24206 14596 27950
rect 15384 27940 15436 27946
rect 15384 27882 15436 27888
rect 14740 26036 14792 26042
rect 14740 25978 14792 25984
rect 14648 24404 14700 24410
rect 14648 24346 14700 24352
rect 14556 24200 14608 24206
rect 14556 24142 14608 24148
rect 14660 23798 14688 24346
rect 14648 23792 14700 23798
rect 14648 23734 14700 23740
rect 14660 22574 14688 23734
rect 14752 23662 14780 25978
rect 15396 25294 15424 27882
rect 15292 25288 15344 25294
rect 15292 25230 15344 25236
rect 15384 25288 15436 25294
rect 15384 25230 15436 25236
rect 15200 25152 15252 25158
rect 15200 25094 15252 25100
rect 15212 24818 15240 25094
rect 15200 24812 15252 24818
rect 15200 24754 15252 24760
rect 15200 24608 15252 24614
rect 15200 24550 15252 24556
rect 14832 24200 14884 24206
rect 14832 24142 14884 24148
rect 14740 23656 14792 23662
rect 14740 23598 14792 23604
rect 14752 23118 14780 23598
rect 14740 23112 14792 23118
rect 14740 23054 14792 23060
rect 14740 22976 14792 22982
rect 14740 22918 14792 22924
rect 14752 22642 14780 22918
rect 14740 22636 14792 22642
rect 14740 22578 14792 22584
rect 14648 22568 14700 22574
rect 14648 22510 14700 22516
rect 14464 20936 14516 20942
rect 14464 20878 14516 20884
rect 14280 20800 14332 20806
rect 14280 20742 14332 20748
rect 14292 20534 14320 20742
rect 14280 20528 14332 20534
rect 14280 20470 14332 20476
rect 13780 20340 14136 20346
rect 13728 20334 14136 20340
rect 13740 20330 14136 20334
rect 14844 20330 14872 24142
rect 15212 23798 15240 24550
rect 15200 23792 15252 23798
rect 15200 23734 15252 23740
rect 15212 23118 15240 23734
rect 15304 23662 15332 25230
rect 15396 25158 15424 25230
rect 15488 25226 15516 28018
rect 15764 26994 15792 28426
rect 15844 27464 15896 27470
rect 15844 27406 15896 27412
rect 15660 26988 15712 26994
rect 15660 26930 15712 26936
rect 15752 26988 15804 26994
rect 15752 26930 15804 26936
rect 15672 26246 15700 26930
rect 15660 26240 15712 26246
rect 15660 26182 15712 26188
rect 15672 25498 15700 26182
rect 15660 25492 15712 25498
rect 15660 25434 15712 25440
rect 15476 25220 15528 25226
rect 15476 25162 15528 25168
rect 15384 25152 15436 25158
rect 15384 25094 15436 25100
rect 15396 24970 15424 25094
rect 15396 24942 15516 24970
rect 15384 24812 15436 24818
rect 15384 24754 15436 24760
rect 15396 23866 15424 24754
rect 15384 23860 15436 23866
rect 15384 23802 15436 23808
rect 15292 23656 15344 23662
rect 15292 23598 15344 23604
rect 15292 23520 15344 23526
rect 15292 23462 15344 23468
rect 15304 23186 15332 23462
rect 15396 23186 15424 23802
rect 15292 23180 15344 23186
rect 15292 23122 15344 23128
rect 15384 23180 15436 23186
rect 15384 23122 15436 23128
rect 15200 23112 15252 23118
rect 15200 23054 15252 23060
rect 15488 22710 15516 24942
rect 15568 24676 15620 24682
rect 15568 24618 15620 24624
rect 15580 24070 15608 24618
rect 15764 24342 15792 26930
rect 15856 26382 15884 27406
rect 15844 26376 15896 26382
rect 15844 26318 15896 26324
rect 15856 24342 15884 26318
rect 15752 24336 15804 24342
rect 15752 24278 15804 24284
rect 15844 24336 15896 24342
rect 15844 24278 15896 24284
rect 15948 24206 15976 28562
rect 16028 28144 16080 28150
rect 16028 28086 16080 28092
rect 16040 27606 16068 28086
rect 16028 27600 16080 27606
rect 16028 27542 16080 27548
rect 16040 27470 16068 27542
rect 16028 27464 16080 27470
rect 16028 27406 16080 27412
rect 15936 24200 15988 24206
rect 15936 24142 15988 24148
rect 15660 24132 15712 24138
rect 15660 24074 15712 24080
rect 15568 24064 15620 24070
rect 15568 24006 15620 24012
rect 15580 23730 15608 24006
rect 15568 23724 15620 23730
rect 15568 23666 15620 23672
rect 15476 22704 15528 22710
rect 15476 22646 15528 22652
rect 15672 22642 15700 24074
rect 15948 23730 15976 24142
rect 15936 23724 15988 23730
rect 15936 23666 15988 23672
rect 15660 22636 15712 22642
rect 15660 22578 15712 22584
rect 15292 21548 15344 21554
rect 15292 21490 15344 21496
rect 15752 21548 15804 21554
rect 15752 21490 15804 21496
rect 15108 20460 15160 20466
rect 15108 20402 15160 20408
rect 13740 20324 14148 20330
rect 13740 20318 14096 20324
rect 14096 20266 14148 20272
rect 14832 20324 14884 20330
rect 14832 20266 14884 20272
rect 13611 20156 13919 20165
rect 13611 20154 13617 20156
rect 13673 20154 13697 20156
rect 13753 20154 13777 20156
rect 13833 20154 13857 20156
rect 13913 20154 13919 20156
rect 13673 20102 13675 20154
rect 13855 20102 13857 20154
rect 13611 20100 13617 20102
rect 13673 20100 13697 20102
rect 13753 20100 13777 20102
rect 13833 20100 13857 20102
rect 13913 20100 13919 20102
rect 13611 20091 13919 20100
rect 15120 19922 15148 20402
rect 15304 20058 15332 21490
rect 15384 21344 15436 21350
rect 15384 21286 15436 21292
rect 15396 20466 15424 21286
rect 15764 20466 15792 21490
rect 15844 21344 15896 21350
rect 15844 21286 15896 21292
rect 15936 21344 15988 21350
rect 15936 21286 15988 21292
rect 15856 20806 15884 21286
rect 15948 20874 15976 21286
rect 15936 20868 15988 20874
rect 15936 20810 15988 20816
rect 15844 20800 15896 20806
rect 15844 20742 15896 20748
rect 15384 20460 15436 20466
rect 15384 20402 15436 20408
rect 15752 20460 15804 20466
rect 15752 20402 15804 20408
rect 15292 20052 15344 20058
rect 15292 19994 15344 20000
rect 15108 19916 15160 19922
rect 15108 19858 15160 19864
rect 13452 19848 13504 19854
rect 13452 19790 13504 19796
rect 14464 19848 14516 19854
rect 14464 19790 14516 19796
rect 13360 17264 13412 17270
rect 13360 17206 13412 17212
rect 13268 16244 13320 16250
rect 13268 16186 13320 16192
rect 13280 15570 13308 16186
rect 13464 16182 13492 19790
rect 13611 19068 13919 19077
rect 13611 19066 13617 19068
rect 13673 19066 13697 19068
rect 13753 19066 13777 19068
rect 13833 19066 13857 19068
rect 13913 19066 13919 19068
rect 13673 19014 13675 19066
rect 13855 19014 13857 19066
rect 13611 19012 13617 19014
rect 13673 19012 13697 19014
rect 13753 19012 13777 19014
rect 13833 19012 13857 19014
rect 13913 19012 13919 19014
rect 13611 19003 13919 19012
rect 13611 17980 13919 17989
rect 13611 17978 13617 17980
rect 13673 17978 13697 17980
rect 13753 17978 13777 17980
rect 13833 17978 13857 17980
rect 13913 17978 13919 17980
rect 13673 17926 13675 17978
rect 13855 17926 13857 17978
rect 13611 17924 13617 17926
rect 13673 17924 13697 17926
rect 13753 17924 13777 17926
rect 13833 17924 13857 17926
rect 13913 17924 13919 17926
rect 13611 17915 13919 17924
rect 13544 17672 13596 17678
rect 13544 17614 13596 17620
rect 13556 17202 13584 17614
rect 14476 17338 14504 19790
rect 14740 19304 14792 19310
rect 14740 19246 14792 19252
rect 14752 18766 14780 19246
rect 14740 18760 14792 18766
rect 14740 18702 14792 18708
rect 14752 18358 14780 18702
rect 14740 18352 14792 18358
rect 14740 18294 14792 18300
rect 14464 17332 14516 17338
rect 14464 17274 14516 17280
rect 13544 17196 13596 17202
rect 13544 17138 13596 17144
rect 13611 16892 13919 16901
rect 13611 16890 13617 16892
rect 13673 16890 13697 16892
rect 13753 16890 13777 16892
rect 13833 16890 13857 16892
rect 13913 16890 13919 16892
rect 13673 16838 13675 16890
rect 13855 16838 13857 16890
rect 13611 16836 13617 16838
rect 13673 16836 13697 16838
rect 13753 16836 13777 16838
rect 13833 16836 13857 16838
rect 13913 16836 13919 16838
rect 13611 16827 13919 16836
rect 14740 16652 14792 16658
rect 14740 16594 14792 16600
rect 14464 16448 14516 16454
rect 14464 16390 14516 16396
rect 13452 16176 13504 16182
rect 13452 16118 13504 16124
rect 14280 16108 14332 16114
rect 14280 16050 14332 16056
rect 13611 15804 13919 15813
rect 13611 15802 13617 15804
rect 13673 15802 13697 15804
rect 13753 15802 13777 15804
rect 13833 15802 13857 15804
rect 13913 15802 13919 15804
rect 13673 15750 13675 15802
rect 13855 15750 13857 15802
rect 13611 15748 13617 15750
rect 13673 15748 13697 15750
rect 13753 15748 13777 15750
rect 13833 15748 13857 15750
rect 13913 15748 13919 15750
rect 13611 15739 13919 15748
rect 13268 15564 13320 15570
rect 13268 15506 13320 15512
rect 13452 14884 13504 14890
rect 13452 14826 13504 14832
rect 13084 14340 13136 14346
rect 13084 14282 13136 14288
rect 13096 14006 13124 14282
rect 13084 14000 13136 14006
rect 13084 13942 13136 13948
rect 13268 13524 13320 13530
rect 13268 13466 13320 13472
rect 13084 13184 13136 13190
rect 13084 13126 13136 13132
rect 12992 12912 13044 12918
rect 12992 12854 13044 12860
rect 12728 12406 12848 12434
rect 12360 11342 12572 11370
rect 12164 11212 12216 11218
rect 12164 11154 12216 11160
rect 12176 10606 12204 11154
rect 12360 10742 12388 11342
rect 12544 11150 12572 11342
rect 12532 11144 12584 11150
rect 12532 11086 12584 11092
rect 12440 11076 12492 11082
rect 12440 11018 12492 11024
rect 12624 11076 12676 11082
rect 12624 11018 12676 11024
rect 12348 10736 12400 10742
rect 12348 10678 12400 10684
rect 12452 10674 12480 11018
rect 12532 10736 12584 10742
rect 12532 10678 12584 10684
rect 12440 10668 12492 10674
rect 12440 10610 12492 10616
rect 12164 10600 12216 10606
rect 12164 10542 12216 10548
rect 12072 9988 12124 9994
rect 12072 9930 12124 9936
rect 12544 9178 12572 10678
rect 12636 10266 12664 11018
rect 12716 11008 12768 11014
rect 12716 10950 12768 10956
rect 12624 10260 12676 10266
rect 12624 10202 12676 10208
rect 12728 9450 12756 10950
rect 12716 9444 12768 9450
rect 12716 9386 12768 9392
rect 12532 9172 12584 9178
rect 12532 9114 12584 9120
rect 11888 7336 11940 7342
rect 11888 7278 11940 7284
rect 11900 5778 11928 7278
rect 12532 7200 12584 7206
rect 12532 7142 12584 7148
rect 12544 6458 12572 7142
rect 12820 6730 12848 12406
rect 13096 11150 13124 13126
rect 12900 11144 12952 11150
rect 12900 11086 12952 11092
rect 13084 11144 13136 11150
rect 13084 11086 13136 11092
rect 12912 10742 12940 11086
rect 12900 10736 12952 10742
rect 12900 10678 12952 10684
rect 13084 7336 13136 7342
rect 13084 7278 13136 7284
rect 13096 7002 13124 7278
rect 13084 6996 13136 7002
rect 13084 6938 13136 6944
rect 12808 6724 12860 6730
rect 12808 6666 12860 6672
rect 12532 6452 12584 6458
rect 12532 6394 12584 6400
rect 12348 6248 12400 6254
rect 12348 6190 12400 6196
rect 11888 5772 11940 5778
rect 11888 5714 11940 5720
rect 11796 5228 11848 5234
rect 11796 5170 11848 5176
rect 11704 5160 11756 5166
rect 11704 5102 11756 5108
rect 10876 4820 10928 4826
rect 10876 4762 10928 4768
rect 10416 4548 10468 4554
rect 10416 4490 10468 4496
rect 10428 4146 10456 4490
rect 11808 4486 11836 5170
rect 11900 4826 11928 5714
rect 12360 5710 12388 6190
rect 12348 5704 12400 5710
rect 12348 5646 12400 5652
rect 12716 5704 12768 5710
rect 12716 5646 12768 5652
rect 11888 4820 11940 4826
rect 11888 4762 11940 4768
rect 11796 4480 11848 4486
rect 11796 4422 11848 4428
rect 10416 4140 10468 4146
rect 10416 4082 10468 4088
rect 10508 4140 10560 4146
rect 10508 4082 10560 4088
rect 10784 4140 10836 4146
rect 10784 4082 10836 4088
rect 10520 3534 10548 4082
rect 10796 3602 10824 4082
rect 11900 4078 11928 4762
rect 12360 4622 12388 5646
rect 12728 5370 12756 5646
rect 12716 5364 12768 5370
rect 12716 5306 12768 5312
rect 13280 4826 13308 13466
rect 13464 11082 13492 14826
rect 13611 14716 13919 14725
rect 13611 14714 13617 14716
rect 13673 14714 13697 14716
rect 13753 14714 13777 14716
rect 13833 14714 13857 14716
rect 13913 14714 13919 14716
rect 13673 14662 13675 14714
rect 13855 14662 13857 14714
rect 13611 14660 13617 14662
rect 13673 14660 13697 14662
rect 13753 14660 13777 14662
rect 13833 14660 13857 14662
rect 13913 14660 13919 14662
rect 13611 14651 13919 14660
rect 14004 13932 14056 13938
rect 14004 13874 14056 13880
rect 13611 13628 13919 13637
rect 13611 13626 13617 13628
rect 13673 13626 13697 13628
rect 13753 13626 13777 13628
rect 13833 13626 13857 13628
rect 13913 13626 13919 13628
rect 13673 13574 13675 13626
rect 13855 13574 13857 13626
rect 13611 13572 13617 13574
rect 13673 13572 13697 13574
rect 13753 13572 13777 13574
rect 13833 13572 13857 13574
rect 13913 13572 13919 13574
rect 13611 13563 13919 13572
rect 14016 13326 14044 13874
rect 14292 13530 14320 16050
rect 14476 15910 14504 16390
rect 14752 16046 14780 16594
rect 14740 16040 14792 16046
rect 14740 15982 14792 15988
rect 14464 15904 14516 15910
rect 14464 15846 14516 15852
rect 14372 14612 14424 14618
rect 14372 14554 14424 14560
rect 14280 13524 14332 13530
rect 14280 13466 14332 13472
rect 14004 13320 14056 13326
rect 14004 13262 14056 13268
rect 13611 12540 13919 12549
rect 13611 12538 13617 12540
rect 13673 12538 13697 12540
rect 13753 12538 13777 12540
rect 13833 12538 13857 12540
rect 13913 12538 13919 12540
rect 13673 12486 13675 12538
rect 13855 12486 13857 12538
rect 13611 12484 13617 12486
rect 13673 12484 13697 12486
rect 13753 12484 13777 12486
rect 13833 12484 13857 12486
rect 13913 12484 13919 12486
rect 13611 12475 13919 12484
rect 14016 12442 14044 13262
rect 14384 13258 14412 14554
rect 14556 13932 14608 13938
rect 14556 13874 14608 13880
rect 14568 13258 14596 13874
rect 14372 13252 14424 13258
rect 14372 13194 14424 13200
rect 14556 13252 14608 13258
rect 14556 13194 14608 13200
rect 14568 12782 14596 13194
rect 14752 12918 14780 15982
rect 15120 14890 15148 19858
rect 15764 19854 15792 20402
rect 15856 19854 15884 20742
rect 16224 20534 16252 32778
rect 16776 32230 16804 32778
rect 17831 32668 18139 32677
rect 17831 32666 17837 32668
rect 17893 32666 17917 32668
rect 17973 32666 17997 32668
rect 18053 32666 18077 32668
rect 18133 32666 18139 32668
rect 17893 32614 17895 32666
rect 18075 32614 18077 32666
rect 17831 32612 17837 32614
rect 17893 32612 17917 32614
rect 17973 32612 17997 32614
rect 18053 32612 18077 32614
rect 18133 32612 18139 32614
rect 17831 32603 18139 32612
rect 17868 32428 17920 32434
rect 17868 32370 17920 32376
rect 18236 32428 18288 32434
rect 18236 32370 18288 32376
rect 17408 32360 17460 32366
rect 17408 32302 17460 32308
rect 16764 32224 16816 32230
rect 16764 32166 16816 32172
rect 16672 31952 16724 31958
rect 16672 31894 16724 31900
rect 16304 31340 16356 31346
rect 16304 31282 16356 31288
rect 16316 30666 16344 31282
rect 16684 30734 16712 31894
rect 16776 31754 16804 32166
rect 17132 31884 17184 31890
rect 17132 31826 17184 31832
rect 16776 31726 16896 31754
rect 16672 30728 16724 30734
rect 16672 30670 16724 30676
rect 16304 30660 16356 30666
rect 16304 30602 16356 30608
rect 16304 25424 16356 25430
rect 16304 25366 16356 25372
rect 16316 24818 16344 25366
rect 16396 25152 16448 25158
rect 16396 25094 16448 25100
rect 16304 24812 16356 24818
rect 16304 24754 16356 24760
rect 16408 24614 16436 25094
rect 16396 24608 16448 24614
rect 16396 24550 16448 24556
rect 16580 23588 16632 23594
rect 16580 23530 16632 23536
rect 16592 23186 16620 23530
rect 16580 23180 16632 23186
rect 16580 23122 16632 23128
rect 16396 22636 16448 22642
rect 16396 22578 16448 22584
rect 16408 22234 16436 22578
rect 16396 22228 16448 22234
rect 16396 22170 16448 22176
rect 16212 20528 16264 20534
rect 16212 20470 16264 20476
rect 15752 19848 15804 19854
rect 15752 19790 15804 19796
rect 15844 19848 15896 19854
rect 15844 19790 15896 19796
rect 15292 19712 15344 19718
rect 15292 19654 15344 19660
rect 15304 18766 15332 19654
rect 15292 18760 15344 18766
rect 15292 18702 15344 18708
rect 16212 18692 16264 18698
rect 16212 18634 16264 18640
rect 15292 18352 15344 18358
rect 15292 18294 15344 18300
rect 15200 16720 15252 16726
rect 15200 16662 15252 16668
rect 15212 16182 15240 16662
rect 15304 16522 15332 18294
rect 15844 18080 15896 18086
rect 15844 18022 15896 18028
rect 15856 16590 15884 18022
rect 16224 17202 16252 18634
rect 16212 17196 16264 17202
rect 16212 17138 16264 17144
rect 16304 17128 16356 17134
rect 16304 17070 16356 17076
rect 16316 16726 16344 17070
rect 16304 16720 16356 16726
rect 16304 16662 16356 16668
rect 15844 16584 15896 16590
rect 15844 16526 15896 16532
rect 16316 16522 16344 16662
rect 15292 16516 15344 16522
rect 15292 16458 15344 16464
rect 16120 16516 16172 16522
rect 16120 16458 16172 16464
rect 16304 16516 16356 16522
rect 16304 16458 16356 16464
rect 15200 16176 15252 16182
rect 15200 16118 15252 16124
rect 15304 15434 15332 16458
rect 15292 15428 15344 15434
rect 15292 15370 15344 15376
rect 15108 14884 15160 14890
rect 15108 14826 15160 14832
rect 15200 13932 15252 13938
rect 15200 13874 15252 13880
rect 15568 13932 15620 13938
rect 15568 13874 15620 13880
rect 15212 13190 15240 13874
rect 15580 13394 15608 13874
rect 15568 13388 15620 13394
rect 15568 13330 15620 13336
rect 15752 13320 15804 13326
rect 15752 13262 15804 13268
rect 15200 13184 15252 13190
rect 15200 13126 15252 13132
rect 14740 12912 14792 12918
rect 14740 12854 14792 12860
rect 15108 12844 15160 12850
rect 15108 12786 15160 12792
rect 14556 12776 14608 12782
rect 14556 12718 14608 12724
rect 14568 12646 14596 12718
rect 14556 12640 14608 12646
rect 14556 12582 14608 12588
rect 14004 12436 14056 12442
rect 14004 12378 14056 12384
rect 13611 11452 13919 11461
rect 13611 11450 13617 11452
rect 13673 11450 13697 11452
rect 13753 11450 13777 11452
rect 13833 11450 13857 11452
rect 13913 11450 13919 11452
rect 13673 11398 13675 11450
rect 13855 11398 13857 11450
rect 13611 11396 13617 11398
rect 13673 11396 13697 11398
rect 13753 11396 13777 11398
rect 13833 11396 13857 11398
rect 13913 11396 13919 11398
rect 13611 11387 13919 11396
rect 13452 11076 13504 11082
rect 13452 11018 13504 11024
rect 14016 10742 14044 12378
rect 14568 12238 14596 12582
rect 15120 12442 15148 12786
rect 15108 12436 15160 12442
rect 15108 12378 15160 12384
rect 15120 12238 15148 12378
rect 14556 12232 14608 12238
rect 14556 12174 14608 12180
rect 15108 12232 15160 12238
rect 15108 12174 15160 12180
rect 15212 11762 15240 13126
rect 15764 12238 15792 13262
rect 16132 12481 16160 16458
rect 16304 16108 16356 16114
rect 16304 16050 16356 16056
rect 16316 15502 16344 16050
rect 16304 15496 16356 15502
rect 16304 15438 16356 15444
rect 16212 15020 16264 15026
rect 16316 15008 16344 15438
rect 16408 15366 16436 22170
rect 16764 19780 16816 19786
rect 16764 19722 16816 19728
rect 16776 19446 16804 19722
rect 16764 19440 16816 19446
rect 16764 19382 16816 19388
rect 16672 18352 16724 18358
rect 16672 18294 16724 18300
rect 16684 16454 16712 18294
rect 16672 16448 16724 16454
rect 16672 16390 16724 16396
rect 16580 15564 16632 15570
rect 16580 15506 16632 15512
rect 16396 15360 16448 15366
rect 16396 15302 16448 15308
rect 16264 14980 16344 15008
rect 16212 14962 16264 14968
rect 16224 13802 16252 14962
rect 16212 13796 16264 13802
rect 16212 13738 16264 13744
rect 16592 12782 16620 15506
rect 16672 15020 16724 15026
rect 16672 14962 16724 14968
rect 16684 14006 16712 14962
rect 16672 14000 16724 14006
rect 16672 13942 16724 13948
rect 16580 12776 16632 12782
rect 16580 12718 16632 12724
rect 16118 12472 16174 12481
rect 16174 12416 16252 12434
rect 16118 12407 16252 12416
rect 16132 12406 16252 12407
rect 15752 12232 15804 12238
rect 15752 12174 15804 12180
rect 15764 11830 15792 12174
rect 15752 11824 15804 11830
rect 15752 11766 15804 11772
rect 15200 11756 15252 11762
rect 15200 11698 15252 11704
rect 15936 11280 15988 11286
rect 15936 11222 15988 11228
rect 14004 10736 14056 10742
rect 14004 10678 14056 10684
rect 14372 10464 14424 10470
rect 14372 10406 14424 10412
rect 13611 10364 13919 10373
rect 13611 10362 13617 10364
rect 13673 10362 13697 10364
rect 13753 10362 13777 10364
rect 13833 10362 13857 10364
rect 13913 10362 13919 10364
rect 13673 10310 13675 10362
rect 13855 10310 13857 10362
rect 13611 10308 13617 10310
rect 13673 10308 13697 10310
rect 13753 10308 13777 10310
rect 13833 10308 13857 10310
rect 13913 10308 13919 10310
rect 13611 10299 13919 10308
rect 13360 9920 13412 9926
rect 13360 9862 13412 9868
rect 13268 4820 13320 4826
rect 13268 4762 13320 4768
rect 12348 4616 12400 4622
rect 12348 4558 12400 4564
rect 13372 4282 13400 9862
rect 13611 9276 13919 9285
rect 13611 9274 13617 9276
rect 13673 9274 13697 9276
rect 13753 9274 13777 9276
rect 13833 9274 13857 9276
rect 13913 9274 13919 9276
rect 13673 9222 13675 9274
rect 13855 9222 13857 9274
rect 13611 9220 13617 9222
rect 13673 9220 13697 9222
rect 13753 9220 13777 9222
rect 13833 9220 13857 9222
rect 13913 9220 13919 9222
rect 13611 9211 13919 9220
rect 13611 8188 13919 8197
rect 13611 8186 13617 8188
rect 13673 8186 13697 8188
rect 13753 8186 13777 8188
rect 13833 8186 13857 8188
rect 13913 8186 13919 8188
rect 13673 8134 13675 8186
rect 13855 8134 13857 8186
rect 13611 8132 13617 8134
rect 13673 8132 13697 8134
rect 13753 8132 13777 8134
rect 13833 8132 13857 8134
rect 13913 8132 13919 8134
rect 13611 8123 13919 8132
rect 13611 7100 13919 7109
rect 13611 7098 13617 7100
rect 13673 7098 13697 7100
rect 13753 7098 13777 7100
rect 13833 7098 13857 7100
rect 13913 7098 13919 7100
rect 13673 7046 13675 7098
rect 13855 7046 13857 7098
rect 13611 7044 13617 7046
rect 13673 7044 13697 7046
rect 13753 7044 13777 7046
rect 13833 7044 13857 7046
rect 13913 7044 13919 7046
rect 13611 7035 13919 7044
rect 13636 6656 13688 6662
rect 13636 6598 13688 6604
rect 13648 6390 13676 6598
rect 13636 6384 13688 6390
rect 13636 6326 13688 6332
rect 13611 6012 13919 6021
rect 13611 6010 13617 6012
rect 13673 6010 13697 6012
rect 13753 6010 13777 6012
rect 13833 6010 13857 6012
rect 13913 6010 13919 6012
rect 13673 5958 13675 6010
rect 13855 5958 13857 6010
rect 13611 5956 13617 5958
rect 13673 5956 13697 5958
rect 13753 5956 13777 5958
rect 13833 5956 13857 5958
rect 13913 5956 13919 5958
rect 13611 5947 13919 5956
rect 14280 5568 14332 5574
rect 14280 5510 14332 5516
rect 13611 4924 13919 4933
rect 13611 4922 13617 4924
rect 13673 4922 13697 4924
rect 13753 4922 13777 4924
rect 13833 4922 13857 4924
rect 13913 4922 13919 4924
rect 13673 4870 13675 4922
rect 13855 4870 13857 4922
rect 13611 4868 13617 4870
rect 13673 4868 13697 4870
rect 13753 4868 13777 4870
rect 13833 4868 13857 4870
rect 13913 4868 13919 4870
rect 13611 4859 13919 4868
rect 14188 4684 14240 4690
rect 14188 4626 14240 4632
rect 13360 4276 13412 4282
rect 13360 4218 13412 4224
rect 14004 4140 14056 4146
rect 14004 4082 14056 4088
rect 11888 4072 11940 4078
rect 11888 4014 11940 4020
rect 12992 3936 13044 3942
rect 12992 3878 13044 3884
rect 10784 3596 10836 3602
rect 10784 3538 10836 3544
rect 10508 3528 10560 3534
rect 10508 3470 10560 3476
rect 10796 3058 10824 3538
rect 13004 3534 13032 3878
rect 13611 3836 13919 3845
rect 13611 3834 13617 3836
rect 13673 3834 13697 3836
rect 13753 3834 13777 3836
rect 13833 3834 13857 3836
rect 13913 3834 13919 3836
rect 13673 3782 13675 3834
rect 13855 3782 13857 3834
rect 13611 3780 13617 3782
rect 13673 3780 13697 3782
rect 13753 3780 13777 3782
rect 13833 3780 13857 3782
rect 13913 3780 13919 3782
rect 13611 3771 13919 3780
rect 14016 3738 14044 4082
rect 14200 4078 14228 4626
rect 14292 4622 14320 5510
rect 14280 4616 14332 4622
rect 14280 4558 14332 4564
rect 14188 4072 14240 4078
rect 14188 4014 14240 4020
rect 14004 3732 14056 3738
rect 14004 3674 14056 3680
rect 12348 3528 12400 3534
rect 12348 3470 12400 3476
rect 12992 3528 13044 3534
rect 12992 3470 13044 3476
rect 12360 3194 12388 3470
rect 12348 3188 12400 3194
rect 12348 3130 12400 3136
rect 10784 3052 10836 3058
rect 10784 2994 10836 3000
rect 13611 2748 13919 2757
rect 13611 2746 13617 2748
rect 13673 2746 13697 2748
rect 13753 2746 13777 2748
rect 13833 2746 13857 2748
rect 13913 2746 13919 2748
rect 13673 2694 13675 2746
rect 13855 2694 13857 2746
rect 13611 2692 13617 2694
rect 13673 2692 13697 2694
rect 13753 2692 13777 2694
rect 13833 2692 13857 2694
rect 13913 2692 13919 2694
rect 13611 2683 13919 2692
rect 10048 2576 10100 2582
rect 10048 2518 10100 2524
rect 14016 2446 14044 3674
rect 14200 2990 14228 4014
rect 14280 3392 14332 3398
rect 14280 3334 14332 3340
rect 14292 2990 14320 3334
rect 14384 3194 14412 10406
rect 15292 9376 15344 9382
rect 15292 9318 15344 9324
rect 15304 8974 15332 9318
rect 15108 8968 15160 8974
rect 15108 8910 15160 8916
rect 15292 8968 15344 8974
rect 15292 8910 15344 8916
rect 15120 7206 15148 8910
rect 15660 8084 15712 8090
rect 15660 8026 15712 8032
rect 15568 7812 15620 7818
rect 15568 7754 15620 7760
rect 15580 7546 15608 7754
rect 15568 7540 15620 7546
rect 15568 7482 15620 7488
rect 15672 7206 15700 8026
rect 15108 7200 15160 7206
rect 15108 7142 15160 7148
rect 15660 7200 15712 7206
rect 15660 7142 15712 7148
rect 15120 6866 15148 7142
rect 15108 6860 15160 6866
rect 15108 6802 15160 6808
rect 15672 6798 15700 7142
rect 15660 6792 15712 6798
rect 15660 6734 15712 6740
rect 15200 5228 15252 5234
rect 15200 5170 15252 5176
rect 14832 5024 14884 5030
rect 14832 4966 14884 4972
rect 14924 5024 14976 5030
rect 14924 4966 14976 4972
rect 14844 4282 14872 4966
rect 14832 4276 14884 4282
rect 14832 4218 14884 4224
rect 14936 4146 14964 4966
rect 14924 4140 14976 4146
rect 14924 4082 14976 4088
rect 14740 3460 14792 3466
rect 14740 3402 14792 3408
rect 14752 3194 14780 3402
rect 14372 3188 14424 3194
rect 14372 3130 14424 3136
rect 14740 3188 14792 3194
rect 14740 3130 14792 3136
rect 14188 2984 14240 2990
rect 14188 2926 14240 2932
rect 14280 2984 14332 2990
rect 14280 2926 14332 2932
rect 8944 2440 8996 2446
rect 8944 2382 8996 2388
rect 10232 2440 10284 2446
rect 10232 2382 10284 2388
rect 11520 2440 11572 2446
rect 11520 2382 11572 2388
rect 12808 2440 12860 2446
rect 12808 2382 12860 2388
rect 14004 2440 14056 2446
rect 14004 2382 14056 2388
rect 7840 2372 7892 2378
rect 7840 2314 7892 2320
rect 8956 800 8984 2382
rect 9390 2204 9698 2213
rect 9390 2202 9396 2204
rect 9452 2202 9476 2204
rect 9532 2202 9556 2204
rect 9612 2202 9636 2204
rect 9692 2202 9698 2204
rect 9452 2150 9454 2202
rect 9634 2150 9636 2202
rect 9390 2148 9396 2150
rect 9452 2148 9476 2150
rect 9532 2148 9556 2150
rect 9612 2148 9636 2150
rect 9692 2148 9698 2150
rect 9390 2139 9698 2148
rect 10244 800 10272 2382
rect 11532 800 11560 2382
rect 12820 800 12848 2382
rect 14096 2372 14148 2378
rect 14096 2314 14148 2320
rect 14108 800 14136 2314
rect 14384 2310 14412 3130
rect 15212 3058 15240 5170
rect 15948 4622 15976 11222
rect 16224 8634 16252 12406
rect 16304 12232 16356 12238
rect 16304 12174 16356 12180
rect 16316 11762 16344 12174
rect 16592 11762 16620 12718
rect 16868 12434 16896 31726
rect 17144 31346 17172 31826
rect 17316 31816 17368 31822
rect 17316 31758 17368 31764
rect 17328 31482 17356 31758
rect 17316 31476 17368 31482
rect 17316 31418 17368 31424
rect 17132 31340 17184 31346
rect 17132 31282 17184 31288
rect 17040 31136 17092 31142
rect 17040 31078 17092 31084
rect 17052 30734 17080 31078
rect 17420 30938 17448 32302
rect 17880 31822 17908 32370
rect 18248 32026 18276 32370
rect 19536 32298 19564 33322
rect 22052 33212 22360 33221
rect 22052 33210 22058 33212
rect 22114 33210 22138 33212
rect 22194 33210 22218 33212
rect 22274 33210 22298 33212
rect 22354 33210 22360 33212
rect 22114 33158 22116 33210
rect 22296 33158 22298 33210
rect 22052 33156 22058 33158
rect 22114 33156 22138 33158
rect 22194 33156 22218 33158
rect 22274 33156 22298 33158
rect 22354 33156 22360 33158
rect 22052 33147 22360 33156
rect 20628 32972 20680 32978
rect 20628 32914 20680 32920
rect 20812 32972 20864 32978
rect 20812 32914 20864 32920
rect 20536 32904 20588 32910
rect 20536 32846 20588 32852
rect 19524 32292 19576 32298
rect 19524 32234 19576 32240
rect 18512 32224 18564 32230
rect 18512 32166 18564 32172
rect 18236 32020 18288 32026
rect 18236 31962 18288 31968
rect 18524 31822 18552 32166
rect 20548 32042 20576 32846
rect 20456 32014 20576 32042
rect 20640 32026 20668 32914
rect 20824 32774 20852 32914
rect 20812 32768 20864 32774
rect 20812 32710 20864 32716
rect 21272 32768 21324 32774
rect 21272 32710 21324 32716
rect 22008 32768 22060 32774
rect 22008 32710 22060 32716
rect 21284 32366 21312 32710
rect 22020 32434 22048 32710
rect 22480 32570 22508 33322
rect 24584 33040 24636 33046
rect 24584 32982 24636 32988
rect 22928 32904 22980 32910
rect 22928 32846 22980 32852
rect 22468 32564 22520 32570
rect 22468 32506 22520 32512
rect 22008 32428 22060 32434
rect 22008 32370 22060 32376
rect 22560 32428 22612 32434
rect 22560 32370 22612 32376
rect 21272 32360 21324 32366
rect 21272 32302 21324 32308
rect 21180 32292 21232 32298
rect 21180 32234 21232 32240
rect 20628 32020 20680 32026
rect 17868 31816 17920 31822
rect 17696 31776 17868 31804
rect 17696 31346 17724 31776
rect 17868 31758 17920 31764
rect 18512 31816 18564 31822
rect 18512 31758 18564 31764
rect 17831 31580 18139 31589
rect 17831 31578 17837 31580
rect 17893 31578 17917 31580
rect 17973 31578 17997 31580
rect 18053 31578 18077 31580
rect 18133 31578 18139 31580
rect 17893 31526 17895 31578
rect 18075 31526 18077 31578
rect 17831 31524 17837 31526
rect 17893 31524 17917 31526
rect 17973 31524 17997 31526
rect 18053 31524 18077 31526
rect 18133 31524 18139 31526
rect 17831 31515 18139 31524
rect 20456 31414 20484 32014
rect 20628 31962 20680 31968
rect 20536 31952 20588 31958
rect 20536 31894 20588 31900
rect 20444 31408 20496 31414
rect 20444 31350 20496 31356
rect 17684 31340 17736 31346
rect 17684 31282 17736 31288
rect 20168 31340 20220 31346
rect 20168 31282 20220 31288
rect 17408 30932 17460 30938
rect 17408 30874 17460 30880
rect 17040 30728 17092 30734
rect 17040 30670 17092 30676
rect 18788 30660 18840 30666
rect 18788 30602 18840 30608
rect 17831 30492 18139 30501
rect 17831 30490 17837 30492
rect 17893 30490 17917 30492
rect 17973 30490 17997 30492
rect 18053 30490 18077 30492
rect 18133 30490 18139 30492
rect 17893 30438 17895 30490
rect 18075 30438 18077 30490
rect 17831 30436 17837 30438
rect 17893 30436 17917 30438
rect 17973 30436 17997 30438
rect 18053 30436 18077 30438
rect 18133 30436 18139 30438
rect 17831 30427 18139 30436
rect 18800 30326 18828 30602
rect 18788 30320 18840 30326
rect 18788 30262 18840 30268
rect 20180 29646 20208 31282
rect 20548 31278 20576 31894
rect 21192 31822 21220 32234
rect 22052 32124 22360 32133
rect 22052 32122 22058 32124
rect 22114 32122 22138 32124
rect 22194 32122 22218 32124
rect 22274 32122 22298 32124
rect 22354 32122 22360 32124
rect 22114 32070 22116 32122
rect 22296 32070 22298 32122
rect 22052 32068 22058 32070
rect 22114 32068 22138 32070
rect 22194 32068 22218 32070
rect 22274 32068 22298 32070
rect 22354 32068 22360 32070
rect 22052 32059 22360 32068
rect 22572 31958 22600 32370
rect 22940 32230 22968 32846
rect 24596 32434 24624 32982
rect 25424 32978 25452 33322
rect 25412 32972 25464 32978
rect 25412 32914 25464 32920
rect 28368 32842 28396 33322
rect 30493 33212 30801 33221
rect 30493 33210 30499 33212
rect 30555 33210 30579 33212
rect 30635 33210 30659 33212
rect 30715 33210 30739 33212
rect 30795 33210 30801 33212
rect 30555 33158 30557 33210
rect 30737 33158 30739 33210
rect 30493 33156 30499 33158
rect 30555 33156 30579 33158
rect 30635 33156 30659 33158
rect 30715 33156 30739 33158
rect 30795 33156 30801 33158
rect 30493 33147 30801 33156
rect 28356 32836 28408 32842
rect 28356 32778 28408 32784
rect 26272 32668 26580 32677
rect 26272 32666 26278 32668
rect 26334 32666 26358 32668
rect 26414 32666 26438 32668
rect 26494 32666 26518 32668
rect 26574 32666 26580 32668
rect 26334 32614 26336 32666
rect 26516 32614 26518 32666
rect 26272 32612 26278 32614
rect 26334 32612 26358 32614
rect 26414 32612 26438 32614
rect 26494 32612 26518 32614
rect 26574 32612 26580 32614
rect 26272 32603 26580 32612
rect 31312 32434 31340 33322
rect 33428 32434 33456 33322
rect 34713 32668 35021 32677
rect 34713 32666 34719 32668
rect 34775 32666 34799 32668
rect 34855 32666 34879 32668
rect 34935 32666 34959 32668
rect 35015 32666 35021 32668
rect 34775 32614 34777 32666
rect 34957 32614 34959 32666
rect 34713 32612 34719 32614
rect 34775 32612 34799 32614
rect 34855 32612 34879 32614
rect 34935 32612 34959 32614
rect 35015 32612 35021 32614
rect 34713 32603 35021 32612
rect 23296 32428 23348 32434
rect 23296 32370 23348 32376
rect 24584 32428 24636 32434
rect 24584 32370 24636 32376
rect 27712 32428 27764 32434
rect 27712 32370 27764 32376
rect 28632 32428 28684 32434
rect 28632 32370 28684 32376
rect 31300 32428 31352 32434
rect 31300 32370 31352 32376
rect 33416 32428 33468 32434
rect 33416 32370 33468 32376
rect 22744 32224 22796 32230
rect 22744 32166 22796 32172
rect 22928 32224 22980 32230
rect 22928 32166 22980 32172
rect 22560 31952 22612 31958
rect 22560 31894 22612 31900
rect 22756 31890 22784 32166
rect 22744 31884 22796 31890
rect 22744 31826 22796 31832
rect 20812 31816 20864 31822
rect 20812 31758 20864 31764
rect 21088 31816 21140 31822
rect 21088 31758 21140 31764
rect 21180 31816 21232 31822
rect 21180 31758 21232 31764
rect 20824 31482 20852 31758
rect 20812 31476 20864 31482
rect 20812 31418 20864 31424
rect 20996 31340 21048 31346
rect 20996 31282 21048 31288
rect 20536 31272 20588 31278
rect 20536 31214 20588 31220
rect 20260 30252 20312 30258
rect 20260 30194 20312 30200
rect 19248 29640 19300 29646
rect 19248 29582 19300 29588
rect 20168 29640 20220 29646
rect 20168 29582 20220 29588
rect 17831 29404 18139 29413
rect 17831 29402 17837 29404
rect 17893 29402 17917 29404
rect 17973 29402 17997 29404
rect 18053 29402 18077 29404
rect 18133 29402 18139 29404
rect 17893 29350 17895 29402
rect 18075 29350 18077 29402
rect 17831 29348 17837 29350
rect 17893 29348 17917 29350
rect 17973 29348 17997 29350
rect 18053 29348 18077 29350
rect 18133 29348 18139 29350
rect 17831 29339 18139 29348
rect 19260 28490 19288 29582
rect 19432 29504 19484 29510
rect 19432 29446 19484 29452
rect 19340 29232 19392 29238
rect 19340 29174 19392 29180
rect 19248 28484 19300 28490
rect 19248 28426 19300 28432
rect 17831 28316 18139 28325
rect 17831 28314 17837 28316
rect 17893 28314 17917 28316
rect 17973 28314 17997 28316
rect 18053 28314 18077 28316
rect 18133 28314 18139 28316
rect 17893 28262 17895 28314
rect 18075 28262 18077 28314
rect 17831 28260 17837 28262
rect 17893 28260 17917 28262
rect 17973 28260 17997 28262
rect 18053 28260 18077 28262
rect 18133 28260 18139 28262
rect 17831 28251 18139 28260
rect 19260 28082 19288 28426
rect 19248 28076 19300 28082
rect 19248 28018 19300 28024
rect 19352 28014 19380 29174
rect 19444 29170 19472 29446
rect 19432 29164 19484 29170
rect 19432 29106 19484 29112
rect 20180 29102 20208 29582
rect 20272 29306 20300 30194
rect 20548 29714 20576 31214
rect 20904 31204 20956 31210
rect 20904 31146 20956 31152
rect 20916 30410 20944 31146
rect 21008 30938 21036 31282
rect 20996 30932 21048 30938
rect 20996 30874 21048 30880
rect 20916 30382 21036 30410
rect 20720 30048 20772 30054
rect 20720 29990 20772 29996
rect 20536 29708 20588 29714
rect 20536 29650 20588 29656
rect 20260 29300 20312 29306
rect 20260 29242 20312 29248
rect 20444 29164 20496 29170
rect 20548 29152 20576 29650
rect 20732 29170 20760 29990
rect 20812 29640 20864 29646
rect 20812 29582 20864 29588
rect 20824 29170 20852 29582
rect 20496 29124 20576 29152
rect 20720 29164 20772 29170
rect 20444 29106 20496 29112
rect 20720 29106 20772 29112
rect 20812 29164 20864 29170
rect 20812 29106 20864 29112
rect 20168 29096 20220 29102
rect 20168 29038 20220 29044
rect 20824 28694 20852 29106
rect 20812 28688 20864 28694
rect 20812 28630 20864 28636
rect 19708 28552 19760 28558
rect 19708 28494 19760 28500
rect 19892 28552 19944 28558
rect 19892 28494 19944 28500
rect 19340 28008 19392 28014
rect 19340 27950 19392 27956
rect 18236 27464 18288 27470
rect 18236 27406 18288 27412
rect 17831 27228 18139 27237
rect 17831 27226 17837 27228
rect 17893 27226 17917 27228
rect 17973 27226 17997 27228
rect 18053 27226 18077 27228
rect 18133 27226 18139 27228
rect 17893 27174 17895 27226
rect 18075 27174 18077 27226
rect 17831 27172 17837 27174
rect 17893 27172 17917 27174
rect 17973 27172 17997 27174
rect 18053 27172 18077 27174
rect 18133 27172 18139 27174
rect 17831 27163 18139 27172
rect 18248 27130 18276 27406
rect 19248 27396 19300 27402
rect 19248 27338 19300 27344
rect 18236 27124 18288 27130
rect 18236 27066 18288 27072
rect 18248 26450 18276 27066
rect 18328 26988 18380 26994
rect 18328 26930 18380 26936
rect 18236 26444 18288 26450
rect 18236 26386 18288 26392
rect 17224 26376 17276 26382
rect 17224 26318 17276 26324
rect 16948 25900 17000 25906
rect 16948 25842 17000 25848
rect 16960 20398 16988 25842
rect 17236 25702 17264 26318
rect 17831 26140 18139 26149
rect 17831 26138 17837 26140
rect 17893 26138 17917 26140
rect 17973 26138 17997 26140
rect 18053 26138 18077 26140
rect 18133 26138 18139 26140
rect 17893 26086 17895 26138
rect 18075 26086 18077 26138
rect 17831 26084 17837 26086
rect 17893 26084 17917 26086
rect 17973 26084 17997 26086
rect 18053 26084 18077 26086
rect 18133 26084 18139 26086
rect 17831 26075 18139 26084
rect 18340 25702 18368 26930
rect 18420 26308 18472 26314
rect 18420 26250 18472 26256
rect 17224 25696 17276 25702
rect 17224 25638 17276 25644
rect 18328 25696 18380 25702
rect 18328 25638 18380 25644
rect 17236 24954 17264 25638
rect 17831 25052 18139 25061
rect 17831 25050 17837 25052
rect 17893 25050 17917 25052
rect 17973 25050 17997 25052
rect 18053 25050 18077 25052
rect 18133 25050 18139 25052
rect 17893 24998 17895 25050
rect 18075 24998 18077 25050
rect 17831 24996 17837 24998
rect 17893 24996 17917 24998
rect 17973 24996 17997 24998
rect 18053 24996 18077 24998
rect 18133 24996 18139 24998
rect 17831 24987 18139 24996
rect 17224 24948 17276 24954
rect 17224 24890 17276 24896
rect 17316 24744 17368 24750
rect 17316 24686 17368 24692
rect 17328 23186 17356 24686
rect 17960 24336 18012 24342
rect 17960 24278 18012 24284
rect 17972 24206 18000 24278
rect 18052 24268 18104 24274
rect 18236 24268 18288 24274
rect 18104 24228 18236 24256
rect 18052 24210 18104 24216
rect 18236 24210 18288 24216
rect 17960 24200 18012 24206
rect 17696 24148 17960 24154
rect 17696 24142 18012 24148
rect 17696 24126 18000 24142
rect 17408 24064 17460 24070
rect 17408 24006 17460 24012
rect 17592 24064 17644 24070
rect 17592 24006 17644 24012
rect 17420 23730 17448 24006
rect 17408 23724 17460 23730
rect 17408 23666 17460 23672
rect 17316 23180 17368 23186
rect 17316 23122 17368 23128
rect 17328 21146 17356 23122
rect 17420 22642 17448 23666
rect 17604 23118 17632 24006
rect 17592 23112 17644 23118
rect 17592 23054 17644 23060
rect 17500 23044 17552 23050
rect 17500 22986 17552 22992
rect 17512 22642 17540 22986
rect 17408 22636 17460 22642
rect 17408 22578 17460 22584
rect 17500 22636 17552 22642
rect 17500 22578 17552 22584
rect 17696 21554 17724 24126
rect 17831 23964 18139 23973
rect 17831 23962 17837 23964
rect 17893 23962 17917 23964
rect 17973 23962 17997 23964
rect 18053 23962 18077 23964
rect 18133 23962 18139 23964
rect 17893 23910 17895 23962
rect 18075 23910 18077 23962
rect 17831 23908 17837 23910
rect 17893 23908 17917 23910
rect 17973 23908 17997 23910
rect 18053 23908 18077 23910
rect 18133 23908 18139 23910
rect 17831 23899 18139 23908
rect 17831 22876 18139 22885
rect 17831 22874 17837 22876
rect 17893 22874 17917 22876
rect 17973 22874 17997 22876
rect 18053 22874 18077 22876
rect 18133 22874 18139 22876
rect 17893 22822 17895 22874
rect 18075 22822 18077 22874
rect 17831 22820 17837 22822
rect 17893 22820 17917 22822
rect 17973 22820 17997 22822
rect 18053 22820 18077 22822
rect 18133 22820 18139 22822
rect 17831 22811 18139 22820
rect 17960 22500 18012 22506
rect 17960 22442 18012 22448
rect 17972 22030 18000 22442
rect 18052 22432 18104 22438
rect 18052 22374 18104 22380
rect 18064 22098 18092 22374
rect 18052 22092 18104 22098
rect 18052 22034 18104 22040
rect 17960 22024 18012 22030
rect 17960 21966 18012 21972
rect 18236 21956 18288 21962
rect 18236 21898 18288 21904
rect 17831 21788 18139 21797
rect 17831 21786 17837 21788
rect 17893 21786 17917 21788
rect 17973 21786 17997 21788
rect 18053 21786 18077 21788
rect 18133 21786 18139 21788
rect 17893 21734 17895 21786
rect 18075 21734 18077 21786
rect 17831 21732 17837 21734
rect 17893 21732 17917 21734
rect 17973 21732 17997 21734
rect 18053 21732 18077 21734
rect 18133 21732 18139 21734
rect 17831 21723 18139 21732
rect 17684 21548 17736 21554
rect 17684 21490 17736 21496
rect 18248 21486 18276 21898
rect 18236 21480 18288 21486
rect 18236 21422 18288 21428
rect 17316 21140 17368 21146
rect 17316 21082 17368 21088
rect 18340 20942 18368 25638
rect 18432 24818 18460 26250
rect 19260 25974 19288 27338
rect 19352 26314 19380 27950
rect 19720 27878 19748 28494
rect 19904 28150 19932 28494
rect 20720 28484 20772 28490
rect 20720 28426 20772 28432
rect 20536 28416 20588 28422
rect 20536 28358 20588 28364
rect 19892 28144 19944 28150
rect 19892 28086 19944 28092
rect 19708 27872 19760 27878
rect 19708 27814 19760 27820
rect 19800 27328 19852 27334
rect 19800 27270 19852 27276
rect 19812 27062 19840 27270
rect 19800 27056 19852 27062
rect 19800 26998 19852 27004
rect 19340 26308 19392 26314
rect 19340 26250 19392 26256
rect 19248 25968 19300 25974
rect 19248 25910 19300 25916
rect 18420 24812 18472 24818
rect 18420 24754 18472 24760
rect 19352 24750 19380 26250
rect 19616 25900 19668 25906
rect 19616 25842 19668 25848
rect 19340 24744 19392 24750
rect 19340 24686 19392 24692
rect 18696 24132 18748 24138
rect 18696 24074 18748 24080
rect 18420 23656 18472 23662
rect 18420 23598 18472 23604
rect 18432 22030 18460 23598
rect 18708 23322 18736 24074
rect 18696 23316 18748 23322
rect 18696 23258 18748 23264
rect 18512 22976 18564 22982
rect 18512 22918 18564 22924
rect 18524 22710 18552 22918
rect 18708 22710 18736 23258
rect 19628 23254 19656 25842
rect 19812 25498 19840 26998
rect 20548 26926 20576 28358
rect 20732 28150 20760 28426
rect 20720 28144 20772 28150
rect 20720 28086 20772 28092
rect 21008 27402 21036 30382
rect 21100 28762 21128 31758
rect 21272 31748 21324 31754
rect 21272 31690 21324 31696
rect 22652 31748 22704 31754
rect 22652 31690 22704 31696
rect 21284 31210 21312 31690
rect 22664 31346 22692 31690
rect 22756 31346 22784 31826
rect 22940 31822 22968 32166
rect 23308 32026 23336 32370
rect 23388 32360 23440 32366
rect 23388 32302 23440 32308
rect 23296 32020 23348 32026
rect 23296 31962 23348 31968
rect 22928 31816 22980 31822
rect 22928 31758 22980 31764
rect 22652 31340 22704 31346
rect 22652 31282 22704 31288
rect 22744 31340 22796 31346
rect 22744 31282 22796 31288
rect 23020 31340 23072 31346
rect 23020 31282 23072 31288
rect 21456 31272 21508 31278
rect 21456 31214 21508 31220
rect 21272 31204 21324 31210
rect 21272 31146 21324 31152
rect 21468 30734 21496 31214
rect 22756 31210 22784 31282
rect 21732 31204 21784 31210
rect 21732 31146 21784 31152
rect 22744 31204 22796 31210
rect 22744 31146 22796 31152
rect 21456 30728 21508 30734
rect 21456 30670 21508 30676
rect 21272 30252 21324 30258
rect 21272 30194 21324 30200
rect 21284 29646 21312 30194
rect 21272 29640 21324 29646
rect 21272 29582 21324 29588
rect 21088 28756 21140 28762
rect 21088 28698 21140 28704
rect 21284 28626 21312 29582
rect 21468 29510 21496 30670
rect 21548 30320 21600 30326
rect 21548 30262 21600 30268
rect 21560 29714 21588 30262
rect 21548 29708 21600 29714
rect 21548 29650 21600 29656
rect 21456 29504 21508 29510
rect 21456 29446 21508 29452
rect 21456 29028 21508 29034
rect 21456 28970 21508 28976
rect 21272 28620 21324 28626
rect 21272 28562 21324 28568
rect 20996 27396 21048 27402
rect 20996 27338 21048 27344
rect 21008 27130 21036 27338
rect 20996 27124 21048 27130
rect 20996 27066 21048 27072
rect 20996 26988 21048 26994
rect 20996 26930 21048 26936
rect 20536 26920 20588 26926
rect 20536 26862 20588 26868
rect 21008 26450 21036 26930
rect 20996 26444 21048 26450
rect 20996 26386 21048 26392
rect 21180 26240 21232 26246
rect 21180 26182 21232 26188
rect 20996 25968 21048 25974
rect 20996 25910 21048 25916
rect 20904 25696 20956 25702
rect 20904 25638 20956 25644
rect 19800 25492 19852 25498
rect 19800 25434 19852 25440
rect 20916 25294 20944 25638
rect 20904 25288 20956 25294
rect 20904 25230 20956 25236
rect 20444 24812 20496 24818
rect 20444 24754 20496 24760
rect 20456 24342 20484 24754
rect 20628 24744 20680 24750
rect 20628 24686 20680 24692
rect 20536 24608 20588 24614
rect 20536 24550 20588 24556
rect 20548 24410 20576 24550
rect 20536 24404 20588 24410
rect 20536 24346 20588 24352
rect 20444 24336 20496 24342
rect 20444 24278 20496 24284
rect 19706 23896 19762 23905
rect 19706 23831 19762 23840
rect 19720 23594 19748 23831
rect 20548 23730 20576 24346
rect 20640 23866 20668 24686
rect 20720 24200 20772 24206
rect 20720 24142 20772 24148
rect 20732 23905 20760 24142
rect 20718 23896 20774 23905
rect 20628 23860 20680 23866
rect 20718 23831 20774 23840
rect 20628 23802 20680 23808
rect 20536 23724 20588 23730
rect 20536 23666 20588 23672
rect 19708 23588 19760 23594
rect 19708 23530 19760 23536
rect 20076 23588 20128 23594
rect 20076 23530 20128 23536
rect 19616 23248 19668 23254
rect 19616 23190 19668 23196
rect 19720 23118 19748 23530
rect 19432 23112 19484 23118
rect 19432 23054 19484 23060
rect 19708 23112 19760 23118
rect 19708 23054 19760 23060
rect 18512 22704 18564 22710
rect 18512 22646 18564 22652
rect 18696 22704 18748 22710
rect 18696 22646 18748 22652
rect 18420 22024 18472 22030
rect 18420 21966 18472 21972
rect 18788 22024 18840 22030
rect 18788 21966 18840 21972
rect 18432 21690 18460 21966
rect 18420 21684 18472 21690
rect 18420 21626 18472 21632
rect 18328 20936 18380 20942
rect 18328 20878 18380 20884
rect 17831 20700 18139 20709
rect 17831 20698 17837 20700
rect 17893 20698 17917 20700
rect 17973 20698 17997 20700
rect 18053 20698 18077 20700
rect 18133 20698 18139 20700
rect 17893 20646 17895 20698
rect 18075 20646 18077 20698
rect 17831 20644 17837 20646
rect 17893 20644 17917 20646
rect 17973 20644 17997 20646
rect 18053 20644 18077 20646
rect 18133 20644 18139 20646
rect 17831 20635 18139 20644
rect 16948 20392 17000 20398
rect 16948 20334 17000 20340
rect 17224 20392 17276 20398
rect 17224 20334 17276 20340
rect 17316 20392 17368 20398
rect 17316 20334 17368 20340
rect 17040 19916 17092 19922
rect 17040 19858 17092 19864
rect 16948 18080 17000 18086
rect 16948 18022 17000 18028
rect 16960 17678 16988 18022
rect 16948 17672 17000 17678
rect 16948 17614 17000 17620
rect 17052 16402 17080 19858
rect 17132 19848 17184 19854
rect 17132 19790 17184 19796
rect 17144 19378 17172 19790
rect 17132 19372 17184 19378
rect 17132 19314 17184 19320
rect 17236 16590 17264 20334
rect 17328 19718 17356 20334
rect 17408 20256 17460 20262
rect 17408 20198 17460 20204
rect 17316 19712 17368 19718
rect 17316 19654 17368 19660
rect 17328 18970 17356 19654
rect 17420 18970 17448 20198
rect 18236 19848 18288 19854
rect 18236 19790 18288 19796
rect 17684 19780 17736 19786
rect 17684 19722 17736 19728
rect 17316 18964 17368 18970
rect 17316 18906 17368 18912
rect 17408 18964 17460 18970
rect 17408 18906 17460 18912
rect 17316 18692 17368 18698
rect 17316 18634 17368 18640
rect 17328 18358 17356 18634
rect 17316 18352 17368 18358
rect 17316 18294 17368 18300
rect 17316 18148 17368 18154
rect 17316 18090 17368 18096
rect 17224 16584 17276 16590
rect 17224 16526 17276 16532
rect 17328 16522 17356 18090
rect 17420 18086 17448 18906
rect 17696 18426 17724 19722
rect 17831 19612 18139 19621
rect 17831 19610 17837 19612
rect 17893 19610 17917 19612
rect 17973 19610 17997 19612
rect 18053 19610 18077 19612
rect 18133 19610 18139 19612
rect 17893 19558 17895 19610
rect 18075 19558 18077 19610
rect 17831 19556 17837 19558
rect 17893 19556 17917 19558
rect 17973 19556 17997 19558
rect 18053 19556 18077 19558
rect 18133 19556 18139 19558
rect 17831 19547 18139 19556
rect 17831 18524 18139 18533
rect 17831 18522 17837 18524
rect 17893 18522 17917 18524
rect 17973 18522 17997 18524
rect 18053 18522 18077 18524
rect 18133 18522 18139 18524
rect 17893 18470 17895 18522
rect 18075 18470 18077 18522
rect 17831 18468 17837 18470
rect 17893 18468 17917 18470
rect 17973 18468 17997 18470
rect 18053 18468 18077 18470
rect 18133 18468 18139 18470
rect 17831 18459 18139 18468
rect 17684 18420 17736 18426
rect 17684 18362 17736 18368
rect 17408 18080 17460 18086
rect 17408 18022 17460 18028
rect 17316 16516 17368 16522
rect 17316 16458 17368 16464
rect 17052 16374 17264 16402
rect 17132 15428 17184 15434
rect 17132 15370 17184 15376
rect 16948 15088 17000 15094
rect 16948 15030 17000 15036
rect 16960 12850 16988 15030
rect 16948 12844 17000 12850
rect 16948 12786 17000 12792
rect 16684 12406 16896 12434
rect 16304 11756 16356 11762
rect 16304 11698 16356 11704
rect 16580 11756 16632 11762
rect 16580 11698 16632 11704
rect 16396 9648 16448 9654
rect 16396 9590 16448 9596
rect 16408 9178 16436 9590
rect 16396 9172 16448 9178
rect 16396 9114 16448 9120
rect 16212 8628 16264 8634
rect 16212 8570 16264 8576
rect 16396 8560 16448 8566
rect 16396 8502 16448 8508
rect 16304 8356 16356 8362
rect 16304 8298 16356 8304
rect 16316 6798 16344 8298
rect 16408 6798 16436 8502
rect 16684 7426 16712 12406
rect 16960 12374 16988 12786
rect 16948 12368 17000 12374
rect 16948 12310 17000 12316
rect 16856 11688 16908 11694
rect 16856 11630 16908 11636
rect 16868 11150 16896 11630
rect 16960 11150 16988 12310
rect 17144 12102 17172 15370
rect 17236 14958 17264 16374
rect 17328 15366 17356 16458
rect 17500 16448 17552 16454
rect 17500 16390 17552 16396
rect 17408 16108 17460 16114
rect 17408 16050 17460 16056
rect 17420 15570 17448 16050
rect 17512 15570 17540 16390
rect 17592 16108 17644 16114
rect 17592 16050 17644 16056
rect 17408 15564 17460 15570
rect 17408 15506 17460 15512
rect 17500 15564 17552 15570
rect 17500 15506 17552 15512
rect 17604 15434 17632 16050
rect 17408 15428 17460 15434
rect 17408 15370 17460 15376
rect 17592 15428 17644 15434
rect 17592 15370 17644 15376
rect 17316 15360 17368 15366
rect 17316 15302 17368 15308
rect 17224 14952 17276 14958
rect 17224 14894 17276 14900
rect 17132 12096 17184 12102
rect 17132 12038 17184 12044
rect 16856 11144 16908 11150
rect 16856 11086 16908 11092
rect 16948 11144 17000 11150
rect 16948 11086 17000 11092
rect 16764 11076 16816 11082
rect 16764 11018 16816 11024
rect 16776 9518 16804 11018
rect 17040 9716 17092 9722
rect 17040 9658 17092 9664
rect 16764 9512 16816 9518
rect 16764 9454 16816 9460
rect 16776 7546 16804 9454
rect 16856 8968 16908 8974
rect 16856 8910 16908 8916
rect 16868 8498 16896 8910
rect 16856 8492 16908 8498
rect 16856 8434 16908 8440
rect 16764 7540 16816 7546
rect 16764 7482 16816 7488
rect 16684 7398 16804 7426
rect 16304 6792 16356 6798
rect 16304 6734 16356 6740
rect 16396 6792 16448 6798
rect 16396 6734 16448 6740
rect 15936 4616 15988 4622
rect 15936 4558 15988 4564
rect 15568 4480 15620 4486
rect 15568 4422 15620 4428
rect 15580 4214 15608 4422
rect 15568 4208 15620 4214
rect 15568 4150 15620 4156
rect 15660 3528 15712 3534
rect 15660 3470 15712 3476
rect 15672 3194 15700 3470
rect 15660 3188 15712 3194
rect 15660 3130 15712 3136
rect 15200 3052 15252 3058
rect 15200 2994 15252 3000
rect 15476 2984 15528 2990
rect 15476 2926 15528 2932
rect 15488 2446 15516 2926
rect 15948 2650 15976 4558
rect 16304 4480 16356 4486
rect 16304 4422 16356 4428
rect 16316 3942 16344 4422
rect 16304 3936 16356 3942
rect 16304 3878 16356 3884
rect 16672 3936 16724 3942
rect 16672 3878 16724 3884
rect 15936 2644 15988 2650
rect 15936 2586 15988 2592
rect 16316 2446 16344 3878
rect 16684 3602 16712 3878
rect 16672 3596 16724 3602
rect 16672 3538 16724 3544
rect 16776 3534 16804 7398
rect 16764 3528 16816 3534
rect 16764 3470 16816 3476
rect 16948 3460 17000 3466
rect 16948 3402 17000 3408
rect 16960 3194 16988 3402
rect 17052 3194 17080 9658
rect 17132 9580 17184 9586
rect 17236 9568 17264 14894
rect 17420 14414 17448 15370
rect 17500 15360 17552 15366
rect 17500 15302 17552 15308
rect 17408 14408 17460 14414
rect 17328 14368 17408 14396
rect 17328 13938 17356 14368
rect 17408 14350 17460 14356
rect 17316 13932 17368 13938
rect 17316 13874 17368 13880
rect 17328 13530 17356 13874
rect 17316 13524 17368 13530
rect 17316 13466 17368 13472
rect 17408 12844 17460 12850
rect 17408 12786 17460 12792
rect 17420 12714 17448 12786
rect 17408 12708 17460 12714
rect 17408 12650 17460 12656
rect 17512 12646 17540 15302
rect 17592 14000 17644 14006
rect 17592 13942 17644 13948
rect 17500 12640 17552 12646
rect 17500 12582 17552 12588
rect 17512 12434 17540 12582
rect 17420 12406 17540 12434
rect 17316 12096 17368 12102
rect 17316 12038 17368 12044
rect 17328 11354 17356 12038
rect 17316 11348 17368 11354
rect 17316 11290 17368 11296
rect 17328 9586 17356 11290
rect 17184 9540 17264 9568
rect 17316 9580 17368 9586
rect 17132 9522 17184 9528
rect 17316 9522 17368 9528
rect 17328 9058 17356 9522
rect 17144 9030 17356 9058
rect 17144 8294 17172 9030
rect 17224 8900 17276 8906
rect 17224 8842 17276 8848
rect 17132 8288 17184 8294
rect 17132 8230 17184 8236
rect 17144 7154 17172 8230
rect 17236 7342 17264 8842
rect 17316 7812 17368 7818
rect 17316 7754 17368 7760
rect 17328 7478 17356 7754
rect 17316 7472 17368 7478
rect 17316 7414 17368 7420
rect 17224 7336 17276 7342
rect 17224 7278 17276 7284
rect 17144 7126 17264 7154
rect 17236 6934 17264 7126
rect 17224 6928 17276 6934
rect 17224 6870 17276 6876
rect 17236 6730 17264 6870
rect 17224 6724 17276 6730
rect 17224 6666 17276 6672
rect 17328 4622 17356 7414
rect 17420 7392 17448 12406
rect 17604 12238 17632 13942
rect 17696 13870 17724 18362
rect 17831 17436 18139 17445
rect 17831 17434 17837 17436
rect 17893 17434 17917 17436
rect 17973 17434 17997 17436
rect 18053 17434 18077 17436
rect 18133 17434 18139 17436
rect 17893 17382 17895 17434
rect 18075 17382 18077 17434
rect 17831 17380 17837 17382
rect 17893 17380 17917 17382
rect 17973 17380 17997 17382
rect 18053 17380 18077 17382
rect 18133 17380 18139 17382
rect 17831 17371 18139 17380
rect 17831 16348 18139 16357
rect 17831 16346 17837 16348
rect 17893 16346 17917 16348
rect 17973 16346 17997 16348
rect 18053 16346 18077 16348
rect 18133 16346 18139 16348
rect 17893 16294 17895 16346
rect 18075 16294 18077 16346
rect 17831 16292 17837 16294
rect 17893 16292 17917 16294
rect 17973 16292 17997 16294
rect 18053 16292 18077 16294
rect 18133 16292 18139 16294
rect 17831 16283 18139 16292
rect 18248 15638 18276 19790
rect 18236 15632 18288 15638
rect 18236 15574 18288 15580
rect 18328 15496 18380 15502
rect 18328 15438 18380 15444
rect 17831 15260 18139 15269
rect 17831 15258 17837 15260
rect 17893 15258 17917 15260
rect 17973 15258 17997 15260
rect 18053 15258 18077 15260
rect 18133 15258 18139 15260
rect 17893 15206 17895 15258
rect 18075 15206 18077 15258
rect 17831 15204 17837 15206
rect 17893 15204 17917 15206
rect 17973 15204 17997 15206
rect 18053 15204 18077 15206
rect 18133 15204 18139 15206
rect 17831 15195 18139 15204
rect 17868 15088 17920 15094
rect 17868 15030 17920 15036
rect 17880 14414 17908 15030
rect 18236 15020 18288 15026
rect 18236 14962 18288 14968
rect 17868 14408 17920 14414
rect 17868 14350 17920 14356
rect 17831 14172 18139 14181
rect 17831 14170 17837 14172
rect 17893 14170 17917 14172
rect 17973 14170 17997 14172
rect 18053 14170 18077 14172
rect 18133 14170 18139 14172
rect 17893 14118 17895 14170
rect 18075 14118 18077 14170
rect 17831 14116 17837 14118
rect 17893 14116 17917 14118
rect 17973 14116 17997 14118
rect 18053 14116 18077 14118
rect 18133 14116 18139 14118
rect 17831 14107 18139 14116
rect 17684 13864 17736 13870
rect 17684 13806 17736 13812
rect 17696 12866 17724 13806
rect 18248 13190 18276 14962
rect 18340 13462 18368 15438
rect 18432 15162 18460 21626
rect 18800 21146 18828 21966
rect 18972 21888 19024 21894
rect 18972 21830 19024 21836
rect 18788 21140 18840 21146
rect 18788 21082 18840 21088
rect 18696 20256 18748 20262
rect 18696 20198 18748 20204
rect 18708 19378 18736 20198
rect 18696 19372 18748 19378
rect 18696 19314 18748 19320
rect 18708 18290 18736 19314
rect 18984 18358 19012 21830
rect 19444 21690 19472 23054
rect 20088 22642 20116 23530
rect 20076 22636 20128 22642
rect 20076 22578 20128 22584
rect 19892 22432 19944 22438
rect 19892 22374 19944 22380
rect 19800 21888 19852 21894
rect 19800 21830 19852 21836
rect 19432 21684 19484 21690
rect 19432 21626 19484 21632
rect 19248 21412 19300 21418
rect 19248 21354 19300 21360
rect 19260 20942 19288 21354
rect 19248 20936 19300 20942
rect 19248 20878 19300 20884
rect 18972 18352 19024 18358
rect 18972 18294 19024 18300
rect 18696 18284 18748 18290
rect 18696 18226 18748 18232
rect 18696 17672 18748 17678
rect 18696 17614 18748 17620
rect 18708 17134 18736 17614
rect 18696 17128 18748 17134
rect 18696 17070 18748 17076
rect 18708 16250 18736 17070
rect 18696 16244 18748 16250
rect 18696 16186 18748 16192
rect 19260 15706 19288 20878
rect 19708 20528 19760 20534
rect 19708 20470 19760 20476
rect 19340 19916 19392 19922
rect 19340 19858 19392 19864
rect 19352 18630 19380 19858
rect 19432 19848 19484 19854
rect 19432 19790 19484 19796
rect 19524 19848 19576 19854
rect 19524 19790 19576 19796
rect 19444 19718 19472 19790
rect 19432 19712 19484 19718
rect 19432 19654 19484 19660
rect 19536 19514 19564 19790
rect 19720 19786 19748 20470
rect 19812 19854 19840 21830
rect 19904 21554 19932 22374
rect 20088 22234 20116 22578
rect 20076 22228 20128 22234
rect 20076 22170 20128 22176
rect 19892 21548 19944 21554
rect 19892 21490 19944 21496
rect 20088 21010 20116 22170
rect 20442 22128 20498 22137
rect 20442 22063 20444 22072
rect 20496 22063 20498 22072
rect 20444 22034 20496 22040
rect 20548 21690 20576 23666
rect 20640 22982 20668 23802
rect 20904 23792 20956 23798
rect 20904 23734 20956 23740
rect 20720 23724 20772 23730
rect 20720 23666 20772 23672
rect 20628 22976 20680 22982
rect 20628 22918 20680 22924
rect 20628 22636 20680 22642
rect 20628 22578 20680 22584
rect 20640 22080 20668 22578
rect 20732 22148 20760 23666
rect 20812 23656 20864 23662
rect 20812 23598 20864 23604
rect 20824 23118 20852 23598
rect 20812 23112 20864 23118
rect 20812 23054 20864 23060
rect 20916 22234 20944 23734
rect 21008 23202 21036 25910
rect 21192 25770 21220 26182
rect 21180 25764 21232 25770
rect 21180 25706 21232 25712
rect 21192 25362 21220 25706
rect 21180 25356 21232 25362
rect 21180 25298 21232 25304
rect 21088 25220 21140 25226
rect 21088 25162 21140 25168
rect 21100 24274 21128 25162
rect 21180 24812 21232 24818
rect 21180 24754 21232 24760
rect 21192 24342 21220 24754
rect 21272 24676 21324 24682
rect 21272 24618 21324 24624
rect 21180 24336 21232 24342
rect 21180 24278 21232 24284
rect 21088 24268 21140 24274
rect 21088 24210 21140 24216
rect 21284 24206 21312 24618
rect 21272 24200 21324 24206
rect 21272 24142 21324 24148
rect 21180 24064 21232 24070
rect 21180 24006 21232 24012
rect 21008 23174 21128 23202
rect 20996 23112 21048 23118
rect 20996 23054 21048 23060
rect 20904 22228 20956 22234
rect 20904 22170 20956 22176
rect 20732 22120 20852 22148
rect 20824 22114 20852 22120
rect 20824 22086 20944 22114
rect 20640 22052 20760 22080
rect 20536 21684 20588 21690
rect 20536 21626 20588 21632
rect 20732 21434 20760 22052
rect 20640 21406 20760 21434
rect 20076 21004 20128 21010
rect 20076 20946 20128 20952
rect 20352 20460 20404 20466
rect 20352 20402 20404 20408
rect 20536 20460 20588 20466
rect 20536 20402 20588 20408
rect 19800 19848 19852 19854
rect 19800 19790 19852 19796
rect 19708 19780 19760 19786
rect 19708 19722 19760 19728
rect 19524 19508 19576 19514
rect 19524 19450 19576 19456
rect 19524 18692 19576 18698
rect 19524 18634 19576 18640
rect 19340 18624 19392 18630
rect 19340 18566 19392 18572
rect 19352 16182 19380 18566
rect 19432 17196 19484 17202
rect 19432 17138 19484 17144
rect 19444 16794 19472 17138
rect 19432 16788 19484 16794
rect 19432 16730 19484 16736
rect 19340 16176 19392 16182
rect 19340 16118 19392 16124
rect 19248 15700 19300 15706
rect 19248 15642 19300 15648
rect 18420 15156 18472 15162
rect 18420 15098 18472 15104
rect 18512 15020 18564 15026
rect 18512 14962 18564 14968
rect 18524 14482 18552 14962
rect 18512 14476 18564 14482
rect 18512 14418 18564 14424
rect 19536 14385 19564 18634
rect 19812 18426 19840 19790
rect 20260 19712 20312 19718
rect 20260 19654 20312 19660
rect 19800 18420 19852 18426
rect 19800 18362 19852 18368
rect 19800 16992 19852 16998
rect 19800 16934 19852 16940
rect 19812 16590 19840 16934
rect 19984 16652 20036 16658
rect 19984 16594 20036 16600
rect 19800 16584 19852 16590
rect 19800 16526 19852 16532
rect 19892 16584 19944 16590
rect 19892 16526 19944 16532
rect 19812 16046 19840 16526
rect 19904 16454 19932 16526
rect 19892 16448 19944 16454
rect 19892 16390 19944 16396
rect 19800 16040 19852 16046
rect 19800 15982 19852 15988
rect 19904 15706 19932 16390
rect 19892 15700 19944 15706
rect 19892 15642 19944 15648
rect 19996 15094 20024 16594
rect 20168 16108 20220 16114
rect 20168 16050 20220 16056
rect 20076 15904 20128 15910
rect 20076 15846 20128 15852
rect 19984 15088 20036 15094
rect 19984 15030 20036 15036
rect 19800 15020 19852 15026
rect 19800 14962 19852 14968
rect 19522 14376 19578 14385
rect 19522 14311 19578 14320
rect 19536 14006 19564 14311
rect 19524 14000 19576 14006
rect 19524 13942 19576 13948
rect 19616 14000 19668 14006
rect 19812 13977 19840 14962
rect 19892 14952 19944 14958
rect 19890 14920 19892 14929
rect 19944 14920 19946 14929
rect 19890 14855 19946 14864
rect 19892 14816 19944 14822
rect 19892 14758 19944 14764
rect 19904 14346 19932 14758
rect 19996 14618 20024 15030
rect 19984 14612 20036 14618
rect 19984 14554 20036 14560
rect 19892 14340 19944 14346
rect 19892 14282 19944 14288
rect 19616 13942 19668 13948
rect 19798 13968 19854 13977
rect 19524 13728 19576 13734
rect 19524 13670 19576 13676
rect 18328 13456 18380 13462
rect 18380 13404 18460 13410
rect 18328 13398 18460 13404
rect 18340 13382 18460 13398
rect 18328 13320 18380 13326
rect 18328 13262 18380 13268
rect 18236 13184 18288 13190
rect 18236 13126 18288 13132
rect 17831 13084 18139 13093
rect 17831 13082 17837 13084
rect 17893 13082 17917 13084
rect 17973 13082 17997 13084
rect 18053 13082 18077 13084
rect 18133 13082 18139 13084
rect 17893 13030 17895 13082
rect 18075 13030 18077 13082
rect 17831 13028 17837 13030
rect 17893 13028 17917 13030
rect 17973 13028 17997 13030
rect 18053 13028 18077 13030
rect 18133 13028 18139 13030
rect 17831 13019 18139 13028
rect 17696 12838 17816 12866
rect 17788 12434 17816 12838
rect 17696 12406 17816 12434
rect 17592 12232 17644 12238
rect 17592 12174 17644 12180
rect 17604 11150 17632 12174
rect 17696 11218 17724 12406
rect 17831 11996 18139 12005
rect 17831 11994 17837 11996
rect 17893 11994 17917 11996
rect 17973 11994 17997 11996
rect 18053 11994 18077 11996
rect 18133 11994 18139 11996
rect 17893 11942 17895 11994
rect 18075 11942 18077 11994
rect 17831 11940 17837 11942
rect 17893 11940 17917 11942
rect 17973 11940 17997 11942
rect 18053 11940 18077 11942
rect 18133 11940 18139 11942
rect 17831 11931 18139 11940
rect 17684 11212 17736 11218
rect 17684 11154 17736 11160
rect 17592 11144 17644 11150
rect 17592 11086 17644 11092
rect 17831 10908 18139 10917
rect 17831 10906 17837 10908
rect 17893 10906 17917 10908
rect 17973 10906 17997 10908
rect 18053 10906 18077 10908
rect 18133 10906 18139 10908
rect 17893 10854 17895 10906
rect 18075 10854 18077 10906
rect 17831 10852 17837 10854
rect 17893 10852 17917 10854
rect 17973 10852 17997 10854
rect 18053 10852 18077 10854
rect 18133 10852 18139 10854
rect 17831 10843 18139 10852
rect 18248 10742 18276 13126
rect 18340 12850 18368 13262
rect 18328 12844 18380 12850
rect 18328 12786 18380 12792
rect 18340 12306 18368 12786
rect 18328 12300 18380 12306
rect 18328 12242 18380 12248
rect 18432 11830 18460 13382
rect 19338 12472 19394 12481
rect 19338 12407 19394 12416
rect 19156 12164 19208 12170
rect 19156 12106 19208 12112
rect 18420 11824 18472 11830
rect 18420 11766 18472 11772
rect 18236 10736 18288 10742
rect 18236 10678 18288 10684
rect 17831 9820 18139 9829
rect 17831 9818 17837 9820
rect 17893 9818 17917 9820
rect 17973 9818 17997 9820
rect 18053 9818 18077 9820
rect 18133 9818 18139 9820
rect 17893 9766 17895 9818
rect 18075 9766 18077 9818
rect 17831 9764 17837 9766
rect 17893 9764 17917 9766
rect 17973 9764 17997 9766
rect 18053 9764 18077 9766
rect 18133 9764 18139 9766
rect 17831 9755 18139 9764
rect 17592 9580 17644 9586
rect 17592 9522 17644 9528
rect 18420 9580 18472 9586
rect 19064 9580 19116 9586
rect 18472 9540 18920 9568
rect 18420 9522 18472 9528
rect 17604 8430 17632 9522
rect 18892 9450 18920 9540
rect 19064 9522 19116 9528
rect 18788 9444 18840 9450
rect 18788 9386 18840 9392
rect 18880 9444 18932 9450
rect 18880 9386 18932 9392
rect 18800 9178 18828 9386
rect 18788 9172 18840 9178
rect 18788 9114 18840 9120
rect 18788 8832 18840 8838
rect 18788 8774 18840 8780
rect 17831 8732 18139 8741
rect 17831 8730 17837 8732
rect 17893 8730 17917 8732
rect 17973 8730 17997 8732
rect 18053 8730 18077 8732
rect 18133 8730 18139 8732
rect 17893 8678 17895 8730
rect 18075 8678 18077 8730
rect 17831 8676 17837 8678
rect 17893 8676 17917 8678
rect 17973 8676 17997 8678
rect 18053 8676 18077 8678
rect 18133 8676 18139 8678
rect 17831 8667 18139 8676
rect 17684 8628 17736 8634
rect 17684 8570 17736 8576
rect 17592 8424 17644 8430
rect 17592 8366 17644 8372
rect 17500 7744 17552 7750
rect 17500 7686 17552 7692
rect 17512 7546 17540 7686
rect 17500 7540 17552 7546
rect 17500 7482 17552 7488
rect 17500 7404 17552 7410
rect 17420 7364 17500 7392
rect 17500 7346 17552 7352
rect 17604 6882 17632 8366
rect 17512 6854 17632 6882
rect 17512 6730 17540 6854
rect 17500 6724 17552 6730
rect 17500 6666 17552 6672
rect 17696 6662 17724 8570
rect 18800 8498 18828 8774
rect 18892 8566 18920 9386
rect 19076 8634 19104 9522
rect 19168 9518 19196 12106
rect 19352 10674 19380 12407
rect 19340 10668 19392 10674
rect 19340 10610 19392 10616
rect 19156 9512 19208 9518
rect 19156 9454 19208 9460
rect 19168 8634 19196 9454
rect 19536 9058 19564 13670
rect 19628 12782 19656 13942
rect 19798 13903 19854 13912
rect 19800 13728 19852 13734
rect 19800 13670 19852 13676
rect 19812 13326 19840 13670
rect 19800 13320 19852 13326
rect 19800 13262 19852 13268
rect 19616 12776 19668 12782
rect 19616 12718 19668 12724
rect 19708 11756 19760 11762
rect 19708 11698 19760 11704
rect 19720 10810 19748 11698
rect 20088 11150 20116 15846
rect 20180 15434 20208 16050
rect 20168 15428 20220 15434
rect 20168 15370 20220 15376
rect 19984 11144 20036 11150
rect 19984 11086 20036 11092
rect 20076 11144 20128 11150
rect 20076 11086 20128 11092
rect 19892 11076 19944 11082
rect 19892 11018 19944 11024
rect 19708 10804 19760 10810
rect 19708 10746 19760 10752
rect 19904 10742 19932 11018
rect 19892 10736 19944 10742
rect 19892 10678 19944 10684
rect 19904 9586 19932 10678
rect 19708 9580 19760 9586
rect 19708 9522 19760 9528
rect 19892 9580 19944 9586
rect 19892 9522 19944 9528
rect 19352 9030 19564 9058
rect 19064 8628 19116 8634
rect 19064 8570 19116 8576
rect 19156 8628 19208 8634
rect 19156 8570 19208 8576
rect 18880 8560 18932 8566
rect 18880 8502 18932 8508
rect 18696 8492 18748 8498
rect 18696 8434 18748 8440
rect 18788 8492 18840 8498
rect 18788 8434 18840 8440
rect 18708 8090 18736 8434
rect 18696 8084 18748 8090
rect 18696 8026 18748 8032
rect 17831 7644 18139 7653
rect 17831 7642 17837 7644
rect 17893 7642 17917 7644
rect 17973 7642 17997 7644
rect 18053 7642 18077 7644
rect 18133 7642 18139 7644
rect 17893 7590 17895 7642
rect 18075 7590 18077 7642
rect 17831 7588 17837 7590
rect 17893 7588 17917 7590
rect 17973 7588 17997 7590
rect 18053 7588 18077 7590
rect 18133 7588 18139 7590
rect 17831 7579 18139 7588
rect 17868 7404 17920 7410
rect 17868 7346 17920 7352
rect 17880 6934 17908 7346
rect 17868 6928 17920 6934
rect 17868 6870 17920 6876
rect 17880 6798 17908 6870
rect 17868 6792 17920 6798
rect 17868 6734 17920 6740
rect 17684 6656 17736 6662
rect 17684 6598 17736 6604
rect 17831 6556 18139 6565
rect 17831 6554 17837 6556
rect 17893 6554 17917 6556
rect 17973 6554 17997 6556
rect 18053 6554 18077 6556
rect 18133 6554 18139 6556
rect 17893 6502 17895 6554
rect 18075 6502 18077 6554
rect 17831 6500 17837 6502
rect 17893 6500 17917 6502
rect 17973 6500 17997 6502
rect 18053 6500 18077 6502
rect 18133 6500 18139 6502
rect 17831 6491 18139 6500
rect 18420 6180 18472 6186
rect 18420 6122 18472 6128
rect 17831 5468 18139 5477
rect 17831 5466 17837 5468
rect 17893 5466 17917 5468
rect 17973 5466 17997 5468
rect 18053 5466 18077 5468
rect 18133 5466 18139 5468
rect 17893 5414 17895 5466
rect 18075 5414 18077 5466
rect 17831 5412 17837 5414
rect 17893 5412 17917 5414
rect 17973 5412 17997 5414
rect 18053 5412 18077 5414
rect 18133 5412 18139 5414
rect 17831 5403 18139 5412
rect 18432 4622 18460 6122
rect 18708 5302 18736 8026
rect 18800 7546 18828 8434
rect 19168 7750 19196 8570
rect 19352 8294 19380 9030
rect 19524 8968 19576 8974
rect 19524 8910 19576 8916
rect 19340 8288 19392 8294
rect 19340 8230 19392 8236
rect 19352 8022 19380 8230
rect 19340 8016 19392 8022
rect 19340 7958 19392 7964
rect 19156 7744 19208 7750
rect 19156 7686 19208 7692
rect 19536 7546 19564 8910
rect 19720 8906 19748 9522
rect 19996 9450 20024 11086
rect 19984 9444 20036 9450
rect 19984 9386 20036 9392
rect 20168 9376 20220 9382
rect 20168 9318 20220 9324
rect 20180 8974 20208 9318
rect 20272 9178 20300 19654
rect 20364 18630 20392 20402
rect 20548 19922 20576 20402
rect 20536 19916 20588 19922
rect 20536 19858 20588 19864
rect 20352 18624 20404 18630
rect 20352 18566 20404 18572
rect 20364 16182 20392 18566
rect 20536 18080 20588 18086
rect 20536 18022 20588 18028
rect 20548 17678 20576 18022
rect 20536 17672 20588 17678
rect 20536 17614 20588 17620
rect 20352 16176 20404 16182
rect 20352 16118 20404 16124
rect 20444 16108 20496 16114
rect 20444 16050 20496 16056
rect 20456 12986 20484 16050
rect 20640 15978 20668 21406
rect 20720 20528 20772 20534
rect 20720 20470 20772 20476
rect 20732 19514 20760 20470
rect 20812 20324 20864 20330
rect 20812 20266 20864 20272
rect 20824 19786 20852 20266
rect 20812 19780 20864 19786
rect 20812 19722 20864 19728
rect 20720 19508 20772 19514
rect 20720 19450 20772 19456
rect 20720 17196 20772 17202
rect 20720 17138 20772 17144
rect 20732 16522 20760 17138
rect 20720 16516 20772 16522
rect 20720 16458 20772 16464
rect 20628 15972 20680 15978
rect 20628 15914 20680 15920
rect 20824 15502 20852 19722
rect 20916 18698 20944 22086
rect 21008 20602 21036 23054
rect 21100 22094 21128 23174
rect 21192 22642 21220 24006
rect 21180 22636 21232 22642
rect 21180 22578 21232 22584
rect 21100 22066 21220 22094
rect 21088 21956 21140 21962
rect 21088 21898 21140 21904
rect 20996 20596 21048 20602
rect 20996 20538 21048 20544
rect 20996 20460 21048 20466
rect 20996 20402 21048 20408
rect 21008 19990 21036 20402
rect 20996 19984 21048 19990
rect 20996 19926 21048 19932
rect 20996 19372 21048 19378
rect 21100 19360 21128 21898
rect 21192 21894 21220 22066
rect 21180 21888 21232 21894
rect 21180 21830 21232 21836
rect 21192 20874 21220 21830
rect 21284 21146 21312 24142
rect 21272 21140 21324 21146
rect 21272 21082 21324 21088
rect 21468 21010 21496 28970
rect 21560 28490 21588 29650
rect 21640 29640 21692 29646
rect 21640 29582 21692 29588
rect 21652 29238 21680 29582
rect 21744 29306 21772 31146
rect 22052 31036 22360 31045
rect 22052 31034 22058 31036
rect 22114 31034 22138 31036
rect 22194 31034 22218 31036
rect 22274 31034 22298 31036
rect 22354 31034 22360 31036
rect 22114 30982 22116 31034
rect 22296 30982 22298 31034
rect 22052 30980 22058 30982
rect 22114 30980 22138 30982
rect 22194 30980 22218 30982
rect 22274 30980 22298 30982
rect 22354 30980 22360 30982
rect 22052 30971 22360 30980
rect 23032 30938 23060 31282
rect 23020 30932 23072 30938
rect 23020 30874 23072 30880
rect 23308 30734 23336 31962
rect 23400 31754 23428 32302
rect 23756 31816 23808 31822
rect 23756 31758 23808 31764
rect 23388 31748 23440 31754
rect 23388 31690 23440 31696
rect 23400 30802 23428 31690
rect 23572 31680 23624 31686
rect 23572 31622 23624 31628
rect 23584 31346 23612 31622
rect 23572 31340 23624 31346
rect 23572 31282 23624 31288
rect 23572 31204 23624 31210
rect 23572 31146 23624 31152
rect 23388 30796 23440 30802
rect 23388 30738 23440 30744
rect 23296 30728 23348 30734
rect 23296 30670 23348 30676
rect 22052 29948 22360 29957
rect 22052 29946 22058 29948
rect 22114 29946 22138 29948
rect 22194 29946 22218 29948
rect 22274 29946 22298 29948
rect 22354 29946 22360 29948
rect 22114 29894 22116 29946
rect 22296 29894 22298 29946
rect 22052 29892 22058 29894
rect 22114 29892 22138 29894
rect 22194 29892 22218 29894
rect 22274 29892 22298 29894
rect 22354 29892 22360 29894
rect 22052 29883 22360 29892
rect 23308 29782 23336 30670
rect 23296 29776 23348 29782
rect 23296 29718 23348 29724
rect 21732 29300 21784 29306
rect 21732 29242 21784 29248
rect 21640 29232 21692 29238
rect 21640 29174 21692 29180
rect 23480 29232 23532 29238
rect 23480 29174 23532 29180
rect 22284 29164 22336 29170
rect 22284 29106 22336 29112
rect 22744 29164 22796 29170
rect 22744 29106 22796 29112
rect 21640 29096 21692 29102
rect 21640 29038 21692 29044
rect 22296 29050 22324 29106
rect 21652 28694 21680 29038
rect 22296 29022 22416 29050
rect 22052 28860 22360 28869
rect 22052 28858 22058 28860
rect 22114 28858 22138 28860
rect 22194 28858 22218 28860
rect 22274 28858 22298 28860
rect 22354 28858 22360 28860
rect 22114 28806 22116 28858
rect 22296 28806 22298 28858
rect 22052 28804 22058 28806
rect 22114 28804 22138 28806
rect 22194 28804 22218 28806
rect 22274 28804 22298 28806
rect 22354 28804 22360 28806
rect 22052 28795 22360 28804
rect 21640 28688 21692 28694
rect 21640 28630 21692 28636
rect 21548 28484 21600 28490
rect 21548 28426 21600 28432
rect 22388 28218 22416 29022
rect 22756 28422 22784 29106
rect 23296 29028 23348 29034
rect 23296 28970 23348 28976
rect 23308 28558 23336 28970
rect 23492 28558 23520 29174
rect 23584 29170 23612 31146
rect 23768 30666 23796 31758
rect 24596 31686 24624 32370
rect 24768 32360 24820 32366
rect 24768 32302 24820 32308
rect 24780 31754 24808 32302
rect 25044 32224 25096 32230
rect 25044 32166 25096 32172
rect 25056 31890 25084 32166
rect 25044 31884 25096 31890
rect 25044 31826 25096 31832
rect 25136 31884 25188 31890
rect 25136 31826 25188 31832
rect 24688 31726 24808 31754
rect 24584 31680 24636 31686
rect 24584 31622 24636 31628
rect 24492 31340 24544 31346
rect 24688 31328 24716 31726
rect 24768 31680 24820 31686
rect 24768 31622 24820 31628
rect 24544 31300 24716 31328
rect 24492 31282 24544 31288
rect 23756 30660 23808 30666
rect 23756 30602 23808 30608
rect 24596 29578 24624 31300
rect 24676 30252 24728 30258
rect 24676 30194 24728 30200
rect 24584 29572 24636 29578
rect 24584 29514 24636 29520
rect 23572 29164 23624 29170
rect 23572 29106 23624 29112
rect 22836 28552 22888 28558
rect 22836 28494 22888 28500
rect 23296 28552 23348 28558
rect 23296 28494 23348 28500
rect 23480 28552 23532 28558
rect 23480 28494 23532 28500
rect 22744 28416 22796 28422
rect 22744 28358 22796 28364
rect 22376 28212 22428 28218
rect 22376 28154 22428 28160
rect 22052 27772 22360 27781
rect 22052 27770 22058 27772
rect 22114 27770 22138 27772
rect 22194 27770 22218 27772
rect 22274 27770 22298 27772
rect 22354 27770 22360 27772
rect 22114 27718 22116 27770
rect 22296 27718 22298 27770
rect 22052 27716 22058 27718
rect 22114 27716 22138 27718
rect 22194 27716 22218 27718
rect 22274 27716 22298 27718
rect 22354 27716 22360 27718
rect 22052 27707 22360 27716
rect 22652 26920 22704 26926
rect 22652 26862 22704 26868
rect 21548 26852 21600 26858
rect 21548 26794 21600 26800
rect 21560 26382 21588 26794
rect 22376 26784 22428 26790
rect 22376 26726 22428 26732
rect 22052 26684 22360 26693
rect 22052 26682 22058 26684
rect 22114 26682 22138 26684
rect 22194 26682 22218 26684
rect 22274 26682 22298 26684
rect 22354 26682 22360 26684
rect 22114 26630 22116 26682
rect 22296 26630 22298 26682
rect 22052 26628 22058 26630
rect 22114 26628 22138 26630
rect 22194 26628 22218 26630
rect 22274 26628 22298 26630
rect 22354 26628 22360 26630
rect 22052 26619 22360 26628
rect 21640 26444 21692 26450
rect 21640 26386 21692 26392
rect 21548 26376 21600 26382
rect 21548 26318 21600 26324
rect 21560 25906 21588 26318
rect 21548 25900 21600 25906
rect 21548 25842 21600 25848
rect 21560 21962 21588 25842
rect 21548 21956 21600 21962
rect 21548 21898 21600 21904
rect 21456 21004 21508 21010
rect 21456 20946 21508 20952
rect 21180 20868 21232 20874
rect 21180 20810 21232 20816
rect 21652 20602 21680 26386
rect 22388 25906 22416 26726
rect 22664 26314 22692 26862
rect 22756 26450 22784 28358
rect 22848 28150 22876 28494
rect 22836 28144 22888 28150
rect 22836 28086 22888 28092
rect 23492 27946 23520 28494
rect 23480 27940 23532 27946
rect 23480 27882 23532 27888
rect 23584 27470 23612 29106
rect 24596 27606 24624 29514
rect 24688 29238 24716 30194
rect 24780 29646 24808 31622
rect 25148 31482 25176 31826
rect 26608 31816 26660 31822
rect 26608 31758 26660 31764
rect 27344 31816 27396 31822
rect 27344 31758 27396 31764
rect 26272 31580 26580 31589
rect 26272 31578 26278 31580
rect 26334 31578 26358 31580
rect 26414 31578 26438 31580
rect 26494 31578 26518 31580
rect 26574 31578 26580 31580
rect 26334 31526 26336 31578
rect 26516 31526 26518 31578
rect 26272 31524 26278 31526
rect 26334 31524 26358 31526
rect 26414 31524 26438 31526
rect 26494 31524 26518 31526
rect 26574 31524 26580 31526
rect 26272 31515 26580 31524
rect 26620 31482 26648 31758
rect 25136 31476 25188 31482
rect 25136 31418 25188 31424
rect 26608 31476 26660 31482
rect 26608 31418 26660 31424
rect 27356 31346 27384 31758
rect 27724 31754 27752 32370
rect 27712 31748 27764 31754
rect 27712 31690 27764 31696
rect 28644 31482 28672 32370
rect 30196 32224 30248 32230
rect 30196 32166 30248 32172
rect 33232 32224 33284 32230
rect 33232 32166 33284 32172
rect 28632 31476 28684 31482
rect 28632 31418 28684 31424
rect 25044 31340 25096 31346
rect 25044 31282 25096 31288
rect 25320 31340 25372 31346
rect 25320 31282 25372 31288
rect 26056 31340 26108 31346
rect 26056 31282 26108 31288
rect 27344 31340 27396 31346
rect 27344 31282 27396 31288
rect 27528 31340 27580 31346
rect 27528 31282 27580 31288
rect 27712 31340 27764 31346
rect 27712 31282 27764 31288
rect 28540 31340 28592 31346
rect 28540 31282 28592 31288
rect 24952 30864 25004 30870
rect 24950 30832 24952 30841
rect 25004 30832 25006 30841
rect 24950 30767 25006 30776
rect 25056 30666 25084 31282
rect 25332 30734 25360 31282
rect 25780 31272 25832 31278
rect 25780 31214 25832 31220
rect 25596 31136 25648 31142
rect 25596 31078 25648 31084
rect 25608 30734 25636 31078
rect 25792 30734 25820 31214
rect 26068 30734 26096 31282
rect 25320 30728 25372 30734
rect 25320 30670 25372 30676
rect 25596 30728 25648 30734
rect 25596 30670 25648 30676
rect 25780 30728 25832 30734
rect 25780 30670 25832 30676
rect 26056 30728 26108 30734
rect 26056 30670 26108 30676
rect 25044 30660 25096 30666
rect 25044 30602 25096 30608
rect 25056 30394 25084 30602
rect 25044 30388 25096 30394
rect 25044 30330 25096 30336
rect 24768 29640 24820 29646
rect 24768 29582 24820 29588
rect 24676 29232 24728 29238
rect 24676 29174 24728 29180
rect 24676 28076 24728 28082
rect 24676 28018 24728 28024
rect 24584 27600 24636 27606
rect 24584 27542 24636 27548
rect 23572 27464 23624 27470
rect 23572 27406 23624 27412
rect 22744 26444 22796 26450
rect 22744 26386 22796 26392
rect 22560 26308 22612 26314
rect 22560 26250 22612 26256
rect 22652 26308 22704 26314
rect 22652 26250 22704 26256
rect 22376 25900 22428 25906
rect 22376 25842 22428 25848
rect 22052 25596 22360 25605
rect 22052 25594 22058 25596
rect 22114 25594 22138 25596
rect 22194 25594 22218 25596
rect 22274 25594 22298 25596
rect 22354 25594 22360 25596
rect 22114 25542 22116 25594
rect 22296 25542 22298 25594
rect 22052 25540 22058 25542
rect 22114 25540 22138 25542
rect 22194 25540 22218 25542
rect 22274 25540 22298 25542
rect 22354 25540 22360 25542
rect 22052 25531 22360 25540
rect 22572 25158 22600 26250
rect 22664 26042 22692 26250
rect 23584 26042 23612 27406
rect 24584 26784 24636 26790
rect 24584 26726 24636 26732
rect 22652 26036 22704 26042
rect 22652 25978 22704 25984
rect 23572 26036 23624 26042
rect 23572 25978 23624 25984
rect 23664 25832 23716 25838
rect 23664 25774 23716 25780
rect 23480 25288 23532 25294
rect 23480 25230 23532 25236
rect 22560 25152 22612 25158
rect 22560 25094 22612 25100
rect 22052 24508 22360 24517
rect 22052 24506 22058 24508
rect 22114 24506 22138 24508
rect 22194 24506 22218 24508
rect 22274 24506 22298 24508
rect 22354 24506 22360 24508
rect 22114 24454 22116 24506
rect 22296 24454 22298 24506
rect 22052 24452 22058 24454
rect 22114 24452 22138 24454
rect 22194 24452 22218 24454
rect 22274 24452 22298 24454
rect 22354 24452 22360 24454
rect 22052 24443 22360 24452
rect 21732 24064 21784 24070
rect 21732 24006 21784 24012
rect 21640 20596 21692 20602
rect 21640 20538 21692 20544
rect 21048 19332 21128 19360
rect 20996 19314 21048 19320
rect 20904 18692 20956 18698
rect 20904 18634 20956 18640
rect 21008 18578 21036 19314
rect 21744 18766 21772 24006
rect 21916 23792 21968 23798
rect 21916 23734 21968 23740
rect 21928 23322 21956 23734
rect 22052 23420 22360 23429
rect 22052 23418 22058 23420
rect 22114 23418 22138 23420
rect 22194 23418 22218 23420
rect 22274 23418 22298 23420
rect 22354 23418 22360 23420
rect 22114 23366 22116 23418
rect 22296 23366 22298 23418
rect 22052 23364 22058 23366
rect 22114 23364 22138 23366
rect 22194 23364 22218 23366
rect 22274 23364 22298 23366
rect 22354 23364 22360 23366
rect 22052 23355 22360 23364
rect 21916 23316 21968 23322
rect 21916 23258 21968 23264
rect 22190 23216 22246 23225
rect 22190 23151 22246 23160
rect 22204 22642 22232 23151
rect 21824 22636 21876 22642
rect 21824 22578 21876 22584
rect 22192 22636 22244 22642
rect 22192 22578 22244 22584
rect 21732 18760 21784 18766
rect 21732 18702 21784 18708
rect 20916 18550 21036 18578
rect 20916 18290 20944 18550
rect 21088 18420 21140 18426
rect 21088 18362 21140 18368
rect 20904 18284 20956 18290
rect 20904 18226 20956 18232
rect 20916 16454 20944 18226
rect 21100 17542 21128 18362
rect 21088 17536 21140 17542
rect 21088 17478 21140 17484
rect 20996 16516 21048 16522
rect 20996 16458 21048 16464
rect 20904 16448 20956 16454
rect 20904 16390 20956 16396
rect 20812 15496 20864 15502
rect 20812 15438 20864 15444
rect 20536 15428 20588 15434
rect 20536 15370 20588 15376
rect 20548 13938 20576 15370
rect 21008 15366 21036 16458
rect 21100 16182 21128 17478
rect 21744 17270 21772 18702
rect 21732 17264 21784 17270
rect 21732 17206 21784 17212
rect 21088 16176 21140 16182
rect 21088 16118 21140 16124
rect 21640 16108 21692 16114
rect 21640 16050 21692 16056
rect 21180 15564 21232 15570
rect 21180 15506 21232 15512
rect 20996 15360 21048 15366
rect 20996 15302 21048 15308
rect 20720 14952 20772 14958
rect 20720 14894 20772 14900
rect 20628 14340 20680 14346
rect 20628 14282 20680 14288
rect 20536 13932 20588 13938
rect 20536 13874 20588 13880
rect 20444 12980 20496 12986
rect 20444 12922 20496 12928
rect 20536 12708 20588 12714
rect 20536 12650 20588 12656
rect 20548 11898 20576 12650
rect 20536 11892 20588 11898
rect 20536 11834 20588 11840
rect 20444 11756 20496 11762
rect 20444 11698 20496 11704
rect 20456 10810 20484 11698
rect 20548 11150 20576 11834
rect 20536 11144 20588 11150
rect 20536 11086 20588 11092
rect 20444 10804 20496 10810
rect 20444 10746 20496 10752
rect 20640 9586 20668 14282
rect 20732 13802 20760 14894
rect 20812 14272 20864 14278
rect 20812 14214 20864 14220
rect 20720 13796 20772 13802
rect 20720 13738 20772 13744
rect 20720 12844 20772 12850
rect 20720 12786 20772 12792
rect 20732 11898 20760 12786
rect 20824 12170 20852 14214
rect 20904 12844 20956 12850
rect 20904 12786 20956 12792
rect 20996 12844 21048 12850
rect 20996 12786 21048 12792
rect 20916 12374 20944 12786
rect 20904 12368 20956 12374
rect 20904 12310 20956 12316
rect 20812 12164 20864 12170
rect 20812 12106 20864 12112
rect 20720 11892 20772 11898
rect 20720 11834 20772 11840
rect 20732 10810 20760 11834
rect 20720 10804 20772 10810
rect 20720 10746 20772 10752
rect 20628 9580 20680 9586
rect 20628 9522 20680 9528
rect 20720 9444 20772 9450
rect 20720 9386 20772 9392
rect 20260 9172 20312 9178
rect 20260 9114 20312 9120
rect 19892 8968 19944 8974
rect 19892 8910 19944 8916
rect 20168 8968 20220 8974
rect 20168 8910 20220 8916
rect 19708 8900 19760 8906
rect 19708 8842 19760 8848
rect 19904 8430 19932 8910
rect 19892 8424 19944 8430
rect 19892 8366 19944 8372
rect 20536 8424 20588 8430
rect 20536 8366 20588 8372
rect 18788 7540 18840 7546
rect 18788 7482 18840 7488
rect 19524 7540 19576 7546
rect 19524 7482 19576 7488
rect 19340 7404 19392 7410
rect 19340 7346 19392 7352
rect 19352 6866 19380 7346
rect 20444 7200 20496 7206
rect 20444 7142 20496 7148
rect 19340 6860 19392 6866
rect 19340 6802 19392 6808
rect 20456 6798 20484 7142
rect 20548 6866 20576 8366
rect 20628 7948 20680 7954
rect 20628 7890 20680 7896
rect 20640 7410 20668 7890
rect 20732 7546 20760 9386
rect 20824 7818 20852 12106
rect 21008 11014 21036 12786
rect 21088 11348 21140 11354
rect 21088 11290 21140 11296
rect 21100 11150 21128 11290
rect 21192 11257 21220 15506
rect 21652 14414 21680 16050
rect 21836 15162 21864 22578
rect 22052 22332 22360 22341
rect 22052 22330 22058 22332
rect 22114 22330 22138 22332
rect 22194 22330 22218 22332
rect 22274 22330 22298 22332
rect 22354 22330 22360 22332
rect 22114 22278 22116 22330
rect 22296 22278 22298 22330
rect 22052 22276 22058 22278
rect 22114 22276 22138 22278
rect 22194 22276 22218 22278
rect 22274 22276 22298 22278
rect 22354 22276 22360 22278
rect 22052 22267 22360 22276
rect 22284 21888 22336 21894
rect 22284 21830 22336 21836
rect 22296 21554 22324 21830
rect 22284 21548 22336 21554
rect 22284 21490 22336 21496
rect 22376 21480 22428 21486
rect 22376 21422 22428 21428
rect 22052 21244 22360 21253
rect 22052 21242 22058 21244
rect 22114 21242 22138 21244
rect 22194 21242 22218 21244
rect 22274 21242 22298 21244
rect 22354 21242 22360 21244
rect 22114 21190 22116 21242
rect 22296 21190 22298 21242
rect 22052 21188 22058 21190
rect 22114 21188 22138 21190
rect 22194 21188 22218 21190
rect 22274 21188 22298 21190
rect 22354 21188 22360 21190
rect 22052 21179 22360 21188
rect 22284 20596 22336 20602
rect 22284 20538 22336 20544
rect 22296 20244 22324 20538
rect 22388 20534 22416 21422
rect 22572 20942 22600 25094
rect 23388 24948 23440 24954
rect 23388 24890 23440 24896
rect 23400 24206 23428 24890
rect 23492 24342 23520 25230
rect 23676 24886 23704 25774
rect 24596 25294 24624 26726
rect 24688 25906 24716 28018
rect 24780 26994 24808 29582
rect 25056 28914 25084 30330
rect 25332 30258 25360 30670
rect 25608 30258 25636 30670
rect 25792 30258 25820 30670
rect 26068 30258 26096 30670
rect 26272 30492 26580 30501
rect 26272 30490 26278 30492
rect 26334 30490 26358 30492
rect 26414 30490 26438 30492
rect 26494 30490 26518 30492
rect 26574 30490 26580 30492
rect 26334 30438 26336 30490
rect 26516 30438 26518 30490
rect 26272 30436 26278 30438
rect 26334 30436 26358 30438
rect 26414 30436 26438 30438
rect 26494 30436 26518 30438
rect 26574 30436 26580 30438
rect 26272 30427 26580 30436
rect 27356 30394 27384 31282
rect 27160 30388 27212 30394
rect 27160 30330 27212 30336
rect 27344 30388 27396 30394
rect 27344 30330 27396 30336
rect 25320 30252 25372 30258
rect 25320 30194 25372 30200
rect 25596 30252 25648 30258
rect 25596 30194 25648 30200
rect 25780 30252 25832 30258
rect 25780 30194 25832 30200
rect 26056 30252 26108 30258
rect 26056 30194 26108 30200
rect 25332 29306 25360 30194
rect 25412 30184 25464 30190
rect 25412 30126 25464 30132
rect 25424 29578 25452 30126
rect 26068 29850 26096 30194
rect 26056 29844 26108 29850
rect 26056 29786 26108 29792
rect 25412 29572 25464 29578
rect 25412 29514 25464 29520
rect 26056 29572 26108 29578
rect 26056 29514 26108 29520
rect 25320 29300 25372 29306
rect 25320 29242 25372 29248
rect 25780 29164 25832 29170
rect 25780 29106 25832 29112
rect 25056 28886 25268 28914
rect 25240 28082 25268 28886
rect 25044 28076 25096 28082
rect 25044 28018 25096 28024
rect 25228 28076 25280 28082
rect 25228 28018 25280 28024
rect 25056 27402 25084 28018
rect 25136 28008 25188 28014
rect 25136 27950 25188 27956
rect 25044 27396 25096 27402
rect 25044 27338 25096 27344
rect 24768 26988 24820 26994
rect 24768 26930 24820 26936
rect 25056 26382 25084 27338
rect 25148 26994 25176 27950
rect 25136 26988 25188 26994
rect 25136 26930 25188 26936
rect 25148 26586 25176 26930
rect 25136 26580 25188 26586
rect 25136 26522 25188 26528
rect 25240 26466 25268 28018
rect 25792 28014 25820 29106
rect 25780 28008 25832 28014
rect 25780 27950 25832 27956
rect 25688 27464 25740 27470
rect 25688 27406 25740 27412
rect 25596 27396 25648 27402
rect 25596 27338 25648 27344
rect 25608 26994 25636 27338
rect 25596 26988 25648 26994
rect 25596 26930 25648 26936
rect 25148 26438 25268 26466
rect 25044 26376 25096 26382
rect 25044 26318 25096 26324
rect 25148 26314 25176 26438
rect 25320 26376 25372 26382
rect 25320 26318 25372 26324
rect 25504 26376 25556 26382
rect 25504 26318 25556 26324
rect 25136 26308 25188 26314
rect 25136 26250 25188 26256
rect 24676 25900 24728 25906
rect 24676 25842 24728 25848
rect 24688 25362 24716 25842
rect 24860 25764 24912 25770
rect 24860 25706 24912 25712
rect 24676 25356 24728 25362
rect 24676 25298 24728 25304
rect 24584 25288 24636 25294
rect 24584 25230 24636 25236
rect 23664 24880 23716 24886
rect 23664 24822 23716 24828
rect 23480 24336 23532 24342
rect 23480 24278 23532 24284
rect 23388 24200 23440 24206
rect 23388 24142 23440 24148
rect 23480 24064 23532 24070
rect 23480 24006 23532 24012
rect 23492 23866 23520 24006
rect 23480 23860 23532 23866
rect 23480 23802 23532 23808
rect 23676 23730 23704 24822
rect 23756 24200 23808 24206
rect 23756 24142 23808 24148
rect 23768 23798 23796 24142
rect 24492 24132 24544 24138
rect 24492 24074 24544 24080
rect 23756 23792 23808 23798
rect 23756 23734 23808 23740
rect 23664 23724 23716 23730
rect 23664 23666 23716 23672
rect 23848 22568 23900 22574
rect 23848 22510 23900 22516
rect 23020 22432 23072 22438
rect 23020 22374 23072 22380
rect 23032 22234 23060 22374
rect 23020 22228 23072 22234
rect 23020 22170 23072 22176
rect 22652 22160 22704 22166
rect 22652 22102 22704 22108
rect 22560 20936 22612 20942
rect 22560 20878 22612 20884
rect 22376 20528 22428 20534
rect 22376 20470 22428 20476
rect 22296 20216 22416 20244
rect 22052 20156 22360 20165
rect 22052 20154 22058 20156
rect 22114 20154 22138 20156
rect 22194 20154 22218 20156
rect 22274 20154 22298 20156
rect 22354 20154 22360 20156
rect 22114 20102 22116 20154
rect 22296 20102 22298 20154
rect 22052 20100 22058 20102
rect 22114 20100 22138 20102
rect 22194 20100 22218 20102
rect 22274 20100 22298 20102
rect 22354 20100 22360 20102
rect 22052 20091 22360 20100
rect 22388 19378 22416 20216
rect 22376 19372 22428 19378
rect 22376 19314 22428 19320
rect 22052 19068 22360 19077
rect 22052 19066 22058 19068
rect 22114 19066 22138 19068
rect 22194 19066 22218 19068
rect 22274 19066 22298 19068
rect 22354 19066 22360 19068
rect 22114 19014 22116 19066
rect 22296 19014 22298 19066
rect 22052 19012 22058 19014
rect 22114 19012 22138 19014
rect 22194 19012 22218 19014
rect 22274 19012 22298 19014
rect 22354 19012 22360 19014
rect 22052 19003 22360 19012
rect 22052 17980 22360 17989
rect 22052 17978 22058 17980
rect 22114 17978 22138 17980
rect 22194 17978 22218 17980
rect 22274 17978 22298 17980
rect 22354 17978 22360 17980
rect 22114 17926 22116 17978
rect 22296 17926 22298 17978
rect 22052 17924 22058 17926
rect 22114 17924 22138 17926
rect 22194 17924 22218 17926
rect 22274 17924 22298 17926
rect 22354 17924 22360 17926
rect 22052 17915 22360 17924
rect 22560 17128 22612 17134
rect 22560 17070 22612 17076
rect 22376 16992 22428 16998
rect 22376 16934 22428 16940
rect 22052 16892 22360 16901
rect 22052 16890 22058 16892
rect 22114 16890 22138 16892
rect 22194 16890 22218 16892
rect 22274 16890 22298 16892
rect 22354 16890 22360 16892
rect 22114 16838 22116 16890
rect 22296 16838 22298 16890
rect 22052 16836 22058 16838
rect 22114 16836 22138 16838
rect 22194 16836 22218 16838
rect 22274 16836 22298 16838
rect 22354 16836 22360 16838
rect 22052 16827 22360 16836
rect 22388 16794 22416 16934
rect 22376 16788 22428 16794
rect 22376 16730 22428 16736
rect 22008 16108 22060 16114
rect 22008 16050 22060 16056
rect 22376 16108 22428 16114
rect 22376 16050 22428 16056
rect 22020 15910 22048 16050
rect 22008 15904 22060 15910
rect 22008 15846 22060 15852
rect 22052 15804 22360 15813
rect 22052 15802 22058 15804
rect 22114 15802 22138 15804
rect 22194 15802 22218 15804
rect 22274 15802 22298 15804
rect 22354 15802 22360 15804
rect 22114 15750 22116 15802
rect 22296 15750 22298 15802
rect 22052 15748 22058 15750
rect 22114 15748 22138 15750
rect 22194 15748 22218 15750
rect 22274 15748 22298 15750
rect 22354 15748 22360 15750
rect 22052 15739 22360 15748
rect 22388 15638 22416 16050
rect 22376 15632 22428 15638
rect 22376 15574 22428 15580
rect 22572 15570 22600 17070
rect 22664 16250 22692 22102
rect 22836 22024 22888 22030
rect 22836 21966 22888 21972
rect 22652 16244 22704 16250
rect 22652 16186 22704 16192
rect 22652 16108 22704 16114
rect 22652 16050 22704 16056
rect 22560 15564 22612 15570
rect 22560 15506 22612 15512
rect 21824 15156 21876 15162
rect 21824 15098 21876 15104
rect 22192 15020 22244 15026
rect 22192 14962 22244 14968
rect 22376 15020 22428 15026
rect 22376 14962 22428 14968
rect 22468 15020 22520 15026
rect 22468 14962 22520 14968
rect 21916 14952 21968 14958
rect 22204 14929 22232 14962
rect 21916 14894 21968 14900
rect 22190 14920 22246 14929
rect 21732 14612 21784 14618
rect 21732 14554 21784 14560
rect 21744 14414 21772 14554
rect 21928 14498 21956 14894
rect 22190 14855 22246 14864
rect 22052 14716 22360 14725
rect 22052 14714 22058 14716
rect 22114 14714 22138 14716
rect 22194 14714 22218 14716
rect 22274 14714 22298 14716
rect 22354 14714 22360 14716
rect 22114 14662 22116 14714
rect 22296 14662 22298 14714
rect 22052 14660 22058 14662
rect 22114 14660 22138 14662
rect 22194 14660 22218 14662
rect 22274 14660 22298 14662
rect 22354 14660 22360 14662
rect 22052 14651 22360 14660
rect 22100 14544 22152 14550
rect 21928 14492 22100 14498
rect 21928 14486 22152 14492
rect 21928 14470 22140 14486
rect 22388 14414 22416 14962
rect 21640 14408 21692 14414
rect 21640 14350 21692 14356
rect 21732 14408 21784 14414
rect 21732 14350 21784 14356
rect 22376 14408 22428 14414
rect 22376 14350 22428 14356
rect 21652 13938 21680 14350
rect 21824 14340 21876 14346
rect 21824 14282 21876 14288
rect 21836 14006 21864 14282
rect 22480 14090 22508 14962
rect 22558 14376 22614 14385
rect 22558 14311 22614 14320
rect 22388 14074 22508 14090
rect 22376 14068 22508 14074
rect 22428 14062 22508 14068
rect 22376 14010 22428 14016
rect 21824 14000 21876 14006
rect 21824 13942 21876 13948
rect 21640 13932 21692 13938
rect 21640 13874 21692 13880
rect 21652 13394 21680 13874
rect 22052 13628 22360 13637
rect 22052 13626 22058 13628
rect 22114 13626 22138 13628
rect 22194 13626 22218 13628
rect 22274 13626 22298 13628
rect 22354 13626 22360 13628
rect 22114 13574 22116 13626
rect 22296 13574 22298 13626
rect 22052 13572 22058 13574
rect 22114 13572 22138 13574
rect 22194 13572 22218 13574
rect 22274 13572 22298 13574
rect 22354 13572 22360 13574
rect 22052 13563 22360 13572
rect 21640 13388 21692 13394
rect 21640 13330 21692 13336
rect 21364 12640 21416 12646
rect 21364 12582 21416 12588
rect 21456 12640 21508 12646
rect 21456 12582 21508 12588
rect 21376 12238 21404 12582
rect 21364 12232 21416 12238
rect 21364 12174 21416 12180
rect 21178 11248 21234 11257
rect 21178 11183 21234 11192
rect 21376 11150 21404 12174
rect 21088 11144 21140 11150
rect 21364 11144 21416 11150
rect 21088 11086 21140 11092
rect 21178 11112 21234 11121
rect 20996 11008 21048 11014
rect 20996 10950 21048 10956
rect 21100 9110 21128 11086
rect 21364 11086 21416 11092
rect 21178 11047 21180 11056
rect 21232 11047 21234 11056
rect 21180 11018 21232 11024
rect 21272 9648 21324 9654
rect 21272 9590 21324 9596
rect 21284 9178 21312 9590
rect 21468 9586 21496 12582
rect 22052 12540 22360 12549
rect 22052 12538 22058 12540
rect 22114 12538 22138 12540
rect 22194 12538 22218 12540
rect 22274 12538 22298 12540
rect 22354 12538 22360 12540
rect 22114 12486 22116 12538
rect 22296 12486 22298 12538
rect 22052 12484 22058 12486
rect 22114 12484 22138 12486
rect 22194 12484 22218 12486
rect 22274 12484 22298 12486
rect 22354 12484 22360 12486
rect 22052 12475 22360 12484
rect 21548 11688 21600 11694
rect 21548 11630 21600 11636
rect 21560 11354 21588 11630
rect 22052 11452 22360 11461
rect 22052 11450 22058 11452
rect 22114 11450 22138 11452
rect 22194 11450 22218 11452
rect 22274 11450 22298 11452
rect 22354 11450 22360 11452
rect 22114 11398 22116 11450
rect 22296 11398 22298 11450
rect 22052 11396 22058 11398
rect 22114 11396 22138 11398
rect 22194 11396 22218 11398
rect 22274 11396 22298 11398
rect 22354 11396 22360 11398
rect 22052 11387 22360 11396
rect 21548 11348 21600 11354
rect 21548 11290 21600 11296
rect 22282 11248 22338 11257
rect 22282 11183 22338 11192
rect 22296 11150 22324 11183
rect 22192 11144 22244 11150
rect 22192 11086 22244 11092
rect 22284 11144 22336 11150
rect 22284 11086 22336 11092
rect 22204 10810 22232 11086
rect 22192 10804 22244 10810
rect 22192 10746 22244 10752
rect 22388 10674 22416 14010
rect 22572 12306 22600 14311
rect 22664 12918 22692 16050
rect 22652 12912 22704 12918
rect 22652 12854 22704 12860
rect 22664 12481 22692 12854
rect 22650 12472 22706 12481
rect 22650 12407 22706 12416
rect 22560 12300 22612 12306
rect 22560 12242 22612 12248
rect 22468 11892 22520 11898
rect 22468 11834 22520 11840
rect 22480 11354 22508 11834
rect 22572 11830 22600 12242
rect 22560 11824 22612 11830
rect 22560 11766 22612 11772
rect 22744 11824 22796 11830
rect 22744 11766 22796 11772
rect 22652 11552 22704 11558
rect 22652 11494 22704 11500
rect 22468 11348 22520 11354
rect 22468 11290 22520 11296
rect 22664 11150 22692 11494
rect 22652 11144 22704 11150
rect 22652 11086 22704 11092
rect 22376 10668 22428 10674
rect 22376 10610 22428 10616
rect 22052 10364 22360 10373
rect 22052 10362 22058 10364
rect 22114 10362 22138 10364
rect 22194 10362 22218 10364
rect 22274 10362 22298 10364
rect 22354 10362 22360 10364
rect 22114 10310 22116 10362
rect 22296 10310 22298 10362
rect 22052 10308 22058 10310
rect 22114 10308 22138 10310
rect 22194 10308 22218 10310
rect 22274 10308 22298 10310
rect 22354 10308 22360 10310
rect 22052 10299 22360 10308
rect 22388 9602 22416 10610
rect 22652 10532 22704 10538
rect 22652 10474 22704 10480
rect 22388 9586 22508 9602
rect 21456 9580 21508 9586
rect 21456 9522 21508 9528
rect 22388 9580 22520 9586
rect 22388 9574 22468 9580
rect 21272 9172 21324 9178
rect 21272 9114 21324 9120
rect 21088 9104 21140 9110
rect 21088 9046 21140 9052
rect 21468 8498 21496 9522
rect 22052 9276 22360 9285
rect 22052 9274 22058 9276
rect 22114 9274 22138 9276
rect 22194 9274 22218 9276
rect 22274 9274 22298 9276
rect 22354 9274 22360 9276
rect 22114 9222 22116 9274
rect 22296 9222 22298 9274
rect 22052 9220 22058 9222
rect 22114 9220 22138 9222
rect 22194 9220 22218 9222
rect 22274 9220 22298 9222
rect 22354 9220 22360 9222
rect 22052 9211 22360 9220
rect 21916 8832 21968 8838
rect 21916 8774 21968 8780
rect 21456 8492 21508 8498
rect 21456 8434 21508 8440
rect 20904 8424 20956 8430
rect 20904 8366 20956 8372
rect 20812 7812 20864 7818
rect 20812 7754 20864 7760
rect 20916 7546 20944 8366
rect 20720 7540 20772 7546
rect 20720 7482 20772 7488
rect 20904 7540 20956 7546
rect 20904 7482 20956 7488
rect 20732 7426 20760 7482
rect 20628 7404 20680 7410
rect 20732 7398 20852 7426
rect 20628 7346 20680 7352
rect 20720 7200 20772 7206
rect 20720 7142 20772 7148
rect 20536 6860 20588 6866
rect 20536 6802 20588 6808
rect 19524 6792 19576 6798
rect 19524 6734 19576 6740
rect 20444 6792 20496 6798
rect 20444 6734 20496 6740
rect 19536 6254 19564 6734
rect 20732 6390 20760 7142
rect 20824 7002 20852 7398
rect 20812 6996 20864 7002
rect 20812 6938 20864 6944
rect 20916 6458 20944 7482
rect 21928 6798 21956 8774
rect 22052 8188 22360 8197
rect 22052 8186 22058 8188
rect 22114 8186 22138 8188
rect 22194 8186 22218 8188
rect 22274 8186 22298 8188
rect 22354 8186 22360 8188
rect 22114 8134 22116 8186
rect 22296 8134 22298 8186
rect 22052 8132 22058 8134
rect 22114 8132 22138 8134
rect 22194 8132 22218 8134
rect 22274 8132 22298 8134
rect 22354 8132 22360 8134
rect 22052 8123 22360 8132
rect 22388 7562 22416 9574
rect 22468 9522 22520 9528
rect 22664 8974 22692 10474
rect 22652 8968 22704 8974
rect 22652 8910 22704 8916
rect 22756 8566 22784 11766
rect 22848 11354 22876 21966
rect 23204 21480 23256 21486
rect 23204 21422 23256 21428
rect 23572 21480 23624 21486
rect 23572 21422 23624 21428
rect 23216 19922 23244 21422
rect 23584 21146 23612 21422
rect 23860 21350 23888 22510
rect 23940 21480 23992 21486
rect 23940 21422 23992 21428
rect 23848 21344 23900 21350
rect 23848 21286 23900 21292
rect 23572 21140 23624 21146
rect 23572 21082 23624 21088
rect 23756 21140 23808 21146
rect 23756 21082 23808 21088
rect 23768 20942 23796 21082
rect 23952 20942 23980 21422
rect 23756 20936 23808 20942
rect 23756 20878 23808 20884
rect 23940 20936 23992 20942
rect 23940 20878 23992 20884
rect 24124 20868 24176 20874
rect 24124 20810 24176 20816
rect 23388 20800 23440 20806
rect 23388 20742 23440 20748
rect 23940 20800 23992 20806
rect 24136 20754 24164 20810
rect 23992 20748 24164 20754
rect 23940 20742 24164 20748
rect 23204 19916 23256 19922
rect 23204 19858 23256 19864
rect 23020 19508 23072 19514
rect 23020 19450 23072 19456
rect 23032 15502 23060 19450
rect 23216 19378 23244 19858
rect 23204 19372 23256 19378
rect 23204 19314 23256 19320
rect 23400 19310 23428 20742
rect 23952 20726 24164 20742
rect 23388 19304 23440 19310
rect 23388 19246 23440 19252
rect 24504 18766 24532 24074
rect 24688 24070 24716 25298
rect 24872 24886 24900 25706
rect 24860 24880 24912 24886
rect 24860 24822 24912 24828
rect 24676 24064 24728 24070
rect 24676 24006 24728 24012
rect 24688 23254 24716 24006
rect 24676 23248 24728 23254
rect 24676 23190 24728 23196
rect 24872 22982 24900 24822
rect 25148 24818 25176 26250
rect 25332 24818 25360 26318
rect 25516 25974 25544 26318
rect 25700 26042 25728 27406
rect 25792 27334 25820 27950
rect 25872 27940 25924 27946
rect 25872 27882 25924 27888
rect 25884 27538 25912 27882
rect 25872 27532 25924 27538
rect 25872 27474 25924 27480
rect 25780 27328 25832 27334
rect 25780 27270 25832 27276
rect 25884 26994 25912 27474
rect 25872 26988 25924 26994
rect 25872 26930 25924 26936
rect 25964 26580 26016 26586
rect 25964 26522 26016 26528
rect 25872 26376 25924 26382
rect 25872 26318 25924 26324
rect 25688 26036 25740 26042
rect 25688 25978 25740 25984
rect 25504 25968 25556 25974
rect 25504 25910 25556 25916
rect 25884 25906 25912 26318
rect 25872 25900 25924 25906
rect 25872 25842 25924 25848
rect 25976 25498 26004 26522
rect 26068 25838 26096 29514
rect 26272 29404 26580 29413
rect 26272 29402 26278 29404
rect 26334 29402 26358 29404
rect 26414 29402 26438 29404
rect 26494 29402 26518 29404
rect 26574 29402 26580 29404
rect 26334 29350 26336 29402
rect 26516 29350 26518 29402
rect 26272 29348 26278 29350
rect 26334 29348 26358 29350
rect 26414 29348 26438 29350
rect 26494 29348 26518 29350
rect 26574 29348 26580 29350
rect 26272 29339 26580 29348
rect 27172 28626 27200 30330
rect 27540 30258 27568 31282
rect 27724 30734 27752 31282
rect 28448 31204 28500 31210
rect 28448 31146 28500 31152
rect 27712 30728 27764 30734
rect 27712 30670 27764 30676
rect 28080 30728 28132 30734
rect 28080 30670 28132 30676
rect 27528 30252 27580 30258
rect 27528 30194 27580 30200
rect 27528 30048 27580 30054
rect 27528 29990 27580 29996
rect 27356 29850 27476 29866
rect 27356 29844 27488 29850
rect 27356 29838 27436 29844
rect 27160 28620 27212 28626
rect 27160 28562 27212 28568
rect 27252 28416 27304 28422
rect 27252 28358 27304 28364
rect 26272 28316 26580 28325
rect 26272 28314 26278 28316
rect 26334 28314 26358 28316
rect 26414 28314 26438 28316
rect 26494 28314 26518 28316
rect 26574 28314 26580 28316
rect 26334 28262 26336 28314
rect 26516 28262 26518 28314
rect 26272 28260 26278 28262
rect 26334 28260 26358 28262
rect 26414 28260 26438 28262
rect 26494 28260 26518 28262
rect 26574 28260 26580 28262
rect 26272 28251 26580 28260
rect 27068 28076 27120 28082
rect 27068 28018 27120 28024
rect 26240 28008 26292 28014
rect 26240 27950 26292 27956
rect 26148 27464 26200 27470
rect 26148 27406 26200 27412
rect 26160 27062 26188 27406
rect 26252 27402 26280 27950
rect 26608 27872 26660 27878
rect 26608 27814 26660 27820
rect 26240 27396 26292 27402
rect 26240 27338 26292 27344
rect 26272 27228 26580 27237
rect 26272 27226 26278 27228
rect 26334 27226 26358 27228
rect 26414 27226 26438 27228
rect 26494 27226 26518 27228
rect 26574 27226 26580 27228
rect 26334 27174 26336 27226
rect 26516 27174 26518 27226
rect 26272 27172 26278 27174
rect 26334 27172 26358 27174
rect 26414 27172 26438 27174
rect 26494 27172 26518 27174
rect 26574 27172 26580 27174
rect 26272 27163 26580 27172
rect 26148 27056 26200 27062
rect 26148 26998 26200 27004
rect 26148 26920 26200 26926
rect 26148 26862 26200 26868
rect 26056 25832 26108 25838
rect 26056 25774 26108 25780
rect 25964 25492 26016 25498
rect 25964 25434 26016 25440
rect 26068 25226 26096 25774
rect 26056 25220 26108 25226
rect 26056 25162 26108 25168
rect 25136 24812 25188 24818
rect 25136 24754 25188 24760
rect 25320 24812 25372 24818
rect 25320 24754 25372 24760
rect 25964 24608 26016 24614
rect 25964 24550 26016 24556
rect 25228 24064 25280 24070
rect 25228 24006 25280 24012
rect 24952 23520 25004 23526
rect 24952 23462 25004 23468
rect 24860 22976 24912 22982
rect 24860 22918 24912 22924
rect 24584 22432 24636 22438
rect 24584 22374 24636 22380
rect 24596 22030 24624 22374
rect 24872 22098 24900 22918
rect 24964 22098 24992 23462
rect 25240 23186 25268 24006
rect 25976 23526 26004 24550
rect 25964 23520 26016 23526
rect 25964 23462 26016 23468
rect 25228 23180 25280 23186
rect 25228 23122 25280 23128
rect 25320 23044 25372 23050
rect 25320 22986 25372 22992
rect 25136 22976 25188 22982
rect 25136 22918 25188 22924
rect 25148 22710 25176 22918
rect 25136 22704 25188 22710
rect 25136 22646 25188 22652
rect 24860 22092 24912 22098
rect 24860 22034 24912 22040
rect 24952 22092 25004 22098
rect 24952 22034 25004 22040
rect 25148 22030 25176 22646
rect 24584 22024 24636 22030
rect 24584 21966 24636 21972
rect 24768 22024 24820 22030
rect 24768 21966 24820 21972
rect 25136 22024 25188 22030
rect 25136 21966 25188 21972
rect 24676 20936 24728 20942
rect 24676 20878 24728 20884
rect 24688 20602 24716 20878
rect 24676 20596 24728 20602
rect 24676 20538 24728 20544
rect 24780 20058 24808 21966
rect 25044 21888 25096 21894
rect 25044 21830 25096 21836
rect 24952 20800 25004 20806
rect 24952 20742 25004 20748
rect 24768 20052 24820 20058
rect 24768 19994 24820 20000
rect 24964 19446 24992 20742
rect 24952 19440 25004 19446
rect 24952 19382 25004 19388
rect 24492 18760 24544 18766
rect 24492 18702 24544 18708
rect 23480 18624 23532 18630
rect 23480 18566 23532 18572
rect 24216 18624 24268 18630
rect 24216 18566 24268 18572
rect 23492 18290 23520 18566
rect 24228 18358 24256 18566
rect 24504 18426 24532 18702
rect 24584 18624 24636 18630
rect 24584 18566 24636 18572
rect 24492 18420 24544 18426
rect 24492 18362 24544 18368
rect 24216 18352 24268 18358
rect 24216 18294 24268 18300
rect 23480 18284 23532 18290
rect 23480 18226 23532 18232
rect 23112 18216 23164 18222
rect 23112 18158 23164 18164
rect 23124 17134 23152 18158
rect 24492 17604 24544 17610
rect 24492 17546 24544 17552
rect 23756 17196 23808 17202
rect 23756 17138 23808 17144
rect 23112 17128 23164 17134
rect 23112 17070 23164 17076
rect 23296 16992 23348 16998
rect 23296 16934 23348 16940
rect 23020 15496 23072 15502
rect 23020 15438 23072 15444
rect 22928 15360 22980 15366
rect 22928 15302 22980 15308
rect 22940 15162 22968 15302
rect 22928 15156 22980 15162
rect 22928 15098 22980 15104
rect 23032 15026 23060 15438
rect 23308 15162 23336 16934
rect 23388 15496 23440 15502
rect 23388 15438 23440 15444
rect 23400 15162 23428 15438
rect 23480 15360 23532 15366
rect 23480 15302 23532 15308
rect 23296 15156 23348 15162
rect 23296 15098 23348 15104
rect 23388 15156 23440 15162
rect 23388 15098 23440 15104
rect 23020 15020 23072 15026
rect 23020 14962 23072 14968
rect 23492 14414 23520 15302
rect 23664 14816 23716 14822
rect 23664 14758 23716 14764
rect 23676 14618 23704 14758
rect 23664 14612 23716 14618
rect 23664 14554 23716 14560
rect 23480 14408 23532 14414
rect 23480 14350 23532 14356
rect 23570 14376 23626 14385
rect 23570 14311 23572 14320
rect 23624 14311 23626 14320
rect 23572 14282 23624 14288
rect 23676 14074 23704 14554
rect 23768 14482 23796 17138
rect 24504 16046 24532 17546
rect 24596 17270 24624 18566
rect 24952 18080 25004 18086
rect 24952 18022 25004 18028
rect 24584 17264 24636 17270
rect 24584 17206 24636 17212
rect 24584 16584 24636 16590
rect 24584 16526 24636 16532
rect 24676 16584 24728 16590
rect 24676 16526 24728 16532
rect 24492 16040 24544 16046
rect 24492 15982 24544 15988
rect 24504 15502 24532 15982
rect 24596 15910 24624 16526
rect 24584 15904 24636 15910
rect 24584 15846 24636 15852
rect 24492 15496 24544 15502
rect 24492 15438 24544 15444
rect 23756 14476 23808 14482
rect 23756 14418 23808 14424
rect 23664 14068 23716 14074
rect 23664 14010 23716 14016
rect 23664 12164 23716 12170
rect 23664 12106 23716 12112
rect 22928 11552 22980 11558
rect 22928 11494 22980 11500
rect 23480 11552 23532 11558
rect 23480 11494 23532 11500
rect 22836 11348 22888 11354
rect 22836 11290 22888 11296
rect 22940 11121 22968 11494
rect 22926 11112 22982 11121
rect 23492 11082 23520 11494
rect 23572 11144 23624 11150
rect 23676 11132 23704 12106
rect 23624 11104 23704 11132
rect 23572 11086 23624 11092
rect 22926 11047 22982 11056
rect 23480 11076 23532 11082
rect 22940 10674 22968 11047
rect 23480 11018 23532 11024
rect 23572 10804 23624 10810
rect 23572 10746 23624 10752
rect 22928 10668 22980 10674
rect 22928 10610 22980 10616
rect 23480 10600 23532 10606
rect 23480 10542 23532 10548
rect 22836 9172 22888 9178
rect 22836 9114 22888 9120
rect 22848 8974 22876 9114
rect 23388 9104 23440 9110
rect 23388 9046 23440 9052
rect 22836 8968 22888 8974
rect 22836 8910 22888 8916
rect 22744 8560 22796 8566
rect 22744 8502 22796 8508
rect 22296 7534 22416 7562
rect 22296 7478 22324 7534
rect 22284 7472 22336 7478
rect 22284 7414 22336 7420
rect 22052 7100 22360 7109
rect 22052 7098 22058 7100
rect 22114 7098 22138 7100
rect 22194 7098 22218 7100
rect 22274 7098 22298 7100
rect 22354 7098 22360 7100
rect 22114 7046 22116 7098
rect 22296 7046 22298 7098
rect 22052 7044 22058 7046
rect 22114 7044 22138 7046
rect 22194 7044 22218 7046
rect 22274 7044 22298 7046
rect 22354 7044 22360 7046
rect 22052 7035 22360 7044
rect 21916 6792 21968 6798
rect 21916 6734 21968 6740
rect 22848 6662 22876 8910
rect 23400 8634 23428 9046
rect 23388 8628 23440 8634
rect 23388 8570 23440 8576
rect 23388 7744 23440 7750
rect 23388 7686 23440 7692
rect 23400 7478 23428 7686
rect 23388 7472 23440 7478
rect 23388 7414 23440 7420
rect 22836 6656 22888 6662
rect 22836 6598 22888 6604
rect 20904 6452 20956 6458
rect 20904 6394 20956 6400
rect 20720 6384 20772 6390
rect 20720 6326 20772 6332
rect 19524 6248 19576 6254
rect 19524 6190 19576 6196
rect 19536 5370 19564 6190
rect 20168 6112 20220 6118
rect 20168 6054 20220 6060
rect 19524 5364 19576 5370
rect 19524 5306 19576 5312
rect 18696 5296 18748 5302
rect 18696 5238 18748 5244
rect 20180 4622 20208 6054
rect 22052 6012 22360 6021
rect 22052 6010 22058 6012
rect 22114 6010 22138 6012
rect 22194 6010 22218 6012
rect 22274 6010 22298 6012
rect 22354 6010 22360 6012
rect 22114 5958 22116 6010
rect 22296 5958 22298 6010
rect 22052 5956 22058 5958
rect 22114 5956 22138 5958
rect 22194 5956 22218 5958
rect 22274 5956 22298 5958
rect 22354 5956 22360 5958
rect 22052 5947 22360 5956
rect 23400 5302 23428 7414
rect 23492 6730 23520 10542
rect 23584 9654 23612 10746
rect 23572 9648 23624 9654
rect 23572 9590 23624 9596
rect 23584 8566 23612 9590
rect 23676 8974 23704 11104
rect 23768 10742 23796 14418
rect 24032 14272 24084 14278
rect 24032 14214 24084 14220
rect 24044 13938 24072 14214
rect 24504 13938 24532 15438
rect 24596 14482 24624 15846
rect 24688 15434 24716 16526
rect 24676 15428 24728 15434
rect 24676 15370 24728 15376
rect 24674 14920 24730 14929
rect 24674 14855 24730 14864
rect 24584 14476 24636 14482
rect 24584 14418 24636 14424
rect 24032 13932 24084 13938
rect 24032 13874 24084 13880
rect 24492 13932 24544 13938
rect 24492 13874 24544 13880
rect 24044 12782 24072 13874
rect 24032 12776 24084 12782
rect 24032 12718 24084 12724
rect 24504 12170 24532 13874
rect 24688 13802 24716 14855
rect 24676 13796 24728 13802
rect 24676 13738 24728 13744
rect 24492 12164 24544 12170
rect 24492 12106 24544 12112
rect 24584 12096 24636 12102
rect 24584 12038 24636 12044
rect 24596 11762 24624 12038
rect 24584 11756 24636 11762
rect 24584 11698 24636 11704
rect 23848 11688 23900 11694
rect 23848 11630 23900 11636
rect 23756 10736 23808 10742
rect 23756 10678 23808 10684
rect 23860 10266 23888 11630
rect 24688 11218 24716 13738
rect 24964 12434 24992 18022
rect 25056 17202 25084 21830
rect 25228 18760 25280 18766
rect 25228 18702 25280 18708
rect 25136 18624 25188 18630
rect 25136 18566 25188 18572
rect 25148 17338 25176 18566
rect 25240 17678 25268 18702
rect 25332 18290 25360 22986
rect 26160 22574 26188 26862
rect 26620 26586 26648 27814
rect 27080 27334 27108 28018
rect 26700 27328 26752 27334
rect 26700 27270 26752 27276
rect 27068 27328 27120 27334
rect 27068 27270 27120 27276
rect 26608 26580 26660 26586
rect 26608 26522 26660 26528
rect 26620 26466 26648 26522
rect 26528 26438 26648 26466
rect 26528 26382 26556 26438
rect 26516 26376 26568 26382
rect 26516 26318 26568 26324
rect 26272 26140 26580 26149
rect 26272 26138 26278 26140
rect 26334 26138 26358 26140
rect 26414 26138 26438 26140
rect 26494 26138 26518 26140
rect 26574 26138 26580 26140
rect 26334 26086 26336 26138
rect 26516 26086 26518 26138
rect 26272 26084 26278 26086
rect 26334 26084 26358 26086
rect 26414 26084 26438 26086
rect 26494 26084 26518 26086
rect 26574 26084 26580 26086
rect 26272 26075 26580 26084
rect 26516 25900 26568 25906
rect 26516 25842 26568 25848
rect 26528 25226 26556 25842
rect 26712 25838 26740 27270
rect 27080 26586 27108 27270
rect 27264 26994 27292 28358
rect 27356 26994 27384 29838
rect 27436 29786 27488 29792
rect 27436 29708 27488 29714
rect 27436 29650 27488 29656
rect 27448 29170 27476 29650
rect 27540 29306 27568 29990
rect 27724 29646 27752 30670
rect 28092 30326 28120 30670
rect 28460 30394 28488 31146
rect 28552 30666 28580 31282
rect 28632 30728 28684 30734
rect 28632 30670 28684 30676
rect 28540 30660 28592 30666
rect 28540 30602 28592 30608
rect 28448 30388 28500 30394
rect 28448 30330 28500 30336
rect 28080 30320 28132 30326
rect 28080 30262 28132 30268
rect 27896 30184 27948 30190
rect 27896 30126 27948 30132
rect 27908 29782 27936 30126
rect 27896 29776 27948 29782
rect 27896 29718 27948 29724
rect 28092 29714 28120 30262
rect 28460 30122 28488 30330
rect 28552 30122 28580 30602
rect 28448 30116 28500 30122
rect 28448 30058 28500 30064
rect 28540 30116 28592 30122
rect 28540 30058 28592 30064
rect 28644 29714 28672 30670
rect 28908 30252 28960 30258
rect 28908 30194 28960 30200
rect 29920 30252 29972 30258
rect 29920 30194 29972 30200
rect 28080 29708 28132 29714
rect 28080 29650 28132 29656
rect 28632 29708 28684 29714
rect 28632 29650 28684 29656
rect 27712 29640 27764 29646
rect 27712 29582 27764 29588
rect 28264 29640 28316 29646
rect 28264 29582 28316 29588
rect 27528 29300 27580 29306
rect 27528 29242 27580 29248
rect 27620 29300 27672 29306
rect 27620 29242 27672 29248
rect 27908 29294 28120 29322
rect 28276 29306 28304 29582
rect 27436 29164 27488 29170
rect 27436 29106 27488 29112
rect 27528 28960 27580 28966
rect 27528 28902 27580 28908
rect 27252 26988 27304 26994
rect 27252 26930 27304 26936
rect 27344 26988 27396 26994
rect 27344 26930 27396 26936
rect 27160 26784 27212 26790
rect 27160 26726 27212 26732
rect 26792 26580 26844 26586
rect 26792 26522 26844 26528
rect 27068 26580 27120 26586
rect 27068 26522 27120 26528
rect 26804 26246 26832 26522
rect 27172 26382 27200 26726
rect 26884 26376 26936 26382
rect 26884 26318 26936 26324
rect 27160 26376 27212 26382
rect 27160 26318 27212 26324
rect 26792 26240 26844 26246
rect 26792 26182 26844 26188
rect 26700 25832 26752 25838
rect 26700 25774 26752 25780
rect 26608 25356 26660 25362
rect 26608 25298 26660 25304
rect 26516 25220 26568 25226
rect 26516 25162 26568 25168
rect 26272 25052 26580 25061
rect 26272 25050 26278 25052
rect 26334 25050 26358 25052
rect 26414 25050 26438 25052
rect 26494 25050 26518 25052
rect 26574 25050 26580 25052
rect 26334 24998 26336 25050
rect 26516 24998 26518 25050
rect 26272 24996 26278 24998
rect 26334 24996 26358 24998
rect 26414 24996 26438 24998
rect 26494 24996 26518 24998
rect 26574 24996 26580 24998
rect 26272 24987 26580 24996
rect 26620 24614 26648 25298
rect 26608 24608 26660 24614
rect 26608 24550 26660 24556
rect 26712 24206 26740 25774
rect 26804 25498 26832 26182
rect 26896 25770 26924 26318
rect 27264 26042 27292 26930
rect 27252 26036 27304 26042
rect 27252 25978 27304 25984
rect 27068 25832 27120 25838
rect 27068 25774 27120 25780
rect 26884 25764 26936 25770
rect 26884 25706 26936 25712
rect 26792 25492 26844 25498
rect 26792 25434 26844 25440
rect 27080 25158 27108 25774
rect 27252 25288 27304 25294
rect 27356 25276 27384 26930
rect 27540 26518 27568 28902
rect 27632 28626 27660 29242
rect 27908 29034 27936 29294
rect 28092 29238 28120 29294
rect 28264 29300 28316 29306
rect 28264 29242 28316 29248
rect 27988 29232 28040 29238
rect 27988 29174 28040 29180
rect 28080 29232 28132 29238
rect 28080 29174 28132 29180
rect 27896 29028 27948 29034
rect 27896 28970 27948 28976
rect 27620 28620 27672 28626
rect 27620 28562 27672 28568
rect 27632 26926 27660 28562
rect 27896 28552 27948 28558
rect 27896 28494 27948 28500
rect 27712 28076 27764 28082
rect 27712 28018 27764 28024
rect 27724 27470 27752 28018
rect 27908 27606 27936 28494
rect 27896 27600 27948 27606
rect 27896 27542 27948 27548
rect 28000 27470 28028 29174
rect 28644 29102 28672 29650
rect 28816 29640 28868 29646
rect 28816 29582 28868 29588
rect 28632 29096 28684 29102
rect 28632 29038 28684 29044
rect 28828 28966 28856 29582
rect 28920 29306 28948 30194
rect 29092 30184 29144 30190
rect 29092 30126 29144 30132
rect 29104 29510 29132 30126
rect 29932 29850 29960 30194
rect 29920 29844 29972 29850
rect 29920 29786 29972 29792
rect 29092 29504 29144 29510
rect 29092 29446 29144 29452
rect 28908 29300 28960 29306
rect 28908 29242 28960 29248
rect 28920 29170 28948 29242
rect 29104 29170 29132 29446
rect 28908 29164 28960 29170
rect 28908 29106 28960 29112
rect 29092 29164 29144 29170
rect 29092 29106 29144 29112
rect 28816 28960 28868 28966
rect 28816 28902 28868 28908
rect 28828 28762 28856 28902
rect 28816 28756 28868 28762
rect 28816 28698 28868 28704
rect 29000 28552 29052 28558
rect 29000 28494 29052 28500
rect 29012 27470 29040 28494
rect 29276 28076 29328 28082
rect 29276 28018 29328 28024
rect 27712 27464 27764 27470
rect 27712 27406 27764 27412
rect 27988 27464 28040 27470
rect 27988 27406 28040 27412
rect 29000 27464 29052 27470
rect 29000 27406 29052 27412
rect 27620 26920 27672 26926
rect 27620 26862 27672 26868
rect 27528 26512 27580 26518
rect 27528 26454 27580 26460
rect 27540 25838 27568 26454
rect 27620 26308 27672 26314
rect 27620 26250 27672 26256
rect 27632 25906 27660 26250
rect 27620 25900 27672 25906
rect 27620 25842 27672 25848
rect 27528 25832 27580 25838
rect 27528 25774 27580 25780
rect 27304 25248 27384 25276
rect 27252 25230 27304 25236
rect 27068 25152 27120 25158
rect 27068 25094 27120 25100
rect 27080 24886 27108 25094
rect 27068 24880 27120 24886
rect 27068 24822 27120 24828
rect 27160 24880 27212 24886
rect 27160 24822 27212 24828
rect 26700 24200 26752 24206
rect 26700 24142 26752 24148
rect 26272 23964 26580 23973
rect 26272 23962 26278 23964
rect 26334 23962 26358 23964
rect 26414 23962 26438 23964
rect 26494 23962 26518 23964
rect 26574 23962 26580 23964
rect 26334 23910 26336 23962
rect 26516 23910 26518 23962
rect 26272 23908 26278 23910
rect 26334 23908 26358 23910
rect 26414 23908 26438 23910
rect 26494 23908 26518 23910
rect 26574 23908 26580 23910
rect 26272 23899 26580 23908
rect 27172 23662 27200 24822
rect 27540 24274 27568 25774
rect 27632 25498 27660 25842
rect 27620 25492 27672 25498
rect 27620 25434 27672 25440
rect 28000 24750 28028 27406
rect 28632 26512 28684 26518
rect 28632 26454 28684 26460
rect 28644 25974 28672 26454
rect 28724 26376 28776 26382
rect 28724 26318 28776 26324
rect 28908 26376 28960 26382
rect 29012 26330 29040 27406
rect 29184 27396 29236 27402
rect 29184 27338 29236 27344
rect 29196 26586 29224 27338
rect 29184 26580 29236 26586
rect 29184 26522 29236 26528
rect 28960 26324 29040 26330
rect 28908 26318 29040 26324
rect 28632 25968 28684 25974
rect 28632 25910 28684 25916
rect 27988 24744 28040 24750
rect 27988 24686 28040 24692
rect 27528 24268 27580 24274
rect 27528 24210 27580 24216
rect 28644 23798 28672 25910
rect 28736 24274 28764 26318
rect 28920 26302 29040 26318
rect 29092 26308 29144 26314
rect 29092 26250 29144 26256
rect 29000 26240 29052 26246
rect 29000 26182 29052 26188
rect 28908 25288 28960 25294
rect 28908 25230 28960 25236
rect 28816 24880 28868 24886
rect 28816 24822 28868 24828
rect 28724 24268 28776 24274
rect 28724 24210 28776 24216
rect 28632 23792 28684 23798
rect 28632 23734 28684 23740
rect 27160 23656 27212 23662
rect 27160 23598 27212 23604
rect 27712 23180 27764 23186
rect 27712 23122 27764 23128
rect 27528 23112 27580 23118
rect 27528 23054 27580 23060
rect 26272 22876 26580 22885
rect 26272 22874 26278 22876
rect 26334 22874 26358 22876
rect 26414 22874 26438 22876
rect 26494 22874 26518 22876
rect 26574 22874 26580 22876
rect 26334 22822 26336 22874
rect 26516 22822 26518 22874
rect 26272 22820 26278 22822
rect 26334 22820 26358 22822
rect 26414 22820 26438 22822
rect 26494 22820 26518 22822
rect 26574 22820 26580 22822
rect 26272 22811 26580 22820
rect 27160 22636 27212 22642
rect 27160 22578 27212 22584
rect 26148 22568 26200 22574
rect 26148 22510 26200 22516
rect 26976 22432 27028 22438
rect 26976 22374 27028 22380
rect 26988 22098 27016 22374
rect 26976 22092 27028 22098
rect 26976 22034 27028 22040
rect 27068 22024 27120 22030
rect 27068 21966 27120 21972
rect 26884 21888 26936 21894
rect 26884 21830 26936 21836
rect 26976 21888 27028 21894
rect 26976 21830 27028 21836
rect 26272 21788 26580 21797
rect 26272 21786 26278 21788
rect 26334 21786 26358 21788
rect 26414 21786 26438 21788
rect 26494 21786 26518 21788
rect 26574 21786 26580 21788
rect 26334 21734 26336 21786
rect 26516 21734 26518 21786
rect 26272 21732 26278 21734
rect 26334 21732 26358 21734
rect 26414 21732 26438 21734
rect 26494 21732 26518 21734
rect 26574 21732 26580 21734
rect 26272 21723 26580 21732
rect 26896 21622 26924 21830
rect 26988 21690 27016 21830
rect 26976 21684 27028 21690
rect 26976 21626 27028 21632
rect 26884 21616 26936 21622
rect 26884 21558 26936 21564
rect 25872 21072 25924 21078
rect 25872 21014 25924 21020
rect 25964 21072 26016 21078
rect 25964 21014 26016 21020
rect 25504 20936 25556 20942
rect 25504 20878 25556 20884
rect 25516 18766 25544 20878
rect 25884 18970 25912 21014
rect 25976 20602 26004 21014
rect 26272 20700 26580 20709
rect 26272 20698 26278 20700
rect 26334 20698 26358 20700
rect 26414 20698 26438 20700
rect 26494 20698 26518 20700
rect 26574 20698 26580 20700
rect 26334 20646 26336 20698
rect 26516 20646 26518 20698
rect 26272 20644 26278 20646
rect 26334 20644 26358 20646
rect 26414 20644 26438 20646
rect 26494 20644 26518 20646
rect 26574 20644 26580 20646
rect 26272 20635 26580 20644
rect 25964 20596 26016 20602
rect 25964 20538 26016 20544
rect 26272 19612 26580 19621
rect 26272 19610 26278 19612
rect 26334 19610 26358 19612
rect 26414 19610 26438 19612
rect 26494 19610 26518 19612
rect 26574 19610 26580 19612
rect 26334 19558 26336 19610
rect 26516 19558 26518 19610
rect 26272 19556 26278 19558
rect 26334 19556 26358 19558
rect 26414 19556 26438 19558
rect 26494 19556 26518 19558
rect 26574 19556 26580 19558
rect 26272 19547 26580 19556
rect 26424 19168 26476 19174
rect 26424 19110 26476 19116
rect 25872 18964 25924 18970
rect 25872 18906 25924 18912
rect 26436 18834 26464 19110
rect 26424 18828 26476 18834
rect 26424 18770 26476 18776
rect 25504 18760 25556 18766
rect 25504 18702 25556 18708
rect 26240 18760 26292 18766
rect 26240 18702 26292 18708
rect 25688 18692 25740 18698
rect 25688 18634 25740 18640
rect 25700 18426 25728 18634
rect 26252 18630 26280 18702
rect 27080 18630 27108 21966
rect 27172 21690 27200 22578
rect 27250 22128 27306 22137
rect 27250 22063 27252 22072
rect 27304 22063 27306 22072
rect 27252 22034 27304 22040
rect 27540 21962 27568 23054
rect 27620 23044 27672 23050
rect 27620 22986 27672 22992
rect 27528 21956 27580 21962
rect 27528 21898 27580 21904
rect 27540 21690 27568 21898
rect 27160 21684 27212 21690
rect 27160 21626 27212 21632
rect 27528 21684 27580 21690
rect 27528 21626 27580 21632
rect 27632 21486 27660 22986
rect 27724 21554 27752 23122
rect 27988 23112 28040 23118
rect 27988 23054 28040 23060
rect 28264 23112 28316 23118
rect 28264 23054 28316 23060
rect 28000 22642 28028 23054
rect 28276 22642 28304 23054
rect 27988 22636 28040 22642
rect 27988 22578 28040 22584
rect 28264 22636 28316 22642
rect 28264 22578 28316 22584
rect 28000 22094 28028 22578
rect 28000 22066 28304 22094
rect 27712 21548 27764 21554
rect 27712 21490 27764 21496
rect 27344 21480 27396 21486
rect 27344 21422 27396 21428
rect 27620 21480 27672 21486
rect 27620 21422 27672 21428
rect 27356 20874 27384 21422
rect 27896 21344 27948 21350
rect 27896 21286 27948 21292
rect 27344 20868 27396 20874
rect 27344 20810 27396 20816
rect 27908 20398 27936 21286
rect 27988 20460 28040 20466
rect 27988 20402 28040 20408
rect 27896 20392 27948 20398
rect 27896 20334 27948 20340
rect 27344 19372 27396 19378
rect 27344 19314 27396 19320
rect 27436 19372 27488 19378
rect 27436 19314 27488 19320
rect 27356 18766 27384 19314
rect 27448 18766 27476 19314
rect 27804 18896 27856 18902
rect 27804 18838 27856 18844
rect 27344 18760 27396 18766
rect 27344 18702 27396 18708
rect 27436 18760 27488 18766
rect 27436 18702 27488 18708
rect 27620 18760 27672 18766
rect 27620 18702 27672 18708
rect 26240 18624 26292 18630
rect 26240 18566 26292 18572
rect 27068 18624 27120 18630
rect 27068 18566 27120 18572
rect 26272 18524 26580 18533
rect 26272 18522 26278 18524
rect 26334 18522 26358 18524
rect 26414 18522 26438 18524
rect 26494 18522 26518 18524
rect 26574 18522 26580 18524
rect 26334 18470 26336 18522
rect 26516 18470 26518 18522
rect 26272 18468 26278 18470
rect 26334 18468 26358 18470
rect 26414 18468 26438 18470
rect 26494 18468 26518 18470
rect 26574 18468 26580 18470
rect 26272 18459 26580 18468
rect 25688 18420 25740 18426
rect 25688 18362 25740 18368
rect 25320 18284 25372 18290
rect 25320 18226 25372 18232
rect 27356 18222 27384 18702
rect 27632 18426 27660 18702
rect 27620 18420 27672 18426
rect 27620 18362 27672 18368
rect 25412 18216 25464 18222
rect 25412 18158 25464 18164
rect 27344 18216 27396 18222
rect 27344 18158 27396 18164
rect 25228 17672 25280 17678
rect 25228 17614 25280 17620
rect 25136 17332 25188 17338
rect 25136 17274 25188 17280
rect 25044 17196 25096 17202
rect 25044 17138 25096 17144
rect 25148 16266 25176 17274
rect 25148 16238 25268 16266
rect 25136 16108 25188 16114
rect 25136 16050 25188 16056
rect 25148 15706 25176 16050
rect 25240 15910 25268 16238
rect 25228 15904 25280 15910
rect 25228 15846 25280 15852
rect 25136 15700 25188 15706
rect 25136 15642 25188 15648
rect 25228 15428 25280 15434
rect 25228 15370 25280 15376
rect 25136 15156 25188 15162
rect 25136 15098 25188 15104
rect 25044 15020 25096 15026
rect 25044 14962 25096 14968
rect 25056 14074 25084 14962
rect 25148 14464 25176 15098
rect 25240 14618 25268 15370
rect 25228 14612 25280 14618
rect 25228 14554 25280 14560
rect 25148 14436 25268 14464
rect 25044 14068 25096 14074
rect 25044 14010 25096 14016
rect 25044 13932 25096 13938
rect 25044 13874 25096 13880
rect 25056 12646 25084 13874
rect 25044 12640 25096 12646
rect 25044 12582 25096 12588
rect 25240 12434 25268 14436
rect 24964 12406 25084 12434
rect 24952 12096 25004 12102
rect 24952 12038 25004 12044
rect 24964 11558 24992 12038
rect 24952 11552 25004 11558
rect 24952 11494 25004 11500
rect 23940 11212 23992 11218
rect 23940 11154 23992 11160
rect 24676 11212 24728 11218
rect 24676 11154 24728 11160
rect 23848 10260 23900 10266
rect 23848 10202 23900 10208
rect 23952 9518 23980 11154
rect 24860 11076 24912 11082
rect 24860 11018 24912 11024
rect 24872 10742 24900 11018
rect 24860 10736 24912 10742
rect 24860 10678 24912 10684
rect 24584 10600 24636 10606
rect 24584 10542 24636 10548
rect 24596 10266 24624 10542
rect 24584 10260 24636 10266
rect 24584 10202 24636 10208
rect 24768 10056 24820 10062
rect 24768 9998 24820 10004
rect 24780 9654 24808 9998
rect 24768 9648 24820 9654
rect 24768 9590 24820 9596
rect 23940 9512 23992 9518
rect 23940 9454 23992 9460
rect 23664 8968 23716 8974
rect 23664 8910 23716 8916
rect 23664 8832 23716 8838
rect 23664 8774 23716 8780
rect 23676 8634 23704 8774
rect 23952 8634 23980 9454
rect 25056 9450 25084 12406
rect 25148 12406 25268 12434
rect 25044 9444 25096 9450
rect 25044 9386 25096 9392
rect 24584 8968 24636 8974
rect 24584 8910 24636 8916
rect 23664 8628 23716 8634
rect 23664 8570 23716 8576
rect 23940 8628 23992 8634
rect 23940 8570 23992 8576
rect 23572 8560 23624 8566
rect 23572 8502 23624 8508
rect 24032 8356 24084 8362
rect 24032 8298 24084 8304
rect 24044 7886 24072 8298
rect 24032 7880 24084 7886
rect 24032 7822 24084 7828
rect 24596 7342 24624 8910
rect 25044 8832 25096 8838
rect 25044 8774 25096 8780
rect 25056 8566 25084 8774
rect 25044 8560 25096 8566
rect 25044 8502 25096 8508
rect 24952 8492 25004 8498
rect 24952 8434 25004 8440
rect 23756 7336 23808 7342
rect 23756 7278 23808 7284
rect 24032 7336 24084 7342
rect 24032 7278 24084 7284
rect 24584 7336 24636 7342
rect 24584 7278 24636 7284
rect 23768 6798 23796 7278
rect 24044 6798 24072 7278
rect 23756 6792 23808 6798
rect 23756 6734 23808 6740
rect 24032 6792 24084 6798
rect 24032 6734 24084 6740
rect 24964 6730 24992 8434
rect 25044 8424 25096 8430
rect 25044 8366 25096 8372
rect 25056 7478 25084 8366
rect 25148 7954 25176 12406
rect 25320 11756 25372 11762
rect 25320 11698 25372 11704
rect 25332 11354 25360 11698
rect 25320 11348 25372 11354
rect 25320 11290 25372 11296
rect 25332 10062 25360 11290
rect 25424 10266 25452 18158
rect 27632 17746 27660 18362
rect 27620 17740 27672 17746
rect 27620 17682 27672 17688
rect 25688 17672 25740 17678
rect 25688 17614 25740 17620
rect 25700 17338 25728 17614
rect 27816 17610 27844 18838
rect 28000 17882 28028 20402
rect 28080 20256 28132 20262
rect 28080 20198 28132 20204
rect 28092 18170 28120 20198
rect 28172 19712 28224 19718
rect 28172 19654 28224 19660
rect 28184 18290 28212 19654
rect 28276 18970 28304 22066
rect 28448 21956 28500 21962
rect 28448 21898 28500 21904
rect 28460 21622 28488 21898
rect 28448 21616 28500 21622
rect 28448 21558 28500 21564
rect 28448 21344 28500 21350
rect 28448 21286 28500 21292
rect 28460 21010 28488 21286
rect 28448 21004 28500 21010
rect 28448 20946 28500 20952
rect 28736 20942 28764 24210
rect 28828 23594 28856 24822
rect 28920 24614 28948 25230
rect 28908 24608 28960 24614
rect 28908 24550 28960 24556
rect 29012 24138 29040 26182
rect 29104 24818 29132 26250
rect 29092 24812 29144 24818
rect 29092 24754 29144 24760
rect 29000 24132 29052 24138
rect 29000 24074 29052 24080
rect 29288 23866 29316 28018
rect 30012 27872 30064 27878
rect 30012 27814 30064 27820
rect 29736 27464 29788 27470
rect 29736 27406 29788 27412
rect 29748 26926 29776 27406
rect 30024 26994 30052 27814
rect 30012 26988 30064 26994
rect 30012 26930 30064 26936
rect 29736 26920 29788 26926
rect 29736 26862 29788 26868
rect 29920 26920 29972 26926
rect 29920 26862 29972 26868
rect 29932 26042 29960 26862
rect 29920 26036 29972 26042
rect 29920 25978 29972 25984
rect 30104 25288 30156 25294
rect 30104 25230 30156 25236
rect 30116 24750 30144 25230
rect 30104 24744 30156 24750
rect 30104 24686 30156 24692
rect 30116 23866 30144 24686
rect 29276 23860 29328 23866
rect 29276 23802 29328 23808
rect 30104 23860 30156 23866
rect 30104 23802 30156 23808
rect 28816 23588 28868 23594
rect 28816 23530 28868 23536
rect 29920 22094 29972 22098
rect 30208 22094 30236 32166
rect 30493 32124 30801 32133
rect 30493 32122 30499 32124
rect 30555 32122 30579 32124
rect 30635 32122 30659 32124
rect 30715 32122 30739 32124
rect 30795 32122 30801 32124
rect 30555 32070 30557 32122
rect 30737 32070 30739 32122
rect 30493 32068 30499 32070
rect 30555 32068 30579 32070
rect 30635 32068 30659 32070
rect 30715 32068 30739 32070
rect 30795 32068 30801 32070
rect 30493 32059 30801 32068
rect 30493 31036 30801 31045
rect 30493 31034 30499 31036
rect 30555 31034 30579 31036
rect 30635 31034 30659 31036
rect 30715 31034 30739 31036
rect 30795 31034 30801 31036
rect 30555 30982 30557 31034
rect 30737 30982 30739 31034
rect 30493 30980 30499 30982
rect 30555 30980 30579 30982
rect 30635 30980 30659 30982
rect 30715 30980 30739 30982
rect 30795 30980 30801 30982
rect 30493 30971 30801 30980
rect 30493 29948 30801 29957
rect 30493 29946 30499 29948
rect 30555 29946 30579 29948
rect 30635 29946 30659 29948
rect 30715 29946 30739 29948
rect 30795 29946 30801 29948
rect 30555 29894 30557 29946
rect 30737 29894 30739 29946
rect 30493 29892 30499 29894
rect 30555 29892 30579 29894
rect 30635 29892 30659 29894
rect 30715 29892 30739 29894
rect 30795 29892 30801 29894
rect 30493 29883 30801 29892
rect 30288 29028 30340 29034
rect 30288 28970 30340 28976
rect 30300 28082 30328 28970
rect 30493 28860 30801 28869
rect 30493 28858 30499 28860
rect 30555 28858 30579 28860
rect 30635 28858 30659 28860
rect 30715 28858 30739 28860
rect 30795 28858 30801 28860
rect 30555 28806 30557 28858
rect 30737 28806 30739 28858
rect 30493 28804 30499 28806
rect 30555 28804 30579 28806
rect 30635 28804 30659 28806
rect 30715 28804 30739 28806
rect 30795 28804 30801 28806
rect 30493 28795 30801 28804
rect 30288 28076 30340 28082
rect 30288 28018 30340 28024
rect 32312 28076 32364 28082
rect 32312 28018 32364 28024
rect 30300 27130 30328 28018
rect 30493 27772 30801 27781
rect 30493 27770 30499 27772
rect 30555 27770 30579 27772
rect 30635 27770 30659 27772
rect 30715 27770 30739 27772
rect 30795 27770 30801 27772
rect 30555 27718 30557 27770
rect 30737 27718 30739 27770
rect 30493 27716 30499 27718
rect 30555 27716 30579 27718
rect 30635 27716 30659 27718
rect 30715 27716 30739 27718
rect 30795 27716 30801 27718
rect 30493 27707 30801 27716
rect 30288 27124 30340 27130
rect 30288 27066 30340 27072
rect 30493 26684 30801 26693
rect 30493 26682 30499 26684
rect 30555 26682 30579 26684
rect 30635 26682 30659 26684
rect 30715 26682 30739 26684
rect 30795 26682 30801 26684
rect 30555 26630 30557 26682
rect 30737 26630 30739 26682
rect 30493 26628 30499 26630
rect 30555 26628 30579 26630
rect 30635 26628 30659 26630
rect 30715 26628 30739 26630
rect 30795 26628 30801 26630
rect 30493 26619 30801 26628
rect 32324 25906 32352 28018
rect 32312 25900 32364 25906
rect 32312 25842 32364 25848
rect 32404 25900 32456 25906
rect 32404 25842 32456 25848
rect 30493 25596 30801 25605
rect 30493 25594 30499 25596
rect 30555 25594 30579 25596
rect 30635 25594 30659 25596
rect 30715 25594 30739 25596
rect 30795 25594 30801 25596
rect 30555 25542 30557 25594
rect 30737 25542 30739 25594
rect 30493 25540 30499 25542
rect 30555 25540 30579 25542
rect 30635 25540 30659 25542
rect 30715 25540 30739 25542
rect 30795 25540 30801 25542
rect 30493 25531 30801 25540
rect 30380 24812 30432 24818
rect 30380 24754 30432 24760
rect 30392 24410 30420 24754
rect 31484 24608 31536 24614
rect 31484 24550 31536 24556
rect 30493 24508 30801 24517
rect 30493 24506 30499 24508
rect 30555 24506 30579 24508
rect 30635 24506 30659 24508
rect 30715 24506 30739 24508
rect 30795 24506 30801 24508
rect 30555 24454 30557 24506
rect 30737 24454 30739 24506
rect 30493 24452 30499 24454
rect 30555 24452 30579 24454
rect 30635 24452 30659 24454
rect 30715 24452 30739 24454
rect 30795 24452 30801 24454
rect 30493 24443 30801 24452
rect 30380 24404 30432 24410
rect 30380 24346 30432 24352
rect 30840 24200 30892 24206
rect 30840 24142 30892 24148
rect 30493 23420 30801 23429
rect 30493 23418 30499 23420
rect 30555 23418 30579 23420
rect 30635 23418 30659 23420
rect 30715 23418 30739 23420
rect 30795 23418 30801 23420
rect 30555 23366 30557 23418
rect 30737 23366 30739 23418
rect 30493 23364 30499 23366
rect 30555 23364 30579 23366
rect 30635 23364 30659 23366
rect 30715 23364 30739 23366
rect 30795 23364 30801 23366
rect 30493 23355 30801 23364
rect 30380 22432 30432 22438
rect 30380 22374 30432 22380
rect 30392 22166 30420 22374
rect 30493 22332 30801 22341
rect 30493 22330 30499 22332
rect 30555 22330 30579 22332
rect 30635 22330 30659 22332
rect 30715 22330 30739 22332
rect 30795 22330 30801 22332
rect 30555 22278 30557 22330
rect 30737 22278 30739 22330
rect 30493 22276 30499 22278
rect 30555 22276 30579 22278
rect 30635 22276 30659 22278
rect 30715 22276 30739 22278
rect 30795 22276 30801 22278
rect 30493 22267 30801 22276
rect 30380 22160 30432 22166
rect 30432 22108 30512 22114
rect 30380 22102 30512 22108
rect 29920 22092 30236 22094
rect 29972 22066 30236 22092
rect 30392 22086 30512 22102
rect 29920 22034 29972 22040
rect 30380 21956 30432 21962
rect 30380 21898 30432 21904
rect 29736 21888 29788 21894
rect 29736 21830 29788 21836
rect 29748 21554 29776 21830
rect 30392 21690 30420 21898
rect 30380 21684 30432 21690
rect 30380 21626 30432 21632
rect 30484 21622 30512 22086
rect 30852 22094 30880 24142
rect 31496 24070 31524 24550
rect 32324 24274 32352 25842
rect 32416 25498 32444 25842
rect 32496 25832 32548 25838
rect 32496 25774 32548 25780
rect 32404 25492 32456 25498
rect 32404 25434 32456 25440
rect 32312 24268 32364 24274
rect 32312 24210 32364 24216
rect 31484 24064 31536 24070
rect 31484 24006 31536 24012
rect 31760 23112 31812 23118
rect 31760 23054 31812 23060
rect 32036 23112 32088 23118
rect 32036 23054 32088 23060
rect 32404 23112 32456 23118
rect 32404 23054 32456 23060
rect 31300 23044 31352 23050
rect 31300 22986 31352 22992
rect 31116 22976 31168 22982
rect 31116 22918 31168 22924
rect 31128 22778 31156 22918
rect 31116 22772 31168 22778
rect 31116 22714 31168 22720
rect 31312 22574 31340 22986
rect 31392 22636 31444 22642
rect 31392 22578 31444 22584
rect 31300 22568 31352 22574
rect 31300 22510 31352 22516
rect 30852 22066 30972 22094
rect 30472 21616 30524 21622
rect 30472 21558 30524 21564
rect 29736 21548 29788 21554
rect 29736 21490 29788 21496
rect 30493 21244 30801 21253
rect 30493 21242 30499 21244
rect 30555 21242 30579 21244
rect 30635 21242 30659 21244
rect 30715 21242 30739 21244
rect 30795 21242 30801 21244
rect 30555 21190 30557 21242
rect 30737 21190 30739 21242
rect 30493 21188 30499 21190
rect 30555 21188 30579 21190
rect 30635 21188 30659 21190
rect 30715 21188 30739 21190
rect 30795 21188 30801 21190
rect 30493 21179 30801 21188
rect 30944 21146 30972 22066
rect 31404 22030 31432 22578
rect 31484 22500 31536 22506
rect 31484 22442 31536 22448
rect 31024 22024 31076 22030
rect 31024 21966 31076 21972
rect 31392 22024 31444 22030
rect 31392 21966 31444 21972
rect 31036 21622 31064 21966
rect 31404 21622 31432 21966
rect 31024 21616 31076 21622
rect 31024 21558 31076 21564
rect 31392 21616 31444 21622
rect 31392 21558 31444 21564
rect 31496 21554 31524 22442
rect 31576 22024 31628 22030
rect 31576 21966 31628 21972
rect 31484 21548 31536 21554
rect 31484 21490 31536 21496
rect 31496 21146 31524 21490
rect 30932 21140 30984 21146
rect 30932 21082 30984 21088
rect 31484 21140 31536 21146
rect 31484 21082 31536 21088
rect 28724 20936 28776 20942
rect 28724 20878 28776 20884
rect 29092 20868 29144 20874
rect 29092 20810 29144 20816
rect 28816 19848 28868 19854
rect 28816 19790 28868 19796
rect 28908 19848 28960 19854
rect 28908 19790 28960 19796
rect 28724 19780 28776 19786
rect 28724 19722 28776 19728
rect 28736 19310 28764 19722
rect 28724 19304 28776 19310
rect 28724 19246 28776 19252
rect 28264 18964 28316 18970
rect 28264 18906 28316 18912
rect 28736 18834 28764 19246
rect 28724 18828 28776 18834
rect 28724 18770 28776 18776
rect 28828 18766 28856 19790
rect 28920 18834 28948 19790
rect 29104 19378 29132 20810
rect 31588 20602 31616 21966
rect 31772 21690 31800 23054
rect 32048 22778 32076 23054
rect 32036 22772 32088 22778
rect 32036 22714 32088 22720
rect 32416 22574 32444 23054
rect 32404 22568 32456 22574
rect 32404 22510 32456 22516
rect 32416 22030 32444 22510
rect 32404 22024 32456 22030
rect 32404 21966 32456 21972
rect 31760 21684 31812 21690
rect 31760 21626 31812 21632
rect 32416 21146 32444 21966
rect 32404 21140 32456 21146
rect 32404 21082 32456 21088
rect 32508 21078 32536 25774
rect 32772 25696 32824 25702
rect 32772 25638 32824 25644
rect 32784 25294 32812 25638
rect 32772 25288 32824 25294
rect 32772 25230 32824 25236
rect 32680 23180 32732 23186
rect 32680 23122 32732 23128
rect 33140 23180 33192 23186
rect 33140 23122 33192 23128
rect 32692 22642 32720 23122
rect 33152 22710 33180 23122
rect 33244 22982 33272 32166
rect 34713 31580 35021 31589
rect 34713 31578 34719 31580
rect 34775 31578 34799 31580
rect 34855 31578 34879 31580
rect 34935 31578 34959 31580
rect 35015 31578 35021 31580
rect 34775 31526 34777 31578
rect 34957 31526 34959 31578
rect 34713 31524 34719 31526
rect 34775 31524 34799 31526
rect 34855 31524 34879 31526
rect 34935 31524 34959 31526
rect 35015 31524 35021 31526
rect 34713 31515 35021 31524
rect 34713 30492 35021 30501
rect 34713 30490 34719 30492
rect 34775 30490 34799 30492
rect 34855 30490 34879 30492
rect 34935 30490 34959 30492
rect 35015 30490 35021 30492
rect 34775 30438 34777 30490
rect 34957 30438 34959 30490
rect 34713 30436 34719 30438
rect 34775 30436 34799 30438
rect 34855 30436 34879 30438
rect 34935 30436 34959 30438
rect 35015 30436 35021 30438
rect 34713 30427 35021 30436
rect 34713 29404 35021 29413
rect 34713 29402 34719 29404
rect 34775 29402 34799 29404
rect 34855 29402 34879 29404
rect 34935 29402 34959 29404
rect 35015 29402 35021 29404
rect 34775 29350 34777 29402
rect 34957 29350 34959 29402
rect 34713 29348 34719 29350
rect 34775 29348 34799 29350
rect 34855 29348 34879 29350
rect 34935 29348 34959 29350
rect 35015 29348 35021 29350
rect 34713 29339 35021 29348
rect 34713 28316 35021 28325
rect 34713 28314 34719 28316
rect 34775 28314 34799 28316
rect 34855 28314 34879 28316
rect 34935 28314 34959 28316
rect 35015 28314 35021 28316
rect 34775 28262 34777 28314
rect 34957 28262 34959 28314
rect 34713 28260 34719 28262
rect 34775 28260 34799 28262
rect 34855 28260 34879 28262
rect 34935 28260 34959 28262
rect 35015 28260 35021 28262
rect 34713 28251 35021 28260
rect 34713 27228 35021 27237
rect 34713 27226 34719 27228
rect 34775 27226 34799 27228
rect 34855 27226 34879 27228
rect 34935 27226 34959 27228
rect 35015 27226 35021 27228
rect 34775 27174 34777 27226
rect 34957 27174 34959 27226
rect 34713 27172 34719 27174
rect 34775 27172 34799 27174
rect 34855 27172 34879 27174
rect 34935 27172 34959 27174
rect 35015 27172 35021 27174
rect 34713 27163 35021 27172
rect 34713 26140 35021 26149
rect 34713 26138 34719 26140
rect 34775 26138 34799 26140
rect 34855 26138 34879 26140
rect 34935 26138 34959 26140
rect 35015 26138 35021 26140
rect 34775 26086 34777 26138
rect 34957 26086 34959 26138
rect 34713 26084 34719 26086
rect 34775 26084 34799 26086
rect 34855 26084 34879 26086
rect 34935 26084 34959 26086
rect 35015 26084 35021 26086
rect 34713 26075 35021 26084
rect 34713 25052 35021 25061
rect 34713 25050 34719 25052
rect 34775 25050 34799 25052
rect 34855 25050 34879 25052
rect 34935 25050 34959 25052
rect 35015 25050 35021 25052
rect 34775 24998 34777 25050
rect 34957 24998 34959 25050
rect 34713 24996 34719 24998
rect 34775 24996 34799 24998
rect 34855 24996 34879 24998
rect 34935 24996 34959 24998
rect 35015 24996 35021 24998
rect 34713 24987 35021 24996
rect 34713 23964 35021 23973
rect 34713 23962 34719 23964
rect 34775 23962 34799 23964
rect 34855 23962 34879 23964
rect 34935 23962 34959 23964
rect 35015 23962 35021 23964
rect 34775 23910 34777 23962
rect 34957 23910 34959 23962
rect 34713 23908 34719 23910
rect 34775 23908 34799 23910
rect 34855 23908 34879 23910
rect 34935 23908 34959 23910
rect 35015 23908 35021 23910
rect 34713 23899 35021 23908
rect 33324 23112 33376 23118
rect 33324 23054 33376 23060
rect 33232 22976 33284 22982
rect 33232 22918 33284 22924
rect 33140 22704 33192 22710
rect 33140 22646 33192 22652
rect 32680 22636 32732 22642
rect 32680 22578 32732 22584
rect 32588 22024 32640 22030
rect 32588 21966 32640 21972
rect 32600 21554 32628 21966
rect 32588 21548 32640 21554
rect 32588 21490 32640 21496
rect 32496 21072 32548 21078
rect 32496 21014 32548 21020
rect 32220 20936 32272 20942
rect 32220 20878 32272 20884
rect 32312 20936 32364 20942
rect 32312 20878 32364 20884
rect 32232 20806 32260 20878
rect 32220 20800 32272 20806
rect 32220 20742 32272 20748
rect 31576 20596 31628 20602
rect 31576 20538 31628 20544
rect 32324 20482 32352 20878
rect 32404 20800 32456 20806
rect 32404 20742 32456 20748
rect 32232 20454 32352 20482
rect 31944 20392 31996 20398
rect 31944 20334 31996 20340
rect 30493 20156 30801 20165
rect 30493 20154 30499 20156
rect 30555 20154 30579 20156
rect 30635 20154 30659 20156
rect 30715 20154 30739 20156
rect 30795 20154 30801 20156
rect 30555 20102 30557 20154
rect 30737 20102 30739 20154
rect 30493 20100 30499 20102
rect 30555 20100 30579 20102
rect 30635 20100 30659 20102
rect 30715 20100 30739 20102
rect 30795 20100 30801 20102
rect 30493 20091 30801 20100
rect 31956 19854 31984 20334
rect 32232 19854 32260 20454
rect 32312 20324 32364 20330
rect 32312 20266 32364 20272
rect 32324 19990 32352 20266
rect 32312 19984 32364 19990
rect 32312 19926 32364 19932
rect 32416 19854 32444 20742
rect 32600 20602 32628 21490
rect 32588 20596 32640 20602
rect 32588 20538 32640 20544
rect 32588 20460 32640 20466
rect 32588 20402 32640 20408
rect 32600 19854 32628 20402
rect 31760 19848 31812 19854
rect 31760 19790 31812 19796
rect 31944 19848 31996 19854
rect 31944 19790 31996 19796
rect 32220 19848 32272 19854
rect 32220 19790 32272 19796
rect 32404 19848 32456 19854
rect 32404 19790 32456 19796
rect 32588 19848 32640 19854
rect 32588 19790 32640 19796
rect 29092 19372 29144 19378
rect 29092 19314 29144 19320
rect 29736 19372 29788 19378
rect 29736 19314 29788 19320
rect 31208 19372 31260 19378
rect 31208 19314 31260 19320
rect 29104 18834 29132 19314
rect 28908 18828 28960 18834
rect 28908 18770 28960 18776
rect 29092 18828 29144 18834
rect 29092 18770 29144 18776
rect 28816 18760 28868 18766
rect 28816 18702 28868 18708
rect 29748 18748 29776 19314
rect 30493 19068 30801 19077
rect 30493 19066 30499 19068
rect 30555 19066 30579 19068
rect 30635 19066 30659 19068
rect 30715 19066 30739 19068
rect 30795 19066 30801 19068
rect 30555 19014 30557 19066
rect 30737 19014 30739 19066
rect 30493 19012 30499 19014
rect 30555 19012 30579 19014
rect 30635 19012 30659 19014
rect 30715 19012 30739 19014
rect 30795 19012 30801 19014
rect 30493 19003 30801 19012
rect 29828 18760 29880 18766
rect 29748 18720 29828 18748
rect 28828 18290 28856 18702
rect 29460 18692 29512 18698
rect 29460 18634 29512 18640
rect 29092 18352 29144 18358
rect 29092 18294 29144 18300
rect 28172 18284 28224 18290
rect 28172 18226 28224 18232
rect 28540 18284 28592 18290
rect 28540 18226 28592 18232
rect 28816 18284 28868 18290
rect 28816 18226 28868 18232
rect 28092 18142 28304 18170
rect 27988 17876 28040 17882
rect 27988 17818 28040 17824
rect 26148 17604 26200 17610
rect 26148 17546 26200 17552
rect 27804 17604 27856 17610
rect 27804 17546 27856 17552
rect 25688 17332 25740 17338
rect 25688 17274 25740 17280
rect 25964 17264 26016 17270
rect 25964 17206 26016 17212
rect 25504 17196 25556 17202
rect 25504 17138 25556 17144
rect 25516 12782 25544 17138
rect 25780 16788 25832 16794
rect 25780 16730 25832 16736
rect 25792 16114 25820 16730
rect 25872 16516 25924 16522
rect 25872 16458 25924 16464
rect 25884 16250 25912 16458
rect 25872 16244 25924 16250
rect 25872 16186 25924 16192
rect 25780 16108 25832 16114
rect 25780 16050 25832 16056
rect 25792 15434 25820 16050
rect 25780 15428 25832 15434
rect 25780 15370 25832 15376
rect 25976 15366 26004 17206
rect 26160 16522 26188 17546
rect 26272 17436 26580 17445
rect 26272 17434 26278 17436
rect 26334 17434 26358 17436
rect 26414 17434 26438 17436
rect 26494 17434 26518 17436
rect 26574 17434 26580 17436
rect 26334 17382 26336 17434
rect 26516 17382 26518 17434
rect 26272 17380 26278 17382
rect 26334 17380 26358 17382
rect 26414 17380 26438 17382
rect 26494 17380 26518 17382
rect 26574 17380 26580 17382
rect 26272 17371 26580 17380
rect 26148 16516 26200 16522
rect 26148 16458 26200 16464
rect 26056 16448 26108 16454
rect 26056 16390 26108 16396
rect 26068 16182 26096 16390
rect 26056 16176 26108 16182
rect 26056 16118 26108 16124
rect 26056 15700 26108 15706
rect 26056 15642 26108 15648
rect 25964 15360 26016 15366
rect 25964 15302 26016 15308
rect 25976 14618 26004 15302
rect 25964 14612 26016 14618
rect 25964 14554 26016 14560
rect 26068 13326 26096 15642
rect 26160 15094 26188 16458
rect 26272 16348 26580 16357
rect 26272 16346 26278 16348
rect 26334 16346 26358 16348
rect 26414 16346 26438 16348
rect 26494 16346 26518 16348
rect 26574 16346 26580 16348
rect 26334 16294 26336 16346
rect 26516 16294 26518 16346
rect 26272 16292 26278 16294
rect 26334 16292 26358 16294
rect 26414 16292 26438 16294
rect 26494 16292 26518 16294
rect 26574 16292 26580 16294
rect 26272 16283 26580 16292
rect 27816 16046 27844 17546
rect 27712 16040 27764 16046
rect 27712 15982 27764 15988
rect 27804 16040 27856 16046
rect 27804 15982 27856 15988
rect 26272 15260 26580 15269
rect 26272 15258 26278 15260
rect 26334 15258 26358 15260
rect 26414 15258 26438 15260
rect 26494 15258 26518 15260
rect 26574 15258 26580 15260
rect 26334 15206 26336 15258
rect 26516 15206 26518 15258
rect 26272 15204 26278 15206
rect 26334 15204 26358 15206
rect 26414 15204 26438 15206
rect 26494 15204 26518 15206
rect 26574 15204 26580 15206
rect 26272 15195 26580 15204
rect 26148 15088 26200 15094
rect 26148 15030 26200 15036
rect 26424 14952 26476 14958
rect 26424 14894 26476 14900
rect 26436 14414 26464 14894
rect 26700 14612 26752 14618
rect 26700 14554 26752 14560
rect 26424 14408 26476 14414
rect 26424 14350 26476 14356
rect 26712 14346 26740 14554
rect 27724 14414 27752 15982
rect 26976 14408 27028 14414
rect 26976 14350 27028 14356
rect 27712 14408 27764 14414
rect 27712 14350 27764 14356
rect 26700 14340 26752 14346
rect 26700 14282 26752 14288
rect 26272 14172 26580 14181
rect 26272 14170 26278 14172
rect 26334 14170 26358 14172
rect 26414 14170 26438 14172
rect 26494 14170 26518 14172
rect 26574 14170 26580 14172
rect 26334 14118 26336 14170
rect 26516 14118 26518 14170
rect 26272 14116 26278 14118
rect 26334 14116 26358 14118
rect 26414 14116 26438 14118
rect 26494 14116 26518 14118
rect 26574 14116 26580 14118
rect 26272 14107 26580 14116
rect 26700 13864 26752 13870
rect 26700 13806 26752 13812
rect 26056 13320 26108 13326
rect 26056 13262 26108 13268
rect 26272 13084 26580 13093
rect 26272 13082 26278 13084
rect 26334 13082 26358 13084
rect 26414 13082 26438 13084
rect 26494 13082 26518 13084
rect 26574 13082 26580 13084
rect 26334 13030 26336 13082
rect 26516 13030 26518 13082
rect 26272 13028 26278 13030
rect 26334 13028 26358 13030
rect 26414 13028 26438 13030
rect 26494 13028 26518 13030
rect 26574 13028 26580 13030
rect 26272 13019 26580 13028
rect 26608 12844 26660 12850
rect 26608 12786 26660 12792
rect 25504 12776 25556 12782
rect 25504 12718 25556 12724
rect 26272 11996 26580 12005
rect 26272 11994 26278 11996
rect 26334 11994 26358 11996
rect 26414 11994 26438 11996
rect 26494 11994 26518 11996
rect 26574 11994 26580 11996
rect 26334 11942 26336 11994
rect 26516 11942 26518 11994
rect 26272 11940 26278 11942
rect 26334 11940 26358 11942
rect 26414 11940 26438 11942
rect 26494 11940 26518 11942
rect 26574 11940 26580 11942
rect 26272 11931 26580 11940
rect 26056 11552 26108 11558
rect 26056 11494 26108 11500
rect 26068 11150 26096 11494
rect 26620 11150 26648 12786
rect 25872 11144 25924 11150
rect 25872 11086 25924 11092
rect 26056 11144 26108 11150
rect 26056 11086 26108 11092
rect 26608 11144 26660 11150
rect 26608 11086 26660 11092
rect 25884 10810 25912 11086
rect 26608 11008 26660 11014
rect 26608 10950 26660 10956
rect 26272 10908 26580 10917
rect 26272 10906 26278 10908
rect 26334 10906 26358 10908
rect 26414 10906 26438 10908
rect 26494 10906 26518 10908
rect 26574 10906 26580 10908
rect 26334 10854 26336 10906
rect 26516 10854 26518 10906
rect 26272 10852 26278 10854
rect 26334 10852 26358 10854
rect 26414 10852 26438 10854
rect 26494 10852 26518 10854
rect 26574 10852 26580 10854
rect 26272 10843 26580 10852
rect 25872 10804 25924 10810
rect 25872 10746 25924 10752
rect 25412 10260 25464 10266
rect 25412 10202 25464 10208
rect 25320 10056 25372 10062
rect 25320 9998 25372 10004
rect 25884 9994 25912 10746
rect 26620 10062 26648 10950
rect 26608 10056 26660 10062
rect 26608 9998 26660 10004
rect 25228 9988 25280 9994
rect 25228 9930 25280 9936
rect 25872 9988 25924 9994
rect 25872 9930 25924 9936
rect 25240 8634 25268 9930
rect 26272 9820 26580 9829
rect 26272 9818 26278 9820
rect 26334 9818 26358 9820
rect 26414 9818 26438 9820
rect 26494 9818 26518 9820
rect 26574 9818 26580 9820
rect 26334 9766 26336 9818
rect 26516 9766 26518 9818
rect 26272 9764 26278 9766
rect 26334 9764 26358 9766
rect 26414 9764 26438 9766
rect 26494 9764 26518 9766
rect 26574 9764 26580 9766
rect 26272 9755 26580 9764
rect 25964 9580 26016 9586
rect 25964 9522 26016 9528
rect 25228 8628 25280 8634
rect 25228 8570 25280 8576
rect 25872 8628 25924 8634
rect 25872 8570 25924 8576
rect 25136 7948 25188 7954
rect 25136 7890 25188 7896
rect 25044 7472 25096 7478
rect 25044 7414 25096 7420
rect 25056 6730 25084 7414
rect 25148 7410 25176 7890
rect 25136 7404 25188 7410
rect 25136 7346 25188 7352
rect 25596 7200 25648 7206
rect 25596 7142 25648 7148
rect 23480 6724 23532 6730
rect 23480 6666 23532 6672
rect 24952 6724 25004 6730
rect 24952 6666 25004 6672
rect 25044 6724 25096 6730
rect 25044 6666 25096 6672
rect 23492 6186 23520 6666
rect 23572 6656 23624 6662
rect 23572 6598 23624 6604
rect 23584 6390 23612 6598
rect 23572 6384 23624 6390
rect 23572 6326 23624 6332
rect 23480 6180 23532 6186
rect 23480 6122 23532 6128
rect 24676 6112 24728 6118
rect 24676 6054 24728 6060
rect 24688 5710 24716 6054
rect 25608 5710 25636 7142
rect 25884 6662 25912 8570
rect 25976 7546 26004 9522
rect 26712 9178 26740 13806
rect 26988 13530 27016 14350
rect 27620 14340 27672 14346
rect 27620 14282 27672 14288
rect 27632 14006 27660 14282
rect 27712 14272 27764 14278
rect 27712 14214 27764 14220
rect 27620 14000 27672 14006
rect 27620 13942 27672 13948
rect 26976 13524 27028 13530
rect 26976 13466 27028 13472
rect 27724 12986 27752 14214
rect 27816 14074 27844 15982
rect 27804 14068 27856 14074
rect 27804 14010 27856 14016
rect 27816 13977 27844 14010
rect 27802 13968 27858 13977
rect 27802 13903 27804 13912
rect 27856 13903 27858 13912
rect 27804 13874 27856 13880
rect 27712 12980 27764 12986
rect 27712 12922 27764 12928
rect 27804 12912 27856 12918
rect 27804 12854 27856 12860
rect 27344 11688 27396 11694
rect 27344 11630 27396 11636
rect 26792 11144 26844 11150
rect 26792 11086 26844 11092
rect 26700 9172 26752 9178
rect 26700 9114 26752 9120
rect 26804 9110 26832 11086
rect 27356 10606 27384 11630
rect 27344 10600 27396 10606
rect 27344 10542 27396 10548
rect 27356 10266 27384 10542
rect 27344 10260 27396 10266
rect 27344 10202 27396 10208
rect 26792 9104 26844 9110
rect 26792 9046 26844 9052
rect 26272 8732 26580 8741
rect 26272 8730 26278 8732
rect 26334 8730 26358 8732
rect 26414 8730 26438 8732
rect 26494 8730 26518 8732
rect 26574 8730 26580 8732
rect 26334 8678 26336 8730
rect 26516 8678 26518 8730
rect 26272 8676 26278 8678
rect 26334 8676 26358 8678
rect 26414 8676 26438 8678
rect 26494 8676 26518 8678
rect 26574 8676 26580 8678
rect 26272 8667 26580 8676
rect 26056 8492 26108 8498
rect 26056 8434 26108 8440
rect 25964 7540 26016 7546
rect 25964 7482 26016 7488
rect 25872 6656 25924 6662
rect 25872 6598 25924 6604
rect 25976 5914 26004 7482
rect 26068 7410 26096 8434
rect 26272 7644 26580 7653
rect 26272 7642 26278 7644
rect 26334 7642 26358 7644
rect 26414 7642 26438 7644
rect 26494 7642 26518 7644
rect 26574 7642 26580 7644
rect 26334 7590 26336 7642
rect 26516 7590 26518 7642
rect 26272 7588 26278 7590
rect 26334 7588 26358 7590
rect 26414 7588 26438 7590
rect 26494 7588 26518 7590
rect 26574 7588 26580 7590
rect 26272 7579 26580 7588
rect 26056 7404 26108 7410
rect 26056 7346 26108 7352
rect 27816 6662 27844 12854
rect 27896 12708 27948 12714
rect 27896 12650 27948 12656
rect 27908 9994 27936 12650
rect 28078 12336 28134 12345
rect 28078 12271 28134 12280
rect 28092 12238 28120 12271
rect 28080 12232 28132 12238
rect 28080 12174 28132 12180
rect 28092 11082 28120 12174
rect 28172 11892 28224 11898
rect 28172 11834 28224 11840
rect 28080 11076 28132 11082
rect 28080 11018 28132 11024
rect 28092 10826 28120 11018
rect 28000 10798 28120 10826
rect 27896 9988 27948 9994
rect 27896 9930 27948 9936
rect 28000 9586 28028 10798
rect 28080 10736 28132 10742
rect 28080 10678 28132 10684
rect 27988 9580 28040 9586
rect 27988 9522 28040 9528
rect 28092 7818 28120 10678
rect 28184 8906 28212 11834
rect 28276 10266 28304 18142
rect 28552 17678 28580 18226
rect 28540 17672 28592 17678
rect 28540 17614 28592 17620
rect 29104 16590 29132 18294
rect 29184 18284 29236 18290
rect 29184 18226 29236 18232
rect 29276 18284 29328 18290
rect 29276 18226 29328 18232
rect 29196 17610 29224 18226
rect 29288 17882 29316 18226
rect 29472 18222 29500 18634
rect 29460 18216 29512 18222
rect 29460 18158 29512 18164
rect 29276 17876 29328 17882
rect 29276 17818 29328 17824
rect 29288 17678 29316 17818
rect 29472 17814 29500 18158
rect 29460 17808 29512 17814
rect 29460 17750 29512 17756
rect 29276 17672 29328 17678
rect 29276 17614 29328 17620
rect 29184 17604 29236 17610
rect 29184 17546 29236 17552
rect 29092 16584 29144 16590
rect 29092 16526 29144 16532
rect 29104 16114 29132 16526
rect 29748 16522 29776 18720
rect 29828 18702 29880 18708
rect 30493 17980 30801 17989
rect 30493 17978 30499 17980
rect 30555 17978 30579 17980
rect 30635 17978 30659 17980
rect 30715 17978 30739 17980
rect 30795 17978 30801 17980
rect 30555 17926 30557 17978
rect 30737 17926 30739 17978
rect 30493 17924 30499 17926
rect 30555 17924 30579 17926
rect 30635 17924 30659 17926
rect 30715 17924 30739 17926
rect 30795 17924 30801 17926
rect 30493 17915 30801 17924
rect 30932 17672 30984 17678
rect 30932 17614 30984 17620
rect 29828 17604 29880 17610
rect 29828 17546 29880 17552
rect 29840 17338 29868 17546
rect 30944 17338 30972 17614
rect 31116 17604 31168 17610
rect 31116 17546 31168 17552
rect 29828 17332 29880 17338
rect 29828 17274 29880 17280
rect 30012 17332 30064 17338
rect 30012 17274 30064 17280
rect 30932 17332 30984 17338
rect 30932 17274 30984 17280
rect 30024 17066 30052 17274
rect 30288 17128 30340 17134
rect 30288 17070 30340 17076
rect 30012 17060 30064 17066
rect 30012 17002 30064 17008
rect 30024 16590 30052 17002
rect 30012 16584 30064 16590
rect 30012 16526 30064 16532
rect 30104 16584 30156 16590
rect 30104 16526 30156 16532
rect 29736 16516 29788 16522
rect 29736 16458 29788 16464
rect 29748 16114 29776 16458
rect 30116 16454 30144 16526
rect 30300 16454 30328 17070
rect 30493 16892 30801 16901
rect 30493 16890 30499 16892
rect 30555 16890 30579 16892
rect 30635 16890 30659 16892
rect 30715 16890 30739 16892
rect 30795 16890 30801 16892
rect 30555 16838 30557 16890
rect 30737 16838 30739 16890
rect 30493 16836 30499 16838
rect 30555 16836 30579 16838
rect 30635 16836 30659 16838
rect 30715 16836 30739 16838
rect 30795 16836 30801 16838
rect 30493 16827 30801 16836
rect 31128 16794 31156 17546
rect 31220 17218 31248 19314
rect 31772 19310 31800 19790
rect 31956 19446 31984 19790
rect 32232 19514 32260 19790
rect 32220 19508 32272 19514
rect 32220 19450 32272 19456
rect 31944 19440 31996 19446
rect 31944 19382 31996 19388
rect 31760 19304 31812 19310
rect 31760 19246 31812 19252
rect 31668 17332 31720 17338
rect 31668 17274 31720 17280
rect 31220 17202 31340 17218
rect 31220 17196 31352 17202
rect 31220 17190 31300 17196
rect 31300 17138 31352 17144
rect 31116 16788 31168 16794
rect 31116 16730 31168 16736
rect 31312 16522 31340 17138
rect 31680 16794 31708 17274
rect 31668 16788 31720 16794
rect 31668 16730 31720 16736
rect 32232 16658 32260 19450
rect 32416 19446 32444 19790
rect 32404 19440 32456 19446
rect 32404 19382 32456 19388
rect 32600 19378 32628 19790
rect 32588 19372 32640 19378
rect 32588 19314 32640 19320
rect 32600 18952 32628 19314
rect 32692 19310 32720 22578
rect 33152 22098 33180 22646
rect 33336 22574 33364 23054
rect 33508 22976 33560 22982
rect 33508 22918 33560 22924
rect 33520 22710 33548 22918
rect 34713 22876 35021 22885
rect 34713 22874 34719 22876
rect 34775 22874 34799 22876
rect 34855 22874 34879 22876
rect 34935 22874 34959 22876
rect 35015 22874 35021 22876
rect 34775 22822 34777 22874
rect 34957 22822 34959 22874
rect 34713 22820 34719 22822
rect 34775 22820 34799 22822
rect 34855 22820 34879 22822
rect 34935 22820 34959 22822
rect 35015 22820 35021 22822
rect 34713 22811 35021 22820
rect 33508 22704 33560 22710
rect 33508 22646 33560 22652
rect 33692 22636 33744 22642
rect 33692 22578 33744 22584
rect 33324 22568 33376 22574
rect 33324 22510 33376 22516
rect 33140 22092 33192 22098
rect 33140 22034 33192 22040
rect 33336 22030 33364 22510
rect 33704 22234 33732 22578
rect 33692 22228 33744 22234
rect 33692 22170 33744 22176
rect 33324 22024 33376 22030
rect 33324 21966 33376 21972
rect 32956 20936 33008 20942
rect 32956 20878 33008 20884
rect 32772 20868 32824 20874
rect 32772 20810 32824 20816
rect 32784 20466 32812 20810
rect 32772 20460 32824 20466
rect 32772 20402 32824 20408
rect 32680 19304 32732 19310
rect 32680 19246 32732 19252
rect 32508 18924 32628 18952
rect 32508 18834 32536 18924
rect 32784 18850 32812 20402
rect 32968 20330 32996 20878
rect 33048 20868 33100 20874
rect 33048 20810 33100 20816
rect 33060 20466 33088 20810
rect 33048 20460 33100 20466
rect 33048 20402 33100 20408
rect 32956 20324 33008 20330
rect 32956 20266 33008 20272
rect 33060 19514 33088 20402
rect 33048 19508 33100 19514
rect 33048 19450 33100 19456
rect 33336 18970 33364 21966
rect 34713 21788 35021 21797
rect 34713 21786 34719 21788
rect 34775 21786 34799 21788
rect 34855 21786 34879 21788
rect 34935 21786 34959 21788
rect 35015 21786 35021 21788
rect 34775 21734 34777 21786
rect 34957 21734 34959 21786
rect 34713 21732 34719 21734
rect 34775 21732 34799 21734
rect 34855 21732 34879 21734
rect 34935 21732 34959 21734
rect 35015 21732 35021 21734
rect 34713 21723 35021 21732
rect 34713 20700 35021 20709
rect 34713 20698 34719 20700
rect 34775 20698 34799 20700
rect 34855 20698 34879 20700
rect 34935 20698 34959 20700
rect 35015 20698 35021 20700
rect 34775 20646 34777 20698
rect 34957 20646 34959 20698
rect 34713 20644 34719 20646
rect 34775 20644 34799 20646
rect 34855 20644 34879 20646
rect 34935 20644 34959 20646
rect 35015 20644 35021 20646
rect 34713 20635 35021 20644
rect 34713 19612 35021 19621
rect 34713 19610 34719 19612
rect 34775 19610 34799 19612
rect 34855 19610 34879 19612
rect 34935 19610 34959 19612
rect 35015 19610 35021 19612
rect 34775 19558 34777 19610
rect 34957 19558 34959 19610
rect 34713 19556 34719 19558
rect 34775 19556 34799 19558
rect 34855 19556 34879 19558
rect 34935 19556 34959 19558
rect 35015 19556 35021 19558
rect 34713 19547 35021 19556
rect 33324 18964 33376 18970
rect 33324 18906 33376 18912
rect 32496 18828 32548 18834
rect 32496 18770 32548 18776
rect 32588 18828 32640 18834
rect 32784 18822 32904 18850
rect 32588 18770 32640 18776
rect 32404 18692 32456 18698
rect 32404 18634 32456 18640
rect 32312 18216 32364 18222
rect 32312 18158 32364 18164
rect 32324 17814 32352 18158
rect 32312 17808 32364 17814
rect 32312 17750 32364 17756
rect 32220 16652 32272 16658
rect 32220 16594 32272 16600
rect 32416 16590 32444 18634
rect 32508 18290 32536 18770
rect 32496 18284 32548 18290
rect 32496 18226 32548 18232
rect 32508 17490 32536 18226
rect 32600 17678 32628 18770
rect 32876 18766 32904 18822
rect 32864 18760 32916 18766
rect 32864 18702 32916 18708
rect 32876 18426 32904 18702
rect 34713 18524 35021 18533
rect 34713 18522 34719 18524
rect 34775 18522 34799 18524
rect 34855 18522 34879 18524
rect 34935 18522 34959 18524
rect 35015 18522 35021 18524
rect 34775 18470 34777 18522
rect 34957 18470 34959 18522
rect 34713 18468 34719 18470
rect 34775 18468 34799 18470
rect 34855 18468 34879 18470
rect 34935 18468 34959 18470
rect 35015 18468 35021 18470
rect 34713 18459 35021 18468
rect 32864 18420 32916 18426
rect 32864 18362 32916 18368
rect 32864 18216 32916 18222
rect 32864 18158 32916 18164
rect 34336 18216 34388 18222
rect 34336 18158 34388 18164
rect 32588 17672 32640 17678
rect 32588 17614 32640 17620
rect 32508 17462 32628 17490
rect 32600 17202 32628 17462
rect 32876 17338 32904 18158
rect 34348 17921 34376 18158
rect 34334 17912 34390 17921
rect 34334 17847 34390 17856
rect 33416 17672 33468 17678
rect 33416 17614 33468 17620
rect 33428 17338 33456 17614
rect 34713 17436 35021 17445
rect 34713 17434 34719 17436
rect 34775 17434 34799 17436
rect 34855 17434 34879 17436
rect 34935 17434 34959 17436
rect 35015 17434 35021 17436
rect 34775 17382 34777 17434
rect 34957 17382 34959 17434
rect 34713 17380 34719 17382
rect 34775 17380 34799 17382
rect 34855 17380 34879 17382
rect 34935 17380 34959 17382
rect 35015 17380 35021 17382
rect 34713 17371 35021 17380
rect 32864 17332 32916 17338
rect 32864 17274 32916 17280
rect 33416 17332 33468 17338
rect 33416 17274 33468 17280
rect 32588 17196 32640 17202
rect 32588 17138 32640 17144
rect 32600 16998 32628 17138
rect 32588 16992 32640 16998
rect 32588 16934 32640 16940
rect 32496 16652 32548 16658
rect 32496 16594 32548 16600
rect 32404 16584 32456 16590
rect 32404 16526 32456 16532
rect 30380 16516 30432 16522
rect 30380 16458 30432 16464
rect 31300 16516 31352 16522
rect 31300 16458 31352 16464
rect 30104 16448 30156 16454
rect 30104 16390 30156 16396
rect 30288 16448 30340 16454
rect 30288 16390 30340 16396
rect 28448 16108 28500 16114
rect 28448 16050 28500 16056
rect 29092 16108 29144 16114
rect 29092 16050 29144 16056
rect 29736 16108 29788 16114
rect 29736 16050 29788 16056
rect 28356 16040 28408 16046
rect 28356 15982 28408 15988
rect 28368 15706 28396 15982
rect 28356 15700 28408 15706
rect 28356 15642 28408 15648
rect 28460 13002 28488 16050
rect 29000 15428 29052 15434
rect 29000 15370 29052 15376
rect 28632 14408 28684 14414
rect 28632 14350 28684 14356
rect 28722 14376 28778 14385
rect 28540 13728 28592 13734
rect 28540 13670 28592 13676
rect 28368 12986 28488 13002
rect 28356 12980 28488 12986
rect 28408 12974 28488 12980
rect 28356 12922 28408 12928
rect 28448 12912 28500 12918
rect 28448 12854 28500 12860
rect 28356 12640 28408 12646
rect 28356 12582 28408 12588
rect 28368 11830 28396 12582
rect 28460 12238 28488 12854
rect 28552 12238 28580 13670
rect 28644 12306 28672 14350
rect 28722 14311 28778 14320
rect 28736 14006 28764 14311
rect 29012 14278 29040 15370
rect 29104 14346 29132 16050
rect 29552 15564 29604 15570
rect 29552 15506 29604 15512
rect 29564 15162 29592 15506
rect 29552 15156 29604 15162
rect 29552 15098 29604 15104
rect 29092 14340 29144 14346
rect 29092 14282 29144 14288
rect 29000 14272 29052 14278
rect 29000 14214 29052 14220
rect 28724 14000 28776 14006
rect 28724 13942 28776 13948
rect 29012 12782 29040 14214
rect 29460 13728 29512 13734
rect 29460 13670 29512 13676
rect 29000 12776 29052 12782
rect 29000 12718 29052 12724
rect 29472 12434 29500 13670
rect 29380 12406 29500 12434
rect 28632 12300 28684 12306
rect 28632 12242 28684 12248
rect 28448 12232 28500 12238
rect 28448 12174 28500 12180
rect 28540 12232 28592 12238
rect 28540 12174 28592 12180
rect 28460 11898 28488 12174
rect 28632 12164 28684 12170
rect 28632 12106 28684 12112
rect 28448 11892 28500 11898
rect 28448 11834 28500 11840
rect 28356 11824 28408 11830
rect 28356 11766 28408 11772
rect 28644 11762 28672 12106
rect 28632 11756 28684 11762
rect 28632 11698 28684 11704
rect 28264 10260 28316 10266
rect 28264 10202 28316 10208
rect 28644 10062 28672 11698
rect 29380 11558 29408 12406
rect 29368 11552 29420 11558
rect 29368 11494 29420 11500
rect 29000 10804 29052 10810
rect 29000 10746 29052 10752
rect 29012 10130 29040 10746
rect 29380 10470 29408 11494
rect 29564 11150 29592 15098
rect 29644 14884 29696 14890
rect 29644 14826 29696 14832
rect 29656 13938 29684 14826
rect 29748 14346 29776 16050
rect 30116 16046 30144 16390
rect 30104 16040 30156 16046
rect 30104 15982 30156 15988
rect 30300 15502 30328 16390
rect 30392 16182 30420 16458
rect 30380 16176 30432 16182
rect 30380 16118 30432 16124
rect 30493 15804 30801 15813
rect 30493 15802 30499 15804
rect 30555 15802 30579 15804
rect 30635 15802 30659 15804
rect 30715 15802 30739 15804
rect 30795 15802 30801 15804
rect 30555 15750 30557 15802
rect 30737 15750 30739 15802
rect 30493 15748 30499 15750
rect 30555 15748 30579 15750
rect 30635 15748 30659 15750
rect 30715 15748 30739 15750
rect 30795 15748 30801 15750
rect 30493 15739 30801 15748
rect 30288 15496 30340 15502
rect 30288 15438 30340 15444
rect 30012 15020 30064 15026
rect 30012 14962 30064 14968
rect 29736 14340 29788 14346
rect 29736 14282 29788 14288
rect 29748 13938 29776 14282
rect 29920 14272 29972 14278
rect 29920 14214 29972 14220
rect 29932 13938 29960 14214
rect 30024 14074 30052 14962
rect 30493 14716 30801 14725
rect 30493 14714 30499 14716
rect 30555 14714 30579 14716
rect 30635 14714 30659 14716
rect 30715 14714 30739 14716
rect 30795 14714 30801 14716
rect 30555 14662 30557 14714
rect 30737 14662 30739 14714
rect 30493 14660 30499 14662
rect 30555 14660 30579 14662
rect 30635 14660 30659 14662
rect 30715 14660 30739 14662
rect 30795 14660 30801 14662
rect 30493 14651 30801 14660
rect 30104 14408 30156 14414
rect 30104 14350 30156 14356
rect 30116 14074 30144 14350
rect 31312 14278 31340 16458
rect 32508 16250 32536 16594
rect 32496 16244 32548 16250
rect 32496 16186 32548 16192
rect 32312 16040 32364 16046
rect 32312 15982 32364 15988
rect 32324 15706 32352 15982
rect 31760 15700 31812 15706
rect 31760 15642 31812 15648
rect 32312 15700 32364 15706
rect 32312 15642 32364 15648
rect 31772 14482 31800 15642
rect 32496 14612 32548 14618
rect 32496 14554 32548 14560
rect 31760 14476 31812 14482
rect 31760 14418 31812 14424
rect 32312 14476 32364 14482
rect 32312 14418 32364 14424
rect 32128 14408 32180 14414
rect 32128 14350 32180 14356
rect 31300 14272 31352 14278
rect 31300 14214 31352 14220
rect 30012 14068 30064 14074
rect 30012 14010 30064 14016
rect 30104 14068 30156 14074
rect 30104 14010 30156 14016
rect 29644 13932 29696 13938
rect 29644 13874 29696 13880
rect 29736 13932 29788 13938
rect 29736 13874 29788 13880
rect 29920 13932 29972 13938
rect 29920 13874 29972 13880
rect 29656 12850 29684 13874
rect 30288 13864 30340 13870
rect 30288 13806 30340 13812
rect 29644 12844 29696 12850
rect 29644 12786 29696 12792
rect 30196 12776 30248 12782
rect 30196 12718 30248 12724
rect 30208 11762 30236 12718
rect 30196 11756 30248 11762
rect 30196 11698 30248 11704
rect 30208 11150 30236 11698
rect 29552 11144 29604 11150
rect 29552 11086 29604 11092
rect 30196 11144 30248 11150
rect 30196 11086 30248 11092
rect 29460 11076 29512 11082
rect 29460 11018 29512 11024
rect 29472 10742 29500 11018
rect 29736 11008 29788 11014
rect 29736 10950 29788 10956
rect 30104 11008 30156 11014
rect 30104 10950 30156 10956
rect 29460 10736 29512 10742
rect 29460 10678 29512 10684
rect 29368 10464 29420 10470
rect 29368 10406 29420 10412
rect 29000 10124 29052 10130
rect 29000 10066 29052 10072
rect 28632 10056 28684 10062
rect 28632 9998 28684 10004
rect 28908 10056 28960 10062
rect 28908 9998 28960 10004
rect 28264 9988 28316 9994
rect 28264 9930 28316 9936
rect 28540 9988 28592 9994
rect 28540 9930 28592 9936
rect 28172 8900 28224 8906
rect 28172 8842 28224 8848
rect 28080 7812 28132 7818
rect 28080 7754 28132 7760
rect 27804 6656 27856 6662
rect 27804 6598 27856 6604
rect 26272 6556 26580 6565
rect 26272 6554 26278 6556
rect 26334 6554 26358 6556
rect 26414 6554 26438 6556
rect 26494 6554 26518 6556
rect 26574 6554 26580 6556
rect 26334 6502 26336 6554
rect 26516 6502 26518 6554
rect 26272 6500 26278 6502
rect 26334 6500 26358 6502
rect 26414 6500 26438 6502
rect 26494 6500 26518 6502
rect 26574 6500 26580 6502
rect 26272 6491 26580 6500
rect 27816 6458 27844 6598
rect 27804 6452 27856 6458
rect 27804 6394 27856 6400
rect 28184 6186 28212 8842
rect 28276 7750 28304 9930
rect 28448 7812 28500 7818
rect 28448 7754 28500 7760
rect 28264 7744 28316 7750
rect 28264 7686 28316 7692
rect 28172 6180 28224 6186
rect 28172 6122 28224 6128
rect 25964 5908 26016 5914
rect 25964 5850 26016 5856
rect 24676 5704 24728 5710
rect 24676 5646 24728 5652
rect 25596 5704 25648 5710
rect 25596 5646 25648 5652
rect 24688 5370 24716 5646
rect 26272 5468 26580 5477
rect 26272 5466 26278 5468
rect 26334 5466 26358 5468
rect 26414 5466 26438 5468
rect 26494 5466 26518 5468
rect 26574 5466 26580 5468
rect 26334 5414 26336 5466
rect 26516 5414 26518 5466
rect 26272 5412 26278 5414
rect 26334 5412 26358 5414
rect 26414 5412 26438 5414
rect 26494 5412 26518 5414
rect 26574 5412 26580 5414
rect 26272 5403 26580 5412
rect 24676 5364 24728 5370
rect 24676 5306 24728 5312
rect 23388 5296 23440 5302
rect 23388 5238 23440 5244
rect 26056 5296 26108 5302
rect 26056 5238 26108 5244
rect 25596 5024 25648 5030
rect 25596 4966 25648 4972
rect 22052 4924 22360 4933
rect 22052 4922 22058 4924
rect 22114 4922 22138 4924
rect 22194 4922 22218 4924
rect 22274 4922 22298 4924
rect 22354 4922 22360 4924
rect 22114 4870 22116 4922
rect 22296 4870 22298 4922
rect 22052 4868 22058 4870
rect 22114 4868 22138 4870
rect 22194 4868 22218 4870
rect 22274 4868 22298 4870
rect 22354 4868 22360 4870
rect 22052 4859 22360 4868
rect 20720 4752 20772 4758
rect 20720 4694 20772 4700
rect 24952 4752 25004 4758
rect 24952 4694 25004 4700
rect 20444 4684 20496 4690
rect 20444 4626 20496 4632
rect 17316 4616 17368 4622
rect 17316 4558 17368 4564
rect 18420 4616 18472 4622
rect 18420 4558 18472 4564
rect 20168 4616 20220 4622
rect 20168 4558 20220 4564
rect 17328 4146 17356 4558
rect 17500 4480 17552 4486
rect 17500 4422 17552 4428
rect 18236 4480 18288 4486
rect 18236 4422 18288 4428
rect 19064 4480 19116 4486
rect 19064 4422 19116 4428
rect 19800 4480 19852 4486
rect 19800 4422 19852 4428
rect 17512 4146 17540 4422
rect 17831 4380 18139 4389
rect 17831 4378 17837 4380
rect 17893 4378 17917 4380
rect 17973 4378 17997 4380
rect 18053 4378 18077 4380
rect 18133 4378 18139 4380
rect 17893 4326 17895 4378
rect 18075 4326 18077 4378
rect 17831 4324 17837 4326
rect 17893 4324 17917 4326
rect 17973 4324 17997 4326
rect 18053 4324 18077 4326
rect 18133 4324 18139 4326
rect 17831 4315 18139 4324
rect 17316 4140 17368 4146
rect 17316 4082 17368 4088
rect 17500 4140 17552 4146
rect 17500 4082 17552 4088
rect 17960 4140 18012 4146
rect 18248 4128 18276 4422
rect 18012 4100 18276 4128
rect 17960 4082 18012 4088
rect 19076 3942 19104 4422
rect 19064 3936 19116 3942
rect 19064 3878 19116 3884
rect 18236 3392 18288 3398
rect 18236 3334 18288 3340
rect 17831 3292 18139 3301
rect 17831 3290 17837 3292
rect 17893 3290 17917 3292
rect 17973 3290 17997 3292
rect 18053 3290 18077 3292
rect 18133 3290 18139 3292
rect 17893 3238 17895 3290
rect 18075 3238 18077 3290
rect 17831 3236 17837 3238
rect 17893 3236 17917 3238
rect 17973 3236 17997 3238
rect 18053 3236 18077 3238
rect 18133 3236 18139 3238
rect 17831 3227 18139 3236
rect 18248 3194 18276 3334
rect 16948 3188 17000 3194
rect 16948 3130 17000 3136
rect 17040 3188 17092 3194
rect 17040 3130 17092 3136
rect 18236 3188 18288 3194
rect 18236 3130 18288 3136
rect 18248 2514 18276 3130
rect 18236 2508 18288 2514
rect 18236 2450 18288 2456
rect 19076 2446 19104 3878
rect 19812 3534 19840 4422
rect 19524 3528 19576 3534
rect 19524 3470 19576 3476
rect 19800 3528 19852 3534
rect 19800 3470 19852 3476
rect 19536 3194 19564 3470
rect 19524 3188 19576 3194
rect 19524 3130 19576 3136
rect 20456 2990 20484 4626
rect 20732 3058 20760 4694
rect 20904 4616 20956 4622
rect 20904 4558 20956 4564
rect 20812 4480 20864 4486
rect 20812 4422 20864 4428
rect 20824 3738 20852 4422
rect 20916 4146 20944 4558
rect 21548 4480 21600 4486
rect 21548 4422 21600 4428
rect 22100 4480 22152 4486
rect 22100 4422 22152 4428
rect 21560 4146 21588 4422
rect 22112 4146 22140 4422
rect 22468 4276 22520 4282
rect 22468 4218 22520 4224
rect 20904 4140 20956 4146
rect 20904 4082 20956 4088
rect 21180 4140 21232 4146
rect 21180 4082 21232 4088
rect 21548 4140 21600 4146
rect 21548 4082 21600 4088
rect 22100 4140 22152 4146
rect 22100 4082 22152 4088
rect 22284 4140 22336 4146
rect 22284 4082 22336 4088
rect 20812 3732 20864 3738
rect 20812 3674 20864 3680
rect 20720 3052 20772 3058
rect 20720 2994 20772 3000
rect 20444 2984 20496 2990
rect 20444 2926 20496 2932
rect 20824 2774 20852 3674
rect 20916 3534 20944 4082
rect 21088 3936 21140 3942
rect 21088 3878 21140 3884
rect 20904 3528 20956 3534
rect 20904 3470 20956 3476
rect 20916 3194 20944 3470
rect 21100 3194 21128 3878
rect 20904 3188 20956 3194
rect 20904 3130 20956 3136
rect 21088 3188 21140 3194
rect 21088 3130 21140 3136
rect 20824 2746 20944 2774
rect 20916 2514 20944 2746
rect 20904 2508 20956 2514
rect 20904 2450 20956 2456
rect 21100 2446 21128 3130
rect 21192 2922 21220 4082
rect 22296 4026 22324 4082
rect 22296 3998 22416 4026
rect 22052 3836 22360 3845
rect 22052 3834 22058 3836
rect 22114 3834 22138 3836
rect 22194 3834 22218 3836
rect 22274 3834 22298 3836
rect 22354 3834 22360 3836
rect 22114 3782 22116 3834
rect 22296 3782 22298 3834
rect 22052 3780 22058 3782
rect 22114 3780 22138 3782
rect 22194 3780 22218 3782
rect 22274 3780 22298 3782
rect 22354 3780 22360 3782
rect 22052 3771 22360 3780
rect 22388 3738 22416 3998
rect 22376 3732 22428 3738
rect 22376 3674 22428 3680
rect 22480 3534 22508 4218
rect 24964 3942 24992 4694
rect 25044 4480 25096 4486
rect 25044 4422 25096 4428
rect 23388 3936 23440 3942
rect 23388 3878 23440 3884
rect 24952 3936 25004 3942
rect 24952 3878 25004 3884
rect 22744 3596 22796 3602
rect 22744 3538 22796 3544
rect 22468 3528 22520 3534
rect 22468 3470 22520 3476
rect 22756 3058 22784 3538
rect 23400 3466 23428 3878
rect 23388 3460 23440 3466
rect 23388 3402 23440 3408
rect 22744 3052 22796 3058
rect 22744 2994 22796 3000
rect 21180 2916 21232 2922
rect 21180 2858 21232 2864
rect 22052 2748 22360 2757
rect 22052 2746 22058 2748
rect 22114 2746 22138 2748
rect 22194 2746 22218 2748
rect 22274 2746 22298 2748
rect 22354 2746 22360 2748
rect 22114 2694 22116 2746
rect 22296 2694 22298 2746
rect 22052 2692 22058 2694
rect 22114 2692 22138 2694
rect 22194 2692 22218 2694
rect 22274 2692 22298 2694
rect 22354 2692 22360 2694
rect 22052 2683 22360 2692
rect 23400 2446 23428 3402
rect 24964 2922 24992 3878
rect 25056 3466 25084 4422
rect 25608 4214 25636 4966
rect 25872 4616 25924 4622
rect 25872 4558 25924 4564
rect 25596 4208 25648 4214
rect 25596 4150 25648 4156
rect 25884 4146 25912 4558
rect 25872 4140 25924 4146
rect 25872 4082 25924 4088
rect 25596 3664 25648 3670
rect 25596 3606 25648 3612
rect 25044 3460 25096 3466
rect 25044 3402 25096 3408
rect 25608 2922 25636 3606
rect 25884 3534 25912 4082
rect 26068 3534 26096 5238
rect 26240 5228 26292 5234
rect 26240 5170 26292 5176
rect 26252 4826 26280 5170
rect 26240 4820 26292 4826
rect 26240 4762 26292 4768
rect 26608 4820 26660 4826
rect 26608 4762 26660 4768
rect 26148 4548 26200 4554
rect 26148 4490 26200 4496
rect 26160 4282 26188 4490
rect 26272 4380 26580 4389
rect 26272 4378 26278 4380
rect 26334 4378 26358 4380
rect 26414 4378 26438 4380
rect 26494 4378 26518 4380
rect 26574 4378 26580 4380
rect 26334 4326 26336 4378
rect 26516 4326 26518 4378
rect 26272 4324 26278 4326
rect 26334 4324 26358 4326
rect 26414 4324 26438 4326
rect 26494 4324 26518 4326
rect 26574 4324 26580 4326
rect 26272 4315 26580 4324
rect 26148 4276 26200 4282
rect 26148 4218 26200 4224
rect 26620 4078 26648 4762
rect 27252 4480 27304 4486
rect 27252 4422 27304 4428
rect 26608 4072 26660 4078
rect 26608 4014 26660 4020
rect 26240 4004 26292 4010
rect 26240 3946 26292 3952
rect 26252 3602 26280 3946
rect 26240 3596 26292 3602
rect 26240 3538 26292 3544
rect 25872 3528 25924 3534
rect 25872 3470 25924 3476
rect 26056 3528 26108 3534
rect 26056 3470 26108 3476
rect 25964 3392 26016 3398
rect 25964 3334 26016 3340
rect 25976 2990 26004 3334
rect 25964 2984 26016 2990
rect 25964 2926 26016 2932
rect 26068 2922 26096 3470
rect 26252 3398 26280 3538
rect 26620 3398 26648 4014
rect 26792 3732 26844 3738
rect 26792 3674 26844 3680
rect 26240 3392 26292 3398
rect 26240 3334 26292 3340
rect 26608 3392 26660 3398
rect 26608 3334 26660 3340
rect 26272 3292 26580 3301
rect 26272 3290 26278 3292
rect 26334 3290 26358 3292
rect 26414 3290 26438 3292
rect 26494 3290 26518 3292
rect 26574 3290 26580 3292
rect 26334 3238 26336 3290
rect 26516 3238 26518 3290
rect 26272 3236 26278 3238
rect 26334 3236 26358 3238
rect 26414 3236 26438 3238
rect 26494 3236 26518 3238
rect 26574 3236 26580 3238
rect 26272 3227 26580 3236
rect 26804 3058 26832 3674
rect 27264 3670 27292 4422
rect 28460 4146 28488 7754
rect 28552 6662 28580 9930
rect 28920 9722 28948 9998
rect 28908 9716 28960 9722
rect 28908 9658 28960 9664
rect 28908 8968 28960 8974
rect 28960 8916 29040 8922
rect 28908 8910 29040 8916
rect 28920 8894 29040 8910
rect 28908 8628 28960 8634
rect 28908 8570 28960 8576
rect 28920 6798 28948 8570
rect 28908 6792 28960 6798
rect 28908 6734 28960 6740
rect 28540 6656 28592 6662
rect 28540 6598 28592 6604
rect 28552 5642 28580 6598
rect 29012 5846 29040 8894
rect 29184 8832 29236 8838
rect 29184 8774 29236 8780
rect 29092 8560 29144 8566
rect 29092 8502 29144 8508
rect 29104 7546 29132 8502
rect 29092 7540 29144 7546
rect 29092 7482 29144 7488
rect 29104 6798 29132 7482
rect 29092 6792 29144 6798
rect 29092 6734 29144 6740
rect 29196 6390 29224 8774
rect 29380 8294 29408 10406
rect 29472 10062 29500 10678
rect 29748 10674 29776 10950
rect 30116 10810 30144 10950
rect 30104 10804 30156 10810
rect 30104 10746 30156 10752
rect 29736 10668 29788 10674
rect 29736 10610 29788 10616
rect 30208 10282 30236 11086
rect 30116 10254 30236 10282
rect 29460 10056 29512 10062
rect 29460 9998 29512 10004
rect 30116 9586 30144 10254
rect 30300 10146 30328 13806
rect 30493 13628 30801 13637
rect 30493 13626 30499 13628
rect 30555 13626 30579 13628
rect 30635 13626 30659 13628
rect 30715 13626 30739 13628
rect 30795 13626 30801 13628
rect 30555 13574 30557 13626
rect 30737 13574 30739 13626
rect 30493 13572 30499 13574
rect 30555 13572 30579 13574
rect 30635 13572 30659 13574
rect 30715 13572 30739 13574
rect 30795 13572 30801 13574
rect 30493 13563 30801 13572
rect 32140 12986 32168 14350
rect 32324 13870 32352 14418
rect 32312 13864 32364 13870
rect 32312 13806 32364 13812
rect 32324 13530 32352 13806
rect 32312 13524 32364 13530
rect 32312 13466 32364 13472
rect 32128 12980 32180 12986
rect 32128 12922 32180 12928
rect 32508 12850 32536 14554
rect 32600 14074 32628 16934
rect 34713 16348 35021 16357
rect 34713 16346 34719 16348
rect 34775 16346 34799 16348
rect 34855 16346 34879 16348
rect 34935 16346 34959 16348
rect 35015 16346 35021 16348
rect 34775 16294 34777 16346
rect 34957 16294 34959 16346
rect 34713 16292 34719 16294
rect 34775 16292 34799 16294
rect 34855 16292 34879 16294
rect 34935 16292 34959 16294
rect 35015 16292 35021 16294
rect 34713 16283 35021 16292
rect 33048 16244 33100 16250
rect 33048 16186 33100 16192
rect 32680 15632 32732 15638
rect 32680 15574 32732 15580
rect 32588 14068 32640 14074
rect 32588 14010 32640 14016
rect 32496 12844 32548 12850
rect 32496 12786 32548 12792
rect 30380 12708 30432 12714
rect 30380 12650 30432 12656
rect 30392 11830 30420 12650
rect 30493 12540 30801 12549
rect 30493 12538 30499 12540
rect 30555 12538 30579 12540
rect 30635 12538 30659 12540
rect 30715 12538 30739 12540
rect 30795 12538 30801 12540
rect 30555 12486 30557 12538
rect 30737 12486 30739 12538
rect 30493 12484 30499 12486
rect 30555 12484 30579 12486
rect 30635 12484 30659 12486
rect 30715 12484 30739 12486
rect 30795 12484 30801 12486
rect 30493 12475 30801 12484
rect 31300 12096 31352 12102
rect 31300 12038 31352 12044
rect 31312 11898 31340 12038
rect 31300 11892 31352 11898
rect 31300 11834 31352 11840
rect 30380 11824 30432 11830
rect 30380 11766 30432 11772
rect 30493 11452 30801 11461
rect 30493 11450 30499 11452
rect 30555 11450 30579 11452
rect 30635 11450 30659 11452
rect 30715 11450 30739 11452
rect 30795 11450 30801 11452
rect 30555 11398 30557 11450
rect 30737 11398 30739 11450
rect 30493 11396 30499 11398
rect 30555 11396 30579 11398
rect 30635 11396 30659 11398
rect 30715 11396 30739 11398
rect 30795 11396 30801 11398
rect 30493 11387 30801 11396
rect 31312 11354 31340 11834
rect 32508 11762 32536 12786
rect 32692 11898 32720 15574
rect 33060 15366 33088 16186
rect 33876 16108 33928 16114
rect 33876 16050 33928 16056
rect 33888 15706 33916 16050
rect 33876 15700 33928 15706
rect 33876 15642 33928 15648
rect 33416 15496 33468 15502
rect 33416 15438 33468 15444
rect 33048 15360 33100 15366
rect 33048 15302 33100 15308
rect 33048 14272 33100 14278
rect 33048 14214 33100 14220
rect 33060 12986 33088 14214
rect 33428 13734 33456 15438
rect 33600 15428 33652 15434
rect 33600 15370 33652 15376
rect 33612 15162 33640 15370
rect 34713 15260 35021 15269
rect 34713 15258 34719 15260
rect 34775 15258 34799 15260
rect 34855 15258 34879 15260
rect 34935 15258 34959 15260
rect 35015 15258 35021 15260
rect 34775 15206 34777 15258
rect 34957 15206 34959 15258
rect 34713 15204 34719 15206
rect 34775 15204 34799 15206
rect 34855 15204 34879 15206
rect 34935 15204 34959 15206
rect 35015 15204 35021 15206
rect 34713 15195 35021 15204
rect 33600 15156 33652 15162
rect 33600 15098 33652 15104
rect 33416 13728 33468 13734
rect 33416 13670 33468 13676
rect 33048 12980 33100 12986
rect 33048 12922 33100 12928
rect 33428 12850 33456 13670
rect 33612 13326 33640 15098
rect 34713 14172 35021 14181
rect 34713 14170 34719 14172
rect 34775 14170 34799 14172
rect 34855 14170 34879 14172
rect 34935 14170 34959 14172
rect 35015 14170 35021 14172
rect 34775 14118 34777 14170
rect 34957 14118 34959 14170
rect 34713 14116 34719 14118
rect 34775 14116 34799 14118
rect 34855 14116 34879 14118
rect 34935 14116 34959 14118
rect 35015 14116 35021 14118
rect 34713 14107 35021 14116
rect 33600 13320 33652 13326
rect 33600 13262 33652 13268
rect 34713 13084 35021 13093
rect 34713 13082 34719 13084
rect 34775 13082 34799 13084
rect 34855 13082 34879 13084
rect 34935 13082 34959 13084
rect 35015 13082 35021 13084
rect 34775 13030 34777 13082
rect 34957 13030 34959 13082
rect 34713 13028 34719 13030
rect 34775 13028 34799 13030
rect 34855 13028 34879 13030
rect 34935 13028 34959 13030
rect 35015 13028 35021 13030
rect 34713 13019 35021 13028
rect 33416 12844 33468 12850
rect 33416 12786 33468 12792
rect 34713 11996 35021 12005
rect 34713 11994 34719 11996
rect 34775 11994 34799 11996
rect 34855 11994 34879 11996
rect 34935 11994 34959 11996
rect 35015 11994 35021 11996
rect 34775 11942 34777 11994
rect 34957 11942 34959 11994
rect 34713 11940 34719 11942
rect 34775 11940 34799 11942
rect 34855 11940 34879 11942
rect 34935 11940 34959 11942
rect 35015 11940 35021 11942
rect 34713 11931 35021 11940
rect 32680 11892 32732 11898
rect 32680 11834 32732 11840
rect 33692 11892 33744 11898
rect 33692 11834 33744 11840
rect 31852 11756 31904 11762
rect 31852 11698 31904 11704
rect 32496 11756 32548 11762
rect 32496 11698 32548 11704
rect 31668 11552 31720 11558
rect 31668 11494 31720 11500
rect 31300 11348 31352 11354
rect 31300 11290 31352 11296
rect 31680 11082 31708 11494
rect 30840 11076 30892 11082
rect 30840 11018 30892 11024
rect 31668 11076 31720 11082
rect 31668 11018 31720 11024
rect 30493 10364 30801 10373
rect 30493 10362 30499 10364
rect 30555 10362 30579 10364
rect 30635 10362 30659 10364
rect 30715 10362 30739 10364
rect 30795 10362 30801 10364
rect 30555 10310 30557 10362
rect 30737 10310 30739 10362
rect 30493 10308 30499 10310
rect 30555 10308 30579 10310
rect 30635 10308 30659 10310
rect 30715 10308 30739 10310
rect 30795 10308 30801 10310
rect 30493 10299 30801 10308
rect 30208 10118 30328 10146
rect 30104 9580 30156 9586
rect 30104 9522 30156 9528
rect 30116 8922 30144 9522
rect 30208 9450 30236 10118
rect 30288 10056 30340 10062
rect 30288 9998 30340 10004
rect 30196 9444 30248 9450
rect 30196 9386 30248 9392
rect 30208 9110 30236 9386
rect 30196 9104 30248 9110
rect 30196 9046 30248 9052
rect 30196 8968 30248 8974
rect 30116 8916 30196 8922
rect 30116 8910 30248 8916
rect 30116 8894 30236 8910
rect 30300 8906 30328 9998
rect 30852 9382 30880 11018
rect 31024 10464 31076 10470
rect 31024 10406 31076 10412
rect 31036 9654 31064 10406
rect 31392 9716 31444 9722
rect 31392 9658 31444 9664
rect 31024 9648 31076 9654
rect 31024 9590 31076 9596
rect 30840 9376 30892 9382
rect 30840 9318 30892 9324
rect 30493 9276 30801 9285
rect 30493 9274 30499 9276
rect 30555 9274 30579 9276
rect 30635 9274 30659 9276
rect 30715 9274 30739 9276
rect 30795 9274 30801 9276
rect 30555 9222 30557 9274
rect 30737 9222 30739 9274
rect 30493 9220 30499 9222
rect 30555 9220 30579 9222
rect 30635 9220 30659 9222
rect 30715 9220 30739 9222
rect 30795 9220 30801 9222
rect 30493 9211 30801 9220
rect 29736 8832 29788 8838
rect 29736 8774 29788 8780
rect 29748 8498 29776 8774
rect 30208 8498 30236 8894
rect 30288 8900 30340 8906
rect 30288 8842 30340 8848
rect 30300 8634 30328 8842
rect 30288 8628 30340 8634
rect 30288 8570 30340 8576
rect 29736 8492 29788 8498
rect 29736 8434 29788 8440
rect 30196 8492 30248 8498
rect 30196 8434 30248 8440
rect 29368 8288 29420 8294
rect 29368 8230 29420 8236
rect 29380 8090 29408 8230
rect 30493 8188 30801 8197
rect 30493 8186 30499 8188
rect 30555 8186 30579 8188
rect 30635 8186 30659 8188
rect 30715 8186 30739 8188
rect 30795 8186 30801 8188
rect 30555 8134 30557 8186
rect 30737 8134 30739 8186
rect 30493 8132 30499 8134
rect 30555 8132 30579 8134
rect 30635 8132 30659 8134
rect 30715 8132 30739 8134
rect 30795 8132 30801 8134
rect 30493 8123 30801 8132
rect 29368 8084 29420 8090
rect 29368 8026 29420 8032
rect 30380 7744 30432 7750
rect 30380 7686 30432 7692
rect 30392 7410 30420 7686
rect 30380 7404 30432 7410
rect 30380 7346 30432 7352
rect 29828 6792 29880 6798
rect 29828 6734 29880 6740
rect 29276 6724 29328 6730
rect 29276 6666 29328 6672
rect 29184 6384 29236 6390
rect 29184 6326 29236 6332
rect 29288 5914 29316 6666
rect 29840 6254 29868 6734
rect 29828 6248 29880 6254
rect 29828 6190 29880 6196
rect 29276 5908 29328 5914
rect 29276 5850 29328 5856
rect 29000 5840 29052 5846
rect 29000 5782 29052 5788
rect 28540 5636 28592 5642
rect 28540 5578 28592 5584
rect 28264 4140 28316 4146
rect 28264 4082 28316 4088
rect 28448 4140 28500 4146
rect 28448 4082 28500 4088
rect 27620 3936 27672 3942
rect 27620 3878 27672 3884
rect 27252 3664 27304 3670
rect 27252 3606 27304 3612
rect 27632 3602 27660 3878
rect 28276 3738 28304 4082
rect 28264 3732 28316 3738
rect 28264 3674 28316 3680
rect 27896 3664 27948 3670
rect 27896 3606 27948 3612
rect 27620 3596 27672 3602
rect 27620 3538 27672 3544
rect 26792 3052 26844 3058
rect 26792 2994 26844 3000
rect 26240 2984 26292 2990
rect 26240 2926 26292 2932
rect 24952 2916 25004 2922
rect 24952 2858 25004 2864
rect 25596 2916 25648 2922
rect 25596 2858 25648 2864
rect 26056 2916 26108 2922
rect 26056 2858 26108 2864
rect 25608 2446 25636 2858
rect 26252 2446 26280 2926
rect 27908 2446 27936 3606
rect 28356 3596 28408 3602
rect 28356 3538 28408 3544
rect 28368 2446 28396 3538
rect 29840 3194 29868 6190
rect 29828 3188 29880 3194
rect 29828 3130 29880 3136
rect 30392 3126 30420 7346
rect 30493 7100 30801 7109
rect 30493 7098 30499 7100
rect 30555 7098 30579 7100
rect 30635 7098 30659 7100
rect 30715 7098 30739 7100
rect 30795 7098 30801 7100
rect 30555 7046 30557 7098
rect 30737 7046 30739 7098
rect 30493 7044 30499 7046
rect 30555 7044 30579 7046
rect 30635 7044 30659 7046
rect 30715 7044 30739 7046
rect 30795 7044 30801 7046
rect 30493 7035 30801 7044
rect 30493 6012 30801 6021
rect 30493 6010 30499 6012
rect 30555 6010 30579 6012
rect 30635 6010 30659 6012
rect 30715 6010 30739 6012
rect 30795 6010 30801 6012
rect 30555 5958 30557 6010
rect 30737 5958 30739 6010
rect 30493 5956 30499 5958
rect 30555 5956 30579 5958
rect 30635 5956 30659 5958
rect 30715 5956 30739 5958
rect 30795 5956 30801 5958
rect 30493 5947 30801 5956
rect 30852 5710 30880 9318
rect 31404 8634 31432 9658
rect 31576 9580 31628 9586
rect 31576 9522 31628 9528
rect 31588 9382 31616 9522
rect 31576 9376 31628 9382
rect 31576 9318 31628 9324
rect 31760 9376 31812 9382
rect 31760 9318 31812 9324
rect 30932 8628 30984 8634
rect 30932 8570 30984 8576
rect 31392 8628 31444 8634
rect 31392 8570 31444 8576
rect 30944 6458 30972 8570
rect 31772 8566 31800 9318
rect 31760 8560 31812 8566
rect 31760 8502 31812 8508
rect 31864 8498 31892 11698
rect 33416 11688 33468 11694
rect 33416 11630 33468 11636
rect 32404 11552 32456 11558
rect 32404 11494 32456 11500
rect 32312 11144 32364 11150
rect 32312 11086 32364 11092
rect 32324 10606 32352 11086
rect 32416 10674 32444 11494
rect 32404 10668 32456 10674
rect 32404 10610 32456 10616
rect 32312 10600 32364 10606
rect 32312 10542 32364 10548
rect 32324 10266 32352 10542
rect 32312 10260 32364 10266
rect 32312 10202 32364 10208
rect 33428 10062 33456 11630
rect 33704 10810 33732 11834
rect 34713 10908 35021 10917
rect 34713 10906 34719 10908
rect 34775 10906 34799 10908
rect 34855 10906 34879 10908
rect 34935 10906 34959 10908
rect 35015 10906 35021 10908
rect 34775 10854 34777 10906
rect 34957 10854 34959 10906
rect 34713 10852 34719 10854
rect 34775 10852 34799 10854
rect 34855 10852 34879 10854
rect 34935 10852 34959 10854
rect 35015 10852 35021 10854
rect 34713 10843 35021 10852
rect 33692 10804 33744 10810
rect 33692 10746 33744 10752
rect 33416 10056 33468 10062
rect 33416 9998 33468 10004
rect 33600 10056 33652 10062
rect 33600 9998 33652 10004
rect 32312 9920 32364 9926
rect 32312 9862 32364 9868
rect 32324 9178 32352 9862
rect 33612 9518 33640 9998
rect 33692 9920 33744 9926
rect 33692 9862 33744 9868
rect 33876 9920 33928 9926
rect 33876 9862 33928 9868
rect 33600 9512 33652 9518
rect 33600 9454 33652 9460
rect 33704 9382 33732 9862
rect 33692 9376 33744 9382
rect 33692 9318 33744 9324
rect 32312 9172 32364 9178
rect 32312 9114 32364 9120
rect 32312 8968 32364 8974
rect 32312 8910 32364 8916
rect 32324 8498 32352 8910
rect 31852 8492 31904 8498
rect 31852 8434 31904 8440
rect 32312 8492 32364 8498
rect 32312 8434 32364 8440
rect 32324 8090 32352 8434
rect 32312 8084 32364 8090
rect 32312 8026 32364 8032
rect 33704 7886 33732 9318
rect 33888 8906 33916 9862
rect 34713 9820 35021 9829
rect 34713 9818 34719 9820
rect 34775 9818 34799 9820
rect 34855 9818 34879 9820
rect 34935 9818 34959 9820
rect 35015 9818 35021 9820
rect 34775 9766 34777 9818
rect 34957 9766 34959 9818
rect 34713 9764 34719 9766
rect 34775 9764 34799 9766
rect 34855 9764 34879 9766
rect 34935 9764 34959 9766
rect 35015 9764 35021 9766
rect 34713 9755 35021 9764
rect 33876 8900 33928 8906
rect 33876 8842 33928 8848
rect 34713 8732 35021 8741
rect 34713 8730 34719 8732
rect 34775 8730 34799 8732
rect 34855 8730 34879 8732
rect 34935 8730 34959 8732
rect 35015 8730 35021 8732
rect 34775 8678 34777 8730
rect 34957 8678 34959 8730
rect 34713 8676 34719 8678
rect 34775 8676 34799 8678
rect 34855 8676 34879 8678
rect 34935 8676 34959 8678
rect 35015 8676 35021 8678
rect 34713 8667 35021 8676
rect 33692 7880 33744 7886
rect 33692 7822 33744 7828
rect 34713 7644 35021 7653
rect 34713 7642 34719 7644
rect 34775 7642 34799 7644
rect 34855 7642 34879 7644
rect 34935 7642 34959 7644
rect 35015 7642 35021 7644
rect 34775 7590 34777 7642
rect 34957 7590 34959 7642
rect 34713 7588 34719 7590
rect 34775 7588 34799 7590
rect 34855 7588 34879 7590
rect 34935 7588 34959 7590
rect 35015 7588 35021 7590
rect 34713 7579 35021 7588
rect 34713 6556 35021 6565
rect 34713 6554 34719 6556
rect 34775 6554 34799 6556
rect 34855 6554 34879 6556
rect 34935 6554 34959 6556
rect 35015 6554 35021 6556
rect 34775 6502 34777 6554
rect 34957 6502 34959 6554
rect 34713 6500 34719 6502
rect 34775 6500 34799 6502
rect 34855 6500 34879 6502
rect 34935 6500 34959 6502
rect 35015 6500 35021 6502
rect 34713 6491 35021 6500
rect 30932 6452 30984 6458
rect 30932 6394 30984 6400
rect 30840 5704 30892 5710
rect 30840 5646 30892 5652
rect 34713 5468 35021 5477
rect 34713 5466 34719 5468
rect 34775 5466 34799 5468
rect 34855 5466 34879 5468
rect 34935 5466 34959 5468
rect 35015 5466 35021 5468
rect 34775 5414 34777 5466
rect 34957 5414 34959 5466
rect 34713 5412 34719 5414
rect 34775 5412 34799 5414
rect 34855 5412 34879 5414
rect 34935 5412 34959 5414
rect 35015 5412 35021 5414
rect 34713 5403 35021 5412
rect 30493 4924 30801 4933
rect 30493 4922 30499 4924
rect 30555 4922 30579 4924
rect 30635 4922 30659 4924
rect 30715 4922 30739 4924
rect 30795 4922 30801 4924
rect 30555 4870 30557 4922
rect 30737 4870 30739 4922
rect 30493 4868 30499 4870
rect 30555 4868 30579 4870
rect 30635 4868 30659 4870
rect 30715 4868 30739 4870
rect 30795 4868 30801 4870
rect 30493 4859 30801 4868
rect 34713 4380 35021 4389
rect 34713 4378 34719 4380
rect 34775 4378 34799 4380
rect 34855 4378 34879 4380
rect 34935 4378 34959 4380
rect 35015 4378 35021 4380
rect 34775 4326 34777 4378
rect 34957 4326 34959 4378
rect 34713 4324 34719 4326
rect 34775 4324 34799 4326
rect 34855 4324 34879 4326
rect 34935 4324 34959 4326
rect 35015 4324 35021 4326
rect 34713 4315 35021 4324
rect 30493 3836 30801 3845
rect 30493 3834 30499 3836
rect 30555 3834 30579 3836
rect 30635 3834 30659 3836
rect 30715 3834 30739 3836
rect 30795 3834 30801 3836
rect 30555 3782 30557 3834
rect 30737 3782 30739 3834
rect 30493 3780 30499 3782
rect 30555 3780 30579 3782
rect 30635 3780 30659 3782
rect 30715 3780 30739 3782
rect 30795 3780 30801 3782
rect 30493 3771 30801 3780
rect 34713 3292 35021 3301
rect 34713 3290 34719 3292
rect 34775 3290 34799 3292
rect 34855 3290 34879 3292
rect 34935 3290 34959 3292
rect 35015 3290 35021 3292
rect 34775 3238 34777 3290
rect 34957 3238 34959 3290
rect 34713 3236 34719 3238
rect 34775 3236 34799 3238
rect 34855 3236 34879 3238
rect 34935 3236 34959 3238
rect 35015 3236 35021 3238
rect 34713 3227 35021 3236
rect 30380 3120 30432 3126
rect 30380 3062 30432 3068
rect 30493 2748 30801 2757
rect 30493 2746 30499 2748
rect 30555 2746 30579 2748
rect 30635 2746 30659 2748
rect 30715 2746 30739 2748
rect 30795 2746 30801 2748
rect 30555 2694 30557 2746
rect 30737 2694 30739 2746
rect 30493 2692 30499 2694
rect 30555 2692 30579 2694
rect 30635 2692 30659 2694
rect 30715 2692 30739 2694
rect 30795 2692 30801 2694
rect 30493 2683 30801 2692
rect 15476 2440 15528 2446
rect 15476 2382 15528 2388
rect 16304 2440 16356 2446
rect 16304 2382 16356 2388
rect 19064 2440 19116 2446
rect 19064 2382 19116 2388
rect 21088 2440 21140 2446
rect 21088 2382 21140 2388
rect 23388 2440 23440 2446
rect 23388 2382 23440 2388
rect 25596 2440 25648 2446
rect 25596 2382 25648 2388
rect 26240 2440 26292 2446
rect 26240 2382 26292 2388
rect 27896 2440 27948 2446
rect 27896 2382 27948 2388
rect 28356 2440 28408 2446
rect 28356 2382 28408 2388
rect 29552 2440 29604 2446
rect 29552 2382 29604 2388
rect 30840 2440 30892 2446
rect 30840 2382 30892 2388
rect 32128 2440 32180 2446
rect 32128 2382 32180 2388
rect 33416 2440 33468 2446
rect 33416 2382 33468 2388
rect 15384 2372 15436 2378
rect 15384 2314 15436 2320
rect 16672 2372 16724 2378
rect 16672 2314 16724 2320
rect 18236 2372 18288 2378
rect 18236 2314 18288 2320
rect 19248 2372 19300 2378
rect 19248 2314 19300 2320
rect 20536 2372 20588 2378
rect 20536 2314 20588 2320
rect 21824 2372 21876 2378
rect 21824 2314 21876 2320
rect 23112 2372 23164 2378
rect 23112 2314 23164 2320
rect 24400 2372 24452 2378
rect 24400 2314 24452 2320
rect 25688 2372 25740 2378
rect 25688 2314 25740 2320
rect 26976 2372 27028 2378
rect 26976 2314 27028 2320
rect 28264 2372 28316 2378
rect 28264 2314 28316 2320
rect 14372 2304 14424 2310
rect 14372 2246 14424 2252
rect 15396 800 15424 2314
rect 16684 800 16712 2314
rect 17831 2204 18139 2213
rect 17831 2202 17837 2204
rect 17893 2202 17917 2204
rect 17973 2202 17997 2204
rect 18053 2202 18077 2204
rect 18133 2202 18139 2204
rect 17893 2150 17895 2202
rect 18075 2150 18077 2202
rect 17831 2148 17837 2150
rect 17893 2148 17917 2150
rect 17973 2148 17997 2150
rect 18053 2148 18077 2150
rect 18133 2148 18139 2150
rect 17831 2139 18139 2148
rect 17972 870 18092 898
rect 17972 800 18000 870
rect 1214 0 1270 800
rect 2502 0 2558 800
rect 3790 0 3846 800
rect 5078 0 5134 800
rect 6366 0 6422 800
rect 7654 0 7710 800
rect 8942 0 8998 800
rect 10230 0 10286 800
rect 11518 0 11574 800
rect 12806 0 12862 800
rect 14094 0 14150 800
rect 15382 0 15438 800
rect 16670 0 16726 800
rect 17958 0 18014 800
rect 18064 762 18092 870
rect 18248 762 18276 2314
rect 19260 800 19288 2314
rect 20548 800 20576 2314
rect 21836 800 21864 2314
rect 23124 800 23152 2314
rect 24412 800 24440 2314
rect 25700 800 25728 2314
rect 26272 2204 26580 2213
rect 26272 2202 26278 2204
rect 26334 2202 26358 2204
rect 26414 2202 26438 2204
rect 26494 2202 26518 2204
rect 26574 2202 26580 2204
rect 26334 2150 26336 2202
rect 26516 2150 26518 2202
rect 26272 2148 26278 2150
rect 26334 2148 26358 2150
rect 26414 2148 26438 2150
rect 26494 2148 26518 2150
rect 26574 2148 26580 2150
rect 26272 2139 26580 2148
rect 26988 800 27016 2314
rect 28276 800 28304 2314
rect 29564 800 29592 2382
rect 30852 800 30880 2382
rect 32140 800 32168 2382
rect 33428 800 33456 2382
rect 34612 2304 34664 2310
rect 34612 2246 34664 2252
rect 34624 1170 34652 2246
rect 34713 2204 35021 2213
rect 34713 2202 34719 2204
rect 34775 2202 34799 2204
rect 34855 2202 34879 2204
rect 34935 2202 34959 2204
rect 35015 2202 35021 2204
rect 34775 2150 34777 2202
rect 34957 2150 34959 2202
rect 34713 2148 34719 2150
rect 34775 2148 34799 2150
rect 34855 2148 34879 2150
rect 34935 2148 34959 2150
rect 35015 2148 35021 2150
rect 34713 2139 35021 2148
rect 34624 1142 34744 1170
rect 34716 800 34744 1142
rect 18064 734 18276 762
rect 19246 0 19302 800
rect 20534 0 20590 800
rect 21822 0 21878 800
rect 23110 0 23166 800
rect 24398 0 24454 800
rect 25686 0 25742 800
rect 26974 0 27030 800
rect 28262 0 28318 800
rect 29550 0 29606 800
rect 30838 0 30894 800
rect 32126 0 32182 800
rect 33414 0 33470 800
rect 34702 0 34758 800
<< via2 >>
rect 9396 33754 9452 33756
rect 9476 33754 9532 33756
rect 9556 33754 9612 33756
rect 9636 33754 9692 33756
rect 9396 33702 9442 33754
rect 9442 33702 9452 33754
rect 9476 33702 9506 33754
rect 9506 33702 9518 33754
rect 9518 33702 9532 33754
rect 9556 33702 9570 33754
rect 9570 33702 9582 33754
rect 9582 33702 9612 33754
rect 9636 33702 9646 33754
rect 9646 33702 9692 33754
rect 9396 33700 9452 33702
rect 9476 33700 9532 33702
rect 9556 33700 9612 33702
rect 9636 33700 9692 33702
rect 17837 33754 17893 33756
rect 17917 33754 17973 33756
rect 17997 33754 18053 33756
rect 18077 33754 18133 33756
rect 17837 33702 17883 33754
rect 17883 33702 17893 33754
rect 17917 33702 17947 33754
rect 17947 33702 17959 33754
rect 17959 33702 17973 33754
rect 17997 33702 18011 33754
rect 18011 33702 18023 33754
rect 18023 33702 18053 33754
rect 18077 33702 18087 33754
rect 18087 33702 18133 33754
rect 17837 33700 17893 33702
rect 17917 33700 17973 33702
rect 17997 33700 18053 33702
rect 18077 33700 18133 33702
rect 26278 33754 26334 33756
rect 26358 33754 26414 33756
rect 26438 33754 26494 33756
rect 26518 33754 26574 33756
rect 26278 33702 26324 33754
rect 26324 33702 26334 33754
rect 26358 33702 26388 33754
rect 26388 33702 26400 33754
rect 26400 33702 26414 33754
rect 26438 33702 26452 33754
rect 26452 33702 26464 33754
rect 26464 33702 26494 33754
rect 26518 33702 26528 33754
rect 26528 33702 26574 33754
rect 26278 33700 26334 33702
rect 26358 33700 26414 33702
rect 26438 33700 26494 33702
rect 26518 33700 26574 33702
rect 34719 33754 34775 33756
rect 34799 33754 34855 33756
rect 34879 33754 34935 33756
rect 34959 33754 35015 33756
rect 34719 33702 34765 33754
rect 34765 33702 34775 33754
rect 34799 33702 34829 33754
rect 34829 33702 34841 33754
rect 34841 33702 34855 33754
rect 34879 33702 34893 33754
rect 34893 33702 34905 33754
rect 34905 33702 34935 33754
rect 34959 33702 34969 33754
rect 34969 33702 35015 33754
rect 34719 33700 34775 33702
rect 34799 33700 34855 33702
rect 34879 33700 34935 33702
rect 34959 33700 35015 33702
rect 5176 33210 5232 33212
rect 5256 33210 5312 33212
rect 5336 33210 5392 33212
rect 5416 33210 5472 33212
rect 5176 33158 5222 33210
rect 5222 33158 5232 33210
rect 5256 33158 5286 33210
rect 5286 33158 5298 33210
rect 5298 33158 5312 33210
rect 5336 33158 5350 33210
rect 5350 33158 5362 33210
rect 5362 33158 5392 33210
rect 5416 33158 5426 33210
rect 5426 33158 5472 33210
rect 5176 33156 5232 33158
rect 5256 33156 5312 33158
rect 5336 33156 5392 33158
rect 5416 33156 5472 33158
rect 5176 32122 5232 32124
rect 5256 32122 5312 32124
rect 5336 32122 5392 32124
rect 5416 32122 5472 32124
rect 5176 32070 5222 32122
rect 5222 32070 5232 32122
rect 5256 32070 5286 32122
rect 5286 32070 5298 32122
rect 5298 32070 5312 32122
rect 5336 32070 5350 32122
rect 5350 32070 5362 32122
rect 5362 32070 5392 32122
rect 5416 32070 5426 32122
rect 5426 32070 5472 32122
rect 5176 32068 5232 32070
rect 5256 32068 5312 32070
rect 5336 32068 5392 32070
rect 5416 32068 5472 32070
rect 9396 32666 9452 32668
rect 9476 32666 9532 32668
rect 9556 32666 9612 32668
rect 9636 32666 9692 32668
rect 9396 32614 9442 32666
rect 9442 32614 9452 32666
rect 9476 32614 9506 32666
rect 9506 32614 9518 32666
rect 9518 32614 9532 32666
rect 9556 32614 9570 32666
rect 9570 32614 9582 32666
rect 9582 32614 9612 32666
rect 9636 32614 9646 32666
rect 9646 32614 9692 32666
rect 9396 32612 9452 32614
rect 9476 32612 9532 32614
rect 9556 32612 9612 32614
rect 9636 32612 9692 32614
rect 5176 31034 5232 31036
rect 5256 31034 5312 31036
rect 5336 31034 5392 31036
rect 5416 31034 5472 31036
rect 5176 30982 5222 31034
rect 5222 30982 5232 31034
rect 5256 30982 5286 31034
rect 5286 30982 5298 31034
rect 5298 30982 5312 31034
rect 5336 30982 5350 31034
rect 5350 30982 5362 31034
rect 5362 30982 5392 31034
rect 5416 30982 5426 31034
rect 5426 30982 5472 31034
rect 5176 30980 5232 30982
rect 5256 30980 5312 30982
rect 5336 30980 5392 30982
rect 5416 30980 5472 30982
rect 5176 29946 5232 29948
rect 5256 29946 5312 29948
rect 5336 29946 5392 29948
rect 5416 29946 5472 29948
rect 5176 29894 5222 29946
rect 5222 29894 5232 29946
rect 5256 29894 5286 29946
rect 5286 29894 5298 29946
rect 5298 29894 5312 29946
rect 5336 29894 5350 29946
rect 5350 29894 5362 29946
rect 5362 29894 5392 29946
rect 5416 29894 5426 29946
rect 5426 29894 5472 29946
rect 5176 29892 5232 29894
rect 5256 29892 5312 29894
rect 5336 29892 5392 29894
rect 5416 29892 5472 29894
rect 5176 28858 5232 28860
rect 5256 28858 5312 28860
rect 5336 28858 5392 28860
rect 5416 28858 5472 28860
rect 5176 28806 5222 28858
rect 5222 28806 5232 28858
rect 5256 28806 5286 28858
rect 5286 28806 5298 28858
rect 5298 28806 5312 28858
rect 5336 28806 5350 28858
rect 5350 28806 5362 28858
rect 5362 28806 5392 28858
rect 5416 28806 5426 28858
rect 5426 28806 5472 28858
rect 5176 28804 5232 28806
rect 5256 28804 5312 28806
rect 5336 28804 5392 28806
rect 5416 28804 5472 28806
rect 9396 31578 9452 31580
rect 9476 31578 9532 31580
rect 9556 31578 9612 31580
rect 9636 31578 9692 31580
rect 9396 31526 9442 31578
rect 9442 31526 9452 31578
rect 9476 31526 9506 31578
rect 9506 31526 9518 31578
rect 9518 31526 9532 31578
rect 9556 31526 9570 31578
rect 9570 31526 9582 31578
rect 9582 31526 9612 31578
rect 9636 31526 9646 31578
rect 9646 31526 9692 31578
rect 9396 31524 9452 31526
rect 9476 31524 9532 31526
rect 9556 31524 9612 31526
rect 9636 31524 9692 31526
rect 13617 33210 13673 33212
rect 13697 33210 13753 33212
rect 13777 33210 13833 33212
rect 13857 33210 13913 33212
rect 13617 33158 13663 33210
rect 13663 33158 13673 33210
rect 13697 33158 13727 33210
rect 13727 33158 13739 33210
rect 13739 33158 13753 33210
rect 13777 33158 13791 33210
rect 13791 33158 13803 33210
rect 13803 33158 13833 33210
rect 13857 33158 13867 33210
rect 13867 33158 13913 33210
rect 13617 33156 13673 33158
rect 13697 33156 13753 33158
rect 13777 33156 13833 33158
rect 13857 33156 13913 33158
rect 9396 30490 9452 30492
rect 9476 30490 9532 30492
rect 9556 30490 9612 30492
rect 9636 30490 9692 30492
rect 9396 30438 9442 30490
rect 9442 30438 9452 30490
rect 9476 30438 9506 30490
rect 9506 30438 9518 30490
rect 9518 30438 9532 30490
rect 9556 30438 9570 30490
rect 9570 30438 9582 30490
rect 9582 30438 9612 30490
rect 9636 30438 9646 30490
rect 9646 30438 9692 30490
rect 9396 30436 9452 30438
rect 9476 30436 9532 30438
rect 9556 30436 9612 30438
rect 9636 30436 9692 30438
rect 9396 29402 9452 29404
rect 9476 29402 9532 29404
rect 9556 29402 9612 29404
rect 9636 29402 9692 29404
rect 9396 29350 9442 29402
rect 9442 29350 9452 29402
rect 9476 29350 9506 29402
rect 9506 29350 9518 29402
rect 9518 29350 9532 29402
rect 9556 29350 9570 29402
rect 9570 29350 9582 29402
rect 9582 29350 9612 29402
rect 9636 29350 9646 29402
rect 9646 29350 9692 29402
rect 9396 29348 9452 29350
rect 9476 29348 9532 29350
rect 9556 29348 9612 29350
rect 9636 29348 9692 29350
rect 5176 27770 5232 27772
rect 5256 27770 5312 27772
rect 5336 27770 5392 27772
rect 5416 27770 5472 27772
rect 5176 27718 5222 27770
rect 5222 27718 5232 27770
rect 5256 27718 5286 27770
rect 5286 27718 5298 27770
rect 5298 27718 5312 27770
rect 5336 27718 5350 27770
rect 5350 27718 5362 27770
rect 5362 27718 5392 27770
rect 5416 27718 5426 27770
rect 5426 27718 5472 27770
rect 5176 27716 5232 27718
rect 5256 27716 5312 27718
rect 5336 27716 5392 27718
rect 5416 27716 5472 27718
rect 9396 28314 9452 28316
rect 9476 28314 9532 28316
rect 9556 28314 9612 28316
rect 9636 28314 9692 28316
rect 9396 28262 9442 28314
rect 9442 28262 9452 28314
rect 9476 28262 9506 28314
rect 9506 28262 9518 28314
rect 9518 28262 9532 28314
rect 9556 28262 9570 28314
rect 9570 28262 9582 28314
rect 9582 28262 9612 28314
rect 9636 28262 9646 28314
rect 9646 28262 9692 28314
rect 9396 28260 9452 28262
rect 9476 28260 9532 28262
rect 9556 28260 9612 28262
rect 9636 28260 9692 28262
rect 5176 26682 5232 26684
rect 5256 26682 5312 26684
rect 5336 26682 5392 26684
rect 5416 26682 5472 26684
rect 5176 26630 5222 26682
rect 5222 26630 5232 26682
rect 5256 26630 5286 26682
rect 5286 26630 5298 26682
rect 5298 26630 5312 26682
rect 5336 26630 5350 26682
rect 5350 26630 5362 26682
rect 5362 26630 5392 26682
rect 5416 26630 5426 26682
rect 5426 26630 5472 26682
rect 5176 26628 5232 26630
rect 5256 26628 5312 26630
rect 5336 26628 5392 26630
rect 5416 26628 5472 26630
rect 9396 27226 9452 27228
rect 9476 27226 9532 27228
rect 9556 27226 9612 27228
rect 9636 27226 9692 27228
rect 9396 27174 9442 27226
rect 9442 27174 9452 27226
rect 9476 27174 9506 27226
rect 9506 27174 9518 27226
rect 9518 27174 9532 27226
rect 9556 27174 9570 27226
rect 9570 27174 9582 27226
rect 9582 27174 9612 27226
rect 9636 27174 9646 27226
rect 9646 27174 9692 27226
rect 9396 27172 9452 27174
rect 9476 27172 9532 27174
rect 9556 27172 9612 27174
rect 9636 27172 9692 27174
rect 9396 26138 9452 26140
rect 9476 26138 9532 26140
rect 9556 26138 9612 26140
rect 9636 26138 9692 26140
rect 9396 26086 9442 26138
rect 9442 26086 9452 26138
rect 9476 26086 9506 26138
rect 9506 26086 9518 26138
rect 9518 26086 9532 26138
rect 9556 26086 9570 26138
rect 9570 26086 9582 26138
rect 9582 26086 9612 26138
rect 9636 26086 9646 26138
rect 9646 26086 9692 26138
rect 9396 26084 9452 26086
rect 9476 26084 9532 26086
rect 9556 26084 9612 26086
rect 9636 26084 9692 26086
rect 5176 25594 5232 25596
rect 5256 25594 5312 25596
rect 5336 25594 5392 25596
rect 5416 25594 5472 25596
rect 5176 25542 5222 25594
rect 5222 25542 5232 25594
rect 5256 25542 5286 25594
rect 5286 25542 5298 25594
rect 5298 25542 5312 25594
rect 5336 25542 5350 25594
rect 5350 25542 5362 25594
rect 5362 25542 5392 25594
rect 5416 25542 5426 25594
rect 5426 25542 5472 25594
rect 5176 25540 5232 25542
rect 5256 25540 5312 25542
rect 5336 25540 5392 25542
rect 5416 25540 5472 25542
rect 9396 25050 9452 25052
rect 9476 25050 9532 25052
rect 9556 25050 9612 25052
rect 9636 25050 9692 25052
rect 9396 24998 9442 25050
rect 9442 24998 9452 25050
rect 9476 24998 9506 25050
rect 9506 24998 9518 25050
rect 9518 24998 9532 25050
rect 9556 24998 9570 25050
rect 9570 24998 9582 25050
rect 9582 24998 9612 25050
rect 9636 24998 9646 25050
rect 9646 24998 9692 25050
rect 9396 24996 9452 24998
rect 9476 24996 9532 24998
rect 9556 24996 9612 24998
rect 9636 24996 9692 24998
rect 5176 24506 5232 24508
rect 5256 24506 5312 24508
rect 5336 24506 5392 24508
rect 5416 24506 5472 24508
rect 5176 24454 5222 24506
rect 5222 24454 5232 24506
rect 5256 24454 5286 24506
rect 5286 24454 5298 24506
rect 5298 24454 5312 24506
rect 5336 24454 5350 24506
rect 5350 24454 5362 24506
rect 5362 24454 5392 24506
rect 5416 24454 5426 24506
rect 5426 24454 5472 24506
rect 5176 24452 5232 24454
rect 5256 24452 5312 24454
rect 5336 24452 5392 24454
rect 5416 24452 5472 24454
rect 5176 23418 5232 23420
rect 5256 23418 5312 23420
rect 5336 23418 5392 23420
rect 5416 23418 5472 23420
rect 5176 23366 5222 23418
rect 5222 23366 5232 23418
rect 5256 23366 5286 23418
rect 5286 23366 5298 23418
rect 5298 23366 5312 23418
rect 5336 23366 5350 23418
rect 5350 23366 5362 23418
rect 5362 23366 5392 23418
rect 5416 23366 5426 23418
rect 5426 23366 5472 23418
rect 5176 23364 5232 23366
rect 5256 23364 5312 23366
rect 5336 23364 5392 23366
rect 5416 23364 5472 23366
rect 5176 22330 5232 22332
rect 5256 22330 5312 22332
rect 5336 22330 5392 22332
rect 5416 22330 5472 22332
rect 5176 22278 5222 22330
rect 5222 22278 5232 22330
rect 5256 22278 5286 22330
rect 5286 22278 5298 22330
rect 5298 22278 5312 22330
rect 5336 22278 5350 22330
rect 5350 22278 5362 22330
rect 5362 22278 5392 22330
rect 5416 22278 5426 22330
rect 5426 22278 5472 22330
rect 5176 22276 5232 22278
rect 5256 22276 5312 22278
rect 5336 22276 5392 22278
rect 5416 22276 5472 22278
rect 5176 21242 5232 21244
rect 5256 21242 5312 21244
rect 5336 21242 5392 21244
rect 5416 21242 5472 21244
rect 5176 21190 5222 21242
rect 5222 21190 5232 21242
rect 5256 21190 5286 21242
rect 5286 21190 5298 21242
rect 5298 21190 5312 21242
rect 5336 21190 5350 21242
rect 5350 21190 5362 21242
rect 5362 21190 5392 21242
rect 5416 21190 5426 21242
rect 5426 21190 5472 21242
rect 5176 21188 5232 21190
rect 5256 21188 5312 21190
rect 5336 21188 5392 21190
rect 5416 21188 5472 21190
rect 5176 20154 5232 20156
rect 5256 20154 5312 20156
rect 5336 20154 5392 20156
rect 5416 20154 5472 20156
rect 5176 20102 5222 20154
rect 5222 20102 5232 20154
rect 5256 20102 5286 20154
rect 5286 20102 5298 20154
rect 5298 20102 5312 20154
rect 5336 20102 5350 20154
rect 5350 20102 5362 20154
rect 5362 20102 5392 20154
rect 5416 20102 5426 20154
rect 5426 20102 5472 20154
rect 5176 20100 5232 20102
rect 5256 20100 5312 20102
rect 5336 20100 5392 20102
rect 5416 20100 5472 20102
rect 5176 19066 5232 19068
rect 5256 19066 5312 19068
rect 5336 19066 5392 19068
rect 5416 19066 5472 19068
rect 5176 19014 5222 19066
rect 5222 19014 5232 19066
rect 5256 19014 5286 19066
rect 5286 19014 5298 19066
rect 5298 19014 5312 19066
rect 5336 19014 5350 19066
rect 5350 19014 5362 19066
rect 5362 19014 5392 19066
rect 5416 19014 5426 19066
rect 5426 19014 5472 19066
rect 5176 19012 5232 19014
rect 5256 19012 5312 19014
rect 5336 19012 5392 19014
rect 5416 19012 5472 19014
rect 5176 17978 5232 17980
rect 5256 17978 5312 17980
rect 5336 17978 5392 17980
rect 5416 17978 5472 17980
rect 5176 17926 5222 17978
rect 5222 17926 5232 17978
rect 5256 17926 5286 17978
rect 5286 17926 5298 17978
rect 5298 17926 5312 17978
rect 5336 17926 5350 17978
rect 5350 17926 5362 17978
rect 5362 17926 5392 17978
rect 5416 17926 5426 17978
rect 5426 17926 5472 17978
rect 5176 17924 5232 17926
rect 5256 17924 5312 17926
rect 5336 17924 5392 17926
rect 5416 17924 5472 17926
rect 5176 16890 5232 16892
rect 5256 16890 5312 16892
rect 5336 16890 5392 16892
rect 5416 16890 5472 16892
rect 5176 16838 5222 16890
rect 5222 16838 5232 16890
rect 5256 16838 5286 16890
rect 5286 16838 5298 16890
rect 5298 16838 5312 16890
rect 5336 16838 5350 16890
rect 5350 16838 5362 16890
rect 5362 16838 5392 16890
rect 5416 16838 5426 16890
rect 5426 16838 5472 16890
rect 5176 16836 5232 16838
rect 5256 16836 5312 16838
rect 5336 16836 5392 16838
rect 5416 16836 5472 16838
rect 5176 15802 5232 15804
rect 5256 15802 5312 15804
rect 5336 15802 5392 15804
rect 5416 15802 5472 15804
rect 5176 15750 5222 15802
rect 5222 15750 5232 15802
rect 5256 15750 5286 15802
rect 5286 15750 5298 15802
rect 5298 15750 5312 15802
rect 5336 15750 5350 15802
rect 5350 15750 5362 15802
rect 5362 15750 5392 15802
rect 5416 15750 5426 15802
rect 5426 15750 5472 15802
rect 5176 15748 5232 15750
rect 5256 15748 5312 15750
rect 5336 15748 5392 15750
rect 5416 15748 5472 15750
rect 9396 23962 9452 23964
rect 9476 23962 9532 23964
rect 9556 23962 9612 23964
rect 9636 23962 9692 23964
rect 9396 23910 9442 23962
rect 9442 23910 9452 23962
rect 9476 23910 9506 23962
rect 9506 23910 9518 23962
rect 9518 23910 9532 23962
rect 9556 23910 9570 23962
rect 9570 23910 9582 23962
rect 9582 23910 9612 23962
rect 9636 23910 9646 23962
rect 9646 23910 9692 23962
rect 9396 23908 9452 23910
rect 9476 23908 9532 23910
rect 9556 23908 9612 23910
rect 9636 23908 9692 23910
rect 9396 22874 9452 22876
rect 9476 22874 9532 22876
rect 9556 22874 9612 22876
rect 9636 22874 9692 22876
rect 9396 22822 9442 22874
rect 9442 22822 9452 22874
rect 9476 22822 9506 22874
rect 9506 22822 9518 22874
rect 9518 22822 9532 22874
rect 9556 22822 9570 22874
rect 9570 22822 9582 22874
rect 9582 22822 9612 22874
rect 9636 22822 9646 22874
rect 9646 22822 9692 22874
rect 9396 22820 9452 22822
rect 9476 22820 9532 22822
rect 9556 22820 9612 22822
rect 9636 22820 9692 22822
rect 5176 14714 5232 14716
rect 5256 14714 5312 14716
rect 5336 14714 5392 14716
rect 5416 14714 5472 14716
rect 5176 14662 5222 14714
rect 5222 14662 5232 14714
rect 5256 14662 5286 14714
rect 5286 14662 5298 14714
rect 5298 14662 5312 14714
rect 5336 14662 5350 14714
rect 5350 14662 5362 14714
rect 5362 14662 5392 14714
rect 5416 14662 5426 14714
rect 5426 14662 5472 14714
rect 5176 14660 5232 14662
rect 5256 14660 5312 14662
rect 5336 14660 5392 14662
rect 5416 14660 5472 14662
rect 5176 13626 5232 13628
rect 5256 13626 5312 13628
rect 5336 13626 5392 13628
rect 5416 13626 5472 13628
rect 5176 13574 5222 13626
rect 5222 13574 5232 13626
rect 5256 13574 5286 13626
rect 5286 13574 5298 13626
rect 5298 13574 5312 13626
rect 5336 13574 5350 13626
rect 5350 13574 5362 13626
rect 5362 13574 5392 13626
rect 5416 13574 5426 13626
rect 5426 13574 5472 13626
rect 5176 13572 5232 13574
rect 5256 13572 5312 13574
rect 5336 13572 5392 13574
rect 5416 13572 5472 13574
rect 5176 12538 5232 12540
rect 5256 12538 5312 12540
rect 5336 12538 5392 12540
rect 5416 12538 5472 12540
rect 5176 12486 5222 12538
rect 5222 12486 5232 12538
rect 5256 12486 5286 12538
rect 5286 12486 5298 12538
rect 5298 12486 5312 12538
rect 5336 12486 5350 12538
rect 5350 12486 5362 12538
rect 5362 12486 5392 12538
rect 5416 12486 5426 12538
rect 5426 12486 5472 12538
rect 5176 12484 5232 12486
rect 5256 12484 5312 12486
rect 5336 12484 5392 12486
rect 5416 12484 5472 12486
rect 9396 21786 9452 21788
rect 9476 21786 9532 21788
rect 9556 21786 9612 21788
rect 9636 21786 9692 21788
rect 9396 21734 9442 21786
rect 9442 21734 9452 21786
rect 9476 21734 9506 21786
rect 9506 21734 9518 21786
rect 9518 21734 9532 21786
rect 9556 21734 9570 21786
rect 9570 21734 9582 21786
rect 9582 21734 9612 21786
rect 9636 21734 9646 21786
rect 9646 21734 9692 21786
rect 9396 21732 9452 21734
rect 9476 21732 9532 21734
rect 9556 21732 9612 21734
rect 9636 21732 9692 21734
rect 9396 20698 9452 20700
rect 9476 20698 9532 20700
rect 9556 20698 9612 20700
rect 9636 20698 9692 20700
rect 9396 20646 9442 20698
rect 9442 20646 9452 20698
rect 9476 20646 9506 20698
rect 9506 20646 9518 20698
rect 9518 20646 9532 20698
rect 9556 20646 9570 20698
rect 9570 20646 9582 20698
rect 9582 20646 9612 20698
rect 9636 20646 9646 20698
rect 9646 20646 9692 20698
rect 9396 20644 9452 20646
rect 9476 20644 9532 20646
rect 9556 20644 9612 20646
rect 9636 20644 9692 20646
rect 9396 19610 9452 19612
rect 9476 19610 9532 19612
rect 9556 19610 9612 19612
rect 9636 19610 9692 19612
rect 9396 19558 9442 19610
rect 9442 19558 9452 19610
rect 9476 19558 9506 19610
rect 9506 19558 9518 19610
rect 9518 19558 9532 19610
rect 9556 19558 9570 19610
rect 9570 19558 9582 19610
rect 9582 19558 9612 19610
rect 9636 19558 9646 19610
rect 9646 19558 9692 19610
rect 9396 19556 9452 19558
rect 9476 19556 9532 19558
rect 9556 19556 9612 19558
rect 9636 19556 9692 19558
rect 9396 18522 9452 18524
rect 9476 18522 9532 18524
rect 9556 18522 9612 18524
rect 9636 18522 9692 18524
rect 9396 18470 9442 18522
rect 9442 18470 9452 18522
rect 9476 18470 9506 18522
rect 9506 18470 9518 18522
rect 9518 18470 9532 18522
rect 9556 18470 9570 18522
rect 9570 18470 9582 18522
rect 9582 18470 9612 18522
rect 9636 18470 9646 18522
rect 9646 18470 9692 18522
rect 9396 18468 9452 18470
rect 9476 18468 9532 18470
rect 9556 18468 9612 18470
rect 9636 18468 9692 18470
rect 9396 17434 9452 17436
rect 9476 17434 9532 17436
rect 9556 17434 9612 17436
rect 9636 17434 9692 17436
rect 9396 17382 9442 17434
rect 9442 17382 9452 17434
rect 9476 17382 9506 17434
rect 9506 17382 9518 17434
rect 9518 17382 9532 17434
rect 9556 17382 9570 17434
rect 9570 17382 9582 17434
rect 9582 17382 9612 17434
rect 9636 17382 9646 17434
rect 9646 17382 9692 17434
rect 9396 17380 9452 17382
rect 9476 17380 9532 17382
rect 9556 17380 9612 17382
rect 9636 17380 9692 17382
rect 9396 16346 9452 16348
rect 9476 16346 9532 16348
rect 9556 16346 9612 16348
rect 9636 16346 9692 16348
rect 9396 16294 9442 16346
rect 9442 16294 9452 16346
rect 9476 16294 9506 16346
rect 9506 16294 9518 16346
rect 9518 16294 9532 16346
rect 9556 16294 9570 16346
rect 9570 16294 9582 16346
rect 9582 16294 9612 16346
rect 9636 16294 9646 16346
rect 9646 16294 9692 16346
rect 9396 16292 9452 16294
rect 9476 16292 9532 16294
rect 9556 16292 9612 16294
rect 9636 16292 9692 16294
rect 9396 15258 9452 15260
rect 9476 15258 9532 15260
rect 9556 15258 9612 15260
rect 9636 15258 9692 15260
rect 9396 15206 9442 15258
rect 9442 15206 9452 15258
rect 9476 15206 9506 15258
rect 9506 15206 9518 15258
rect 9518 15206 9532 15258
rect 9556 15206 9570 15258
rect 9570 15206 9582 15258
rect 9582 15206 9612 15258
rect 9636 15206 9646 15258
rect 9646 15206 9692 15258
rect 9396 15204 9452 15206
rect 9476 15204 9532 15206
rect 9556 15204 9612 15206
rect 9636 15204 9692 15206
rect 5176 11450 5232 11452
rect 5256 11450 5312 11452
rect 5336 11450 5392 11452
rect 5416 11450 5472 11452
rect 5176 11398 5222 11450
rect 5222 11398 5232 11450
rect 5256 11398 5286 11450
rect 5286 11398 5298 11450
rect 5298 11398 5312 11450
rect 5336 11398 5350 11450
rect 5350 11398 5362 11450
rect 5362 11398 5392 11450
rect 5416 11398 5426 11450
rect 5426 11398 5472 11450
rect 5176 11396 5232 11398
rect 5256 11396 5312 11398
rect 5336 11396 5392 11398
rect 5416 11396 5472 11398
rect 5176 10362 5232 10364
rect 5256 10362 5312 10364
rect 5336 10362 5392 10364
rect 5416 10362 5472 10364
rect 5176 10310 5222 10362
rect 5222 10310 5232 10362
rect 5256 10310 5286 10362
rect 5286 10310 5298 10362
rect 5298 10310 5312 10362
rect 5336 10310 5350 10362
rect 5350 10310 5362 10362
rect 5362 10310 5392 10362
rect 5416 10310 5426 10362
rect 5426 10310 5472 10362
rect 5176 10308 5232 10310
rect 5256 10308 5312 10310
rect 5336 10308 5392 10310
rect 5416 10308 5472 10310
rect 5176 9274 5232 9276
rect 5256 9274 5312 9276
rect 5336 9274 5392 9276
rect 5416 9274 5472 9276
rect 5176 9222 5222 9274
rect 5222 9222 5232 9274
rect 5256 9222 5286 9274
rect 5286 9222 5298 9274
rect 5298 9222 5312 9274
rect 5336 9222 5350 9274
rect 5350 9222 5362 9274
rect 5362 9222 5392 9274
rect 5416 9222 5426 9274
rect 5426 9222 5472 9274
rect 5176 9220 5232 9222
rect 5256 9220 5312 9222
rect 5336 9220 5392 9222
rect 5416 9220 5472 9222
rect 5176 8186 5232 8188
rect 5256 8186 5312 8188
rect 5336 8186 5392 8188
rect 5416 8186 5472 8188
rect 5176 8134 5222 8186
rect 5222 8134 5232 8186
rect 5256 8134 5286 8186
rect 5286 8134 5298 8186
rect 5298 8134 5312 8186
rect 5336 8134 5350 8186
rect 5350 8134 5362 8186
rect 5362 8134 5392 8186
rect 5416 8134 5426 8186
rect 5426 8134 5472 8186
rect 5176 8132 5232 8134
rect 5256 8132 5312 8134
rect 5336 8132 5392 8134
rect 5416 8132 5472 8134
rect 5176 7098 5232 7100
rect 5256 7098 5312 7100
rect 5336 7098 5392 7100
rect 5416 7098 5472 7100
rect 5176 7046 5222 7098
rect 5222 7046 5232 7098
rect 5256 7046 5286 7098
rect 5286 7046 5298 7098
rect 5298 7046 5312 7098
rect 5336 7046 5350 7098
rect 5350 7046 5362 7098
rect 5362 7046 5392 7098
rect 5416 7046 5426 7098
rect 5426 7046 5472 7098
rect 5176 7044 5232 7046
rect 5256 7044 5312 7046
rect 5336 7044 5392 7046
rect 5416 7044 5472 7046
rect 5176 6010 5232 6012
rect 5256 6010 5312 6012
rect 5336 6010 5392 6012
rect 5416 6010 5472 6012
rect 5176 5958 5222 6010
rect 5222 5958 5232 6010
rect 5256 5958 5286 6010
rect 5286 5958 5298 6010
rect 5298 5958 5312 6010
rect 5336 5958 5350 6010
rect 5350 5958 5362 6010
rect 5362 5958 5392 6010
rect 5416 5958 5426 6010
rect 5426 5958 5472 6010
rect 5176 5956 5232 5958
rect 5256 5956 5312 5958
rect 5336 5956 5392 5958
rect 5416 5956 5472 5958
rect 5176 4922 5232 4924
rect 5256 4922 5312 4924
rect 5336 4922 5392 4924
rect 5416 4922 5472 4924
rect 5176 4870 5222 4922
rect 5222 4870 5232 4922
rect 5256 4870 5286 4922
rect 5286 4870 5298 4922
rect 5298 4870 5312 4922
rect 5336 4870 5350 4922
rect 5350 4870 5362 4922
rect 5362 4870 5392 4922
rect 5416 4870 5426 4922
rect 5426 4870 5472 4922
rect 5176 4868 5232 4870
rect 5256 4868 5312 4870
rect 5336 4868 5392 4870
rect 5416 4868 5472 4870
rect 5176 3834 5232 3836
rect 5256 3834 5312 3836
rect 5336 3834 5392 3836
rect 5416 3834 5472 3836
rect 5176 3782 5222 3834
rect 5222 3782 5232 3834
rect 5256 3782 5286 3834
rect 5286 3782 5298 3834
rect 5298 3782 5312 3834
rect 5336 3782 5350 3834
rect 5350 3782 5362 3834
rect 5362 3782 5392 3834
rect 5416 3782 5426 3834
rect 5426 3782 5472 3834
rect 5176 3780 5232 3782
rect 5256 3780 5312 3782
rect 5336 3780 5392 3782
rect 5416 3780 5472 3782
rect 5176 2746 5232 2748
rect 5256 2746 5312 2748
rect 5336 2746 5392 2748
rect 5416 2746 5472 2748
rect 5176 2694 5222 2746
rect 5222 2694 5232 2746
rect 5256 2694 5286 2746
rect 5286 2694 5298 2746
rect 5298 2694 5312 2746
rect 5336 2694 5350 2746
rect 5350 2694 5362 2746
rect 5362 2694 5392 2746
rect 5416 2694 5426 2746
rect 5426 2694 5472 2746
rect 5176 2692 5232 2694
rect 5256 2692 5312 2694
rect 5336 2692 5392 2694
rect 5416 2692 5472 2694
rect 9396 14170 9452 14172
rect 9476 14170 9532 14172
rect 9556 14170 9612 14172
rect 9636 14170 9692 14172
rect 9396 14118 9442 14170
rect 9442 14118 9452 14170
rect 9476 14118 9506 14170
rect 9506 14118 9518 14170
rect 9518 14118 9532 14170
rect 9556 14118 9570 14170
rect 9570 14118 9582 14170
rect 9582 14118 9612 14170
rect 9636 14118 9646 14170
rect 9646 14118 9692 14170
rect 9396 14116 9452 14118
rect 9476 14116 9532 14118
rect 9556 14116 9612 14118
rect 9636 14116 9692 14118
rect 9396 13082 9452 13084
rect 9476 13082 9532 13084
rect 9556 13082 9612 13084
rect 9636 13082 9692 13084
rect 9396 13030 9442 13082
rect 9442 13030 9452 13082
rect 9476 13030 9506 13082
rect 9506 13030 9518 13082
rect 9518 13030 9532 13082
rect 9556 13030 9570 13082
rect 9570 13030 9582 13082
rect 9582 13030 9612 13082
rect 9636 13030 9646 13082
rect 9646 13030 9692 13082
rect 9396 13028 9452 13030
rect 9476 13028 9532 13030
rect 9556 13028 9612 13030
rect 9636 13028 9692 13030
rect 9396 11994 9452 11996
rect 9476 11994 9532 11996
rect 9556 11994 9612 11996
rect 9636 11994 9692 11996
rect 9396 11942 9442 11994
rect 9442 11942 9452 11994
rect 9476 11942 9506 11994
rect 9506 11942 9518 11994
rect 9518 11942 9532 11994
rect 9556 11942 9570 11994
rect 9570 11942 9582 11994
rect 9582 11942 9612 11994
rect 9636 11942 9646 11994
rect 9646 11942 9692 11994
rect 9396 11940 9452 11942
rect 9476 11940 9532 11942
rect 9556 11940 9612 11942
rect 9636 11940 9692 11942
rect 9396 10906 9452 10908
rect 9476 10906 9532 10908
rect 9556 10906 9612 10908
rect 9636 10906 9692 10908
rect 9396 10854 9442 10906
rect 9442 10854 9452 10906
rect 9476 10854 9506 10906
rect 9506 10854 9518 10906
rect 9518 10854 9532 10906
rect 9556 10854 9570 10906
rect 9570 10854 9582 10906
rect 9582 10854 9612 10906
rect 9636 10854 9646 10906
rect 9646 10854 9692 10906
rect 9396 10852 9452 10854
rect 9476 10852 9532 10854
rect 9556 10852 9612 10854
rect 9636 10852 9692 10854
rect 9396 9818 9452 9820
rect 9476 9818 9532 9820
rect 9556 9818 9612 9820
rect 9636 9818 9692 9820
rect 9396 9766 9442 9818
rect 9442 9766 9452 9818
rect 9476 9766 9506 9818
rect 9506 9766 9518 9818
rect 9518 9766 9532 9818
rect 9556 9766 9570 9818
rect 9570 9766 9582 9818
rect 9582 9766 9612 9818
rect 9636 9766 9646 9818
rect 9646 9766 9692 9818
rect 9396 9764 9452 9766
rect 9476 9764 9532 9766
rect 9556 9764 9612 9766
rect 9636 9764 9692 9766
rect 9396 8730 9452 8732
rect 9476 8730 9532 8732
rect 9556 8730 9612 8732
rect 9636 8730 9692 8732
rect 9396 8678 9442 8730
rect 9442 8678 9452 8730
rect 9476 8678 9506 8730
rect 9506 8678 9518 8730
rect 9518 8678 9532 8730
rect 9556 8678 9570 8730
rect 9570 8678 9582 8730
rect 9582 8678 9612 8730
rect 9636 8678 9646 8730
rect 9646 8678 9692 8730
rect 9396 8676 9452 8678
rect 9476 8676 9532 8678
rect 9556 8676 9612 8678
rect 9636 8676 9692 8678
rect 9396 7642 9452 7644
rect 9476 7642 9532 7644
rect 9556 7642 9612 7644
rect 9636 7642 9692 7644
rect 9396 7590 9442 7642
rect 9442 7590 9452 7642
rect 9476 7590 9506 7642
rect 9506 7590 9518 7642
rect 9518 7590 9532 7642
rect 9556 7590 9570 7642
rect 9570 7590 9582 7642
rect 9582 7590 9612 7642
rect 9636 7590 9646 7642
rect 9646 7590 9692 7642
rect 9396 7588 9452 7590
rect 9476 7588 9532 7590
rect 9556 7588 9612 7590
rect 9636 7588 9692 7590
rect 9396 6554 9452 6556
rect 9476 6554 9532 6556
rect 9556 6554 9612 6556
rect 9636 6554 9692 6556
rect 9396 6502 9442 6554
rect 9442 6502 9452 6554
rect 9476 6502 9506 6554
rect 9506 6502 9518 6554
rect 9518 6502 9532 6554
rect 9556 6502 9570 6554
rect 9570 6502 9582 6554
rect 9582 6502 9612 6554
rect 9636 6502 9646 6554
rect 9646 6502 9692 6554
rect 9396 6500 9452 6502
rect 9476 6500 9532 6502
rect 9556 6500 9612 6502
rect 9636 6500 9692 6502
rect 9396 5466 9452 5468
rect 9476 5466 9532 5468
rect 9556 5466 9612 5468
rect 9636 5466 9692 5468
rect 9396 5414 9442 5466
rect 9442 5414 9452 5466
rect 9476 5414 9506 5466
rect 9506 5414 9518 5466
rect 9518 5414 9532 5466
rect 9556 5414 9570 5466
rect 9570 5414 9582 5466
rect 9582 5414 9612 5466
rect 9636 5414 9646 5466
rect 9646 5414 9692 5466
rect 9396 5412 9452 5414
rect 9476 5412 9532 5414
rect 9556 5412 9612 5414
rect 9636 5412 9692 5414
rect 9396 4378 9452 4380
rect 9476 4378 9532 4380
rect 9556 4378 9612 4380
rect 9636 4378 9692 4380
rect 9396 4326 9442 4378
rect 9442 4326 9452 4378
rect 9476 4326 9506 4378
rect 9506 4326 9518 4378
rect 9518 4326 9532 4378
rect 9556 4326 9570 4378
rect 9570 4326 9582 4378
rect 9582 4326 9612 4378
rect 9636 4326 9646 4378
rect 9646 4326 9692 4378
rect 9396 4324 9452 4326
rect 9476 4324 9532 4326
rect 9556 4324 9612 4326
rect 9636 4324 9692 4326
rect 9396 3290 9452 3292
rect 9476 3290 9532 3292
rect 9556 3290 9612 3292
rect 9636 3290 9692 3292
rect 9396 3238 9442 3290
rect 9442 3238 9452 3290
rect 9476 3238 9506 3290
rect 9506 3238 9518 3290
rect 9518 3238 9532 3290
rect 9556 3238 9570 3290
rect 9570 3238 9582 3290
rect 9582 3238 9612 3290
rect 9636 3238 9646 3290
rect 9646 3238 9692 3290
rect 9396 3236 9452 3238
rect 9476 3236 9532 3238
rect 9556 3236 9612 3238
rect 9636 3236 9692 3238
rect 13617 32122 13673 32124
rect 13697 32122 13753 32124
rect 13777 32122 13833 32124
rect 13857 32122 13913 32124
rect 13617 32070 13663 32122
rect 13663 32070 13673 32122
rect 13697 32070 13727 32122
rect 13727 32070 13739 32122
rect 13739 32070 13753 32122
rect 13777 32070 13791 32122
rect 13791 32070 13803 32122
rect 13803 32070 13833 32122
rect 13857 32070 13867 32122
rect 13867 32070 13913 32122
rect 13617 32068 13673 32070
rect 13697 32068 13753 32070
rect 13777 32068 13833 32070
rect 13857 32068 13913 32070
rect 13617 31034 13673 31036
rect 13697 31034 13753 31036
rect 13777 31034 13833 31036
rect 13857 31034 13913 31036
rect 13617 30982 13663 31034
rect 13663 30982 13673 31034
rect 13697 30982 13727 31034
rect 13727 30982 13739 31034
rect 13739 30982 13753 31034
rect 13777 30982 13791 31034
rect 13791 30982 13803 31034
rect 13803 30982 13833 31034
rect 13857 30982 13867 31034
rect 13867 30982 13913 31034
rect 13617 30980 13673 30982
rect 13697 30980 13753 30982
rect 13777 30980 13833 30982
rect 13857 30980 13913 30982
rect 13617 29946 13673 29948
rect 13697 29946 13753 29948
rect 13777 29946 13833 29948
rect 13857 29946 13913 29948
rect 13617 29894 13663 29946
rect 13663 29894 13673 29946
rect 13697 29894 13727 29946
rect 13727 29894 13739 29946
rect 13739 29894 13753 29946
rect 13777 29894 13791 29946
rect 13791 29894 13803 29946
rect 13803 29894 13833 29946
rect 13857 29894 13867 29946
rect 13867 29894 13913 29946
rect 13617 29892 13673 29894
rect 13697 29892 13753 29894
rect 13777 29892 13833 29894
rect 13857 29892 13913 29894
rect 13617 28858 13673 28860
rect 13697 28858 13753 28860
rect 13777 28858 13833 28860
rect 13857 28858 13913 28860
rect 13617 28806 13663 28858
rect 13663 28806 13673 28858
rect 13697 28806 13727 28858
rect 13727 28806 13739 28858
rect 13739 28806 13753 28858
rect 13777 28806 13791 28858
rect 13791 28806 13803 28858
rect 13803 28806 13833 28858
rect 13857 28806 13867 28858
rect 13867 28806 13913 28858
rect 13617 28804 13673 28806
rect 13697 28804 13753 28806
rect 13777 28804 13833 28806
rect 13857 28804 13913 28806
rect 13617 27770 13673 27772
rect 13697 27770 13753 27772
rect 13777 27770 13833 27772
rect 13857 27770 13913 27772
rect 13617 27718 13663 27770
rect 13663 27718 13673 27770
rect 13697 27718 13727 27770
rect 13727 27718 13739 27770
rect 13739 27718 13753 27770
rect 13777 27718 13791 27770
rect 13791 27718 13803 27770
rect 13803 27718 13833 27770
rect 13857 27718 13867 27770
rect 13867 27718 13913 27770
rect 13617 27716 13673 27718
rect 13697 27716 13753 27718
rect 13777 27716 13833 27718
rect 13857 27716 13913 27718
rect 13617 26682 13673 26684
rect 13697 26682 13753 26684
rect 13777 26682 13833 26684
rect 13857 26682 13913 26684
rect 13617 26630 13663 26682
rect 13663 26630 13673 26682
rect 13697 26630 13727 26682
rect 13727 26630 13739 26682
rect 13739 26630 13753 26682
rect 13777 26630 13791 26682
rect 13791 26630 13803 26682
rect 13803 26630 13833 26682
rect 13857 26630 13867 26682
rect 13867 26630 13913 26682
rect 13617 26628 13673 26630
rect 13697 26628 13753 26630
rect 13777 26628 13833 26630
rect 13857 26628 13913 26630
rect 13617 25594 13673 25596
rect 13697 25594 13753 25596
rect 13777 25594 13833 25596
rect 13857 25594 13913 25596
rect 13617 25542 13663 25594
rect 13663 25542 13673 25594
rect 13697 25542 13727 25594
rect 13727 25542 13739 25594
rect 13739 25542 13753 25594
rect 13777 25542 13791 25594
rect 13791 25542 13803 25594
rect 13803 25542 13833 25594
rect 13857 25542 13867 25594
rect 13867 25542 13913 25594
rect 13617 25540 13673 25542
rect 13697 25540 13753 25542
rect 13777 25540 13833 25542
rect 13857 25540 13913 25542
rect 13617 24506 13673 24508
rect 13697 24506 13753 24508
rect 13777 24506 13833 24508
rect 13857 24506 13913 24508
rect 13617 24454 13663 24506
rect 13663 24454 13673 24506
rect 13697 24454 13727 24506
rect 13727 24454 13739 24506
rect 13739 24454 13753 24506
rect 13777 24454 13791 24506
rect 13791 24454 13803 24506
rect 13803 24454 13833 24506
rect 13857 24454 13867 24506
rect 13867 24454 13913 24506
rect 13617 24452 13673 24454
rect 13697 24452 13753 24454
rect 13777 24452 13833 24454
rect 13857 24452 13913 24454
rect 13617 23418 13673 23420
rect 13697 23418 13753 23420
rect 13777 23418 13833 23420
rect 13857 23418 13913 23420
rect 13617 23366 13663 23418
rect 13663 23366 13673 23418
rect 13697 23366 13727 23418
rect 13727 23366 13739 23418
rect 13739 23366 13753 23418
rect 13777 23366 13791 23418
rect 13791 23366 13803 23418
rect 13803 23366 13833 23418
rect 13857 23366 13867 23418
rect 13867 23366 13913 23418
rect 13617 23364 13673 23366
rect 13697 23364 13753 23366
rect 13777 23364 13833 23366
rect 13857 23364 13913 23366
rect 13617 22330 13673 22332
rect 13697 22330 13753 22332
rect 13777 22330 13833 22332
rect 13857 22330 13913 22332
rect 13617 22278 13663 22330
rect 13663 22278 13673 22330
rect 13697 22278 13727 22330
rect 13727 22278 13739 22330
rect 13739 22278 13753 22330
rect 13777 22278 13791 22330
rect 13791 22278 13803 22330
rect 13803 22278 13833 22330
rect 13857 22278 13867 22330
rect 13867 22278 13913 22330
rect 13617 22276 13673 22278
rect 13697 22276 13753 22278
rect 13777 22276 13833 22278
rect 13857 22276 13913 22278
rect 13617 21242 13673 21244
rect 13697 21242 13753 21244
rect 13777 21242 13833 21244
rect 13857 21242 13913 21244
rect 13617 21190 13663 21242
rect 13663 21190 13673 21242
rect 13697 21190 13727 21242
rect 13727 21190 13739 21242
rect 13739 21190 13753 21242
rect 13777 21190 13791 21242
rect 13791 21190 13803 21242
rect 13803 21190 13833 21242
rect 13857 21190 13867 21242
rect 13867 21190 13913 21242
rect 13617 21188 13673 21190
rect 13697 21188 13753 21190
rect 13777 21188 13833 21190
rect 13857 21188 13913 21190
rect 13617 20154 13673 20156
rect 13697 20154 13753 20156
rect 13777 20154 13833 20156
rect 13857 20154 13913 20156
rect 13617 20102 13663 20154
rect 13663 20102 13673 20154
rect 13697 20102 13727 20154
rect 13727 20102 13739 20154
rect 13739 20102 13753 20154
rect 13777 20102 13791 20154
rect 13791 20102 13803 20154
rect 13803 20102 13833 20154
rect 13857 20102 13867 20154
rect 13867 20102 13913 20154
rect 13617 20100 13673 20102
rect 13697 20100 13753 20102
rect 13777 20100 13833 20102
rect 13857 20100 13913 20102
rect 13617 19066 13673 19068
rect 13697 19066 13753 19068
rect 13777 19066 13833 19068
rect 13857 19066 13913 19068
rect 13617 19014 13663 19066
rect 13663 19014 13673 19066
rect 13697 19014 13727 19066
rect 13727 19014 13739 19066
rect 13739 19014 13753 19066
rect 13777 19014 13791 19066
rect 13791 19014 13803 19066
rect 13803 19014 13833 19066
rect 13857 19014 13867 19066
rect 13867 19014 13913 19066
rect 13617 19012 13673 19014
rect 13697 19012 13753 19014
rect 13777 19012 13833 19014
rect 13857 19012 13913 19014
rect 13617 17978 13673 17980
rect 13697 17978 13753 17980
rect 13777 17978 13833 17980
rect 13857 17978 13913 17980
rect 13617 17926 13663 17978
rect 13663 17926 13673 17978
rect 13697 17926 13727 17978
rect 13727 17926 13739 17978
rect 13739 17926 13753 17978
rect 13777 17926 13791 17978
rect 13791 17926 13803 17978
rect 13803 17926 13833 17978
rect 13857 17926 13867 17978
rect 13867 17926 13913 17978
rect 13617 17924 13673 17926
rect 13697 17924 13753 17926
rect 13777 17924 13833 17926
rect 13857 17924 13913 17926
rect 13617 16890 13673 16892
rect 13697 16890 13753 16892
rect 13777 16890 13833 16892
rect 13857 16890 13913 16892
rect 13617 16838 13663 16890
rect 13663 16838 13673 16890
rect 13697 16838 13727 16890
rect 13727 16838 13739 16890
rect 13739 16838 13753 16890
rect 13777 16838 13791 16890
rect 13791 16838 13803 16890
rect 13803 16838 13833 16890
rect 13857 16838 13867 16890
rect 13867 16838 13913 16890
rect 13617 16836 13673 16838
rect 13697 16836 13753 16838
rect 13777 16836 13833 16838
rect 13857 16836 13913 16838
rect 13617 15802 13673 15804
rect 13697 15802 13753 15804
rect 13777 15802 13833 15804
rect 13857 15802 13913 15804
rect 13617 15750 13663 15802
rect 13663 15750 13673 15802
rect 13697 15750 13727 15802
rect 13727 15750 13739 15802
rect 13739 15750 13753 15802
rect 13777 15750 13791 15802
rect 13791 15750 13803 15802
rect 13803 15750 13833 15802
rect 13857 15750 13867 15802
rect 13867 15750 13913 15802
rect 13617 15748 13673 15750
rect 13697 15748 13753 15750
rect 13777 15748 13833 15750
rect 13857 15748 13913 15750
rect 13617 14714 13673 14716
rect 13697 14714 13753 14716
rect 13777 14714 13833 14716
rect 13857 14714 13913 14716
rect 13617 14662 13663 14714
rect 13663 14662 13673 14714
rect 13697 14662 13727 14714
rect 13727 14662 13739 14714
rect 13739 14662 13753 14714
rect 13777 14662 13791 14714
rect 13791 14662 13803 14714
rect 13803 14662 13833 14714
rect 13857 14662 13867 14714
rect 13867 14662 13913 14714
rect 13617 14660 13673 14662
rect 13697 14660 13753 14662
rect 13777 14660 13833 14662
rect 13857 14660 13913 14662
rect 13617 13626 13673 13628
rect 13697 13626 13753 13628
rect 13777 13626 13833 13628
rect 13857 13626 13913 13628
rect 13617 13574 13663 13626
rect 13663 13574 13673 13626
rect 13697 13574 13727 13626
rect 13727 13574 13739 13626
rect 13739 13574 13753 13626
rect 13777 13574 13791 13626
rect 13791 13574 13803 13626
rect 13803 13574 13833 13626
rect 13857 13574 13867 13626
rect 13867 13574 13913 13626
rect 13617 13572 13673 13574
rect 13697 13572 13753 13574
rect 13777 13572 13833 13574
rect 13857 13572 13913 13574
rect 13617 12538 13673 12540
rect 13697 12538 13753 12540
rect 13777 12538 13833 12540
rect 13857 12538 13913 12540
rect 13617 12486 13663 12538
rect 13663 12486 13673 12538
rect 13697 12486 13727 12538
rect 13727 12486 13739 12538
rect 13739 12486 13753 12538
rect 13777 12486 13791 12538
rect 13791 12486 13803 12538
rect 13803 12486 13833 12538
rect 13857 12486 13867 12538
rect 13867 12486 13913 12538
rect 13617 12484 13673 12486
rect 13697 12484 13753 12486
rect 13777 12484 13833 12486
rect 13857 12484 13913 12486
rect 17837 32666 17893 32668
rect 17917 32666 17973 32668
rect 17997 32666 18053 32668
rect 18077 32666 18133 32668
rect 17837 32614 17883 32666
rect 17883 32614 17893 32666
rect 17917 32614 17947 32666
rect 17947 32614 17959 32666
rect 17959 32614 17973 32666
rect 17997 32614 18011 32666
rect 18011 32614 18023 32666
rect 18023 32614 18053 32666
rect 18077 32614 18087 32666
rect 18087 32614 18133 32666
rect 17837 32612 17893 32614
rect 17917 32612 17973 32614
rect 17997 32612 18053 32614
rect 18077 32612 18133 32614
rect 13617 11450 13673 11452
rect 13697 11450 13753 11452
rect 13777 11450 13833 11452
rect 13857 11450 13913 11452
rect 13617 11398 13663 11450
rect 13663 11398 13673 11450
rect 13697 11398 13727 11450
rect 13727 11398 13739 11450
rect 13739 11398 13753 11450
rect 13777 11398 13791 11450
rect 13791 11398 13803 11450
rect 13803 11398 13833 11450
rect 13857 11398 13867 11450
rect 13867 11398 13913 11450
rect 13617 11396 13673 11398
rect 13697 11396 13753 11398
rect 13777 11396 13833 11398
rect 13857 11396 13913 11398
rect 16118 12416 16174 12472
rect 13617 10362 13673 10364
rect 13697 10362 13753 10364
rect 13777 10362 13833 10364
rect 13857 10362 13913 10364
rect 13617 10310 13663 10362
rect 13663 10310 13673 10362
rect 13697 10310 13727 10362
rect 13727 10310 13739 10362
rect 13739 10310 13753 10362
rect 13777 10310 13791 10362
rect 13791 10310 13803 10362
rect 13803 10310 13833 10362
rect 13857 10310 13867 10362
rect 13867 10310 13913 10362
rect 13617 10308 13673 10310
rect 13697 10308 13753 10310
rect 13777 10308 13833 10310
rect 13857 10308 13913 10310
rect 13617 9274 13673 9276
rect 13697 9274 13753 9276
rect 13777 9274 13833 9276
rect 13857 9274 13913 9276
rect 13617 9222 13663 9274
rect 13663 9222 13673 9274
rect 13697 9222 13727 9274
rect 13727 9222 13739 9274
rect 13739 9222 13753 9274
rect 13777 9222 13791 9274
rect 13791 9222 13803 9274
rect 13803 9222 13833 9274
rect 13857 9222 13867 9274
rect 13867 9222 13913 9274
rect 13617 9220 13673 9222
rect 13697 9220 13753 9222
rect 13777 9220 13833 9222
rect 13857 9220 13913 9222
rect 13617 8186 13673 8188
rect 13697 8186 13753 8188
rect 13777 8186 13833 8188
rect 13857 8186 13913 8188
rect 13617 8134 13663 8186
rect 13663 8134 13673 8186
rect 13697 8134 13727 8186
rect 13727 8134 13739 8186
rect 13739 8134 13753 8186
rect 13777 8134 13791 8186
rect 13791 8134 13803 8186
rect 13803 8134 13833 8186
rect 13857 8134 13867 8186
rect 13867 8134 13913 8186
rect 13617 8132 13673 8134
rect 13697 8132 13753 8134
rect 13777 8132 13833 8134
rect 13857 8132 13913 8134
rect 13617 7098 13673 7100
rect 13697 7098 13753 7100
rect 13777 7098 13833 7100
rect 13857 7098 13913 7100
rect 13617 7046 13663 7098
rect 13663 7046 13673 7098
rect 13697 7046 13727 7098
rect 13727 7046 13739 7098
rect 13739 7046 13753 7098
rect 13777 7046 13791 7098
rect 13791 7046 13803 7098
rect 13803 7046 13833 7098
rect 13857 7046 13867 7098
rect 13867 7046 13913 7098
rect 13617 7044 13673 7046
rect 13697 7044 13753 7046
rect 13777 7044 13833 7046
rect 13857 7044 13913 7046
rect 13617 6010 13673 6012
rect 13697 6010 13753 6012
rect 13777 6010 13833 6012
rect 13857 6010 13913 6012
rect 13617 5958 13663 6010
rect 13663 5958 13673 6010
rect 13697 5958 13727 6010
rect 13727 5958 13739 6010
rect 13739 5958 13753 6010
rect 13777 5958 13791 6010
rect 13791 5958 13803 6010
rect 13803 5958 13833 6010
rect 13857 5958 13867 6010
rect 13867 5958 13913 6010
rect 13617 5956 13673 5958
rect 13697 5956 13753 5958
rect 13777 5956 13833 5958
rect 13857 5956 13913 5958
rect 13617 4922 13673 4924
rect 13697 4922 13753 4924
rect 13777 4922 13833 4924
rect 13857 4922 13913 4924
rect 13617 4870 13663 4922
rect 13663 4870 13673 4922
rect 13697 4870 13727 4922
rect 13727 4870 13739 4922
rect 13739 4870 13753 4922
rect 13777 4870 13791 4922
rect 13791 4870 13803 4922
rect 13803 4870 13833 4922
rect 13857 4870 13867 4922
rect 13867 4870 13913 4922
rect 13617 4868 13673 4870
rect 13697 4868 13753 4870
rect 13777 4868 13833 4870
rect 13857 4868 13913 4870
rect 13617 3834 13673 3836
rect 13697 3834 13753 3836
rect 13777 3834 13833 3836
rect 13857 3834 13913 3836
rect 13617 3782 13663 3834
rect 13663 3782 13673 3834
rect 13697 3782 13727 3834
rect 13727 3782 13739 3834
rect 13739 3782 13753 3834
rect 13777 3782 13791 3834
rect 13791 3782 13803 3834
rect 13803 3782 13833 3834
rect 13857 3782 13867 3834
rect 13867 3782 13913 3834
rect 13617 3780 13673 3782
rect 13697 3780 13753 3782
rect 13777 3780 13833 3782
rect 13857 3780 13913 3782
rect 13617 2746 13673 2748
rect 13697 2746 13753 2748
rect 13777 2746 13833 2748
rect 13857 2746 13913 2748
rect 13617 2694 13663 2746
rect 13663 2694 13673 2746
rect 13697 2694 13727 2746
rect 13727 2694 13739 2746
rect 13739 2694 13753 2746
rect 13777 2694 13791 2746
rect 13791 2694 13803 2746
rect 13803 2694 13833 2746
rect 13857 2694 13867 2746
rect 13867 2694 13913 2746
rect 13617 2692 13673 2694
rect 13697 2692 13753 2694
rect 13777 2692 13833 2694
rect 13857 2692 13913 2694
rect 9396 2202 9452 2204
rect 9476 2202 9532 2204
rect 9556 2202 9612 2204
rect 9636 2202 9692 2204
rect 9396 2150 9442 2202
rect 9442 2150 9452 2202
rect 9476 2150 9506 2202
rect 9506 2150 9518 2202
rect 9518 2150 9532 2202
rect 9556 2150 9570 2202
rect 9570 2150 9582 2202
rect 9582 2150 9612 2202
rect 9636 2150 9646 2202
rect 9646 2150 9692 2202
rect 9396 2148 9452 2150
rect 9476 2148 9532 2150
rect 9556 2148 9612 2150
rect 9636 2148 9692 2150
rect 22058 33210 22114 33212
rect 22138 33210 22194 33212
rect 22218 33210 22274 33212
rect 22298 33210 22354 33212
rect 22058 33158 22104 33210
rect 22104 33158 22114 33210
rect 22138 33158 22168 33210
rect 22168 33158 22180 33210
rect 22180 33158 22194 33210
rect 22218 33158 22232 33210
rect 22232 33158 22244 33210
rect 22244 33158 22274 33210
rect 22298 33158 22308 33210
rect 22308 33158 22354 33210
rect 22058 33156 22114 33158
rect 22138 33156 22194 33158
rect 22218 33156 22274 33158
rect 22298 33156 22354 33158
rect 17837 31578 17893 31580
rect 17917 31578 17973 31580
rect 17997 31578 18053 31580
rect 18077 31578 18133 31580
rect 17837 31526 17883 31578
rect 17883 31526 17893 31578
rect 17917 31526 17947 31578
rect 17947 31526 17959 31578
rect 17959 31526 17973 31578
rect 17997 31526 18011 31578
rect 18011 31526 18023 31578
rect 18023 31526 18053 31578
rect 18077 31526 18087 31578
rect 18087 31526 18133 31578
rect 17837 31524 17893 31526
rect 17917 31524 17973 31526
rect 17997 31524 18053 31526
rect 18077 31524 18133 31526
rect 17837 30490 17893 30492
rect 17917 30490 17973 30492
rect 17997 30490 18053 30492
rect 18077 30490 18133 30492
rect 17837 30438 17883 30490
rect 17883 30438 17893 30490
rect 17917 30438 17947 30490
rect 17947 30438 17959 30490
rect 17959 30438 17973 30490
rect 17997 30438 18011 30490
rect 18011 30438 18023 30490
rect 18023 30438 18053 30490
rect 18077 30438 18087 30490
rect 18087 30438 18133 30490
rect 17837 30436 17893 30438
rect 17917 30436 17973 30438
rect 17997 30436 18053 30438
rect 18077 30436 18133 30438
rect 22058 32122 22114 32124
rect 22138 32122 22194 32124
rect 22218 32122 22274 32124
rect 22298 32122 22354 32124
rect 22058 32070 22104 32122
rect 22104 32070 22114 32122
rect 22138 32070 22168 32122
rect 22168 32070 22180 32122
rect 22180 32070 22194 32122
rect 22218 32070 22232 32122
rect 22232 32070 22244 32122
rect 22244 32070 22274 32122
rect 22298 32070 22308 32122
rect 22308 32070 22354 32122
rect 22058 32068 22114 32070
rect 22138 32068 22194 32070
rect 22218 32068 22274 32070
rect 22298 32068 22354 32070
rect 30499 33210 30555 33212
rect 30579 33210 30635 33212
rect 30659 33210 30715 33212
rect 30739 33210 30795 33212
rect 30499 33158 30545 33210
rect 30545 33158 30555 33210
rect 30579 33158 30609 33210
rect 30609 33158 30621 33210
rect 30621 33158 30635 33210
rect 30659 33158 30673 33210
rect 30673 33158 30685 33210
rect 30685 33158 30715 33210
rect 30739 33158 30749 33210
rect 30749 33158 30795 33210
rect 30499 33156 30555 33158
rect 30579 33156 30635 33158
rect 30659 33156 30715 33158
rect 30739 33156 30795 33158
rect 26278 32666 26334 32668
rect 26358 32666 26414 32668
rect 26438 32666 26494 32668
rect 26518 32666 26574 32668
rect 26278 32614 26324 32666
rect 26324 32614 26334 32666
rect 26358 32614 26388 32666
rect 26388 32614 26400 32666
rect 26400 32614 26414 32666
rect 26438 32614 26452 32666
rect 26452 32614 26464 32666
rect 26464 32614 26494 32666
rect 26518 32614 26528 32666
rect 26528 32614 26574 32666
rect 26278 32612 26334 32614
rect 26358 32612 26414 32614
rect 26438 32612 26494 32614
rect 26518 32612 26574 32614
rect 34719 32666 34775 32668
rect 34799 32666 34855 32668
rect 34879 32666 34935 32668
rect 34959 32666 35015 32668
rect 34719 32614 34765 32666
rect 34765 32614 34775 32666
rect 34799 32614 34829 32666
rect 34829 32614 34841 32666
rect 34841 32614 34855 32666
rect 34879 32614 34893 32666
rect 34893 32614 34905 32666
rect 34905 32614 34935 32666
rect 34959 32614 34969 32666
rect 34969 32614 35015 32666
rect 34719 32612 34775 32614
rect 34799 32612 34855 32614
rect 34879 32612 34935 32614
rect 34959 32612 35015 32614
rect 17837 29402 17893 29404
rect 17917 29402 17973 29404
rect 17997 29402 18053 29404
rect 18077 29402 18133 29404
rect 17837 29350 17883 29402
rect 17883 29350 17893 29402
rect 17917 29350 17947 29402
rect 17947 29350 17959 29402
rect 17959 29350 17973 29402
rect 17997 29350 18011 29402
rect 18011 29350 18023 29402
rect 18023 29350 18053 29402
rect 18077 29350 18087 29402
rect 18087 29350 18133 29402
rect 17837 29348 17893 29350
rect 17917 29348 17973 29350
rect 17997 29348 18053 29350
rect 18077 29348 18133 29350
rect 17837 28314 17893 28316
rect 17917 28314 17973 28316
rect 17997 28314 18053 28316
rect 18077 28314 18133 28316
rect 17837 28262 17883 28314
rect 17883 28262 17893 28314
rect 17917 28262 17947 28314
rect 17947 28262 17959 28314
rect 17959 28262 17973 28314
rect 17997 28262 18011 28314
rect 18011 28262 18023 28314
rect 18023 28262 18053 28314
rect 18077 28262 18087 28314
rect 18087 28262 18133 28314
rect 17837 28260 17893 28262
rect 17917 28260 17973 28262
rect 17997 28260 18053 28262
rect 18077 28260 18133 28262
rect 17837 27226 17893 27228
rect 17917 27226 17973 27228
rect 17997 27226 18053 27228
rect 18077 27226 18133 27228
rect 17837 27174 17883 27226
rect 17883 27174 17893 27226
rect 17917 27174 17947 27226
rect 17947 27174 17959 27226
rect 17959 27174 17973 27226
rect 17997 27174 18011 27226
rect 18011 27174 18023 27226
rect 18023 27174 18053 27226
rect 18077 27174 18087 27226
rect 18087 27174 18133 27226
rect 17837 27172 17893 27174
rect 17917 27172 17973 27174
rect 17997 27172 18053 27174
rect 18077 27172 18133 27174
rect 17837 26138 17893 26140
rect 17917 26138 17973 26140
rect 17997 26138 18053 26140
rect 18077 26138 18133 26140
rect 17837 26086 17883 26138
rect 17883 26086 17893 26138
rect 17917 26086 17947 26138
rect 17947 26086 17959 26138
rect 17959 26086 17973 26138
rect 17997 26086 18011 26138
rect 18011 26086 18023 26138
rect 18023 26086 18053 26138
rect 18077 26086 18087 26138
rect 18087 26086 18133 26138
rect 17837 26084 17893 26086
rect 17917 26084 17973 26086
rect 17997 26084 18053 26086
rect 18077 26084 18133 26086
rect 17837 25050 17893 25052
rect 17917 25050 17973 25052
rect 17997 25050 18053 25052
rect 18077 25050 18133 25052
rect 17837 24998 17883 25050
rect 17883 24998 17893 25050
rect 17917 24998 17947 25050
rect 17947 24998 17959 25050
rect 17959 24998 17973 25050
rect 17997 24998 18011 25050
rect 18011 24998 18023 25050
rect 18023 24998 18053 25050
rect 18077 24998 18087 25050
rect 18087 24998 18133 25050
rect 17837 24996 17893 24998
rect 17917 24996 17973 24998
rect 17997 24996 18053 24998
rect 18077 24996 18133 24998
rect 17837 23962 17893 23964
rect 17917 23962 17973 23964
rect 17997 23962 18053 23964
rect 18077 23962 18133 23964
rect 17837 23910 17883 23962
rect 17883 23910 17893 23962
rect 17917 23910 17947 23962
rect 17947 23910 17959 23962
rect 17959 23910 17973 23962
rect 17997 23910 18011 23962
rect 18011 23910 18023 23962
rect 18023 23910 18053 23962
rect 18077 23910 18087 23962
rect 18087 23910 18133 23962
rect 17837 23908 17893 23910
rect 17917 23908 17973 23910
rect 17997 23908 18053 23910
rect 18077 23908 18133 23910
rect 17837 22874 17893 22876
rect 17917 22874 17973 22876
rect 17997 22874 18053 22876
rect 18077 22874 18133 22876
rect 17837 22822 17883 22874
rect 17883 22822 17893 22874
rect 17917 22822 17947 22874
rect 17947 22822 17959 22874
rect 17959 22822 17973 22874
rect 17997 22822 18011 22874
rect 18011 22822 18023 22874
rect 18023 22822 18053 22874
rect 18077 22822 18087 22874
rect 18087 22822 18133 22874
rect 17837 22820 17893 22822
rect 17917 22820 17973 22822
rect 17997 22820 18053 22822
rect 18077 22820 18133 22822
rect 17837 21786 17893 21788
rect 17917 21786 17973 21788
rect 17997 21786 18053 21788
rect 18077 21786 18133 21788
rect 17837 21734 17883 21786
rect 17883 21734 17893 21786
rect 17917 21734 17947 21786
rect 17947 21734 17959 21786
rect 17959 21734 17973 21786
rect 17997 21734 18011 21786
rect 18011 21734 18023 21786
rect 18023 21734 18053 21786
rect 18077 21734 18087 21786
rect 18087 21734 18133 21786
rect 17837 21732 17893 21734
rect 17917 21732 17973 21734
rect 17997 21732 18053 21734
rect 18077 21732 18133 21734
rect 19706 23840 19762 23896
rect 20718 23840 20774 23896
rect 17837 20698 17893 20700
rect 17917 20698 17973 20700
rect 17997 20698 18053 20700
rect 18077 20698 18133 20700
rect 17837 20646 17883 20698
rect 17883 20646 17893 20698
rect 17917 20646 17947 20698
rect 17947 20646 17959 20698
rect 17959 20646 17973 20698
rect 17997 20646 18011 20698
rect 18011 20646 18023 20698
rect 18023 20646 18053 20698
rect 18077 20646 18087 20698
rect 18087 20646 18133 20698
rect 17837 20644 17893 20646
rect 17917 20644 17973 20646
rect 17997 20644 18053 20646
rect 18077 20644 18133 20646
rect 17837 19610 17893 19612
rect 17917 19610 17973 19612
rect 17997 19610 18053 19612
rect 18077 19610 18133 19612
rect 17837 19558 17883 19610
rect 17883 19558 17893 19610
rect 17917 19558 17947 19610
rect 17947 19558 17959 19610
rect 17959 19558 17973 19610
rect 17997 19558 18011 19610
rect 18011 19558 18023 19610
rect 18023 19558 18053 19610
rect 18077 19558 18087 19610
rect 18087 19558 18133 19610
rect 17837 19556 17893 19558
rect 17917 19556 17973 19558
rect 17997 19556 18053 19558
rect 18077 19556 18133 19558
rect 17837 18522 17893 18524
rect 17917 18522 17973 18524
rect 17997 18522 18053 18524
rect 18077 18522 18133 18524
rect 17837 18470 17883 18522
rect 17883 18470 17893 18522
rect 17917 18470 17947 18522
rect 17947 18470 17959 18522
rect 17959 18470 17973 18522
rect 17997 18470 18011 18522
rect 18011 18470 18023 18522
rect 18023 18470 18053 18522
rect 18077 18470 18087 18522
rect 18087 18470 18133 18522
rect 17837 18468 17893 18470
rect 17917 18468 17973 18470
rect 17997 18468 18053 18470
rect 18077 18468 18133 18470
rect 17837 17434 17893 17436
rect 17917 17434 17973 17436
rect 17997 17434 18053 17436
rect 18077 17434 18133 17436
rect 17837 17382 17883 17434
rect 17883 17382 17893 17434
rect 17917 17382 17947 17434
rect 17947 17382 17959 17434
rect 17959 17382 17973 17434
rect 17997 17382 18011 17434
rect 18011 17382 18023 17434
rect 18023 17382 18053 17434
rect 18077 17382 18087 17434
rect 18087 17382 18133 17434
rect 17837 17380 17893 17382
rect 17917 17380 17973 17382
rect 17997 17380 18053 17382
rect 18077 17380 18133 17382
rect 17837 16346 17893 16348
rect 17917 16346 17973 16348
rect 17997 16346 18053 16348
rect 18077 16346 18133 16348
rect 17837 16294 17883 16346
rect 17883 16294 17893 16346
rect 17917 16294 17947 16346
rect 17947 16294 17959 16346
rect 17959 16294 17973 16346
rect 17997 16294 18011 16346
rect 18011 16294 18023 16346
rect 18023 16294 18053 16346
rect 18077 16294 18087 16346
rect 18087 16294 18133 16346
rect 17837 16292 17893 16294
rect 17917 16292 17973 16294
rect 17997 16292 18053 16294
rect 18077 16292 18133 16294
rect 17837 15258 17893 15260
rect 17917 15258 17973 15260
rect 17997 15258 18053 15260
rect 18077 15258 18133 15260
rect 17837 15206 17883 15258
rect 17883 15206 17893 15258
rect 17917 15206 17947 15258
rect 17947 15206 17959 15258
rect 17959 15206 17973 15258
rect 17997 15206 18011 15258
rect 18011 15206 18023 15258
rect 18023 15206 18053 15258
rect 18077 15206 18087 15258
rect 18087 15206 18133 15258
rect 17837 15204 17893 15206
rect 17917 15204 17973 15206
rect 17997 15204 18053 15206
rect 18077 15204 18133 15206
rect 17837 14170 17893 14172
rect 17917 14170 17973 14172
rect 17997 14170 18053 14172
rect 18077 14170 18133 14172
rect 17837 14118 17883 14170
rect 17883 14118 17893 14170
rect 17917 14118 17947 14170
rect 17947 14118 17959 14170
rect 17959 14118 17973 14170
rect 17997 14118 18011 14170
rect 18011 14118 18023 14170
rect 18023 14118 18053 14170
rect 18077 14118 18087 14170
rect 18087 14118 18133 14170
rect 17837 14116 17893 14118
rect 17917 14116 17973 14118
rect 17997 14116 18053 14118
rect 18077 14116 18133 14118
rect 20442 22092 20498 22128
rect 20442 22072 20444 22092
rect 20444 22072 20496 22092
rect 20496 22072 20498 22092
rect 19522 14320 19578 14376
rect 19890 14900 19892 14920
rect 19892 14900 19944 14920
rect 19944 14900 19946 14920
rect 19890 14864 19946 14900
rect 17837 13082 17893 13084
rect 17917 13082 17973 13084
rect 17997 13082 18053 13084
rect 18077 13082 18133 13084
rect 17837 13030 17883 13082
rect 17883 13030 17893 13082
rect 17917 13030 17947 13082
rect 17947 13030 17959 13082
rect 17959 13030 17973 13082
rect 17997 13030 18011 13082
rect 18011 13030 18023 13082
rect 18023 13030 18053 13082
rect 18077 13030 18087 13082
rect 18087 13030 18133 13082
rect 17837 13028 17893 13030
rect 17917 13028 17973 13030
rect 17997 13028 18053 13030
rect 18077 13028 18133 13030
rect 17837 11994 17893 11996
rect 17917 11994 17973 11996
rect 17997 11994 18053 11996
rect 18077 11994 18133 11996
rect 17837 11942 17883 11994
rect 17883 11942 17893 11994
rect 17917 11942 17947 11994
rect 17947 11942 17959 11994
rect 17959 11942 17973 11994
rect 17997 11942 18011 11994
rect 18011 11942 18023 11994
rect 18023 11942 18053 11994
rect 18077 11942 18087 11994
rect 18087 11942 18133 11994
rect 17837 11940 17893 11942
rect 17917 11940 17973 11942
rect 17997 11940 18053 11942
rect 18077 11940 18133 11942
rect 17837 10906 17893 10908
rect 17917 10906 17973 10908
rect 17997 10906 18053 10908
rect 18077 10906 18133 10908
rect 17837 10854 17883 10906
rect 17883 10854 17893 10906
rect 17917 10854 17947 10906
rect 17947 10854 17959 10906
rect 17959 10854 17973 10906
rect 17997 10854 18011 10906
rect 18011 10854 18023 10906
rect 18023 10854 18053 10906
rect 18077 10854 18087 10906
rect 18087 10854 18133 10906
rect 17837 10852 17893 10854
rect 17917 10852 17973 10854
rect 17997 10852 18053 10854
rect 18077 10852 18133 10854
rect 19338 12416 19394 12472
rect 17837 9818 17893 9820
rect 17917 9818 17973 9820
rect 17997 9818 18053 9820
rect 18077 9818 18133 9820
rect 17837 9766 17883 9818
rect 17883 9766 17893 9818
rect 17917 9766 17947 9818
rect 17947 9766 17959 9818
rect 17959 9766 17973 9818
rect 17997 9766 18011 9818
rect 18011 9766 18023 9818
rect 18023 9766 18053 9818
rect 18077 9766 18087 9818
rect 18087 9766 18133 9818
rect 17837 9764 17893 9766
rect 17917 9764 17973 9766
rect 17997 9764 18053 9766
rect 18077 9764 18133 9766
rect 17837 8730 17893 8732
rect 17917 8730 17973 8732
rect 17997 8730 18053 8732
rect 18077 8730 18133 8732
rect 17837 8678 17883 8730
rect 17883 8678 17893 8730
rect 17917 8678 17947 8730
rect 17947 8678 17959 8730
rect 17959 8678 17973 8730
rect 17997 8678 18011 8730
rect 18011 8678 18023 8730
rect 18023 8678 18053 8730
rect 18077 8678 18087 8730
rect 18087 8678 18133 8730
rect 17837 8676 17893 8678
rect 17917 8676 17973 8678
rect 17997 8676 18053 8678
rect 18077 8676 18133 8678
rect 19798 13912 19854 13968
rect 17837 7642 17893 7644
rect 17917 7642 17973 7644
rect 17997 7642 18053 7644
rect 18077 7642 18133 7644
rect 17837 7590 17883 7642
rect 17883 7590 17893 7642
rect 17917 7590 17947 7642
rect 17947 7590 17959 7642
rect 17959 7590 17973 7642
rect 17997 7590 18011 7642
rect 18011 7590 18023 7642
rect 18023 7590 18053 7642
rect 18077 7590 18087 7642
rect 18087 7590 18133 7642
rect 17837 7588 17893 7590
rect 17917 7588 17973 7590
rect 17997 7588 18053 7590
rect 18077 7588 18133 7590
rect 17837 6554 17893 6556
rect 17917 6554 17973 6556
rect 17997 6554 18053 6556
rect 18077 6554 18133 6556
rect 17837 6502 17883 6554
rect 17883 6502 17893 6554
rect 17917 6502 17947 6554
rect 17947 6502 17959 6554
rect 17959 6502 17973 6554
rect 17997 6502 18011 6554
rect 18011 6502 18023 6554
rect 18023 6502 18053 6554
rect 18077 6502 18087 6554
rect 18087 6502 18133 6554
rect 17837 6500 17893 6502
rect 17917 6500 17973 6502
rect 17997 6500 18053 6502
rect 18077 6500 18133 6502
rect 17837 5466 17893 5468
rect 17917 5466 17973 5468
rect 17997 5466 18053 5468
rect 18077 5466 18133 5468
rect 17837 5414 17883 5466
rect 17883 5414 17893 5466
rect 17917 5414 17947 5466
rect 17947 5414 17959 5466
rect 17959 5414 17973 5466
rect 17997 5414 18011 5466
rect 18011 5414 18023 5466
rect 18023 5414 18053 5466
rect 18077 5414 18087 5466
rect 18087 5414 18133 5466
rect 17837 5412 17893 5414
rect 17917 5412 17973 5414
rect 17997 5412 18053 5414
rect 18077 5412 18133 5414
rect 22058 31034 22114 31036
rect 22138 31034 22194 31036
rect 22218 31034 22274 31036
rect 22298 31034 22354 31036
rect 22058 30982 22104 31034
rect 22104 30982 22114 31034
rect 22138 30982 22168 31034
rect 22168 30982 22180 31034
rect 22180 30982 22194 31034
rect 22218 30982 22232 31034
rect 22232 30982 22244 31034
rect 22244 30982 22274 31034
rect 22298 30982 22308 31034
rect 22308 30982 22354 31034
rect 22058 30980 22114 30982
rect 22138 30980 22194 30982
rect 22218 30980 22274 30982
rect 22298 30980 22354 30982
rect 22058 29946 22114 29948
rect 22138 29946 22194 29948
rect 22218 29946 22274 29948
rect 22298 29946 22354 29948
rect 22058 29894 22104 29946
rect 22104 29894 22114 29946
rect 22138 29894 22168 29946
rect 22168 29894 22180 29946
rect 22180 29894 22194 29946
rect 22218 29894 22232 29946
rect 22232 29894 22244 29946
rect 22244 29894 22274 29946
rect 22298 29894 22308 29946
rect 22308 29894 22354 29946
rect 22058 29892 22114 29894
rect 22138 29892 22194 29894
rect 22218 29892 22274 29894
rect 22298 29892 22354 29894
rect 22058 28858 22114 28860
rect 22138 28858 22194 28860
rect 22218 28858 22274 28860
rect 22298 28858 22354 28860
rect 22058 28806 22104 28858
rect 22104 28806 22114 28858
rect 22138 28806 22168 28858
rect 22168 28806 22180 28858
rect 22180 28806 22194 28858
rect 22218 28806 22232 28858
rect 22232 28806 22244 28858
rect 22244 28806 22274 28858
rect 22298 28806 22308 28858
rect 22308 28806 22354 28858
rect 22058 28804 22114 28806
rect 22138 28804 22194 28806
rect 22218 28804 22274 28806
rect 22298 28804 22354 28806
rect 22058 27770 22114 27772
rect 22138 27770 22194 27772
rect 22218 27770 22274 27772
rect 22298 27770 22354 27772
rect 22058 27718 22104 27770
rect 22104 27718 22114 27770
rect 22138 27718 22168 27770
rect 22168 27718 22180 27770
rect 22180 27718 22194 27770
rect 22218 27718 22232 27770
rect 22232 27718 22244 27770
rect 22244 27718 22274 27770
rect 22298 27718 22308 27770
rect 22308 27718 22354 27770
rect 22058 27716 22114 27718
rect 22138 27716 22194 27718
rect 22218 27716 22274 27718
rect 22298 27716 22354 27718
rect 22058 26682 22114 26684
rect 22138 26682 22194 26684
rect 22218 26682 22274 26684
rect 22298 26682 22354 26684
rect 22058 26630 22104 26682
rect 22104 26630 22114 26682
rect 22138 26630 22168 26682
rect 22168 26630 22180 26682
rect 22180 26630 22194 26682
rect 22218 26630 22232 26682
rect 22232 26630 22244 26682
rect 22244 26630 22274 26682
rect 22298 26630 22308 26682
rect 22308 26630 22354 26682
rect 22058 26628 22114 26630
rect 22138 26628 22194 26630
rect 22218 26628 22274 26630
rect 22298 26628 22354 26630
rect 26278 31578 26334 31580
rect 26358 31578 26414 31580
rect 26438 31578 26494 31580
rect 26518 31578 26574 31580
rect 26278 31526 26324 31578
rect 26324 31526 26334 31578
rect 26358 31526 26388 31578
rect 26388 31526 26400 31578
rect 26400 31526 26414 31578
rect 26438 31526 26452 31578
rect 26452 31526 26464 31578
rect 26464 31526 26494 31578
rect 26518 31526 26528 31578
rect 26528 31526 26574 31578
rect 26278 31524 26334 31526
rect 26358 31524 26414 31526
rect 26438 31524 26494 31526
rect 26518 31524 26574 31526
rect 24950 30812 24952 30832
rect 24952 30812 25004 30832
rect 25004 30812 25006 30832
rect 24950 30776 25006 30812
rect 22058 25594 22114 25596
rect 22138 25594 22194 25596
rect 22218 25594 22274 25596
rect 22298 25594 22354 25596
rect 22058 25542 22104 25594
rect 22104 25542 22114 25594
rect 22138 25542 22168 25594
rect 22168 25542 22180 25594
rect 22180 25542 22194 25594
rect 22218 25542 22232 25594
rect 22232 25542 22244 25594
rect 22244 25542 22274 25594
rect 22298 25542 22308 25594
rect 22308 25542 22354 25594
rect 22058 25540 22114 25542
rect 22138 25540 22194 25542
rect 22218 25540 22274 25542
rect 22298 25540 22354 25542
rect 22058 24506 22114 24508
rect 22138 24506 22194 24508
rect 22218 24506 22274 24508
rect 22298 24506 22354 24508
rect 22058 24454 22104 24506
rect 22104 24454 22114 24506
rect 22138 24454 22168 24506
rect 22168 24454 22180 24506
rect 22180 24454 22194 24506
rect 22218 24454 22232 24506
rect 22232 24454 22244 24506
rect 22244 24454 22274 24506
rect 22298 24454 22308 24506
rect 22308 24454 22354 24506
rect 22058 24452 22114 24454
rect 22138 24452 22194 24454
rect 22218 24452 22274 24454
rect 22298 24452 22354 24454
rect 22058 23418 22114 23420
rect 22138 23418 22194 23420
rect 22218 23418 22274 23420
rect 22298 23418 22354 23420
rect 22058 23366 22104 23418
rect 22104 23366 22114 23418
rect 22138 23366 22168 23418
rect 22168 23366 22180 23418
rect 22180 23366 22194 23418
rect 22218 23366 22232 23418
rect 22232 23366 22244 23418
rect 22244 23366 22274 23418
rect 22298 23366 22308 23418
rect 22308 23366 22354 23418
rect 22058 23364 22114 23366
rect 22138 23364 22194 23366
rect 22218 23364 22274 23366
rect 22298 23364 22354 23366
rect 22190 23160 22246 23216
rect 22058 22330 22114 22332
rect 22138 22330 22194 22332
rect 22218 22330 22274 22332
rect 22298 22330 22354 22332
rect 22058 22278 22104 22330
rect 22104 22278 22114 22330
rect 22138 22278 22168 22330
rect 22168 22278 22180 22330
rect 22180 22278 22194 22330
rect 22218 22278 22232 22330
rect 22232 22278 22244 22330
rect 22244 22278 22274 22330
rect 22298 22278 22308 22330
rect 22308 22278 22354 22330
rect 22058 22276 22114 22278
rect 22138 22276 22194 22278
rect 22218 22276 22274 22278
rect 22298 22276 22354 22278
rect 22058 21242 22114 21244
rect 22138 21242 22194 21244
rect 22218 21242 22274 21244
rect 22298 21242 22354 21244
rect 22058 21190 22104 21242
rect 22104 21190 22114 21242
rect 22138 21190 22168 21242
rect 22168 21190 22180 21242
rect 22180 21190 22194 21242
rect 22218 21190 22232 21242
rect 22232 21190 22244 21242
rect 22244 21190 22274 21242
rect 22298 21190 22308 21242
rect 22308 21190 22354 21242
rect 22058 21188 22114 21190
rect 22138 21188 22194 21190
rect 22218 21188 22274 21190
rect 22298 21188 22354 21190
rect 26278 30490 26334 30492
rect 26358 30490 26414 30492
rect 26438 30490 26494 30492
rect 26518 30490 26574 30492
rect 26278 30438 26324 30490
rect 26324 30438 26334 30490
rect 26358 30438 26388 30490
rect 26388 30438 26400 30490
rect 26400 30438 26414 30490
rect 26438 30438 26452 30490
rect 26452 30438 26464 30490
rect 26464 30438 26494 30490
rect 26518 30438 26528 30490
rect 26528 30438 26574 30490
rect 26278 30436 26334 30438
rect 26358 30436 26414 30438
rect 26438 30436 26494 30438
rect 26518 30436 26574 30438
rect 22058 20154 22114 20156
rect 22138 20154 22194 20156
rect 22218 20154 22274 20156
rect 22298 20154 22354 20156
rect 22058 20102 22104 20154
rect 22104 20102 22114 20154
rect 22138 20102 22168 20154
rect 22168 20102 22180 20154
rect 22180 20102 22194 20154
rect 22218 20102 22232 20154
rect 22232 20102 22244 20154
rect 22244 20102 22274 20154
rect 22298 20102 22308 20154
rect 22308 20102 22354 20154
rect 22058 20100 22114 20102
rect 22138 20100 22194 20102
rect 22218 20100 22274 20102
rect 22298 20100 22354 20102
rect 22058 19066 22114 19068
rect 22138 19066 22194 19068
rect 22218 19066 22274 19068
rect 22298 19066 22354 19068
rect 22058 19014 22104 19066
rect 22104 19014 22114 19066
rect 22138 19014 22168 19066
rect 22168 19014 22180 19066
rect 22180 19014 22194 19066
rect 22218 19014 22232 19066
rect 22232 19014 22244 19066
rect 22244 19014 22274 19066
rect 22298 19014 22308 19066
rect 22308 19014 22354 19066
rect 22058 19012 22114 19014
rect 22138 19012 22194 19014
rect 22218 19012 22274 19014
rect 22298 19012 22354 19014
rect 22058 17978 22114 17980
rect 22138 17978 22194 17980
rect 22218 17978 22274 17980
rect 22298 17978 22354 17980
rect 22058 17926 22104 17978
rect 22104 17926 22114 17978
rect 22138 17926 22168 17978
rect 22168 17926 22180 17978
rect 22180 17926 22194 17978
rect 22218 17926 22232 17978
rect 22232 17926 22244 17978
rect 22244 17926 22274 17978
rect 22298 17926 22308 17978
rect 22308 17926 22354 17978
rect 22058 17924 22114 17926
rect 22138 17924 22194 17926
rect 22218 17924 22274 17926
rect 22298 17924 22354 17926
rect 22058 16890 22114 16892
rect 22138 16890 22194 16892
rect 22218 16890 22274 16892
rect 22298 16890 22354 16892
rect 22058 16838 22104 16890
rect 22104 16838 22114 16890
rect 22138 16838 22168 16890
rect 22168 16838 22180 16890
rect 22180 16838 22194 16890
rect 22218 16838 22232 16890
rect 22232 16838 22244 16890
rect 22244 16838 22274 16890
rect 22298 16838 22308 16890
rect 22308 16838 22354 16890
rect 22058 16836 22114 16838
rect 22138 16836 22194 16838
rect 22218 16836 22274 16838
rect 22298 16836 22354 16838
rect 22058 15802 22114 15804
rect 22138 15802 22194 15804
rect 22218 15802 22274 15804
rect 22298 15802 22354 15804
rect 22058 15750 22104 15802
rect 22104 15750 22114 15802
rect 22138 15750 22168 15802
rect 22168 15750 22180 15802
rect 22180 15750 22194 15802
rect 22218 15750 22232 15802
rect 22232 15750 22244 15802
rect 22244 15750 22274 15802
rect 22298 15750 22308 15802
rect 22308 15750 22354 15802
rect 22058 15748 22114 15750
rect 22138 15748 22194 15750
rect 22218 15748 22274 15750
rect 22298 15748 22354 15750
rect 22190 14864 22246 14920
rect 22058 14714 22114 14716
rect 22138 14714 22194 14716
rect 22218 14714 22274 14716
rect 22298 14714 22354 14716
rect 22058 14662 22104 14714
rect 22104 14662 22114 14714
rect 22138 14662 22168 14714
rect 22168 14662 22180 14714
rect 22180 14662 22194 14714
rect 22218 14662 22232 14714
rect 22232 14662 22244 14714
rect 22244 14662 22274 14714
rect 22298 14662 22308 14714
rect 22308 14662 22354 14714
rect 22058 14660 22114 14662
rect 22138 14660 22194 14662
rect 22218 14660 22274 14662
rect 22298 14660 22354 14662
rect 22558 14320 22614 14376
rect 22058 13626 22114 13628
rect 22138 13626 22194 13628
rect 22218 13626 22274 13628
rect 22298 13626 22354 13628
rect 22058 13574 22104 13626
rect 22104 13574 22114 13626
rect 22138 13574 22168 13626
rect 22168 13574 22180 13626
rect 22180 13574 22194 13626
rect 22218 13574 22232 13626
rect 22232 13574 22244 13626
rect 22244 13574 22274 13626
rect 22298 13574 22308 13626
rect 22308 13574 22354 13626
rect 22058 13572 22114 13574
rect 22138 13572 22194 13574
rect 22218 13572 22274 13574
rect 22298 13572 22354 13574
rect 21178 11192 21234 11248
rect 21178 11076 21234 11112
rect 21178 11056 21180 11076
rect 21180 11056 21232 11076
rect 21232 11056 21234 11076
rect 22058 12538 22114 12540
rect 22138 12538 22194 12540
rect 22218 12538 22274 12540
rect 22298 12538 22354 12540
rect 22058 12486 22104 12538
rect 22104 12486 22114 12538
rect 22138 12486 22168 12538
rect 22168 12486 22180 12538
rect 22180 12486 22194 12538
rect 22218 12486 22232 12538
rect 22232 12486 22244 12538
rect 22244 12486 22274 12538
rect 22298 12486 22308 12538
rect 22308 12486 22354 12538
rect 22058 12484 22114 12486
rect 22138 12484 22194 12486
rect 22218 12484 22274 12486
rect 22298 12484 22354 12486
rect 22058 11450 22114 11452
rect 22138 11450 22194 11452
rect 22218 11450 22274 11452
rect 22298 11450 22354 11452
rect 22058 11398 22104 11450
rect 22104 11398 22114 11450
rect 22138 11398 22168 11450
rect 22168 11398 22180 11450
rect 22180 11398 22194 11450
rect 22218 11398 22232 11450
rect 22232 11398 22244 11450
rect 22244 11398 22274 11450
rect 22298 11398 22308 11450
rect 22308 11398 22354 11450
rect 22058 11396 22114 11398
rect 22138 11396 22194 11398
rect 22218 11396 22274 11398
rect 22298 11396 22354 11398
rect 22282 11192 22338 11248
rect 22650 12416 22706 12472
rect 22058 10362 22114 10364
rect 22138 10362 22194 10364
rect 22218 10362 22274 10364
rect 22298 10362 22354 10364
rect 22058 10310 22104 10362
rect 22104 10310 22114 10362
rect 22138 10310 22168 10362
rect 22168 10310 22180 10362
rect 22180 10310 22194 10362
rect 22218 10310 22232 10362
rect 22232 10310 22244 10362
rect 22244 10310 22274 10362
rect 22298 10310 22308 10362
rect 22308 10310 22354 10362
rect 22058 10308 22114 10310
rect 22138 10308 22194 10310
rect 22218 10308 22274 10310
rect 22298 10308 22354 10310
rect 22058 9274 22114 9276
rect 22138 9274 22194 9276
rect 22218 9274 22274 9276
rect 22298 9274 22354 9276
rect 22058 9222 22104 9274
rect 22104 9222 22114 9274
rect 22138 9222 22168 9274
rect 22168 9222 22180 9274
rect 22180 9222 22194 9274
rect 22218 9222 22232 9274
rect 22232 9222 22244 9274
rect 22244 9222 22274 9274
rect 22298 9222 22308 9274
rect 22308 9222 22354 9274
rect 22058 9220 22114 9222
rect 22138 9220 22194 9222
rect 22218 9220 22274 9222
rect 22298 9220 22354 9222
rect 22058 8186 22114 8188
rect 22138 8186 22194 8188
rect 22218 8186 22274 8188
rect 22298 8186 22354 8188
rect 22058 8134 22104 8186
rect 22104 8134 22114 8186
rect 22138 8134 22168 8186
rect 22168 8134 22180 8186
rect 22180 8134 22194 8186
rect 22218 8134 22232 8186
rect 22232 8134 22244 8186
rect 22244 8134 22274 8186
rect 22298 8134 22308 8186
rect 22308 8134 22354 8186
rect 22058 8132 22114 8134
rect 22138 8132 22194 8134
rect 22218 8132 22274 8134
rect 22298 8132 22354 8134
rect 26278 29402 26334 29404
rect 26358 29402 26414 29404
rect 26438 29402 26494 29404
rect 26518 29402 26574 29404
rect 26278 29350 26324 29402
rect 26324 29350 26334 29402
rect 26358 29350 26388 29402
rect 26388 29350 26400 29402
rect 26400 29350 26414 29402
rect 26438 29350 26452 29402
rect 26452 29350 26464 29402
rect 26464 29350 26494 29402
rect 26518 29350 26528 29402
rect 26528 29350 26574 29402
rect 26278 29348 26334 29350
rect 26358 29348 26414 29350
rect 26438 29348 26494 29350
rect 26518 29348 26574 29350
rect 26278 28314 26334 28316
rect 26358 28314 26414 28316
rect 26438 28314 26494 28316
rect 26518 28314 26574 28316
rect 26278 28262 26324 28314
rect 26324 28262 26334 28314
rect 26358 28262 26388 28314
rect 26388 28262 26400 28314
rect 26400 28262 26414 28314
rect 26438 28262 26452 28314
rect 26452 28262 26464 28314
rect 26464 28262 26494 28314
rect 26518 28262 26528 28314
rect 26528 28262 26574 28314
rect 26278 28260 26334 28262
rect 26358 28260 26414 28262
rect 26438 28260 26494 28262
rect 26518 28260 26574 28262
rect 26278 27226 26334 27228
rect 26358 27226 26414 27228
rect 26438 27226 26494 27228
rect 26518 27226 26574 27228
rect 26278 27174 26324 27226
rect 26324 27174 26334 27226
rect 26358 27174 26388 27226
rect 26388 27174 26400 27226
rect 26400 27174 26414 27226
rect 26438 27174 26452 27226
rect 26452 27174 26464 27226
rect 26464 27174 26494 27226
rect 26518 27174 26528 27226
rect 26528 27174 26574 27226
rect 26278 27172 26334 27174
rect 26358 27172 26414 27174
rect 26438 27172 26494 27174
rect 26518 27172 26574 27174
rect 23570 14340 23626 14376
rect 23570 14320 23572 14340
rect 23572 14320 23624 14340
rect 23624 14320 23626 14340
rect 22926 11056 22982 11112
rect 22058 7098 22114 7100
rect 22138 7098 22194 7100
rect 22218 7098 22274 7100
rect 22298 7098 22354 7100
rect 22058 7046 22104 7098
rect 22104 7046 22114 7098
rect 22138 7046 22168 7098
rect 22168 7046 22180 7098
rect 22180 7046 22194 7098
rect 22218 7046 22232 7098
rect 22232 7046 22244 7098
rect 22244 7046 22274 7098
rect 22298 7046 22308 7098
rect 22308 7046 22354 7098
rect 22058 7044 22114 7046
rect 22138 7044 22194 7046
rect 22218 7044 22274 7046
rect 22298 7044 22354 7046
rect 22058 6010 22114 6012
rect 22138 6010 22194 6012
rect 22218 6010 22274 6012
rect 22298 6010 22354 6012
rect 22058 5958 22104 6010
rect 22104 5958 22114 6010
rect 22138 5958 22168 6010
rect 22168 5958 22180 6010
rect 22180 5958 22194 6010
rect 22218 5958 22232 6010
rect 22232 5958 22244 6010
rect 22244 5958 22274 6010
rect 22298 5958 22308 6010
rect 22308 5958 22354 6010
rect 22058 5956 22114 5958
rect 22138 5956 22194 5958
rect 22218 5956 22274 5958
rect 22298 5956 22354 5958
rect 24674 14864 24730 14920
rect 26278 26138 26334 26140
rect 26358 26138 26414 26140
rect 26438 26138 26494 26140
rect 26518 26138 26574 26140
rect 26278 26086 26324 26138
rect 26324 26086 26334 26138
rect 26358 26086 26388 26138
rect 26388 26086 26400 26138
rect 26400 26086 26414 26138
rect 26438 26086 26452 26138
rect 26452 26086 26464 26138
rect 26464 26086 26494 26138
rect 26518 26086 26528 26138
rect 26528 26086 26574 26138
rect 26278 26084 26334 26086
rect 26358 26084 26414 26086
rect 26438 26084 26494 26086
rect 26518 26084 26574 26086
rect 26278 25050 26334 25052
rect 26358 25050 26414 25052
rect 26438 25050 26494 25052
rect 26518 25050 26574 25052
rect 26278 24998 26324 25050
rect 26324 24998 26334 25050
rect 26358 24998 26388 25050
rect 26388 24998 26400 25050
rect 26400 24998 26414 25050
rect 26438 24998 26452 25050
rect 26452 24998 26464 25050
rect 26464 24998 26494 25050
rect 26518 24998 26528 25050
rect 26528 24998 26574 25050
rect 26278 24996 26334 24998
rect 26358 24996 26414 24998
rect 26438 24996 26494 24998
rect 26518 24996 26574 24998
rect 26278 23962 26334 23964
rect 26358 23962 26414 23964
rect 26438 23962 26494 23964
rect 26518 23962 26574 23964
rect 26278 23910 26324 23962
rect 26324 23910 26334 23962
rect 26358 23910 26388 23962
rect 26388 23910 26400 23962
rect 26400 23910 26414 23962
rect 26438 23910 26452 23962
rect 26452 23910 26464 23962
rect 26464 23910 26494 23962
rect 26518 23910 26528 23962
rect 26528 23910 26574 23962
rect 26278 23908 26334 23910
rect 26358 23908 26414 23910
rect 26438 23908 26494 23910
rect 26518 23908 26574 23910
rect 26278 22874 26334 22876
rect 26358 22874 26414 22876
rect 26438 22874 26494 22876
rect 26518 22874 26574 22876
rect 26278 22822 26324 22874
rect 26324 22822 26334 22874
rect 26358 22822 26388 22874
rect 26388 22822 26400 22874
rect 26400 22822 26414 22874
rect 26438 22822 26452 22874
rect 26452 22822 26464 22874
rect 26464 22822 26494 22874
rect 26518 22822 26528 22874
rect 26528 22822 26574 22874
rect 26278 22820 26334 22822
rect 26358 22820 26414 22822
rect 26438 22820 26494 22822
rect 26518 22820 26574 22822
rect 26278 21786 26334 21788
rect 26358 21786 26414 21788
rect 26438 21786 26494 21788
rect 26518 21786 26574 21788
rect 26278 21734 26324 21786
rect 26324 21734 26334 21786
rect 26358 21734 26388 21786
rect 26388 21734 26400 21786
rect 26400 21734 26414 21786
rect 26438 21734 26452 21786
rect 26452 21734 26464 21786
rect 26464 21734 26494 21786
rect 26518 21734 26528 21786
rect 26528 21734 26574 21786
rect 26278 21732 26334 21734
rect 26358 21732 26414 21734
rect 26438 21732 26494 21734
rect 26518 21732 26574 21734
rect 26278 20698 26334 20700
rect 26358 20698 26414 20700
rect 26438 20698 26494 20700
rect 26518 20698 26574 20700
rect 26278 20646 26324 20698
rect 26324 20646 26334 20698
rect 26358 20646 26388 20698
rect 26388 20646 26400 20698
rect 26400 20646 26414 20698
rect 26438 20646 26452 20698
rect 26452 20646 26464 20698
rect 26464 20646 26494 20698
rect 26518 20646 26528 20698
rect 26528 20646 26574 20698
rect 26278 20644 26334 20646
rect 26358 20644 26414 20646
rect 26438 20644 26494 20646
rect 26518 20644 26574 20646
rect 26278 19610 26334 19612
rect 26358 19610 26414 19612
rect 26438 19610 26494 19612
rect 26518 19610 26574 19612
rect 26278 19558 26324 19610
rect 26324 19558 26334 19610
rect 26358 19558 26388 19610
rect 26388 19558 26400 19610
rect 26400 19558 26414 19610
rect 26438 19558 26452 19610
rect 26452 19558 26464 19610
rect 26464 19558 26494 19610
rect 26518 19558 26528 19610
rect 26528 19558 26574 19610
rect 26278 19556 26334 19558
rect 26358 19556 26414 19558
rect 26438 19556 26494 19558
rect 26518 19556 26574 19558
rect 27250 22092 27306 22128
rect 27250 22072 27252 22092
rect 27252 22072 27304 22092
rect 27304 22072 27306 22092
rect 26278 18522 26334 18524
rect 26358 18522 26414 18524
rect 26438 18522 26494 18524
rect 26518 18522 26574 18524
rect 26278 18470 26324 18522
rect 26324 18470 26334 18522
rect 26358 18470 26388 18522
rect 26388 18470 26400 18522
rect 26400 18470 26414 18522
rect 26438 18470 26452 18522
rect 26452 18470 26464 18522
rect 26464 18470 26494 18522
rect 26518 18470 26528 18522
rect 26528 18470 26574 18522
rect 26278 18468 26334 18470
rect 26358 18468 26414 18470
rect 26438 18468 26494 18470
rect 26518 18468 26574 18470
rect 30499 32122 30555 32124
rect 30579 32122 30635 32124
rect 30659 32122 30715 32124
rect 30739 32122 30795 32124
rect 30499 32070 30545 32122
rect 30545 32070 30555 32122
rect 30579 32070 30609 32122
rect 30609 32070 30621 32122
rect 30621 32070 30635 32122
rect 30659 32070 30673 32122
rect 30673 32070 30685 32122
rect 30685 32070 30715 32122
rect 30739 32070 30749 32122
rect 30749 32070 30795 32122
rect 30499 32068 30555 32070
rect 30579 32068 30635 32070
rect 30659 32068 30715 32070
rect 30739 32068 30795 32070
rect 30499 31034 30555 31036
rect 30579 31034 30635 31036
rect 30659 31034 30715 31036
rect 30739 31034 30795 31036
rect 30499 30982 30545 31034
rect 30545 30982 30555 31034
rect 30579 30982 30609 31034
rect 30609 30982 30621 31034
rect 30621 30982 30635 31034
rect 30659 30982 30673 31034
rect 30673 30982 30685 31034
rect 30685 30982 30715 31034
rect 30739 30982 30749 31034
rect 30749 30982 30795 31034
rect 30499 30980 30555 30982
rect 30579 30980 30635 30982
rect 30659 30980 30715 30982
rect 30739 30980 30795 30982
rect 30499 29946 30555 29948
rect 30579 29946 30635 29948
rect 30659 29946 30715 29948
rect 30739 29946 30795 29948
rect 30499 29894 30545 29946
rect 30545 29894 30555 29946
rect 30579 29894 30609 29946
rect 30609 29894 30621 29946
rect 30621 29894 30635 29946
rect 30659 29894 30673 29946
rect 30673 29894 30685 29946
rect 30685 29894 30715 29946
rect 30739 29894 30749 29946
rect 30749 29894 30795 29946
rect 30499 29892 30555 29894
rect 30579 29892 30635 29894
rect 30659 29892 30715 29894
rect 30739 29892 30795 29894
rect 30499 28858 30555 28860
rect 30579 28858 30635 28860
rect 30659 28858 30715 28860
rect 30739 28858 30795 28860
rect 30499 28806 30545 28858
rect 30545 28806 30555 28858
rect 30579 28806 30609 28858
rect 30609 28806 30621 28858
rect 30621 28806 30635 28858
rect 30659 28806 30673 28858
rect 30673 28806 30685 28858
rect 30685 28806 30715 28858
rect 30739 28806 30749 28858
rect 30749 28806 30795 28858
rect 30499 28804 30555 28806
rect 30579 28804 30635 28806
rect 30659 28804 30715 28806
rect 30739 28804 30795 28806
rect 30499 27770 30555 27772
rect 30579 27770 30635 27772
rect 30659 27770 30715 27772
rect 30739 27770 30795 27772
rect 30499 27718 30545 27770
rect 30545 27718 30555 27770
rect 30579 27718 30609 27770
rect 30609 27718 30621 27770
rect 30621 27718 30635 27770
rect 30659 27718 30673 27770
rect 30673 27718 30685 27770
rect 30685 27718 30715 27770
rect 30739 27718 30749 27770
rect 30749 27718 30795 27770
rect 30499 27716 30555 27718
rect 30579 27716 30635 27718
rect 30659 27716 30715 27718
rect 30739 27716 30795 27718
rect 30499 26682 30555 26684
rect 30579 26682 30635 26684
rect 30659 26682 30715 26684
rect 30739 26682 30795 26684
rect 30499 26630 30545 26682
rect 30545 26630 30555 26682
rect 30579 26630 30609 26682
rect 30609 26630 30621 26682
rect 30621 26630 30635 26682
rect 30659 26630 30673 26682
rect 30673 26630 30685 26682
rect 30685 26630 30715 26682
rect 30739 26630 30749 26682
rect 30749 26630 30795 26682
rect 30499 26628 30555 26630
rect 30579 26628 30635 26630
rect 30659 26628 30715 26630
rect 30739 26628 30795 26630
rect 30499 25594 30555 25596
rect 30579 25594 30635 25596
rect 30659 25594 30715 25596
rect 30739 25594 30795 25596
rect 30499 25542 30545 25594
rect 30545 25542 30555 25594
rect 30579 25542 30609 25594
rect 30609 25542 30621 25594
rect 30621 25542 30635 25594
rect 30659 25542 30673 25594
rect 30673 25542 30685 25594
rect 30685 25542 30715 25594
rect 30739 25542 30749 25594
rect 30749 25542 30795 25594
rect 30499 25540 30555 25542
rect 30579 25540 30635 25542
rect 30659 25540 30715 25542
rect 30739 25540 30795 25542
rect 30499 24506 30555 24508
rect 30579 24506 30635 24508
rect 30659 24506 30715 24508
rect 30739 24506 30795 24508
rect 30499 24454 30545 24506
rect 30545 24454 30555 24506
rect 30579 24454 30609 24506
rect 30609 24454 30621 24506
rect 30621 24454 30635 24506
rect 30659 24454 30673 24506
rect 30673 24454 30685 24506
rect 30685 24454 30715 24506
rect 30739 24454 30749 24506
rect 30749 24454 30795 24506
rect 30499 24452 30555 24454
rect 30579 24452 30635 24454
rect 30659 24452 30715 24454
rect 30739 24452 30795 24454
rect 30499 23418 30555 23420
rect 30579 23418 30635 23420
rect 30659 23418 30715 23420
rect 30739 23418 30795 23420
rect 30499 23366 30545 23418
rect 30545 23366 30555 23418
rect 30579 23366 30609 23418
rect 30609 23366 30621 23418
rect 30621 23366 30635 23418
rect 30659 23366 30673 23418
rect 30673 23366 30685 23418
rect 30685 23366 30715 23418
rect 30739 23366 30749 23418
rect 30749 23366 30795 23418
rect 30499 23364 30555 23366
rect 30579 23364 30635 23366
rect 30659 23364 30715 23366
rect 30739 23364 30795 23366
rect 30499 22330 30555 22332
rect 30579 22330 30635 22332
rect 30659 22330 30715 22332
rect 30739 22330 30795 22332
rect 30499 22278 30545 22330
rect 30545 22278 30555 22330
rect 30579 22278 30609 22330
rect 30609 22278 30621 22330
rect 30621 22278 30635 22330
rect 30659 22278 30673 22330
rect 30673 22278 30685 22330
rect 30685 22278 30715 22330
rect 30739 22278 30749 22330
rect 30749 22278 30795 22330
rect 30499 22276 30555 22278
rect 30579 22276 30635 22278
rect 30659 22276 30715 22278
rect 30739 22276 30795 22278
rect 30499 21242 30555 21244
rect 30579 21242 30635 21244
rect 30659 21242 30715 21244
rect 30739 21242 30795 21244
rect 30499 21190 30545 21242
rect 30545 21190 30555 21242
rect 30579 21190 30609 21242
rect 30609 21190 30621 21242
rect 30621 21190 30635 21242
rect 30659 21190 30673 21242
rect 30673 21190 30685 21242
rect 30685 21190 30715 21242
rect 30739 21190 30749 21242
rect 30749 21190 30795 21242
rect 30499 21188 30555 21190
rect 30579 21188 30635 21190
rect 30659 21188 30715 21190
rect 30739 21188 30795 21190
rect 34719 31578 34775 31580
rect 34799 31578 34855 31580
rect 34879 31578 34935 31580
rect 34959 31578 35015 31580
rect 34719 31526 34765 31578
rect 34765 31526 34775 31578
rect 34799 31526 34829 31578
rect 34829 31526 34841 31578
rect 34841 31526 34855 31578
rect 34879 31526 34893 31578
rect 34893 31526 34905 31578
rect 34905 31526 34935 31578
rect 34959 31526 34969 31578
rect 34969 31526 35015 31578
rect 34719 31524 34775 31526
rect 34799 31524 34855 31526
rect 34879 31524 34935 31526
rect 34959 31524 35015 31526
rect 34719 30490 34775 30492
rect 34799 30490 34855 30492
rect 34879 30490 34935 30492
rect 34959 30490 35015 30492
rect 34719 30438 34765 30490
rect 34765 30438 34775 30490
rect 34799 30438 34829 30490
rect 34829 30438 34841 30490
rect 34841 30438 34855 30490
rect 34879 30438 34893 30490
rect 34893 30438 34905 30490
rect 34905 30438 34935 30490
rect 34959 30438 34969 30490
rect 34969 30438 35015 30490
rect 34719 30436 34775 30438
rect 34799 30436 34855 30438
rect 34879 30436 34935 30438
rect 34959 30436 35015 30438
rect 34719 29402 34775 29404
rect 34799 29402 34855 29404
rect 34879 29402 34935 29404
rect 34959 29402 35015 29404
rect 34719 29350 34765 29402
rect 34765 29350 34775 29402
rect 34799 29350 34829 29402
rect 34829 29350 34841 29402
rect 34841 29350 34855 29402
rect 34879 29350 34893 29402
rect 34893 29350 34905 29402
rect 34905 29350 34935 29402
rect 34959 29350 34969 29402
rect 34969 29350 35015 29402
rect 34719 29348 34775 29350
rect 34799 29348 34855 29350
rect 34879 29348 34935 29350
rect 34959 29348 35015 29350
rect 34719 28314 34775 28316
rect 34799 28314 34855 28316
rect 34879 28314 34935 28316
rect 34959 28314 35015 28316
rect 34719 28262 34765 28314
rect 34765 28262 34775 28314
rect 34799 28262 34829 28314
rect 34829 28262 34841 28314
rect 34841 28262 34855 28314
rect 34879 28262 34893 28314
rect 34893 28262 34905 28314
rect 34905 28262 34935 28314
rect 34959 28262 34969 28314
rect 34969 28262 35015 28314
rect 34719 28260 34775 28262
rect 34799 28260 34855 28262
rect 34879 28260 34935 28262
rect 34959 28260 35015 28262
rect 34719 27226 34775 27228
rect 34799 27226 34855 27228
rect 34879 27226 34935 27228
rect 34959 27226 35015 27228
rect 34719 27174 34765 27226
rect 34765 27174 34775 27226
rect 34799 27174 34829 27226
rect 34829 27174 34841 27226
rect 34841 27174 34855 27226
rect 34879 27174 34893 27226
rect 34893 27174 34905 27226
rect 34905 27174 34935 27226
rect 34959 27174 34969 27226
rect 34969 27174 35015 27226
rect 34719 27172 34775 27174
rect 34799 27172 34855 27174
rect 34879 27172 34935 27174
rect 34959 27172 35015 27174
rect 34719 26138 34775 26140
rect 34799 26138 34855 26140
rect 34879 26138 34935 26140
rect 34959 26138 35015 26140
rect 34719 26086 34765 26138
rect 34765 26086 34775 26138
rect 34799 26086 34829 26138
rect 34829 26086 34841 26138
rect 34841 26086 34855 26138
rect 34879 26086 34893 26138
rect 34893 26086 34905 26138
rect 34905 26086 34935 26138
rect 34959 26086 34969 26138
rect 34969 26086 35015 26138
rect 34719 26084 34775 26086
rect 34799 26084 34855 26086
rect 34879 26084 34935 26086
rect 34959 26084 35015 26086
rect 34719 25050 34775 25052
rect 34799 25050 34855 25052
rect 34879 25050 34935 25052
rect 34959 25050 35015 25052
rect 34719 24998 34765 25050
rect 34765 24998 34775 25050
rect 34799 24998 34829 25050
rect 34829 24998 34841 25050
rect 34841 24998 34855 25050
rect 34879 24998 34893 25050
rect 34893 24998 34905 25050
rect 34905 24998 34935 25050
rect 34959 24998 34969 25050
rect 34969 24998 35015 25050
rect 34719 24996 34775 24998
rect 34799 24996 34855 24998
rect 34879 24996 34935 24998
rect 34959 24996 35015 24998
rect 34719 23962 34775 23964
rect 34799 23962 34855 23964
rect 34879 23962 34935 23964
rect 34959 23962 35015 23964
rect 34719 23910 34765 23962
rect 34765 23910 34775 23962
rect 34799 23910 34829 23962
rect 34829 23910 34841 23962
rect 34841 23910 34855 23962
rect 34879 23910 34893 23962
rect 34893 23910 34905 23962
rect 34905 23910 34935 23962
rect 34959 23910 34969 23962
rect 34969 23910 35015 23962
rect 34719 23908 34775 23910
rect 34799 23908 34855 23910
rect 34879 23908 34935 23910
rect 34959 23908 35015 23910
rect 30499 20154 30555 20156
rect 30579 20154 30635 20156
rect 30659 20154 30715 20156
rect 30739 20154 30795 20156
rect 30499 20102 30545 20154
rect 30545 20102 30555 20154
rect 30579 20102 30609 20154
rect 30609 20102 30621 20154
rect 30621 20102 30635 20154
rect 30659 20102 30673 20154
rect 30673 20102 30685 20154
rect 30685 20102 30715 20154
rect 30739 20102 30749 20154
rect 30749 20102 30795 20154
rect 30499 20100 30555 20102
rect 30579 20100 30635 20102
rect 30659 20100 30715 20102
rect 30739 20100 30795 20102
rect 30499 19066 30555 19068
rect 30579 19066 30635 19068
rect 30659 19066 30715 19068
rect 30739 19066 30795 19068
rect 30499 19014 30545 19066
rect 30545 19014 30555 19066
rect 30579 19014 30609 19066
rect 30609 19014 30621 19066
rect 30621 19014 30635 19066
rect 30659 19014 30673 19066
rect 30673 19014 30685 19066
rect 30685 19014 30715 19066
rect 30739 19014 30749 19066
rect 30749 19014 30795 19066
rect 30499 19012 30555 19014
rect 30579 19012 30635 19014
rect 30659 19012 30715 19014
rect 30739 19012 30795 19014
rect 26278 17434 26334 17436
rect 26358 17434 26414 17436
rect 26438 17434 26494 17436
rect 26518 17434 26574 17436
rect 26278 17382 26324 17434
rect 26324 17382 26334 17434
rect 26358 17382 26388 17434
rect 26388 17382 26400 17434
rect 26400 17382 26414 17434
rect 26438 17382 26452 17434
rect 26452 17382 26464 17434
rect 26464 17382 26494 17434
rect 26518 17382 26528 17434
rect 26528 17382 26574 17434
rect 26278 17380 26334 17382
rect 26358 17380 26414 17382
rect 26438 17380 26494 17382
rect 26518 17380 26574 17382
rect 26278 16346 26334 16348
rect 26358 16346 26414 16348
rect 26438 16346 26494 16348
rect 26518 16346 26574 16348
rect 26278 16294 26324 16346
rect 26324 16294 26334 16346
rect 26358 16294 26388 16346
rect 26388 16294 26400 16346
rect 26400 16294 26414 16346
rect 26438 16294 26452 16346
rect 26452 16294 26464 16346
rect 26464 16294 26494 16346
rect 26518 16294 26528 16346
rect 26528 16294 26574 16346
rect 26278 16292 26334 16294
rect 26358 16292 26414 16294
rect 26438 16292 26494 16294
rect 26518 16292 26574 16294
rect 26278 15258 26334 15260
rect 26358 15258 26414 15260
rect 26438 15258 26494 15260
rect 26518 15258 26574 15260
rect 26278 15206 26324 15258
rect 26324 15206 26334 15258
rect 26358 15206 26388 15258
rect 26388 15206 26400 15258
rect 26400 15206 26414 15258
rect 26438 15206 26452 15258
rect 26452 15206 26464 15258
rect 26464 15206 26494 15258
rect 26518 15206 26528 15258
rect 26528 15206 26574 15258
rect 26278 15204 26334 15206
rect 26358 15204 26414 15206
rect 26438 15204 26494 15206
rect 26518 15204 26574 15206
rect 26278 14170 26334 14172
rect 26358 14170 26414 14172
rect 26438 14170 26494 14172
rect 26518 14170 26574 14172
rect 26278 14118 26324 14170
rect 26324 14118 26334 14170
rect 26358 14118 26388 14170
rect 26388 14118 26400 14170
rect 26400 14118 26414 14170
rect 26438 14118 26452 14170
rect 26452 14118 26464 14170
rect 26464 14118 26494 14170
rect 26518 14118 26528 14170
rect 26528 14118 26574 14170
rect 26278 14116 26334 14118
rect 26358 14116 26414 14118
rect 26438 14116 26494 14118
rect 26518 14116 26574 14118
rect 26278 13082 26334 13084
rect 26358 13082 26414 13084
rect 26438 13082 26494 13084
rect 26518 13082 26574 13084
rect 26278 13030 26324 13082
rect 26324 13030 26334 13082
rect 26358 13030 26388 13082
rect 26388 13030 26400 13082
rect 26400 13030 26414 13082
rect 26438 13030 26452 13082
rect 26452 13030 26464 13082
rect 26464 13030 26494 13082
rect 26518 13030 26528 13082
rect 26528 13030 26574 13082
rect 26278 13028 26334 13030
rect 26358 13028 26414 13030
rect 26438 13028 26494 13030
rect 26518 13028 26574 13030
rect 26278 11994 26334 11996
rect 26358 11994 26414 11996
rect 26438 11994 26494 11996
rect 26518 11994 26574 11996
rect 26278 11942 26324 11994
rect 26324 11942 26334 11994
rect 26358 11942 26388 11994
rect 26388 11942 26400 11994
rect 26400 11942 26414 11994
rect 26438 11942 26452 11994
rect 26452 11942 26464 11994
rect 26464 11942 26494 11994
rect 26518 11942 26528 11994
rect 26528 11942 26574 11994
rect 26278 11940 26334 11942
rect 26358 11940 26414 11942
rect 26438 11940 26494 11942
rect 26518 11940 26574 11942
rect 26278 10906 26334 10908
rect 26358 10906 26414 10908
rect 26438 10906 26494 10908
rect 26518 10906 26574 10908
rect 26278 10854 26324 10906
rect 26324 10854 26334 10906
rect 26358 10854 26388 10906
rect 26388 10854 26400 10906
rect 26400 10854 26414 10906
rect 26438 10854 26452 10906
rect 26452 10854 26464 10906
rect 26464 10854 26494 10906
rect 26518 10854 26528 10906
rect 26528 10854 26574 10906
rect 26278 10852 26334 10854
rect 26358 10852 26414 10854
rect 26438 10852 26494 10854
rect 26518 10852 26574 10854
rect 26278 9818 26334 9820
rect 26358 9818 26414 9820
rect 26438 9818 26494 9820
rect 26518 9818 26574 9820
rect 26278 9766 26324 9818
rect 26324 9766 26334 9818
rect 26358 9766 26388 9818
rect 26388 9766 26400 9818
rect 26400 9766 26414 9818
rect 26438 9766 26452 9818
rect 26452 9766 26464 9818
rect 26464 9766 26494 9818
rect 26518 9766 26528 9818
rect 26528 9766 26574 9818
rect 26278 9764 26334 9766
rect 26358 9764 26414 9766
rect 26438 9764 26494 9766
rect 26518 9764 26574 9766
rect 27802 13932 27858 13968
rect 27802 13912 27804 13932
rect 27804 13912 27856 13932
rect 27856 13912 27858 13932
rect 26278 8730 26334 8732
rect 26358 8730 26414 8732
rect 26438 8730 26494 8732
rect 26518 8730 26574 8732
rect 26278 8678 26324 8730
rect 26324 8678 26334 8730
rect 26358 8678 26388 8730
rect 26388 8678 26400 8730
rect 26400 8678 26414 8730
rect 26438 8678 26452 8730
rect 26452 8678 26464 8730
rect 26464 8678 26494 8730
rect 26518 8678 26528 8730
rect 26528 8678 26574 8730
rect 26278 8676 26334 8678
rect 26358 8676 26414 8678
rect 26438 8676 26494 8678
rect 26518 8676 26574 8678
rect 26278 7642 26334 7644
rect 26358 7642 26414 7644
rect 26438 7642 26494 7644
rect 26518 7642 26574 7644
rect 26278 7590 26324 7642
rect 26324 7590 26334 7642
rect 26358 7590 26388 7642
rect 26388 7590 26400 7642
rect 26400 7590 26414 7642
rect 26438 7590 26452 7642
rect 26452 7590 26464 7642
rect 26464 7590 26494 7642
rect 26518 7590 26528 7642
rect 26528 7590 26574 7642
rect 26278 7588 26334 7590
rect 26358 7588 26414 7590
rect 26438 7588 26494 7590
rect 26518 7588 26574 7590
rect 28078 12280 28134 12336
rect 30499 17978 30555 17980
rect 30579 17978 30635 17980
rect 30659 17978 30715 17980
rect 30739 17978 30795 17980
rect 30499 17926 30545 17978
rect 30545 17926 30555 17978
rect 30579 17926 30609 17978
rect 30609 17926 30621 17978
rect 30621 17926 30635 17978
rect 30659 17926 30673 17978
rect 30673 17926 30685 17978
rect 30685 17926 30715 17978
rect 30739 17926 30749 17978
rect 30749 17926 30795 17978
rect 30499 17924 30555 17926
rect 30579 17924 30635 17926
rect 30659 17924 30715 17926
rect 30739 17924 30795 17926
rect 30499 16890 30555 16892
rect 30579 16890 30635 16892
rect 30659 16890 30715 16892
rect 30739 16890 30795 16892
rect 30499 16838 30545 16890
rect 30545 16838 30555 16890
rect 30579 16838 30609 16890
rect 30609 16838 30621 16890
rect 30621 16838 30635 16890
rect 30659 16838 30673 16890
rect 30673 16838 30685 16890
rect 30685 16838 30715 16890
rect 30739 16838 30749 16890
rect 30749 16838 30795 16890
rect 30499 16836 30555 16838
rect 30579 16836 30635 16838
rect 30659 16836 30715 16838
rect 30739 16836 30795 16838
rect 34719 22874 34775 22876
rect 34799 22874 34855 22876
rect 34879 22874 34935 22876
rect 34959 22874 35015 22876
rect 34719 22822 34765 22874
rect 34765 22822 34775 22874
rect 34799 22822 34829 22874
rect 34829 22822 34841 22874
rect 34841 22822 34855 22874
rect 34879 22822 34893 22874
rect 34893 22822 34905 22874
rect 34905 22822 34935 22874
rect 34959 22822 34969 22874
rect 34969 22822 35015 22874
rect 34719 22820 34775 22822
rect 34799 22820 34855 22822
rect 34879 22820 34935 22822
rect 34959 22820 35015 22822
rect 34719 21786 34775 21788
rect 34799 21786 34855 21788
rect 34879 21786 34935 21788
rect 34959 21786 35015 21788
rect 34719 21734 34765 21786
rect 34765 21734 34775 21786
rect 34799 21734 34829 21786
rect 34829 21734 34841 21786
rect 34841 21734 34855 21786
rect 34879 21734 34893 21786
rect 34893 21734 34905 21786
rect 34905 21734 34935 21786
rect 34959 21734 34969 21786
rect 34969 21734 35015 21786
rect 34719 21732 34775 21734
rect 34799 21732 34855 21734
rect 34879 21732 34935 21734
rect 34959 21732 35015 21734
rect 34719 20698 34775 20700
rect 34799 20698 34855 20700
rect 34879 20698 34935 20700
rect 34959 20698 35015 20700
rect 34719 20646 34765 20698
rect 34765 20646 34775 20698
rect 34799 20646 34829 20698
rect 34829 20646 34841 20698
rect 34841 20646 34855 20698
rect 34879 20646 34893 20698
rect 34893 20646 34905 20698
rect 34905 20646 34935 20698
rect 34959 20646 34969 20698
rect 34969 20646 35015 20698
rect 34719 20644 34775 20646
rect 34799 20644 34855 20646
rect 34879 20644 34935 20646
rect 34959 20644 35015 20646
rect 34719 19610 34775 19612
rect 34799 19610 34855 19612
rect 34879 19610 34935 19612
rect 34959 19610 35015 19612
rect 34719 19558 34765 19610
rect 34765 19558 34775 19610
rect 34799 19558 34829 19610
rect 34829 19558 34841 19610
rect 34841 19558 34855 19610
rect 34879 19558 34893 19610
rect 34893 19558 34905 19610
rect 34905 19558 34935 19610
rect 34959 19558 34969 19610
rect 34969 19558 35015 19610
rect 34719 19556 34775 19558
rect 34799 19556 34855 19558
rect 34879 19556 34935 19558
rect 34959 19556 35015 19558
rect 34719 18522 34775 18524
rect 34799 18522 34855 18524
rect 34879 18522 34935 18524
rect 34959 18522 35015 18524
rect 34719 18470 34765 18522
rect 34765 18470 34775 18522
rect 34799 18470 34829 18522
rect 34829 18470 34841 18522
rect 34841 18470 34855 18522
rect 34879 18470 34893 18522
rect 34893 18470 34905 18522
rect 34905 18470 34935 18522
rect 34959 18470 34969 18522
rect 34969 18470 35015 18522
rect 34719 18468 34775 18470
rect 34799 18468 34855 18470
rect 34879 18468 34935 18470
rect 34959 18468 35015 18470
rect 34334 17856 34390 17912
rect 34719 17434 34775 17436
rect 34799 17434 34855 17436
rect 34879 17434 34935 17436
rect 34959 17434 35015 17436
rect 34719 17382 34765 17434
rect 34765 17382 34775 17434
rect 34799 17382 34829 17434
rect 34829 17382 34841 17434
rect 34841 17382 34855 17434
rect 34879 17382 34893 17434
rect 34893 17382 34905 17434
rect 34905 17382 34935 17434
rect 34959 17382 34969 17434
rect 34969 17382 35015 17434
rect 34719 17380 34775 17382
rect 34799 17380 34855 17382
rect 34879 17380 34935 17382
rect 34959 17380 35015 17382
rect 28722 14320 28778 14376
rect 30499 15802 30555 15804
rect 30579 15802 30635 15804
rect 30659 15802 30715 15804
rect 30739 15802 30795 15804
rect 30499 15750 30545 15802
rect 30545 15750 30555 15802
rect 30579 15750 30609 15802
rect 30609 15750 30621 15802
rect 30621 15750 30635 15802
rect 30659 15750 30673 15802
rect 30673 15750 30685 15802
rect 30685 15750 30715 15802
rect 30739 15750 30749 15802
rect 30749 15750 30795 15802
rect 30499 15748 30555 15750
rect 30579 15748 30635 15750
rect 30659 15748 30715 15750
rect 30739 15748 30795 15750
rect 30499 14714 30555 14716
rect 30579 14714 30635 14716
rect 30659 14714 30715 14716
rect 30739 14714 30795 14716
rect 30499 14662 30545 14714
rect 30545 14662 30555 14714
rect 30579 14662 30609 14714
rect 30609 14662 30621 14714
rect 30621 14662 30635 14714
rect 30659 14662 30673 14714
rect 30673 14662 30685 14714
rect 30685 14662 30715 14714
rect 30739 14662 30749 14714
rect 30749 14662 30795 14714
rect 30499 14660 30555 14662
rect 30579 14660 30635 14662
rect 30659 14660 30715 14662
rect 30739 14660 30795 14662
rect 26278 6554 26334 6556
rect 26358 6554 26414 6556
rect 26438 6554 26494 6556
rect 26518 6554 26574 6556
rect 26278 6502 26324 6554
rect 26324 6502 26334 6554
rect 26358 6502 26388 6554
rect 26388 6502 26400 6554
rect 26400 6502 26414 6554
rect 26438 6502 26452 6554
rect 26452 6502 26464 6554
rect 26464 6502 26494 6554
rect 26518 6502 26528 6554
rect 26528 6502 26574 6554
rect 26278 6500 26334 6502
rect 26358 6500 26414 6502
rect 26438 6500 26494 6502
rect 26518 6500 26574 6502
rect 26278 5466 26334 5468
rect 26358 5466 26414 5468
rect 26438 5466 26494 5468
rect 26518 5466 26574 5468
rect 26278 5414 26324 5466
rect 26324 5414 26334 5466
rect 26358 5414 26388 5466
rect 26388 5414 26400 5466
rect 26400 5414 26414 5466
rect 26438 5414 26452 5466
rect 26452 5414 26464 5466
rect 26464 5414 26494 5466
rect 26518 5414 26528 5466
rect 26528 5414 26574 5466
rect 26278 5412 26334 5414
rect 26358 5412 26414 5414
rect 26438 5412 26494 5414
rect 26518 5412 26574 5414
rect 22058 4922 22114 4924
rect 22138 4922 22194 4924
rect 22218 4922 22274 4924
rect 22298 4922 22354 4924
rect 22058 4870 22104 4922
rect 22104 4870 22114 4922
rect 22138 4870 22168 4922
rect 22168 4870 22180 4922
rect 22180 4870 22194 4922
rect 22218 4870 22232 4922
rect 22232 4870 22244 4922
rect 22244 4870 22274 4922
rect 22298 4870 22308 4922
rect 22308 4870 22354 4922
rect 22058 4868 22114 4870
rect 22138 4868 22194 4870
rect 22218 4868 22274 4870
rect 22298 4868 22354 4870
rect 17837 4378 17893 4380
rect 17917 4378 17973 4380
rect 17997 4378 18053 4380
rect 18077 4378 18133 4380
rect 17837 4326 17883 4378
rect 17883 4326 17893 4378
rect 17917 4326 17947 4378
rect 17947 4326 17959 4378
rect 17959 4326 17973 4378
rect 17997 4326 18011 4378
rect 18011 4326 18023 4378
rect 18023 4326 18053 4378
rect 18077 4326 18087 4378
rect 18087 4326 18133 4378
rect 17837 4324 17893 4326
rect 17917 4324 17973 4326
rect 17997 4324 18053 4326
rect 18077 4324 18133 4326
rect 17837 3290 17893 3292
rect 17917 3290 17973 3292
rect 17997 3290 18053 3292
rect 18077 3290 18133 3292
rect 17837 3238 17883 3290
rect 17883 3238 17893 3290
rect 17917 3238 17947 3290
rect 17947 3238 17959 3290
rect 17959 3238 17973 3290
rect 17997 3238 18011 3290
rect 18011 3238 18023 3290
rect 18023 3238 18053 3290
rect 18077 3238 18087 3290
rect 18087 3238 18133 3290
rect 17837 3236 17893 3238
rect 17917 3236 17973 3238
rect 17997 3236 18053 3238
rect 18077 3236 18133 3238
rect 22058 3834 22114 3836
rect 22138 3834 22194 3836
rect 22218 3834 22274 3836
rect 22298 3834 22354 3836
rect 22058 3782 22104 3834
rect 22104 3782 22114 3834
rect 22138 3782 22168 3834
rect 22168 3782 22180 3834
rect 22180 3782 22194 3834
rect 22218 3782 22232 3834
rect 22232 3782 22244 3834
rect 22244 3782 22274 3834
rect 22298 3782 22308 3834
rect 22308 3782 22354 3834
rect 22058 3780 22114 3782
rect 22138 3780 22194 3782
rect 22218 3780 22274 3782
rect 22298 3780 22354 3782
rect 22058 2746 22114 2748
rect 22138 2746 22194 2748
rect 22218 2746 22274 2748
rect 22298 2746 22354 2748
rect 22058 2694 22104 2746
rect 22104 2694 22114 2746
rect 22138 2694 22168 2746
rect 22168 2694 22180 2746
rect 22180 2694 22194 2746
rect 22218 2694 22232 2746
rect 22232 2694 22244 2746
rect 22244 2694 22274 2746
rect 22298 2694 22308 2746
rect 22308 2694 22354 2746
rect 22058 2692 22114 2694
rect 22138 2692 22194 2694
rect 22218 2692 22274 2694
rect 22298 2692 22354 2694
rect 26278 4378 26334 4380
rect 26358 4378 26414 4380
rect 26438 4378 26494 4380
rect 26518 4378 26574 4380
rect 26278 4326 26324 4378
rect 26324 4326 26334 4378
rect 26358 4326 26388 4378
rect 26388 4326 26400 4378
rect 26400 4326 26414 4378
rect 26438 4326 26452 4378
rect 26452 4326 26464 4378
rect 26464 4326 26494 4378
rect 26518 4326 26528 4378
rect 26528 4326 26574 4378
rect 26278 4324 26334 4326
rect 26358 4324 26414 4326
rect 26438 4324 26494 4326
rect 26518 4324 26574 4326
rect 26278 3290 26334 3292
rect 26358 3290 26414 3292
rect 26438 3290 26494 3292
rect 26518 3290 26574 3292
rect 26278 3238 26324 3290
rect 26324 3238 26334 3290
rect 26358 3238 26388 3290
rect 26388 3238 26400 3290
rect 26400 3238 26414 3290
rect 26438 3238 26452 3290
rect 26452 3238 26464 3290
rect 26464 3238 26494 3290
rect 26518 3238 26528 3290
rect 26528 3238 26574 3290
rect 26278 3236 26334 3238
rect 26358 3236 26414 3238
rect 26438 3236 26494 3238
rect 26518 3236 26574 3238
rect 30499 13626 30555 13628
rect 30579 13626 30635 13628
rect 30659 13626 30715 13628
rect 30739 13626 30795 13628
rect 30499 13574 30545 13626
rect 30545 13574 30555 13626
rect 30579 13574 30609 13626
rect 30609 13574 30621 13626
rect 30621 13574 30635 13626
rect 30659 13574 30673 13626
rect 30673 13574 30685 13626
rect 30685 13574 30715 13626
rect 30739 13574 30749 13626
rect 30749 13574 30795 13626
rect 30499 13572 30555 13574
rect 30579 13572 30635 13574
rect 30659 13572 30715 13574
rect 30739 13572 30795 13574
rect 34719 16346 34775 16348
rect 34799 16346 34855 16348
rect 34879 16346 34935 16348
rect 34959 16346 35015 16348
rect 34719 16294 34765 16346
rect 34765 16294 34775 16346
rect 34799 16294 34829 16346
rect 34829 16294 34841 16346
rect 34841 16294 34855 16346
rect 34879 16294 34893 16346
rect 34893 16294 34905 16346
rect 34905 16294 34935 16346
rect 34959 16294 34969 16346
rect 34969 16294 35015 16346
rect 34719 16292 34775 16294
rect 34799 16292 34855 16294
rect 34879 16292 34935 16294
rect 34959 16292 35015 16294
rect 30499 12538 30555 12540
rect 30579 12538 30635 12540
rect 30659 12538 30715 12540
rect 30739 12538 30795 12540
rect 30499 12486 30545 12538
rect 30545 12486 30555 12538
rect 30579 12486 30609 12538
rect 30609 12486 30621 12538
rect 30621 12486 30635 12538
rect 30659 12486 30673 12538
rect 30673 12486 30685 12538
rect 30685 12486 30715 12538
rect 30739 12486 30749 12538
rect 30749 12486 30795 12538
rect 30499 12484 30555 12486
rect 30579 12484 30635 12486
rect 30659 12484 30715 12486
rect 30739 12484 30795 12486
rect 30499 11450 30555 11452
rect 30579 11450 30635 11452
rect 30659 11450 30715 11452
rect 30739 11450 30795 11452
rect 30499 11398 30545 11450
rect 30545 11398 30555 11450
rect 30579 11398 30609 11450
rect 30609 11398 30621 11450
rect 30621 11398 30635 11450
rect 30659 11398 30673 11450
rect 30673 11398 30685 11450
rect 30685 11398 30715 11450
rect 30739 11398 30749 11450
rect 30749 11398 30795 11450
rect 30499 11396 30555 11398
rect 30579 11396 30635 11398
rect 30659 11396 30715 11398
rect 30739 11396 30795 11398
rect 34719 15258 34775 15260
rect 34799 15258 34855 15260
rect 34879 15258 34935 15260
rect 34959 15258 35015 15260
rect 34719 15206 34765 15258
rect 34765 15206 34775 15258
rect 34799 15206 34829 15258
rect 34829 15206 34841 15258
rect 34841 15206 34855 15258
rect 34879 15206 34893 15258
rect 34893 15206 34905 15258
rect 34905 15206 34935 15258
rect 34959 15206 34969 15258
rect 34969 15206 35015 15258
rect 34719 15204 34775 15206
rect 34799 15204 34855 15206
rect 34879 15204 34935 15206
rect 34959 15204 35015 15206
rect 34719 14170 34775 14172
rect 34799 14170 34855 14172
rect 34879 14170 34935 14172
rect 34959 14170 35015 14172
rect 34719 14118 34765 14170
rect 34765 14118 34775 14170
rect 34799 14118 34829 14170
rect 34829 14118 34841 14170
rect 34841 14118 34855 14170
rect 34879 14118 34893 14170
rect 34893 14118 34905 14170
rect 34905 14118 34935 14170
rect 34959 14118 34969 14170
rect 34969 14118 35015 14170
rect 34719 14116 34775 14118
rect 34799 14116 34855 14118
rect 34879 14116 34935 14118
rect 34959 14116 35015 14118
rect 34719 13082 34775 13084
rect 34799 13082 34855 13084
rect 34879 13082 34935 13084
rect 34959 13082 35015 13084
rect 34719 13030 34765 13082
rect 34765 13030 34775 13082
rect 34799 13030 34829 13082
rect 34829 13030 34841 13082
rect 34841 13030 34855 13082
rect 34879 13030 34893 13082
rect 34893 13030 34905 13082
rect 34905 13030 34935 13082
rect 34959 13030 34969 13082
rect 34969 13030 35015 13082
rect 34719 13028 34775 13030
rect 34799 13028 34855 13030
rect 34879 13028 34935 13030
rect 34959 13028 35015 13030
rect 34719 11994 34775 11996
rect 34799 11994 34855 11996
rect 34879 11994 34935 11996
rect 34959 11994 35015 11996
rect 34719 11942 34765 11994
rect 34765 11942 34775 11994
rect 34799 11942 34829 11994
rect 34829 11942 34841 11994
rect 34841 11942 34855 11994
rect 34879 11942 34893 11994
rect 34893 11942 34905 11994
rect 34905 11942 34935 11994
rect 34959 11942 34969 11994
rect 34969 11942 35015 11994
rect 34719 11940 34775 11942
rect 34799 11940 34855 11942
rect 34879 11940 34935 11942
rect 34959 11940 35015 11942
rect 30499 10362 30555 10364
rect 30579 10362 30635 10364
rect 30659 10362 30715 10364
rect 30739 10362 30795 10364
rect 30499 10310 30545 10362
rect 30545 10310 30555 10362
rect 30579 10310 30609 10362
rect 30609 10310 30621 10362
rect 30621 10310 30635 10362
rect 30659 10310 30673 10362
rect 30673 10310 30685 10362
rect 30685 10310 30715 10362
rect 30739 10310 30749 10362
rect 30749 10310 30795 10362
rect 30499 10308 30555 10310
rect 30579 10308 30635 10310
rect 30659 10308 30715 10310
rect 30739 10308 30795 10310
rect 30499 9274 30555 9276
rect 30579 9274 30635 9276
rect 30659 9274 30715 9276
rect 30739 9274 30795 9276
rect 30499 9222 30545 9274
rect 30545 9222 30555 9274
rect 30579 9222 30609 9274
rect 30609 9222 30621 9274
rect 30621 9222 30635 9274
rect 30659 9222 30673 9274
rect 30673 9222 30685 9274
rect 30685 9222 30715 9274
rect 30739 9222 30749 9274
rect 30749 9222 30795 9274
rect 30499 9220 30555 9222
rect 30579 9220 30635 9222
rect 30659 9220 30715 9222
rect 30739 9220 30795 9222
rect 30499 8186 30555 8188
rect 30579 8186 30635 8188
rect 30659 8186 30715 8188
rect 30739 8186 30795 8188
rect 30499 8134 30545 8186
rect 30545 8134 30555 8186
rect 30579 8134 30609 8186
rect 30609 8134 30621 8186
rect 30621 8134 30635 8186
rect 30659 8134 30673 8186
rect 30673 8134 30685 8186
rect 30685 8134 30715 8186
rect 30739 8134 30749 8186
rect 30749 8134 30795 8186
rect 30499 8132 30555 8134
rect 30579 8132 30635 8134
rect 30659 8132 30715 8134
rect 30739 8132 30795 8134
rect 30499 7098 30555 7100
rect 30579 7098 30635 7100
rect 30659 7098 30715 7100
rect 30739 7098 30795 7100
rect 30499 7046 30545 7098
rect 30545 7046 30555 7098
rect 30579 7046 30609 7098
rect 30609 7046 30621 7098
rect 30621 7046 30635 7098
rect 30659 7046 30673 7098
rect 30673 7046 30685 7098
rect 30685 7046 30715 7098
rect 30739 7046 30749 7098
rect 30749 7046 30795 7098
rect 30499 7044 30555 7046
rect 30579 7044 30635 7046
rect 30659 7044 30715 7046
rect 30739 7044 30795 7046
rect 30499 6010 30555 6012
rect 30579 6010 30635 6012
rect 30659 6010 30715 6012
rect 30739 6010 30795 6012
rect 30499 5958 30545 6010
rect 30545 5958 30555 6010
rect 30579 5958 30609 6010
rect 30609 5958 30621 6010
rect 30621 5958 30635 6010
rect 30659 5958 30673 6010
rect 30673 5958 30685 6010
rect 30685 5958 30715 6010
rect 30739 5958 30749 6010
rect 30749 5958 30795 6010
rect 30499 5956 30555 5958
rect 30579 5956 30635 5958
rect 30659 5956 30715 5958
rect 30739 5956 30795 5958
rect 34719 10906 34775 10908
rect 34799 10906 34855 10908
rect 34879 10906 34935 10908
rect 34959 10906 35015 10908
rect 34719 10854 34765 10906
rect 34765 10854 34775 10906
rect 34799 10854 34829 10906
rect 34829 10854 34841 10906
rect 34841 10854 34855 10906
rect 34879 10854 34893 10906
rect 34893 10854 34905 10906
rect 34905 10854 34935 10906
rect 34959 10854 34969 10906
rect 34969 10854 35015 10906
rect 34719 10852 34775 10854
rect 34799 10852 34855 10854
rect 34879 10852 34935 10854
rect 34959 10852 35015 10854
rect 34719 9818 34775 9820
rect 34799 9818 34855 9820
rect 34879 9818 34935 9820
rect 34959 9818 35015 9820
rect 34719 9766 34765 9818
rect 34765 9766 34775 9818
rect 34799 9766 34829 9818
rect 34829 9766 34841 9818
rect 34841 9766 34855 9818
rect 34879 9766 34893 9818
rect 34893 9766 34905 9818
rect 34905 9766 34935 9818
rect 34959 9766 34969 9818
rect 34969 9766 35015 9818
rect 34719 9764 34775 9766
rect 34799 9764 34855 9766
rect 34879 9764 34935 9766
rect 34959 9764 35015 9766
rect 34719 8730 34775 8732
rect 34799 8730 34855 8732
rect 34879 8730 34935 8732
rect 34959 8730 35015 8732
rect 34719 8678 34765 8730
rect 34765 8678 34775 8730
rect 34799 8678 34829 8730
rect 34829 8678 34841 8730
rect 34841 8678 34855 8730
rect 34879 8678 34893 8730
rect 34893 8678 34905 8730
rect 34905 8678 34935 8730
rect 34959 8678 34969 8730
rect 34969 8678 35015 8730
rect 34719 8676 34775 8678
rect 34799 8676 34855 8678
rect 34879 8676 34935 8678
rect 34959 8676 35015 8678
rect 34719 7642 34775 7644
rect 34799 7642 34855 7644
rect 34879 7642 34935 7644
rect 34959 7642 35015 7644
rect 34719 7590 34765 7642
rect 34765 7590 34775 7642
rect 34799 7590 34829 7642
rect 34829 7590 34841 7642
rect 34841 7590 34855 7642
rect 34879 7590 34893 7642
rect 34893 7590 34905 7642
rect 34905 7590 34935 7642
rect 34959 7590 34969 7642
rect 34969 7590 35015 7642
rect 34719 7588 34775 7590
rect 34799 7588 34855 7590
rect 34879 7588 34935 7590
rect 34959 7588 35015 7590
rect 34719 6554 34775 6556
rect 34799 6554 34855 6556
rect 34879 6554 34935 6556
rect 34959 6554 35015 6556
rect 34719 6502 34765 6554
rect 34765 6502 34775 6554
rect 34799 6502 34829 6554
rect 34829 6502 34841 6554
rect 34841 6502 34855 6554
rect 34879 6502 34893 6554
rect 34893 6502 34905 6554
rect 34905 6502 34935 6554
rect 34959 6502 34969 6554
rect 34969 6502 35015 6554
rect 34719 6500 34775 6502
rect 34799 6500 34855 6502
rect 34879 6500 34935 6502
rect 34959 6500 35015 6502
rect 34719 5466 34775 5468
rect 34799 5466 34855 5468
rect 34879 5466 34935 5468
rect 34959 5466 35015 5468
rect 34719 5414 34765 5466
rect 34765 5414 34775 5466
rect 34799 5414 34829 5466
rect 34829 5414 34841 5466
rect 34841 5414 34855 5466
rect 34879 5414 34893 5466
rect 34893 5414 34905 5466
rect 34905 5414 34935 5466
rect 34959 5414 34969 5466
rect 34969 5414 35015 5466
rect 34719 5412 34775 5414
rect 34799 5412 34855 5414
rect 34879 5412 34935 5414
rect 34959 5412 35015 5414
rect 30499 4922 30555 4924
rect 30579 4922 30635 4924
rect 30659 4922 30715 4924
rect 30739 4922 30795 4924
rect 30499 4870 30545 4922
rect 30545 4870 30555 4922
rect 30579 4870 30609 4922
rect 30609 4870 30621 4922
rect 30621 4870 30635 4922
rect 30659 4870 30673 4922
rect 30673 4870 30685 4922
rect 30685 4870 30715 4922
rect 30739 4870 30749 4922
rect 30749 4870 30795 4922
rect 30499 4868 30555 4870
rect 30579 4868 30635 4870
rect 30659 4868 30715 4870
rect 30739 4868 30795 4870
rect 34719 4378 34775 4380
rect 34799 4378 34855 4380
rect 34879 4378 34935 4380
rect 34959 4378 35015 4380
rect 34719 4326 34765 4378
rect 34765 4326 34775 4378
rect 34799 4326 34829 4378
rect 34829 4326 34841 4378
rect 34841 4326 34855 4378
rect 34879 4326 34893 4378
rect 34893 4326 34905 4378
rect 34905 4326 34935 4378
rect 34959 4326 34969 4378
rect 34969 4326 35015 4378
rect 34719 4324 34775 4326
rect 34799 4324 34855 4326
rect 34879 4324 34935 4326
rect 34959 4324 35015 4326
rect 30499 3834 30555 3836
rect 30579 3834 30635 3836
rect 30659 3834 30715 3836
rect 30739 3834 30795 3836
rect 30499 3782 30545 3834
rect 30545 3782 30555 3834
rect 30579 3782 30609 3834
rect 30609 3782 30621 3834
rect 30621 3782 30635 3834
rect 30659 3782 30673 3834
rect 30673 3782 30685 3834
rect 30685 3782 30715 3834
rect 30739 3782 30749 3834
rect 30749 3782 30795 3834
rect 30499 3780 30555 3782
rect 30579 3780 30635 3782
rect 30659 3780 30715 3782
rect 30739 3780 30795 3782
rect 34719 3290 34775 3292
rect 34799 3290 34855 3292
rect 34879 3290 34935 3292
rect 34959 3290 35015 3292
rect 34719 3238 34765 3290
rect 34765 3238 34775 3290
rect 34799 3238 34829 3290
rect 34829 3238 34841 3290
rect 34841 3238 34855 3290
rect 34879 3238 34893 3290
rect 34893 3238 34905 3290
rect 34905 3238 34935 3290
rect 34959 3238 34969 3290
rect 34969 3238 35015 3290
rect 34719 3236 34775 3238
rect 34799 3236 34855 3238
rect 34879 3236 34935 3238
rect 34959 3236 35015 3238
rect 30499 2746 30555 2748
rect 30579 2746 30635 2748
rect 30659 2746 30715 2748
rect 30739 2746 30795 2748
rect 30499 2694 30545 2746
rect 30545 2694 30555 2746
rect 30579 2694 30609 2746
rect 30609 2694 30621 2746
rect 30621 2694 30635 2746
rect 30659 2694 30673 2746
rect 30673 2694 30685 2746
rect 30685 2694 30715 2746
rect 30739 2694 30749 2746
rect 30749 2694 30795 2746
rect 30499 2692 30555 2694
rect 30579 2692 30635 2694
rect 30659 2692 30715 2694
rect 30739 2692 30795 2694
rect 17837 2202 17893 2204
rect 17917 2202 17973 2204
rect 17997 2202 18053 2204
rect 18077 2202 18133 2204
rect 17837 2150 17883 2202
rect 17883 2150 17893 2202
rect 17917 2150 17947 2202
rect 17947 2150 17959 2202
rect 17959 2150 17973 2202
rect 17997 2150 18011 2202
rect 18011 2150 18023 2202
rect 18023 2150 18053 2202
rect 18077 2150 18087 2202
rect 18087 2150 18133 2202
rect 17837 2148 17893 2150
rect 17917 2148 17973 2150
rect 17997 2148 18053 2150
rect 18077 2148 18133 2150
rect 26278 2202 26334 2204
rect 26358 2202 26414 2204
rect 26438 2202 26494 2204
rect 26518 2202 26574 2204
rect 26278 2150 26324 2202
rect 26324 2150 26334 2202
rect 26358 2150 26388 2202
rect 26388 2150 26400 2202
rect 26400 2150 26414 2202
rect 26438 2150 26452 2202
rect 26452 2150 26464 2202
rect 26464 2150 26494 2202
rect 26518 2150 26528 2202
rect 26528 2150 26574 2202
rect 26278 2148 26334 2150
rect 26358 2148 26414 2150
rect 26438 2148 26494 2150
rect 26518 2148 26574 2150
rect 34719 2202 34775 2204
rect 34799 2202 34855 2204
rect 34879 2202 34935 2204
rect 34959 2202 35015 2204
rect 34719 2150 34765 2202
rect 34765 2150 34775 2202
rect 34799 2150 34829 2202
rect 34829 2150 34841 2202
rect 34841 2150 34855 2202
rect 34879 2150 34893 2202
rect 34893 2150 34905 2202
rect 34905 2150 34935 2202
rect 34959 2150 34969 2202
rect 34969 2150 35015 2202
rect 34719 2148 34775 2150
rect 34799 2148 34855 2150
rect 34879 2148 34935 2150
rect 34959 2148 35015 2150
<< metal3 >>
rect 9386 33760 9702 33761
rect 9386 33696 9392 33760
rect 9456 33696 9472 33760
rect 9536 33696 9552 33760
rect 9616 33696 9632 33760
rect 9696 33696 9702 33760
rect 9386 33695 9702 33696
rect 17827 33760 18143 33761
rect 17827 33696 17833 33760
rect 17897 33696 17913 33760
rect 17977 33696 17993 33760
rect 18057 33696 18073 33760
rect 18137 33696 18143 33760
rect 17827 33695 18143 33696
rect 26268 33760 26584 33761
rect 26268 33696 26274 33760
rect 26338 33696 26354 33760
rect 26418 33696 26434 33760
rect 26498 33696 26514 33760
rect 26578 33696 26584 33760
rect 26268 33695 26584 33696
rect 34709 33760 35025 33761
rect 34709 33696 34715 33760
rect 34779 33696 34795 33760
rect 34859 33696 34875 33760
rect 34939 33696 34955 33760
rect 35019 33696 35025 33760
rect 34709 33695 35025 33696
rect 5166 33216 5482 33217
rect 5166 33152 5172 33216
rect 5236 33152 5252 33216
rect 5316 33152 5332 33216
rect 5396 33152 5412 33216
rect 5476 33152 5482 33216
rect 5166 33151 5482 33152
rect 13607 33216 13923 33217
rect 13607 33152 13613 33216
rect 13677 33152 13693 33216
rect 13757 33152 13773 33216
rect 13837 33152 13853 33216
rect 13917 33152 13923 33216
rect 13607 33151 13923 33152
rect 22048 33216 22364 33217
rect 22048 33152 22054 33216
rect 22118 33152 22134 33216
rect 22198 33152 22214 33216
rect 22278 33152 22294 33216
rect 22358 33152 22364 33216
rect 22048 33151 22364 33152
rect 30489 33216 30805 33217
rect 30489 33152 30495 33216
rect 30559 33152 30575 33216
rect 30639 33152 30655 33216
rect 30719 33152 30735 33216
rect 30799 33152 30805 33216
rect 30489 33151 30805 33152
rect 9386 32672 9702 32673
rect 9386 32608 9392 32672
rect 9456 32608 9472 32672
rect 9536 32608 9552 32672
rect 9616 32608 9632 32672
rect 9696 32608 9702 32672
rect 9386 32607 9702 32608
rect 17827 32672 18143 32673
rect 17827 32608 17833 32672
rect 17897 32608 17913 32672
rect 17977 32608 17993 32672
rect 18057 32608 18073 32672
rect 18137 32608 18143 32672
rect 17827 32607 18143 32608
rect 26268 32672 26584 32673
rect 26268 32608 26274 32672
rect 26338 32608 26354 32672
rect 26418 32608 26434 32672
rect 26498 32608 26514 32672
rect 26578 32608 26584 32672
rect 26268 32607 26584 32608
rect 34709 32672 35025 32673
rect 34709 32608 34715 32672
rect 34779 32608 34795 32672
rect 34859 32608 34875 32672
rect 34939 32608 34955 32672
rect 35019 32608 35025 32672
rect 34709 32607 35025 32608
rect 5166 32128 5482 32129
rect 5166 32064 5172 32128
rect 5236 32064 5252 32128
rect 5316 32064 5332 32128
rect 5396 32064 5412 32128
rect 5476 32064 5482 32128
rect 5166 32063 5482 32064
rect 13607 32128 13923 32129
rect 13607 32064 13613 32128
rect 13677 32064 13693 32128
rect 13757 32064 13773 32128
rect 13837 32064 13853 32128
rect 13917 32064 13923 32128
rect 13607 32063 13923 32064
rect 22048 32128 22364 32129
rect 22048 32064 22054 32128
rect 22118 32064 22134 32128
rect 22198 32064 22214 32128
rect 22278 32064 22294 32128
rect 22358 32064 22364 32128
rect 22048 32063 22364 32064
rect 30489 32128 30805 32129
rect 30489 32064 30495 32128
rect 30559 32064 30575 32128
rect 30639 32064 30655 32128
rect 30719 32064 30735 32128
rect 30799 32064 30805 32128
rect 30489 32063 30805 32064
rect 9386 31584 9702 31585
rect 9386 31520 9392 31584
rect 9456 31520 9472 31584
rect 9536 31520 9552 31584
rect 9616 31520 9632 31584
rect 9696 31520 9702 31584
rect 9386 31519 9702 31520
rect 17827 31584 18143 31585
rect 17827 31520 17833 31584
rect 17897 31520 17913 31584
rect 17977 31520 17993 31584
rect 18057 31520 18073 31584
rect 18137 31520 18143 31584
rect 17827 31519 18143 31520
rect 26268 31584 26584 31585
rect 26268 31520 26274 31584
rect 26338 31520 26354 31584
rect 26418 31520 26434 31584
rect 26498 31520 26514 31584
rect 26578 31520 26584 31584
rect 26268 31519 26584 31520
rect 34709 31584 35025 31585
rect 34709 31520 34715 31584
rect 34779 31520 34795 31584
rect 34859 31520 34875 31584
rect 34939 31520 34955 31584
rect 35019 31520 35025 31584
rect 34709 31519 35025 31520
rect 5166 31040 5482 31041
rect 5166 30976 5172 31040
rect 5236 30976 5252 31040
rect 5316 30976 5332 31040
rect 5396 30976 5412 31040
rect 5476 30976 5482 31040
rect 5166 30975 5482 30976
rect 13607 31040 13923 31041
rect 13607 30976 13613 31040
rect 13677 30976 13693 31040
rect 13757 30976 13773 31040
rect 13837 30976 13853 31040
rect 13917 30976 13923 31040
rect 13607 30975 13923 30976
rect 22048 31040 22364 31041
rect 22048 30976 22054 31040
rect 22118 30976 22134 31040
rect 22198 30976 22214 31040
rect 22278 30976 22294 31040
rect 22358 30976 22364 31040
rect 22048 30975 22364 30976
rect 30489 31040 30805 31041
rect 30489 30976 30495 31040
rect 30559 30976 30575 31040
rect 30639 30976 30655 31040
rect 30719 30976 30735 31040
rect 30799 30976 30805 31040
rect 30489 30975 30805 30976
rect 24945 30836 25011 30837
rect 24894 30772 24900 30836
rect 24964 30834 25011 30836
rect 24964 30832 25056 30834
rect 25006 30776 25056 30832
rect 24964 30774 25056 30776
rect 24964 30772 25011 30774
rect 24945 30771 25011 30772
rect 9386 30496 9702 30497
rect 9386 30432 9392 30496
rect 9456 30432 9472 30496
rect 9536 30432 9552 30496
rect 9616 30432 9632 30496
rect 9696 30432 9702 30496
rect 9386 30431 9702 30432
rect 17827 30496 18143 30497
rect 17827 30432 17833 30496
rect 17897 30432 17913 30496
rect 17977 30432 17993 30496
rect 18057 30432 18073 30496
rect 18137 30432 18143 30496
rect 17827 30431 18143 30432
rect 26268 30496 26584 30497
rect 26268 30432 26274 30496
rect 26338 30432 26354 30496
rect 26418 30432 26434 30496
rect 26498 30432 26514 30496
rect 26578 30432 26584 30496
rect 26268 30431 26584 30432
rect 34709 30496 35025 30497
rect 34709 30432 34715 30496
rect 34779 30432 34795 30496
rect 34859 30432 34875 30496
rect 34939 30432 34955 30496
rect 35019 30432 35025 30496
rect 34709 30431 35025 30432
rect 5166 29952 5482 29953
rect 5166 29888 5172 29952
rect 5236 29888 5252 29952
rect 5316 29888 5332 29952
rect 5396 29888 5412 29952
rect 5476 29888 5482 29952
rect 5166 29887 5482 29888
rect 13607 29952 13923 29953
rect 13607 29888 13613 29952
rect 13677 29888 13693 29952
rect 13757 29888 13773 29952
rect 13837 29888 13853 29952
rect 13917 29888 13923 29952
rect 13607 29887 13923 29888
rect 22048 29952 22364 29953
rect 22048 29888 22054 29952
rect 22118 29888 22134 29952
rect 22198 29888 22214 29952
rect 22278 29888 22294 29952
rect 22358 29888 22364 29952
rect 22048 29887 22364 29888
rect 30489 29952 30805 29953
rect 30489 29888 30495 29952
rect 30559 29888 30575 29952
rect 30639 29888 30655 29952
rect 30719 29888 30735 29952
rect 30799 29888 30805 29952
rect 30489 29887 30805 29888
rect 9386 29408 9702 29409
rect 9386 29344 9392 29408
rect 9456 29344 9472 29408
rect 9536 29344 9552 29408
rect 9616 29344 9632 29408
rect 9696 29344 9702 29408
rect 9386 29343 9702 29344
rect 17827 29408 18143 29409
rect 17827 29344 17833 29408
rect 17897 29344 17913 29408
rect 17977 29344 17993 29408
rect 18057 29344 18073 29408
rect 18137 29344 18143 29408
rect 17827 29343 18143 29344
rect 26268 29408 26584 29409
rect 26268 29344 26274 29408
rect 26338 29344 26354 29408
rect 26418 29344 26434 29408
rect 26498 29344 26514 29408
rect 26578 29344 26584 29408
rect 26268 29343 26584 29344
rect 34709 29408 35025 29409
rect 34709 29344 34715 29408
rect 34779 29344 34795 29408
rect 34859 29344 34875 29408
rect 34939 29344 34955 29408
rect 35019 29344 35025 29408
rect 34709 29343 35025 29344
rect 5166 28864 5482 28865
rect 5166 28800 5172 28864
rect 5236 28800 5252 28864
rect 5316 28800 5332 28864
rect 5396 28800 5412 28864
rect 5476 28800 5482 28864
rect 5166 28799 5482 28800
rect 13607 28864 13923 28865
rect 13607 28800 13613 28864
rect 13677 28800 13693 28864
rect 13757 28800 13773 28864
rect 13837 28800 13853 28864
rect 13917 28800 13923 28864
rect 13607 28799 13923 28800
rect 22048 28864 22364 28865
rect 22048 28800 22054 28864
rect 22118 28800 22134 28864
rect 22198 28800 22214 28864
rect 22278 28800 22294 28864
rect 22358 28800 22364 28864
rect 22048 28799 22364 28800
rect 30489 28864 30805 28865
rect 30489 28800 30495 28864
rect 30559 28800 30575 28864
rect 30639 28800 30655 28864
rect 30719 28800 30735 28864
rect 30799 28800 30805 28864
rect 30489 28799 30805 28800
rect 9386 28320 9702 28321
rect 9386 28256 9392 28320
rect 9456 28256 9472 28320
rect 9536 28256 9552 28320
rect 9616 28256 9632 28320
rect 9696 28256 9702 28320
rect 9386 28255 9702 28256
rect 17827 28320 18143 28321
rect 17827 28256 17833 28320
rect 17897 28256 17913 28320
rect 17977 28256 17993 28320
rect 18057 28256 18073 28320
rect 18137 28256 18143 28320
rect 17827 28255 18143 28256
rect 26268 28320 26584 28321
rect 26268 28256 26274 28320
rect 26338 28256 26354 28320
rect 26418 28256 26434 28320
rect 26498 28256 26514 28320
rect 26578 28256 26584 28320
rect 26268 28255 26584 28256
rect 34709 28320 35025 28321
rect 34709 28256 34715 28320
rect 34779 28256 34795 28320
rect 34859 28256 34875 28320
rect 34939 28256 34955 28320
rect 35019 28256 35025 28320
rect 34709 28255 35025 28256
rect 5166 27776 5482 27777
rect 5166 27712 5172 27776
rect 5236 27712 5252 27776
rect 5316 27712 5332 27776
rect 5396 27712 5412 27776
rect 5476 27712 5482 27776
rect 5166 27711 5482 27712
rect 13607 27776 13923 27777
rect 13607 27712 13613 27776
rect 13677 27712 13693 27776
rect 13757 27712 13773 27776
rect 13837 27712 13853 27776
rect 13917 27712 13923 27776
rect 13607 27711 13923 27712
rect 22048 27776 22364 27777
rect 22048 27712 22054 27776
rect 22118 27712 22134 27776
rect 22198 27712 22214 27776
rect 22278 27712 22294 27776
rect 22358 27712 22364 27776
rect 22048 27711 22364 27712
rect 30489 27776 30805 27777
rect 30489 27712 30495 27776
rect 30559 27712 30575 27776
rect 30639 27712 30655 27776
rect 30719 27712 30735 27776
rect 30799 27712 30805 27776
rect 30489 27711 30805 27712
rect 9386 27232 9702 27233
rect 9386 27168 9392 27232
rect 9456 27168 9472 27232
rect 9536 27168 9552 27232
rect 9616 27168 9632 27232
rect 9696 27168 9702 27232
rect 9386 27167 9702 27168
rect 17827 27232 18143 27233
rect 17827 27168 17833 27232
rect 17897 27168 17913 27232
rect 17977 27168 17993 27232
rect 18057 27168 18073 27232
rect 18137 27168 18143 27232
rect 17827 27167 18143 27168
rect 26268 27232 26584 27233
rect 26268 27168 26274 27232
rect 26338 27168 26354 27232
rect 26418 27168 26434 27232
rect 26498 27168 26514 27232
rect 26578 27168 26584 27232
rect 26268 27167 26584 27168
rect 34709 27232 35025 27233
rect 34709 27168 34715 27232
rect 34779 27168 34795 27232
rect 34859 27168 34875 27232
rect 34939 27168 34955 27232
rect 35019 27168 35025 27232
rect 34709 27167 35025 27168
rect 5166 26688 5482 26689
rect 5166 26624 5172 26688
rect 5236 26624 5252 26688
rect 5316 26624 5332 26688
rect 5396 26624 5412 26688
rect 5476 26624 5482 26688
rect 5166 26623 5482 26624
rect 13607 26688 13923 26689
rect 13607 26624 13613 26688
rect 13677 26624 13693 26688
rect 13757 26624 13773 26688
rect 13837 26624 13853 26688
rect 13917 26624 13923 26688
rect 13607 26623 13923 26624
rect 22048 26688 22364 26689
rect 22048 26624 22054 26688
rect 22118 26624 22134 26688
rect 22198 26624 22214 26688
rect 22278 26624 22294 26688
rect 22358 26624 22364 26688
rect 22048 26623 22364 26624
rect 30489 26688 30805 26689
rect 30489 26624 30495 26688
rect 30559 26624 30575 26688
rect 30639 26624 30655 26688
rect 30719 26624 30735 26688
rect 30799 26624 30805 26688
rect 30489 26623 30805 26624
rect 9386 26144 9702 26145
rect 9386 26080 9392 26144
rect 9456 26080 9472 26144
rect 9536 26080 9552 26144
rect 9616 26080 9632 26144
rect 9696 26080 9702 26144
rect 9386 26079 9702 26080
rect 17827 26144 18143 26145
rect 17827 26080 17833 26144
rect 17897 26080 17913 26144
rect 17977 26080 17993 26144
rect 18057 26080 18073 26144
rect 18137 26080 18143 26144
rect 17827 26079 18143 26080
rect 26268 26144 26584 26145
rect 26268 26080 26274 26144
rect 26338 26080 26354 26144
rect 26418 26080 26434 26144
rect 26498 26080 26514 26144
rect 26578 26080 26584 26144
rect 26268 26079 26584 26080
rect 34709 26144 35025 26145
rect 34709 26080 34715 26144
rect 34779 26080 34795 26144
rect 34859 26080 34875 26144
rect 34939 26080 34955 26144
rect 35019 26080 35025 26144
rect 34709 26079 35025 26080
rect 5166 25600 5482 25601
rect 5166 25536 5172 25600
rect 5236 25536 5252 25600
rect 5316 25536 5332 25600
rect 5396 25536 5412 25600
rect 5476 25536 5482 25600
rect 5166 25535 5482 25536
rect 13607 25600 13923 25601
rect 13607 25536 13613 25600
rect 13677 25536 13693 25600
rect 13757 25536 13773 25600
rect 13837 25536 13853 25600
rect 13917 25536 13923 25600
rect 13607 25535 13923 25536
rect 22048 25600 22364 25601
rect 22048 25536 22054 25600
rect 22118 25536 22134 25600
rect 22198 25536 22214 25600
rect 22278 25536 22294 25600
rect 22358 25536 22364 25600
rect 22048 25535 22364 25536
rect 30489 25600 30805 25601
rect 30489 25536 30495 25600
rect 30559 25536 30575 25600
rect 30639 25536 30655 25600
rect 30719 25536 30735 25600
rect 30799 25536 30805 25600
rect 30489 25535 30805 25536
rect 9386 25056 9702 25057
rect 9386 24992 9392 25056
rect 9456 24992 9472 25056
rect 9536 24992 9552 25056
rect 9616 24992 9632 25056
rect 9696 24992 9702 25056
rect 9386 24991 9702 24992
rect 17827 25056 18143 25057
rect 17827 24992 17833 25056
rect 17897 24992 17913 25056
rect 17977 24992 17993 25056
rect 18057 24992 18073 25056
rect 18137 24992 18143 25056
rect 17827 24991 18143 24992
rect 26268 25056 26584 25057
rect 26268 24992 26274 25056
rect 26338 24992 26354 25056
rect 26418 24992 26434 25056
rect 26498 24992 26514 25056
rect 26578 24992 26584 25056
rect 26268 24991 26584 24992
rect 34709 25056 35025 25057
rect 34709 24992 34715 25056
rect 34779 24992 34795 25056
rect 34859 24992 34875 25056
rect 34939 24992 34955 25056
rect 35019 24992 35025 25056
rect 34709 24991 35025 24992
rect 5166 24512 5482 24513
rect 5166 24448 5172 24512
rect 5236 24448 5252 24512
rect 5316 24448 5332 24512
rect 5396 24448 5412 24512
rect 5476 24448 5482 24512
rect 5166 24447 5482 24448
rect 13607 24512 13923 24513
rect 13607 24448 13613 24512
rect 13677 24448 13693 24512
rect 13757 24448 13773 24512
rect 13837 24448 13853 24512
rect 13917 24448 13923 24512
rect 13607 24447 13923 24448
rect 22048 24512 22364 24513
rect 22048 24448 22054 24512
rect 22118 24448 22134 24512
rect 22198 24448 22214 24512
rect 22278 24448 22294 24512
rect 22358 24448 22364 24512
rect 22048 24447 22364 24448
rect 30489 24512 30805 24513
rect 30489 24448 30495 24512
rect 30559 24448 30575 24512
rect 30639 24448 30655 24512
rect 30719 24448 30735 24512
rect 30799 24448 30805 24512
rect 30489 24447 30805 24448
rect 9386 23968 9702 23969
rect 9386 23904 9392 23968
rect 9456 23904 9472 23968
rect 9536 23904 9552 23968
rect 9616 23904 9632 23968
rect 9696 23904 9702 23968
rect 9386 23903 9702 23904
rect 17827 23968 18143 23969
rect 17827 23904 17833 23968
rect 17897 23904 17913 23968
rect 17977 23904 17993 23968
rect 18057 23904 18073 23968
rect 18137 23904 18143 23968
rect 17827 23903 18143 23904
rect 26268 23968 26584 23969
rect 26268 23904 26274 23968
rect 26338 23904 26354 23968
rect 26418 23904 26434 23968
rect 26498 23904 26514 23968
rect 26578 23904 26584 23968
rect 26268 23903 26584 23904
rect 34709 23968 35025 23969
rect 34709 23904 34715 23968
rect 34779 23904 34795 23968
rect 34859 23904 34875 23968
rect 34939 23904 34955 23968
rect 35019 23904 35025 23968
rect 34709 23903 35025 23904
rect 19701 23898 19767 23901
rect 20713 23898 20779 23901
rect 19701 23896 20779 23898
rect 19701 23840 19706 23896
rect 19762 23840 20718 23896
rect 20774 23840 20779 23896
rect 19701 23838 20779 23840
rect 19701 23835 19767 23838
rect 20713 23835 20779 23838
rect 5166 23424 5482 23425
rect 5166 23360 5172 23424
rect 5236 23360 5252 23424
rect 5316 23360 5332 23424
rect 5396 23360 5412 23424
rect 5476 23360 5482 23424
rect 5166 23359 5482 23360
rect 13607 23424 13923 23425
rect 13607 23360 13613 23424
rect 13677 23360 13693 23424
rect 13757 23360 13773 23424
rect 13837 23360 13853 23424
rect 13917 23360 13923 23424
rect 13607 23359 13923 23360
rect 22048 23424 22364 23425
rect 22048 23360 22054 23424
rect 22118 23360 22134 23424
rect 22198 23360 22214 23424
rect 22278 23360 22294 23424
rect 22358 23360 22364 23424
rect 22048 23359 22364 23360
rect 30489 23424 30805 23425
rect 30489 23360 30495 23424
rect 30559 23360 30575 23424
rect 30639 23360 30655 23424
rect 30719 23360 30735 23424
rect 30799 23360 30805 23424
rect 30489 23359 30805 23360
rect 22185 23218 22251 23221
rect 24894 23218 24900 23220
rect 22185 23216 24900 23218
rect 22185 23160 22190 23216
rect 22246 23160 24900 23216
rect 22185 23158 24900 23160
rect 22185 23155 22251 23158
rect 24894 23156 24900 23158
rect 24964 23156 24970 23220
rect 9386 22880 9702 22881
rect 9386 22816 9392 22880
rect 9456 22816 9472 22880
rect 9536 22816 9552 22880
rect 9616 22816 9632 22880
rect 9696 22816 9702 22880
rect 9386 22815 9702 22816
rect 17827 22880 18143 22881
rect 17827 22816 17833 22880
rect 17897 22816 17913 22880
rect 17977 22816 17993 22880
rect 18057 22816 18073 22880
rect 18137 22816 18143 22880
rect 17827 22815 18143 22816
rect 26268 22880 26584 22881
rect 26268 22816 26274 22880
rect 26338 22816 26354 22880
rect 26418 22816 26434 22880
rect 26498 22816 26514 22880
rect 26578 22816 26584 22880
rect 26268 22815 26584 22816
rect 34709 22880 35025 22881
rect 34709 22816 34715 22880
rect 34779 22816 34795 22880
rect 34859 22816 34875 22880
rect 34939 22816 34955 22880
rect 35019 22816 35025 22880
rect 34709 22815 35025 22816
rect 5166 22336 5482 22337
rect 5166 22272 5172 22336
rect 5236 22272 5252 22336
rect 5316 22272 5332 22336
rect 5396 22272 5412 22336
rect 5476 22272 5482 22336
rect 5166 22271 5482 22272
rect 13607 22336 13923 22337
rect 13607 22272 13613 22336
rect 13677 22272 13693 22336
rect 13757 22272 13773 22336
rect 13837 22272 13853 22336
rect 13917 22272 13923 22336
rect 13607 22271 13923 22272
rect 22048 22336 22364 22337
rect 22048 22272 22054 22336
rect 22118 22272 22134 22336
rect 22198 22272 22214 22336
rect 22278 22272 22294 22336
rect 22358 22272 22364 22336
rect 22048 22271 22364 22272
rect 30489 22336 30805 22337
rect 30489 22272 30495 22336
rect 30559 22272 30575 22336
rect 30639 22272 30655 22336
rect 30719 22272 30735 22336
rect 30799 22272 30805 22336
rect 30489 22271 30805 22272
rect 20437 22130 20503 22133
rect 27245 22130 27311 22133
rect 20437 22128 27311 22130
rect 20437 22072 20442 22128
rect 20498 22072 27250 22128
rect 27306 22072 27311 22128
rect 20437 22070 27311 22072
rect 20437 22067 20503 22070
rect 27245 22067 27311 22070
rect 9386 21792 9702 21793
rect 9386 21728 9392 21792
rect 9456 21728 9472 21792
rect 9536 21728 9552 21792
rect 9616 21728 9632 21792
rect 9696 21728 9702 21792
rect 9386 21727 9702 21728
rect 17827 21792 18143 21793
rect 17827 21728 17833 21792
rect 17897 21728 17913 21792
rect 17977 21728 17993 21792
rect 18057 21728 18073 21792
rect 18137 21728 18143 21792
rect 17827 21727 18143 21728
rect 26268 21792 26584 21793
rect 26268 21728 26274 21792
rect 26338 21728 26354 21792
rect 26418 21728 26434 21792
rect 26498 21728 26514 21792
rect 26578 21728 26584 21792
rect 26268 21727 26584 21728
rect 34709 21792 35025 21793
rect 34709 21728 34715 21792
rect 34779 21728 34795 21792
rect 34859 21728 34875 21792
rect 34939 21728 34955 21792
rect 35019 21728 35025 21792
rect 34709 21727 35025 21728
rect 5166 21248 5482 21249
rect 5166 21184 5172 21248
rect 5236 21184 5252 21248
rect 5316 21184 5332 21248
rect 5396 21184 5412 21248
rect 5476 21184 5482 21248
rect 5166 21183 5482 21184
rect 13607 21248 13923 21249
rect 13607 21184 13613 21248
rect 13677 21184 13693 21248
rect 13757 21184 13773 21248
rect 13837 21184 13853 21248
rect 13917 21184 13923 21248
rect 13607 21183 13923 21184
rect 22048 21248 22364 21249
rect 22048 21184 22054 21248
rect 22118 21184 22134 21248
rect 22198 21184 22214 21248
rect 22278 21184 22294 21248
rect 22358 21184 22364 21248
rect 22048 21183 22364 21184
rect 30489 21248 30805 21249
rect 30489 21184 30495 21248
rect 30559 21184 30575 21248
rect 30639 21184 30655 21248
rect 30719 21184 30735 21248
rect 30799 21184 30805 21248
rect 30489 21183 30805 21184
rect 9386 20704 9702 20705
rect 9386 20640 9392 20704
rect 9456 20640 9472 20704
rect 9536 20640 9552 20704
rect 9616 20640 9632 20704
rect 9696 20640 9702 20704
rect 9386 20639 9702 20640
rect 17827 20704 18143 20705
rect 17827 20640 17833 20704
rect 17897 20640 17913 20704
rect 17977 20640 17993 20704
rect 18057 20640 18073 20704
rect 18137 20640 18143 20704
rect 17827 20639 18143 20640
rect 26268 20704 26584 20705
rect 26268 20640 26274 20704
rect 26338 20640 26354 20704
rect 26418 20640 26434 20704
rect 26498 20640 26514 20704
rect 26578 20640 26584 20704
rect 26268 20639 26584 20640
rect 34709 20704 35025 20705
rect 34709 20640 34715 20704
rect 34779 20640 34795 20704
rect 34859 20640 34875 20704
rect 34939 20640 34955 20704
rect 35019 20640 35025 20704
rect 34709 20639 35025 20640
rect 5166 20160 5482 20161
rect 5166 20096 5172 20160
rect 5236 20096 5252 20160
rect 5316 20096 5332 20160
rect 5396 20096 5412 20160
rect 5476 20096 5482 20160
rect 5166 20095 5482 20096
rect 13607 20160 13923 20161
rect 13607 20096 13613 20160
rect 13677 20096 13693 20160
rect 13757 20096 13773 20160
rect 13837 20096 13853 20160
rect 13917 20096 13923 20160
rect 13607 20095 13923 20096
rect 22048 20160 22364 20161
rect 22048 20096 22054 20160
rect 22118 20096 22134 20160
rect 22198 20096 22214 20160
rect 22278 20096 22294 20160
rect 22358 20096 22364 20160
rect 22048 20095 22364 20096
rect 30489 20160 30805 20161
rect 30489 20096 30495 20160
rect 30559 20096 30575 20160
rect 30639 20096 30655 20160
rect 30719 20096 30735 20160
rect 30799 20096 30805 20160
rect 30489 20095 30805 20096
rect 9386 19616 9702 19617
rect 9386 19552 9392 19616
rect 9456 19552 9472 19616
rect 9536 19552 9552 19616
rect 9616 19552 9632 19616
rect 9696 19552 9702 19616
rect 9386 19551 9702 19552
rect 17827 19616 18143 19617
rect 17827 19552 17833 19616
rect 17897 19552 17913 19616
rect 17977 19552 17993 19616
rect 18057 19552 18073 19616
rect 18137 19552 18143 19616
rect 17827 19551 18143 19552
rect 26268 19616 26584 19617
rect 26268 19552 26274 19616
rect 26338 19552 26354 19616
rect 26418 19552 26434 19616
rect 26498 19552 26514 19616
rect 26578 19552 26584 19616
rect 26268 19551 26584 19552
rect 34709 19616 35025 19617
rect 34709 19552 34715 19616
rect 34779 19552 34795 19616
rect 34859 19552 34875 19616
rect 34939 19552 34955 19616
rect 35019 19552 35025 19616
rect 34709 19551 35025 19552
rect 5166 19072 5482 19073
rect 5166 19008 5172 19072
rect 5236 19008 5252 19072
rect 5316 19008 5332 19072
rect 5396 19008 5412 19072
rect 5476 19008 5482 19072
rect 5166 19007 5482 19008
rect 13607 19072 13923 19073
rect 13607 19008 13613 19072
rect 13677 19008 13693 19072
rect 13757 19008 13773 19072
rect 13837 19008 13853 19072
rect 13917 19008 13923 19072
rect 13607 19007 13923 19008
rect 22048 19072 22364 19073
rect 22048 19008 22054 19072
rect 22118 19008 22134 19072
rect 22198 19008 22214 19072
rect 22278 19008 22294 19072
rect 22358 19008 22364 19072
rect 22048 19007 22364 19008
rect 30489 19072 30805 19073
rect 30489 19008 30495 19072
rect 30559 19008 30575 19072
rect 30639 19008 30655 19072
rect 30719 19008 30735 19072
rect 30799 19008 30805 19072
rect 30489 19007 30805 19008
rect 9386 18528 9702 18529
rect 9386 18464 9392 18528
rect 9456 18464 9472 18528
rect 9536 18464 9552 18528
rect 9616 18464 9632 18528
rect 9696 18464 9702 18528
rect 9386 18463 9702 18464
rect 17827 18528 18143 18529
rect 17827 18464 17833 18528
rect 17897 18464 17913 18528
rect 17977 18464 17993 18528
rect 18057 18464 18073 18528
rect 18137 18464 18143 18528
rect 17827 18463 18143 18464
rect 26268 18528 26584 18529
rect 26268 18464 26274 18528
rect 26338 18464 26354 18528
rect 26418 18464 26434 18528
rect 26498 18464 26514 18528
rect 26578 18464 26584 18528
rect 26268 18463 26584 18464
rect 34709 18528 35025 18529
rect 34709 18464 34715 18528
rect 34779 18464 34795 18528
rect 34859 18464 34875 18528
rect 34939 18464 34955 18528
rect 35019 18464 35025 18528
rect 34709 18463 35025 18464
rect 5166 17984 5482 17985
rect 5166 17920 5172 17984
rect 5236 17920 5252 17984
rect 5316 17920 5332 17984
rect 5396 17920 5412 17984
rect 5476 17920 5482 17984
rect 5166 17919 5482 17920
rect 13607 17984 13923 17985
rect 13607 17920 13613 17984
rect 13677 17920 13693 17984
rect 13757 17920 13773 17984
rect 13837 17920 13853 17984
rect 13917 17920 13923 17984
rect 13607 17919 13923 17920
rect 22048 17984 22364 17985
rect 22048 17920 22054 17984
rect 22118 17920 22134 17984
rect 22198 17920 22214 17984
rect 22278 17920 22294 17984
rect 22358 17920 22364 17984
rect 22048 17919 22364 17920
rect 30489 17984 30805 17985
rect 30489 17920 30495 17984
rect 30559 17920 30575 17984
rect 30639 17920 30655 17984
rect 30719 17920 30735 17984
rect 30799 17920 30805 17984
rect 30489 17919 30805 17920
rect 34329 17914 34395 17917
rect 35200 17914 36000 17944
rect 34329 17912 36000 17914
rect 34329 17856 34334 17912
rect 34390 17856 36000 17912
rect 34329 17854 36000 17856
rect 34329 17851 34395 17854
rect 35200 17824 36000 17854
rect 9386 17440 9702 17441
rect 9386 17376 9392 17440
rect 9456 17376 9472 17440
rect 9536 17376 9552 17440
rect 9616 17376 9632 17440
rect 9696 17376 9702 17440
rect 9386 17375 9702 17376
rect 17827 17440 18143 17441
rect 17827 17376 17833 17440
rect 17897 17376 17913 17440
rect 17977 17376 17993 17440
rect 18057 17376 18073 17440
rect 18137 17376 18143 17440
rect 17827 17375 18143 17376
rect 26268 17440 26584 17441
rect 26268 17376 26274 17440
rect 26338 17376 26354 17440
rect 26418 17376 26434 17440
rect 26498 17376 26514 17440
rect 26578 17376 26584 17440
rect 26268 17375 26584 17376
rect 34709 17440 35025 17441
rect 34709 17376 34715 17440
rect 34779 17376 34795 17440
rect 34859 17376 34875 17440
rect 34939 17376 34955 17440
rect 35019 17376 35025 17440
rect 34709 17375 35025 17376
rect 5166 16896 5482 16897
rect 5166 16832 5172 16896
rect 5236 16832 5252 16896
rect 5316 16832 5332 16896
rect 5396 16832 5412 16896
rect 5476 16832 5482 16896
rect 5166 16831 5482 16832
rect 13607 16896 13923 16897
rect 13607 16832 13613 16896
rect 13677 16832 13693 16896
rect 13757 16832 13773 16896
rect 13837 16832 13853 16896
rect 13917 16832 13923 16896
rect 13607 16831 13923 16832
rect 22048 16896 22364 16897
rect 22048 16832 22054 16896
rect 22118 16832 22134 16896
rect 22198 16832 22214 16896
rect 22278 16832 22294 16896
rect 22358 16832 22364 16896
rect 22048 16831 22364 16832
rect 30489 16896 30805 16897
rect 30489 16832 30495 16896
rect 30559 16832 30575 16896
rect 30639 16832 30655 16896
rect 30719 16832 30735 16896
rect 30799 16832 30805 16896
rect 30489 16831 30805 16832
rect 9386 16352 9702 16353
rect 9386 16288 9392 16352
rect 9456 16288 9472 16352
rect 9536 16288 9552 16352
rect 9616 16288 9632 16352
rect 9696 16288 9702 16352
rect 9386 16287 9702 16288
rect 17827 16352 18143 16353
rect 17827 16288 17833 16352
rect 17897 16288 17913 16352
rect 17977 16288 17993 16352
rect 18057 16288 18073 16352
rect 18137 16288 18143 16352
rect 17827 16287 18143 16288
rect 26268 16352 26584 16353
rect 26268 16288 26274 16352
rect 26338 16288 26354 16352
rect 26418 16288 26434 16352
rect 26498 16288 26514 16352
rect 26578 16288 26584 16352
rect 26268 16287 26584 16288
rect 34709 16352 35025 16353
rect 34709 16288 34715 16352
rect 34779 16288 34795 16352
rect 34859 16288 34875 16352
rect 34939 16288 34955 16352
rect 35019 16288 35025 16352
rect 34709 16287 35025 16288
rect 5166 15808 5482 15809
rect 5166 15744 5172 15808
rect 5236 15744 5252 15808
rect 5316 15744 5332 15808
rect 5396 15744 5412 15808
rect 5476 15744 5482 15808
rect 5166 15743 5482 15744
rect 13607 15808 13923 15809
rect 13607 15744 13613 15808
rect 13677 15744 13693 15808
rect 13757 15744 13773 15808
rect 13837 15744 13853 15808
rect 13917 15744 13923 15808
rect 13607 15743 13923 15744
rect 22048 15808 22364 15809
rect 22048 15744 22054 15808
rect 22118 15744 22134 15808
rect 22198 15744 22214 15808
rect 22278 15744 22294 15808
rect 22358 15744 22364 15808
rect 22048 15743 22364 15744
rect 30489 15808 30805 15809
rect 30489 15744 30495 15808
rect 30559 15744 30575 15808
rect 30639 15744 30655 15808
rect 30719 15744 30735 15808
rect 30799 15744 30805 15808
rect 30489 15743 30805 15744
rect 9386 15264 9702 15265
rect 9386 15200 9392 15264
rect 9456 15200 9472 15264
rect 9536 15200 9552 15264
rect 9616 15200 9632 15264
rect 9696 15200 9702 15264
rect 9386 15199 9702 15200
rect 17827 15264 18143 15265
rect 17827 15200 17833 15264
rect 17897 15200 17913 15264
rect 17977 15200 17993 15264
rect 18057 15200 18073 15264
rect 18137 15200 18143 15264
rect 17827 15199 18143 15200
rect 26268 15264 26584 15265
rect 26268 15200 26274 15264
rect 26338 15200 26354 15264
rect 26418 15200 26434 15264
rect 26498 15200 26514 15264
rect 26578 15200 26584 15264
rect 26268 15199 26584 15200
rect 34709 15264 35025 15265
rect 34709 15200 34715 15264
rect 34779 15200 34795 15264
rect 34859 15200 34875 15264
rect 34939 15200 34955 15264
rect 35019 15200 35025 15264
rect 34709 15199 35025 15200
rect 19885 14922 19951 14925
rect 22185 14922 22251 14925
rect 24669 14922 24735 14925
rect 19885 14920 24735 14922
rect 19885 14864 19890 14920
rect 19946 14864 22190 14920
rect 22246 14864 24674 14920
rect 24730 14864 24735 14920
rect 19885 14862 24735 14864
rect 19885 14859 19951 14862
rect 22185 14859 22251 14862
rect 24669 14859 24735 14862
rect 5166 14720 5482 14721
rect 5166 14656 5172 14720
rect 5236 14656 5252 14720
rect 5316 14656 5332 14720
rect 5396 14656 5412 14720
rect 5476 14656 5482 14720
rect 5166 14655 5482 14656
rect 13607 14720 13923 14721
rect 13607 14656 13613 14720
rect 13677 14656 13693 14720
rect 13757 14656 13773 14720
rect 13837 14656 13853 14720
rect 13917 14656 13923 14720
rect 13607 14655 13923 14656
rect 22048 14720 22364 14721
rect 22048 14656 22054 14720
rect 22118 14656 22134 14720
rect 22198 14656 22214 14720
rect 22278 14656 22294 14720
rect 22358 14656 22364 14720
rect 22048 14655 22364 14656
rect 30489 14720 30805 14721
rect 30489 14656 30495 14720
rect 30559 14656 30575 14720
rect 30639 14656 30655 14720
rect 30719 14656 30735 14720
rect 30799 14656 30805 14720
rect 30489 14655 30805 14656
rect 19517 14378 19583 14381
rect 22553 14378 22619 14381
rect 23565 14378 23631 14381
rect 28717 14378 28783 14381
rect 19517 14376 28783 14378
rect 19517 14320 19522 14376
rect 19578 14320 22558 14376
rect 22614 14320 23570 14376
rect 23626 14320 28722 14376
rect 28778 14320 28783 14376
rect 19517 14318 28783 14320
rect 19517 14315 19583 14318
rect 22553 14315 22619 14318
rect 23565 14315 23631 14318
rect 28717 14315 28783 14318
rect 9386 14176 9702 14177
rect 9386 14112 9392 14176
rect 9456 14112 9472 14176
rect 9536 14112 9552 14176
rect 9616 14112 9632 14176
rect 9696 14112 9702 14176
rect 9386 14111 9702 14112
rect 17827 14176 18143 14177
rect 17827 14112 17833 14176
rect 17897 14112 17913 14176
rect 17977 14112 17993 14176
rect 18057 14112 18073 14176
rect 18137 14112 18143 14176
rect 17827 14111 18143 14112
rect 26268 14176 26584 14177
rect 26268 14112 26274 14176
rect 26338 14112 26354 14176
rect 26418 14112 26434 14176
rect 26498 14112 26514 14176
rect 26578 14112 26584 14176
rect 26268 14111 26584 14112
rect 34709 14176 35025 14177
rect 34709 14112 34715 14176
rect 34779 14112 34795 14176
rect 34859 14112 34875 14176
rect 34939 14112 34955 14176
rect 35019 14112 35025 14176
rect 34709 14111 35025 14112
rect 19793 13970 19859 13973
rect 27797 13970 27863 13973
rect 19793 13968 27863 13970
rect 19793 13912 19798 13968
rect 19854 13912 27802 13968
rect 27858 13912 27863 13968
rect 19793 13910 27863 13912
rect 19793 13907 19859 13910
rect 27797 13907 27863 13910
rect 5166 13632 5482 13633
rect 5166 13568 5172 13632
rect 5236 13568 5252 13632
rect 5316 13568 5332 13632
rect 5396 13568 5412 13632
rect 5476 13568 5482 13632
rect 5166 13567 5482 13568
rect 13607 13632 13923 13633
rect 13607 13568 13613 13632
rect 13677 13568 13693 13632
rect 13757 13568 13773 13632
rect 13837 13568 13853 13632
rect 13917 13568 13923 13632
rect 13607 13567 13923 13568
rect 22048 13632 22364 13633
rect 22048 13568 22054 13632
rect 22118 13568 22134 13632
rect 22198 13568 22214 13632
rect 22278 13568 22294 13632
rect 22358 13568 22364 13632
rect 22048 13567 22364 13568
rect 30489 13632 30805 13633
rect 30489 13568 30495 13632
rect 30559 13568 30575 13632
rect 30639 13568 30655 13632
rect 30719 13568 30735 13632
rect 30799 13568 30805 13632
rect 30489 13567 30805 13568
rect 9386 13088 9702 13089
rect 9386 13024 9392 13088
rect 9456 13024 9472 13088
rect 9536 13024 9552 13088
rect 9616 13024 9632 13088
rect 9696 13024 9702 13088
rect 9386 13023 9702 13024
rect 17827 13088 18143 13089
rect 17827 13024 17833 13088
rect 17897 13024 17913 13088
rect 17977 13024 17993 13088
rect 18057 13024 18073 13088
rect 18137 13024 18143 13088
rect 17827 13023 18143 13024
rect 26268 13088 26584 13089
rect 26268 13024 26274 13088
rect 26338 13024 26354 13088
rect 26418 13024 26434 13088
rect 26498 13024 26514 13088
rect 26578 13024 26584 13088
rect 26268 13023 26584 13024
rect 34709 13088 35025 13089
rect 34709 13024 34715 13088
rect 34779 13024 34795 13088
rect 34859 13024 34875 13088
rect 34939 13024 34955 13088
rect 35019 13024 35025 13088
rect 34709 13023 35025 13024
rect 5166 12544 5482 12545
rect 5166 12480 5172 12544
rect 5236 12480 5252 12544
rect 5316 12480 5332 12544
rect 5396 12480 5412 12544
rect 5476 12480 5482 12544
rect 5166 12479 5482 12480
rect 13607 12544 13923 12545
rect 13607 12480 13613 12544
rect 13677 12480 13693 12544
rect 13757 12480 13773 12544
rect 13837 12480 13853 12544
rect 13917 12480 13923 12544
rect 13607 12479 13923 12480
rect 22048 12544 22364 12545
rect 22048 12480 22054 12544
rect 22118 12480 22134 12544
rect 22198 12480 22214 12544
rect 22278 12480 22294 12544
rect 22358 12480 22364 12544
rect 22048 12479 22364 12480
rect 30489 12544 30805 12545
rect 30489 12480 30495 12544
rect 30559 12480 30575 12544
rect 30639 12480 30655 12544
rect 30719 12480 30735 12544
rect 30799 12480 30805 12544
rect 30489 12479 30805 12480
rect 16113 12474 16179 12477
rect 19333 12474 19399 12477
rect 16113 12472 19399 12474
rect 16113 12416 16118 12472
rect 16174 12416 19338 12472
rect 19394 12416 19399 12472
rect 16113 12414 19399 12416
rect 16113 12411 16179 12414
rect 19333 12411 19399 12414
rect 22645 12474 22711 12477
rect 22645 12472 22754 12474
rect 22645 12416 22650 12472
rect 22706 12416 22754 12472
rect 22645 12411 22754 12416
rect 22694 12338 22754 12411
rect 28073 12338 28139 12341
rect 22694 12336 28139 12338
rect 22694 12280 28078 12336
rect 28134 12280 28139 12336
rect 22694 12278 28139 12280
rect 28073 12275 28139 12278
rect 9386 12000 9702 12001
rect 9386 11936 9392 12000
rect 9456 11936 9472 12000
rect 9536 11936 9552 12000
rect 9616 11936 9632 12000
rect 9696 11936 9702 12000
rect 9386 11935 9702 11936
rect 17827 12000 18143 12001
rect 17827 11936 17833 12000
rect 17897 11936 17913 12000
rect 17977 11936 17993 12000
rect 18057 11936 18073 12000
rect 18137 11936 18143 12000
rect 17827 11935 18143 11936
rect 26268 12000 26584 12001
rect 26268 11936 26274 12000
rect 26338 11936 26354 12000
rect 26418 11936 26434 12000
rect 26498 11936 26514 12000
rect 26578 11936 26584 12000
rect 26268 11935 26584 11936
rect 34709 12000 35025 12001
rect 34709 11936 34715 12000
rect 34779 11936 34795 12000
rect 34859 11936 34875 12000
rect 34939 11936 34955 12000
rect 35019 11936 35025 12000
rect 34709 11935 35025 11936
rect 5166 11456 5482 11457
rect 5166 11392 5172 11456
rect 5236 11392 5252 11456
rect 5316 11392 5332 11456
rect 5396 11392 5412 11456
rect 5476 11392 5482 11456
rect 5166 11391 5482 11392
rect 13607 11456 13923 11457
rect 13607 11392 13613 11456
rect 13677 11392 13693 11456
rect 13757 11392 13773 11456
rect 13837 11392 13853 11456
rect 13917 11392 13923 11456
rect 13607 11391 13923 11392
rect 22048 11456 22364 11457
rect 22048 11392 22054 11456
rect 22118 11392 22134 11456
rect 22198 11392 22214 11456
rect 22278 11392 22294 11456
rect 22358 11392 22364 11456
rect 22048 11391 22364 11392
rect 30489 11456 30805 11457
rect 30489 11392 30495 11456
rect 30559 11392 30575 11456
rect 30639 11392 30655 11456
rect 30719 11392 30735 11456
rect 30799 11392 30805 11456
rect 30489 11391 30805 11392
rect 21173 11250 21239 11253
rect 22277 11250 22343 11253
rect 21173 11248 22343 11250
rect 21173 11192 21178 11248
rect 21234 11192 22282 11248
rect 22338 11192 22343 11248
rect 21173 11190 22343 11192
rect 21173 11187 21239 11190
rect 22277 11187 22343 11190
rect 21173 11114 21239 11117
rect 22921 11114 22987 11117
rect 21173 11112 22987 11114
rect 21173 11056 21178 11112
rect 21234 11056 22926 11112
rect 22982 11056 22987 11112
rect 21173 11054 22987 11056
rect 21173 11051 21239 11054
rect 22921 11051 22987 11054
rect 9386 10912 9702 10913
rect 9386 10848 9392 10912
rect 9456 10848 9472 10912
rect 9536 10848 9552 10912
rect 9616 10848 9632 10912
rect 9696 10848 9702 10912
rect 9386 10847 9702 10848
rect 17827 10912 18143 10913
rect 17827 10848 17833 10912
rect 17897 10848 17913 10912
rect 17977 10848 17993 10912
rect 18057 10848 18073 10912
rect 18137 10848 18143 10912
rect 17827 10847 18143 10848
rect 26268 10912 26584 10913
rect 26268 10848 26274 10912
rect 26338 10848 26354 10912
rect 26418 10848 26434 10912
rect 26498 10848 26514 10912
rect 26578 10848 26584 10912
rect 26268 10847 26584 10848
rect 34709 10912 35025 10913
rect 34709 10848 34715 10912
rect 34779 10848 34795 10912
rect 34859 10848 34875 10912
rect 34939 10848 34955 10912
rect 35019 10848 35025 10912
rect 34709 10847 35025 10848
rect 5166 10368 5482 10369
rect 5166 10304 5172 10368
rect 5236 10304 5252 10368
rect 5316 10304 5332 10368
rect 5396 10304 5412 10368
rect 5476 10304 5482 10368
rect 5166 10303 5482 10304
rect 13607 10368 13923 10369
rect 13607 10304 13613 10368
rect 13677 10304 13693 10368
rect 13757 10304 13773 10368
rect 13837 10304 13853 10368
rect 13917 10304 13923 10368
rect 13607 10303 13923 10304
rect 22048 10368 22364 10369
rect 22048 10304 22054 10368
rect 22118 10304 22134 10368
rect 22198 10304 22214 10368
rect 22278 10304 22294 10368
rect 22358 10304 22364 10368
rect 22048 10303 22364 10304
rect 30489 10368 30805 10369
rect 30489 10304 30495 10368
rect 30559 10304 30575 10368
rect 30639 10304 30655 10368
rect 30719 10304 30735 10368
rect 30799 10304 30805 10368
rect 30489 10303 30805 10304
rect 9386 9824 9702 9825
rect 9386 9760 9392 9824
rect 9456 9760 9472 9824
rect 9536 9760 9552 9824
rect 9616 9760 9632 9824
rect 9696 9760 9702 9824
rect 9386 9759 9702 9760
rect 17827 9824 18143 9825
rect 17827 9760 17833 9824
rect 17897 9760 17913 9824
rect 17977 9760 17993 9824
rect 18057 9760 18073 9824
rect 18137 9760 18143 9824
rect 17827 9759 18143 9760
rect 26268 9824 26584 9825
rect 26268 9760 26274 9824
rect 26338 9760 26354 9824
rect 26418 9760 26434 9824
rect 26498 9760 26514 9824
rect 26578 9760 26584 9824
rect 26268 9759 26584 9760
rect 34709 9824 35025 9825
rect 34709 9760 34715 9824
rect 34779 9760 34795 9824
rect 34859 9760 34875 9824
rect 34939 9760 34955 9824
rect 35019 9760 35025 9824
rect 34709 9759 35025 9760
rect 5166 9280 5482 9281
rect 5166 9216 5172 9280
rect 5236 9216 5252 9280
rect 5316 9216 5332 9280
rect 5396 9216 5412 9280
rect 5476 9216 5482 9280
rect 5166 9215 5482 9216
rect 13607 9280 13923 9281
rect 13607 9216 13613 9280
rect 13677 9216 13693 9280
rect 13757 9216 13773 9280
rect 13837 9216 13853 9280
rect 13917 9216 13923 9280
rect 13607 9215 13923 9216
rect 22048 9280 22364 9281
rect 22048 9216 22054 9280
rect 22118 9216 22134 9280
rect 22198 9216 22214 9280
rect 22278 9216 22294 9280
rect 22358 9216 22364 9280
rect 22048 9215 22364 9216
rect 30489 9280 30805 9281
rect 30489 9216 30495 9280
rect 30559 9216 30575 9280
rect 30639 9216 30655 9280
rect 30719 9216 30735 9280
rect 30799 9216 30805 9280
rect 30489 9215 30805 9216
rect 9386 8736 9702 8737
rect 9386 8672 9392 8736
rect 9456 8672 9472 8736
rect 9536 8672 9552 8736
rect 9616 8672 9632 8736
rect 9696 8672 9702 8736
rect 9386 8671 9702 8672
rect 17827 8736 18143 8737
rect 17827 8672 17833 8736
rect 17897 8672 17913 8736
rect 17977 8672 17993 8736
rect 18057 8672 18073 8736
rect 18137 8672 18143 8736
rect 17827 8671 18143 8672
rect 26268 8736 26584 8737
rect 26268 8672 26274 8736
rect 26338 8672 26354 8736
rect 26418 8672 26434 8736
rect 26498 8672 26514 8736
rect 26578 8672 26584 8736
rect 26268 8671 26584 8672
rect 34709 8736 35025 8737
rect 34709 8672 34715 8736
rect 34779 8672 34795 8736
rect 34859 8672 34875 8736
rect 34939 8672 34955 8736
rect 35019 8672 35025 8736
rect 34709 8671 35025 8672
rect 5166 8192 5482 8193
rect 5166 8128 5172 8192
rect 5236 8128 5252 8192
rect 5316 8128 5332 8192
rect 5396 8128 5412 8192
rect 5476 8128 5482 8192
rect 5166 8127 5482 8128
rect 13607 8192 13923 8193
rect 13607 8128 13613 8192
rect 13677 8128 13693 8192
rect 13757 8128 13773 8192
rect 13837 8128 13853 8192
rect 13917 8128 13923 8192
rect 13607 8127 13923 8128
rect 22048 8192 22364 8193
rect 22048 8128 22054 8192
rect 22118 8128 22134 8192
rect 22198 8128 22214 8192
rect 22278 8128 22294 8192
rect 22358 8128 22364 8192
rect 22048 8127 22364 8128
rect 30489 8192 30805 8193
rect 30489 8128 30495 8192
rect 30559 8128 30575 8192
rect 30639 8128 30655 8192
rect 30719 8128 30735 8192
rect 30799 8128 30805 8192
rect 30489 8127 30805 8128
rect 9386 7648 9702 7649
rect 9386 7584 9392 7648
rect 9456 7584 9472 7648
rect 9536 7584 9552 7648
rect 9616 7584 9632 7648
rect 9696 7584 9702 7648
rect 9386 7583 9702 7584
rect 17827 7648 18143 7649
rect 17827 7584 17833 7648
rect 17897 7584 17913 7648
rect 17977 7584 17993 7648
rect 18057 7584 18073 7648
rect 18137 7584 18143 7648
rect 17827 7583 18143 7584
rect 26268 7648 26584 7649
rect 26268 7584 26274 7648
rect 26338 7584 26354 7648
rect 26418 7584 26434 7648
rect 26498 7584 26514 7648
rect 26578 7584 26584 7648
rect 26268 7583 26584 7584
rect 34709 7648 35025 7649
rect 34709 7584 34715 7648
rect 34779 7584 34795 7648
rect 34859 7584 34875 7648
rect 34939 7584 34955 7648
rect 35019 7584 35025 7648
rect 34709 7583 35025 7584
rect 5166 7104 5482 7105
rect 5166 7040 5172 7104
rect 5236 7040 5252 7104
rect 5316 7040 5332 7104
rect 5396 7040 5412 7104
rect 5476 7040 5482 7104
rect 5166 7039 5482 7040
rect 13607 7104 13923 7105
rect 13607 7040 13613 7104
rect 13677 7040 13693 7104
rect 13757 7040 13773 7104
rect 13837 7040 13853 7104
rect 13917 7040 13923 7104
rect 13607 7039 13923 7040
rect 22048 7104 22364 7105
rect 22048 7040 22054 7104
rect 22118 7040 22134 7104
rect 22198 7040 22214 7104
rect 22278 7040 22294 7104
rect 22358 7040 22364 7104
rect 22048 7039 22364 7040
rect 30489 7104 30805 7105
rect 30489 7040 30495 7104
rect 30559 7040 30575 7104
rect 30639 7040 30655 7104
rect 30719 7040 30735 7104
rect 30799 7040 30805 7104
rect 30489 7039 30805 7040
rect 9386 6560 9702 6561
rect 9386 6496 9392 6560
rect 9456 6496 9472 6560
rect 9536 6496 9552 6560
rect 9616 6496 9632 6560
rect 9696 6496 9702 6560
rect 9386 6495 9702 6496
rect 17827 6560 18143 6561
rect 17827 6496 17833 6560
rect 17897 6496 17913 6560
rect 17977 6496 17993 6560
rect 18057 6496 18073 6560
rect 18137 6496 18143 6560
rect 17827 6495 18143 6496
rect 26268 6560 26584 6561
rect 26268 6496 26274 6560
rect 26338 6496 26354 6560
rect 26418 6496 26434 6560
rect 26498 6496 26514 6560
rect 26578 6496 26584 6560
rect 26268 6495 26584 6496
rect 34709 6560 35025 6561
rect 34709 6496 34715 6560
rect 34779 6496 34795 6560
rect 34859 6496 34875 6560
rect 34939 6496 34955 6560
rect 35019 6496 35025 6560
rect 34709 6495 35025 6496
rect 5166 6016 5482 6017
rect 5166 5952 5172 6016
rect 5236 5952 5252 6016
rect 5316 5952 5332 6016
rect 5396 5952 5412 6016
rect 5476 5952 5482 6016
rect 5166 5951 5482 5952
rect 13607 6016 13923 6017
rect 13607 5952 13613 6016
rect 13677 5952 13693 6016
rect 13757 5952 13773 6016
rect 13837 5952 13853 6016
rect 13917 5952 13923 6016
rect 13607 5951 13923 5952
rect 22048 6016 22364 6017
rect 22048 5952 22054 6016
rect 22118 5952 22134 6016
rect 22198 5952 22214 6016
rect 22278 5952 22294 6016
rect 22358 5952 22364 6016
rect 22048 5951 22364 5952
rect 30489 6016 30805 6017
rect 30489 5952 30495 6016
rect 30559 5952 30575 6016
rect 30639 5952 30655 6016
rect 30719 5952 30735 6016
rect 30799 5952 30805 6016
rect 30489 5951 30805 5952
rect 9386 5472 9702 5473
rect 9386 5408 9392 5472
rect 9456 5408 9472 5472
rect 9536 5408 9552 5472
rect 9616 5408 9632 5472
rect 9696 5408 9702 5472
rect 9386 5407 9702 5408
rect 17827 5472 18143 5473
rect 17827 5408 17833 5472
rect 17897 5408 17913 5472
rect 17977 5408 17993 5472
rect 18057 5408 18073 5472
rect 18137 5408 18143 5472
rect 17827 5407 18143 5408
rect 26268 5472 26584 5473
rect 26268 5408 26274 5472
rect 26338 5408 26354 5472
rect 26418 5408 26434 5472
rect 26498 5408 26514 5472
rect 26578 5408 26584 5472
rect 26268 5407 26584 5408
rect 34709 5472 35025 5473
rect 34709 5408 34715 5472
rect 34779 5408 34795 5472
rect 34859 5408 34875 5472
rect 34939 5408 34955 5472
rect 35019 5408 35025 5472
rect 34709 5407 35025 5408
rect 5166 4928 5482 4929
rect 5166 4864 5172 4928
rect 5236 4864 5252 4928
rect 5316 4864 5332 4928
rect 5396 4864 5412 4928
rect 5476 4864 5482 4928
rect 5166 4863 5482 4864
rect 13607 4928 13923 4929
rect 13607 4864 13613 4928
rect 13677 4864 13693 4928
rect 13757 4864 13773 4928
rect 13837 4864 13853 4928
rect 13917 4864 13923 4928
rect 13607 4863 13923 4864
rect 22048 4928 22364 4929
rect 22048 4864 22054 4928
rect 22118 4864 22134 4928
rect 22198 4864 22214 4928
rect 22278 4864 22294 4928
rect 22358 4864 22364 4928
rect 22048 4863 22364 4864
rect 30489 4928 30805 4929
rect 30489 4864 30495 4928
rect 30559 4864 30575 4928
rect 30639 4864 30655 4928
rect 30719 4864 30735 4928
rect 30799 4864 30805 4928
rect 30489 4863 30805 4864
rect 9386 4384 9702 4385
rect 9386 4320 9392 4384
rect 9456 4320 9472 4384
rect 9536 4320 9552 4384
rect 9616 4320 9632 4384
rect 9696 4320 9702 4384
rect 9386 4319 9702 4320
rect 17827 4384 18143 4385
rect 17827 4320 17833 4384
rect 17897 4320 17913 4384
rect 17977 4320 17993 4384
rect 18057 4320 18073 4384
rect 18137 4320 18143 4384
rect 17827 4319 18143 4320
rect 26268 4384 26584 4385
rect 26268 4320 26274 4384
rect 26338 4320 26354 4384
rect 26418 4320 26434 4384
rect 26498 4320 26514 4384
rect 26578 4320 26584 4384
rect 26268 4319 26584 4320
rect 34709 4384 35025 4385
rect 34709 4320 34715 4384
rect 34779 4320 34795 4384
rect 34859 4320 34875 4384
rect 34939 4320 34955 4384
rect 35019 4320 35025 4384
rect 34709 4319 35025 4320
rect 5166 3840 5482 3841
rect 5166 3776 5172 3840
rect 5236 3776 5252 3840
rect 5316 3776 5332 3840
rect 5396 3776 5412 3840
rect 5476 3776 5482 3840
rect 5166 3775 5482 3776
rect 13607 3840 13923 3841
rect 13607 3776 13613 3840
rect 13677 3776 13693 3840
rect 13757 3776 13773 3840
rect 13837 3776 13853 3840
rect 13917 3776 13923 3840
rect 13607 3775 13923 3776
rect 22048 3840 22364 3841
rect 22048 3776 22054 3840
rect 22118 3776 22134 3840
rect 22198 3776 22214 3840
rect 22278 3776 22294 3840
rect 22358 3776 22364 3840
rect 22048 3775 22364 3776
rect 30489 3840 30805 3841
rect 30489 3776 30495 3840
rect 30559 3776 30575 3840
rect 30639 3776 30655 3840
rect 30719 3776 30735 3840
rect 30799 3776 30805 3840
rect 30489 3775 30805 3776
rect 9386 3296 9702 3297
rect 9386 3232 9392 3296
rect 9456 3232 9472 3296
rect 9536 3232 9552 3296
rect 9616 3232 9632 3296
rect 9696 3232 9702 3296
rect 9386 3231 9702 3232
rect 17827 3296 18143 3297
rect 17827 3232 17833 3296
rect 17897 3232 17913 3296
rect 17977 3232 17993 3296
rect 18057 3232 18073 3296
rect 18137 3232 18143 3296
rect 17827 3231 18143 3232
rect 26268 3296 26584 3297
rect 26268 3232 26274 3296
rect 26338 3232 26354 3296
rect 26418 3232 26434 3296
rect 26498 3232 26514 3296
rect 26578 3232 26584 3296
rect 26268 3231 26584 3232
rect 34709 3296 35025 3297
rect 34709 3232 34715 3296
rect 34779 3232 34795 3296
rect 34859 3232 34875 3296
rect 34939 3232 34955 3296
rect 35019 3232 35025 3296
rect 34709 3231 35025 3232
rect 5166 2752 5482 2753
rect 5166 2688 5172 2752
rect 5236 2688 5252 2752
rect 5316 2688 5332 2752
rect 5396 2688 5412 2752
rect 5476 2688 5482 2752
rect 5166 2687 5482 2688
rect 13607 2752 13923 2753
rect 13607 2688 13613 2752
rect 13677 2688 13693 2752
rect 13757 2688 13773 2752
rect 13837 2688 13853 2752
rect 13917 2688 13923 2752
rect 13607 2687 13923 2688
rect 22048 2752 22364 2753
rect 22048 2688 22054 2752
rect 22118 2688 22134 2752
rect 22198 2688 22214 2752
rect 22278 2688 22294 2752
rect 22358 2688 22364 2752
rect 22048 2687 22364 2688
rect 30489 2752 30805 2753
rect 30489 2688 30495 2752
rect 30559 2688 30575 2752
rect 30639 2688 30655 2752
rect 30719 2688 30735 2752
rect 30799 2688 30805 2752
rect 30489 2687 30805 2688
rect 9386 2208 9702 2209
rect 9386 2144 9392 2208
rect 9456 2144 9472 2208
rect 9536 2144 9552 2208
rect 9616 2144 9632 2208
rect 9696 2144 9702 2208
rect 9386 2143 9702 2144
rect 17827 2208 18143 2209
rect 17827 2144 17833 2208
rect 17897 2144 17913 2208
rect 17977 2144 17993 2208
rect 18057 2144 18073 2208
rect 18137 2144 18143 2208
rect 17827 2143 18143 2144
rect 26268 2208 26584 2209
rect 26268 2144 26274 2208
rect 26338 2144 26354 2208
rect 26418 2144 26434 2208
rect 26498 2144 26514 2208
rect 26578 2144 26584 2208
rect 26268 2143 26584 2144
rect 34709 2208 35025 2209
rect 34709 2144 34715 2208
rect 34779 2144 34795 2208
rect 34859 2144 34875 2208
rect 34939 2144 34955 2208
rect 35019 2144 35025 2208
rect 34709 2143 35025 2144
<< via3 >>
rect 9392 33756 9456 33760
rect 9392 33700 9396 33756
rect 9396 33700 9452 33756
rect 9452 33700 9456 33756
rect 9392 33696 9456 33700
rect 9472 33756 9536 33760
rect 9472 33700 9476 33756
rect 9476 33700 9532 33756
rect 9532 33700 9536 33756
rect 9472 33696 9536 33700
rect 9552 33756 9616 33760
rect 9552 33700 9556 33756
rect 9556 33700 9612 33756
rect 9612 33700 9616 33756
rect 9552 33696 9616 33700
rect 9632 33756 9696 33760
rect 9632 33700 9636 33756
rect 9636 33700 9692 33756
rect 9692 33700 9696 33756
rect 9632 33696 9696 33700
rect 17833 33756 17897 33760
rect 17833 33700 17837 33756
rect 17837 33700 17893 33756
rect 17893 33700 17897 33756
rect 17833 33696 17897 33700
rect 17913 33756 17977 33760
rect 17913 33700 17917 33756
rect 17917 33700 17973 33756
rect 17973 33700 17977 33756
rect 17913 33696 17977 33700
rect 17993 33756 18057 33760
rect 17993 33700 17997 33756
rect 17997 33700 18053 33756
rect 18053 33700 18057 33756
rect 17993 33696 18057 33700
rect 18073 33756 18137 33760
rect 18073 33700 18077 33756
rect 18077 33700 18133 33756
rect 18133 33700 18137 33756
rect 18073 33696 18137 33700
rect 26274 33756 26338 33760
rect 26274 33700 26278 33756
rect 26278 33700 26334 33756
rect 26334 33700 26338 33756
rect 26274 33696 26338 33700
rect 26354 33756 26418 33760
rect 26354 33700 26358 33756
rect 26358 33700 26414 33756
rect 26414 33700 26418 33756
rect 26354 33696 26418 33700
rect 26434 33756 26498 33760
rect 26434 33700 26438 33756
rect 26438 33700 26494 33756
rect 26494 33700 26498 33756
rect 26434 33696 26498 33700
rect 26514 33756 26578 33760
rect 26514 33700 26518 33756
rect 26518 33700 26574 33756
rect 26574 33700 26578 33756
rect 26514 33696 26578 33700
rect 34715 33756 34779 33760
rect 34715 33700 34719 33756
rect 34719 33700 34775 33756
rect 34775 33700 34779 33756
rect 34715 33696 34779 33700
rect 34795 33756 34859 33760
rect 34795 33700 34799 33756
rect 34799 33700 34855 33756
rect 34855 33700 34859 33756
rect 34795 33696 34859 33700
rect 34875 33756 34939 33760
rect 34875 33700 34879 33756
rect 34879 33700 34935 33756
rect 34935 33700 34939 33756
rect 34875 33696 34939 33700
rect 34955 33756 35019 33760
rect 34955 33700 34959 33756
rect 34959 33700 35015 33756
rect 35015 33700 35019 33756
rect 34955 33696 35019 33700
rect 5172 33212 5236 33216
rect 5172 33156 5176 33212
rect 5176 33156 5232 33212
rect 5232 33156 5236 33212
rect 5172 33152 5236 33156
rect 5252 33212 5316 33216
rect 5252 33156 5256 33212
rect 5256 33156 5312 33212
rect 5312 33156 5316 33212
rect 5252 33152 5316 33156
rect 5332 33212 5396 33216
rect 5332 33156 5336 33212
rect 5336 33156 5392 33212
rect 5392 33156 5396 33212
rect 5332 33152 5396 33156
rect 5412 33212 5476 33216
rect 5412 33156 5416 33212
rect 5416 33156 5472 33212
rect 5472 33156 5476 33212
rect 5412 33152 5476 33156
rect 13613 33212 13677 33216
rect 13613 33156 13617 33212
rect 13617 33156 13673 33212
rect 13673 33156 13677 33212
rect 13613 33152 13677 33156
rect 13693 33212 13757 33216
rect 13693 33156 13697 33212
rect 13697 33156 13753 33212
rect 13753 33156 13757 33212
rect 13693 33152 13757 33156
rect 13773 33212 13837 33216
rect 13773 33156 13777 33212
rect 13777 33156 13833 33212
rect 13833 33156 13837 33212
rect 13773 33152 13837 33156
rect 13853 33212 13917 33216
rect 13853 33156 13857 33212
rect 13857 33156 13913 33212
rect 13913 33156 13917 33212
rect 13853 33152 13917 33156
rect 22054 33212 22118 33216
rect 22054 33156 22058 33212
rect 22058 33156 22114 33212
rect 22114 33156 22118 33212
rect 22054 33152 22118 33156
rect 22134 33212 22198 33216
rect 22134 33156 22138 33212
rect 22138 33156 22194 33212
rect 22194 33156 22198 33212
rect 22134 33152 22198 33156
rect 22214 33212 22278 33216
rect 22214 33156 22218 33212
rect 22218 33156 22274 33212
rect 22274 33156 22278 33212
rect 22214 33152 22278 33156
rect 22294 33212 22358 33216
rect 22294 33156 22298 33212
rect 22298 33156 22354 33212
rect 22354 33156 22358 33212
rect 22294 33152 22358 33156
rect 30495 33212 30559 33216
rect 30495 33156 30499 33212
rect 30499 33156 30555 33212
rect 30555 33156 30559 33212
rect 30495 33152 30559 33156
rect 30575 33212 30639 33216
rect 30575 33156 30579 33212
rect 30579 33156 30635 33212
rect 30635 33156 30639 33212
rect 30575 33152 30639 33156
rect 30655 33212 30719 33216
rect 30655 33156 30659 33212
rect 30659 33156 30715 33212
rect 30715 33156 30719 33212
rect 30655 33152 30719 33156
rect 30735 33212 30799 33216
rect 30735 33156 30739 33212
rect 30739 33156 30795 33212
rect 30795 33156 30799 33212
rect 30735 33152 30799 33156
rect 9392 32668 9456 32672
rect 9392 32612 9396 32668
rect 9396 32612 9452 32668
rect 9452 32612 9456 32668
rect 9392 32608 9456 32612
rect 9472 32668 9536 32672
rect 9472 32612 9476 32668
rect 9476 32612 9532 32668
rect 9532 32612 9536 32668
rect 9472 32608 9536 32612
rect 9552 32668 9616 32672
rect 9552 32612 9556 32668
rect 9556 32612 9612 32668
rect 9612 32612 9616 32668
rect 9552 32608 9616 32612
rect 9632 32668 9696 32672
rect 9632 32612 9636 32668
rect 9636 32612 9692 32668
rect 9692 32612 9696 32668
rect 9632 32608 9696 32612
rect 17833 32668 17897 32672
rect 17833 32612 17837 32668
rect 17837 32612 17893 32668
rect 17893 32612 17897 32668
rect 17833 32608 17897 32612
rect 17913 32668 17977 32672
rect 17913 32612 17917 32668
rect 17917 32612 17973 32668
rect 17973 32612 17977 32668
rect 17913 32608 17977 32612
rect 17993 32668 18057 32672
rect 17993 32612 17997 32668
rect 17997 32612 18053 32668
rect 18053 32612 18057 32668
rect 17993 32608 18057 32612
rect 18073 32668 18137 32672
rect 18073 32612 18077 32668
rect 18077 32612 18133 32668
rect 18133 32612 18137 32668
rect 18073 32608 18137 32612
rect 26274 32668 26338 32672
rect 26274 32612 26278 32668
rect 26278 32612 26334 32668
rect 26334 32612 26338 32668
rect 26274 32608 26338 32612
rect 26354 32668 26418 32672
rect 26354 32612 26358 32668
rect 26358 32612 26414 32668
rect 26414 32612 26418 32668
rect 26354 32608 26418 32612
rect 26434 32668 26498 32672
rect 26434 32612 26438 32668
rect 26438 32612 26494 32668
rect 26494 32612 26498 32668
rect 26434 32608 26498 32612
rect 26514 32668 26578 32672
rect 26514 32612 26518 32668
rect 26518 32612 26574 32668
rect 26574 32612 26578 32668
rect 26514 32608 26578 32612
rect 34715 32668 34779 32672
rect 34715 32612 34719 32668
rect 34719 32612 34775 32668
rect 34775 32612 34779 32668
rect 34715 32608 34779 32612
rect 34795 32668 34859 32672
rect 34795 32612 34799 32668
rect 34799 32612 34855 32668
rect 34855 32612 34859 32668
rect 34795 32608 34859 32612
rect 34875 32668 34939 32672
rect 34875 32612 34879 32668
rect 34879 32612 34935 32668
rect 34935 32612 34939 32668
rect 34875 32608 34939 32612
rect 34955 32668 35019 32672
rect 34955 32612 34959 32668
rect 34959 32612 35015 32668
rect 35015 32612 35019 32668
rect 34955 32608 35019 32612
rect 5172 32124 5236 32128
rect 5172 32068 5176 32124
rect 5176 32068 5232 32124
rect 5232 32068 5236 32124
rect 5172 32064 5236 32068
rect 5252 32124 5316 32128
rect 5252 32068 5256 32124
rect 5256 32068 5312 32124
rect 5312 32068 5316 32124
rect 5252 32064 5316 32068
rect 5332 32124 5396 32128
rect 5332 32068 5336 32124
rect 5336 32068 5392 32124
rect 5392 32068 5396 32124
rect 5332 32064 5396 32068
rect 5412 32124 5476 32128
rect 5412 32068 5416 32124
rect 5416 32068 5472 32124
rect 5472 32068 5476 32124
rect 5412 32064 5476 32068
rect 13613 32124 13677 32128
rect 13613 32068 13617 32124
rect 13617 32068 13673 32124
rect 13673 32068 13677 32124
rect 13613 32064 13677 32068
rect 13693 32124 13757 32128
rect 13693 32068 13697 32124
rect 13697 32068 13753 32124
rect 13753 32068 13757 32124
rect 13693 32064 13757 32068
rect 13773 32124 13837 32128
rect 13773 32068 13777 32124
rect 13777 32068 13833 32124
rect 13833 32068 13837 32124
rect 13773 32064 13837 32068
rect 13853 32124 13917 32128
rect 13853 32068 13857 32124
rect 13857 32068 13913 32124
rect 13913 32068 13917 32124
rect 13853 32064 13917 32068
rect 22054 32124 22118 32128
rect 22054 32068 22058 32124
rect 22058 32068 22114 32124
rect 22114 32068 22118 32124
rect 22054 32064 22118 32068
rect 22134 32124 22198 32128
rect 22134 32068 22138 32124
rect 22138 32068 22194 32124
rect 22194 32068 22198 32124
rect 22134 32064 22198 32068
rect 22214 32124 22278 32128
rect 22214 32068 22218 32124
rect 22218 32068 22274 32124
rect 22274 32068 22278 32124
rect 22214 32064 22278 32068
rect 22294 32124 22358 32128
rect 22294 32068 22298 32124
rect 22298 32068 22354 32124
rect 22354 32068 22358 32124
rect 22294 32064 22358 32068
rect 30495 32124 30559 32128
rect 30495 32068 30499 32124
rect 30499 32068 30555 32124
rect 30555 32068 30559 32124
rect 30495 32064 30559 32068
rect 30575 32124 30639 32128
rect 30575 32068 30579 32124
rect 30579 32068 30635 32124
rect 30635 32068 30639 32124
rect 30575 32064 30639 32068
rect 30655 32124 30719 32128
rect 30655 32068 30659 32124
rect 30659 32068 30715 32124
rect 30715 32068 30719 32124
rect 30655 32064 30719 32068
rect 30735 32124 30799 32128
rect 30735 32068 30739 32124
rect 30739 32068 30795 32124
rect 30795 32068 30799 32124
rect 30735 32064 30799 32068
rect 9392 31580 9456 31584
rect 9392 31524 9396 31580
rect 9396 31524 9452 31580
rect 9452 31524 9456 31580
rect 9392 31520 9456 31524
rect 9472 31580 9536 31584
rect 9472 31524 9476 31580
rect 9476 31524 9532 31580
rect 9532 31524 9536 31580
rect 9472 31520 9536 31524
rect 9552 31580 9616 31584
rect 9552 31524 9556 31580
rect 9556 31524 9612 31580
rect 9612 31524 9616 31580
rect 9552 31520 9616 31524
rect 9632 31580 9696 31584
rect 9632 31524 9636 31580
rect 9636 31524 9692 31580
rect 9692 31524 9696 31580
rect 9632 31520 9696 31524
rect 17833 31580 17897 31584
rect 17833 31524 17837 31580
rect 17837 31524 17893 31580
rect 17893 31524 17897 31580
rect 17833 31520 17897 31524
rect 17913 31580 17977 31584
rect 17913 31524 17917 31580
rect 17917 31524 17973 31580
rect 17973 31524 17977 31580
rect 17913 31520 17977 31524
rect 17993 31580 18057 31584
rect 17993 31524 17997 31580
rect 17997 31524 18053 31580
rect 18053 31524 18057 31580
rect 17993 31520 18057 31524
rect 18073 31580 18137 31584
rect 18073 31524 18077 31580
rect 18077 31524 18133 31580
rect 18133 31524 18137 31580
rect 18073 31520 18137 31524
rect 26274 31580 26338 31584
rect 26274 31524 26278 31580
rect 26278 31524 26334 31580
rect 26334 31524 26338 31580
rect 26274 31520 26338 31524
rect 26354 31580 26418 31584
rect 26354 31524 26358 31580
rect 26358 31524 26414 31580
rect 26414 31524 26418 31580
rect 26354 31520 26418 31524
rect 26434 31580 26498 31584
rect 26434 31524 26438 31580
rect 26438 31524 26494 31580
rect 26494 31524 26498 31580
rect 26434 31520 26498 31524
rect 26514 31580 26578 31584
rect 26514 31524 26518 31580
rect 26518 31524 26574 31580
rect 26574 31524 26578 31580
rect 26514 31520 26578 31524
rect 34715 31580 34779 31584
rect 34715 31524 34719 31580
rect 34719 31524 34775 31580
rect 34775 31524 34779 31580
rect 34715 31520 34779 31524
rect 34795 31580 34859 31584
rect 34795 31524 34799 31580
rect 34799 31524 34855 31580
rect 34855 31524 34859 31580
rect 34795 31520 34859 31524
rect 34875 31580 34939 31584
rect 34875 31524 34879 31580
rect 34879 31524 34935 31580
rect 34935 31524 34939 31580
rect 34875 31520 34939 31524
rect 34955 31580 35019 31584
rect 34955 31524 34959 31580
rect 34959 31524 35015 31580
rect 35015 31524 35019 31580
rect 34955 31520 35019 31524
rect 5172 31036 5236 31040
rect 5172 30980 5176 31036
rect 5176 30980 5232 31036
rect 5232 30980 5236 31036
rect 5172 30976 5236 30980
rect 5252 31036 5316 31040
rect 5252 30980 5256 31036
rect 5256 30980 5312 31036
rect 5312 30980 5316 31036
rect 5252 30976 5316 30980
rect 5332 31036 5396 31040
rect 5332 30980 5336 31036
rect 5336 30980 5392 31036
rect 5392 30980 5396 31036
rect 5332 30976 5396 30980
rect 5412 31036 5476 31040
rect 5412 30980 5416 31036
rect 5416 30980 5472 31036
rect 5472 30980 5476 31036
rect 5412 30976 5476 30980
rect 13613 31036 13677 31040
rect 13613 30980 13617 31036
rect 13617 30980 13673 31036
rect 13673 30980 13677 31036
rect 13613 30976 13677 30980
rect 13693 31036 13757 31040
rect 13693 30980 13697 31036
rect 13697 30980 13753 31036
rect 13753 30980 13757 31036
rect 13693 30976 13757 30980
rect 13773 31036 13837 31040
rect 13773 30980 13777 31036
rect 13777 30980 13833 31036
rect 13833 30980 13837 31036
rect 13773 30976 13837 30980
rect 13853 31036 13917 31040
rect 13853 30980 13857 31036
rect 13857 30980 13913 31036
rect 13913 30980 13917 31036
rect 13853 30976 13917 30980
rect 22054 31036 22118 31040
rect 22054 30980 22058 31036
rect 22058 30980 22114 31036
rect 22114 30980 22118 31036
rect 22054 30976 22118 30980
rect 22134 31036 22198 31040
rect 22134 30980 22138 31036
rect 22138 30980 22194 31036
rect 22194 30980 22198 31036
rect 22134 30976 22198 30980
rect 22214 31036 22278 31040
rect 22214 30980 22218 31036
rect 22218 30980 22274 31036
rect 22274 30980 22278 31036
rect 22214 30976 22278 30980
rect 22294 31036 22358 31040
rect 22294 30980 22298 31036
rect 22298 30980 22354 31036
rect 22354 30980 22358 31036
rect 22294 30976 22358 30980
rect 30495 31036 30559 31040
rect 30495 30980 30499 31036
rect 30499 30980 30555 31036
rect 30555 30980 30559 31036
rect 30495 30976 30559 30980
rect 30575 31036 30639 31040
rect 30575 30980 30579 31036
rect 30579 30980 30635 31036
rect 30635 30980 30639 31036
rect 30575 30976 30639 30980
rect 30655 31036 30719 31040
rect 30655 30980 30659 31036
rect 30659 30980 30715 31036
rect 30715 30980 30719 31036
rect 30655 30976 30719 30980
rect 30735 31036 30799 31040
rect 30735 30980 30739 31036
rect 30739 30980 30795 31036
rect 30795 30980 30799 31036
rect 30735 30976 30799 30980
rect 24900 30832 24964 30836
rect 24900 30776 24950 30832
rect 24950 30776 24964 30832
rect 24900 30772 24964 30776
rect 9392 30492 9456 30496
rect 9392 30436 9396 30492
rect 9396 30436 9452 30492
rect 9452 30436 9456 30492
rect 9392 30432 9456 30436
rect 9472 30492 9536 30496
rect 9472 30436 9476 30492
rect 9476 30436 9532 30492
rect 9532 30436 9536 30492
rect 9472 30432 9536 30436
rect 9552 30492 9616 30496
rect 9552 30436 9556 30492
rect 9556 30436 9612 30492
rect 9612 30436 9616 30492
rect 9552 30432 9616 30436
rect 9632 30492 9696 30496
rect 9632 30436 9636 30492
rect 9636 30436 9692 30492
rect 9692 30436 9696 30492
rect 9632 30432 9696 30436
rect 17833 30492 17897 30496
rect 17833 30436 17837 30492
rect 17837 30436 17893 30492
rect 17893 30436 17897 30492
rect 17833 30432 17897 30436
rect 17913 30492 17977 30496
rect 17913 30436 17917 30492
rect 17917 30436 17973 30492
rect 17973 30436 17977 30492
rect 17913 30432 17977 30436
rect 17993 30492 18057 30496
rect 17993 30436 17997 30492
rect 17997 30436 18053 30492
rect 18053 30436 18057 30492
rect 17993 30432 18057 30436
rect 18073 30492 18137 30496
rect 18073 30436 18077 30492
rect 18077 30436 18133 30492
rect 18133 30436 18137 30492
rect 18073 30432 18137 30436
rect 26274 30492 26338 30496
rect 26274 30436 26278 30492
rect 26278 30436 26334 30492
rect 26334 30436 26338 30492
rect 26274 30432 26338 30436
rect 26354 30492 26418 30496
rect 26354 30436 26358 30492
rect 26358 30436 26414 30492
rect 26414 30436 26418 30492
rect 26354 30432 26418 30436
rect 26434 30492 26498 30496
rect 26434 30436 26438 30492
rect 26438 30436 26494 30492
rect 26494 30436 26498 30492
rect 26434 30432 26498 30436
rect 26514 30492 26578 30496
rect 26514 30436 26518 30492
rect 26518 30436 26574 30492
rect 26574 30436 26578 30492
rect 26514 30432 26578 30436
rect 34715 30492 34779 30496
rect 34715 30436 34719 30492
rect 34719 30436 34775 30492
rect 34775 30436 34779 30492
rect 34715 30432 34779 30436
rect 34795 30492 34859 30496
rect 34795 30436 34799 30492
rect 34799 30436 34855 30492
rect 34855 30436 34859 30492
rect 34795 30432 34859 30436
rect 34875 30492 34939 30496
rect 34875 30436 34879 30492
rect 34879 30436 34935 30492
rect 34935 30436 34939 30492
rect 34875 30432 34939 30436
rect 34955 30492 35019 30496
rect 34955 30436 34959 30492
rect 34959 30436 35015 30492
rect 35015 30436 35019 30492
rect 34955 30432 35019 30436
rect 5172 29948 5236 29952
rect 5172 29892 5176 29948
rect 5176 29892 5232 29948
rect 5232 29892 5236 29948
rect 5172 29888 5236 29892
rect 5252 29948 5316 29952
rect 5252 29892 5256 29948
rect 5256 29892 5312 29948
rect 5312 29892 5316 29948
rect 5252 29888 5316 29892
rect 5332 29948 5396 29952
rect 5332 29892 5336 29948
rect 5336 29892 5392 29948
rect 5392 29892 5396 29948
rect 5332 29888 5396 29892
rect 5412 29948 5476 29952
rect 5412 29892 5416 29948
rect 5416 29892 5472 29948
rect 5472 29892 5476 29948
rect 5412 29888 5476 29892
rect 13613 29948 13677 29952
rect 13613 29892 13617 29948
rect 13617 29892 13673 29948
rect 13673 29892 13677 29948
rect 13613 29888 13677 29892
rect 13693 29948 13757 29952
rect 13693 29892 13697 29948
rect 13697 29892 13753 29948
rect 13753 29892 13757 29948
rect 13693 29888 13757 29892
rect 13773 29948 13837 29952
rect 13773 29892 13777 29948
rect 13777 29892 13833 29948
rect 13833 29892 13837 29948
rect 13773 29888 13837 29892
rect 13853 29948 13917 29952
rect 13853 29892 13857 29948
rect 13857 29892 13913 29948
rect 13913 29892 13917 29948
rect 13853 29888 13917 29892
rect 22054 29948 22118 29952
rect 22054 29892 22058 29948
rect 22058 29892 22114 29948
rect 22114 29892 22118 29948
rect 22054 29888 22118 29892
rect 22134 29948 22198 29952
rect 22134 29892 22138 29948
rect 22138 29892 22194 29948
rect 22194 29892 22198 29948
rect 22134 29888 22198 29892
rect 22214 29948 22278 29952
rect 22214 29892 22218 29948
rect 22218 29892 22274 29948
rect 22274 29892 22278 29948
rect 22214 29888 22278 29892
rect 22294 29948 22358 29952
rect 22294 29892 22298 29948
rect 22298 29892 22354 29948
rect 22354 29892 22358 29948
rect 22294 29888 22358 29892
rect 30495 29948 30559 29952
rect 30495 29892 30499 29948
rect 30499 29892 30555 29948
rect 30555 29892 30559 29948
rect 30495 29888 30559 29892
rect 30575 29948 30639 29952
rect 30575 29892 30579 29948
rect 30579 29892 30635 29948
rect 30635 29892 30639 29948
rect 30575 29888 30639 29892
rect 30655 29948 30719 29952
rect 30655 29892 30659 29948
rect 30659 29892 30715 29948
rect 30715 29892 30719 29948
rect 30655 29888 30719 29892
rect 30735 29948 30799 29952
rect 30735 29892 30739 29948
rect 30739 29892 30795 29948
rect 30795 29892 30799 29948
rect 30735 29888 30799 29892
rect 9392 29404 9456 29408
rect 9392 29348 9396 29404
rect 9396 29348 9452 29404
rect 9452 29348 9456 29404
rect 9392 29344 9456 29348
rect 9472 29404 9536 29408
rect 9472 29348 9476 29404
rect 9476 29348 9532 29404
rect 9532 29348 9536 29404
rect 9472 29344 9536 29348
rect 9552 29404 9616 29408
rect 9552 29348 9556 29404
rect 9556 29348 9612 29404
rect 9612 29348 9616 29404
rect 9552 29344 9616 29348
rect 9632 29404 9696 29408
rect 9632 29348 9636 29404
rect 9636 29348 9692 29404
rect 9692 29348 9696 29404
rect 9632 29344 9696 29348
rect 17833 29404 17897 29408
rect 17833 29348 17837 29404
rect 17837 29348 17893 29404
rect 17893 29348 17897 29404
rect 17833 29344 17897 29348
rect 17913 29404 17977 29408
rect 17913 29348 17917 29404
rect 17917 29348 17973 29404
rect 17973 29348 17977 29404
rect 17913 29344 17977 29348
rect 17993 29404 18057 29408
rect 17993 29348 17997 29404
rect 17997 29348 18053 29404
rect 18053 29348 18057 29404
rect 17993 29344 18057 29348
rect 18073 29404 18137 29408
rect 18073 29348 18077 29404
rect 18077 29348 18133 29404
rect 18133 29348 18137 29404
rect 18073 29344 18137 29348
rect 26274 29404 26338 29408
rect 26274 29348 26278 29404
rect 26278 29348 26334 29404
rect 26334 29348 26338 29404
rect 26274 29344 26338 29348
rect 26354 29404 26418 29408
rect 26354 29348 26358 29404
rect 26358 29348 26414 29404
rect 26414 29348 26418 29404
rect 26354 29344 26418 29348
rect 26434 29404 26498 29408
rect 26434 29348 26438 29404
rect 26438 29348 26494 29404
rect 26494 29348 26498 29404
rect 26434 29344 26498 29348
rect 26514 29404 26578 29408
rect 26514 29348 26518 29404
rect 26518 29348 26574 29404
rect 26574 29348 26578 29404
rect 26514 29344 26578 29348
rect 34715 29404 34779 29408
rect 34715 29348 34719 29404
rect 34719 29348 34775 29404
rect 34775 29348 34779 29404
rect 34715 29344 34779 29348
rect 34795 29404 34859 29408
rect 34795 29348 34799 29404
rect 34799 29348 34855 29404
rect 34855 29348 34859 29404
rect 34795 29344 34859 29348
rect 34875 29404 34939 29408
rect 34875 29348 34879 29404
rect 34879 29348 34935 29404
rect 34935 29348 34939 29404
rect 34875 29344 34939 29348
rect 34955 29404 35019 29408
rect 34955 29348 34959 29404
rect 34959 29348 35015 29404
rect 35015 29348 35019 29404
rect 34955 29344 35019 29348
rect 5172 28860 5236 28864
rect 5172 28804 5176 28860
rect 5176 28804 5232 28860
rect 5232 28804 5236 28860
rect 5172 28800 5236 28804
rect 5252 28860 5316 28864
rect 5252 28804 5256 28860
rect 5256 28804 5312 28860
rect 5312 28804 5316 28860
rect 5252 28800 5316 28804
rect 5332 28860 5396 28864
rect 5332 28804 5336 28860
rect 5336 28804 5392 28860
rect 5392 28804 5396 28860
rect 5332 28800 5396 28804
rect 5412 28860 5476 28864
rect 5412 28804 5416 28860
rect 5416 28804 5472 28860
rect 5472 28804 5476 28860
rect 5412 28800 5476 28804
rect 13613 28860 13677 28864
rect 13613 28804 13617 28860
rect 13617 28804 13673 28860
rect 13673 28804 13677 28860
rect 13613 28800 13677 28804
rect 13693 28860 13757 28864
rect 13693 28804 13697 28860
rect 13697 28804 13753 28860
rect 13753 28804 13757 28860
rect 13693 28800 13757 28804
rect 13773 28860 13837 28864
rect 13773 28804 13777 28860
rect 13777 28804 13833 28860
rect 13833 28804 13837 28860
rect 13773 28800 13837 28804
rect 13853 28860 13917 28864
rect 13853 28804 13857 28860
rect 13857 28804 13913 28860
rect 13913 28804 13917 28860
rect 13853 28800 13917 28804
rect 22054 28860 22118 28864
rect 22054 28804 22058 28860
rect 22058 28804 22114 28860
rect 22114 28804 22118 28860
rect 22054 28800 22118 28804
rect 22134 28860 22198 28864
rect 22134 28804 22138 28860
rect 22138 28804 22194 28860
rect 22194 28804 22198 28860
rect 22134 28800 22198 28804
rect 22214 28860 22278 28864
rect 22214 28804 22218 28860
rect 22218 28804 22274 28860
rect 22274 28804 22278 28860
rect 22214 28800 22278 28804
rect 22294 28860 22358 28864
rect 22294 28804 22298 28860
rect 22298 28804 22354 28860
rect 22354 28804 22358 28860
rect 22294 28800 22358 28804
rect 30495 28860 30559 28864
rect 30495 28804 30499 28860
rect 30499 28804 30555 28860
rect 30555 28804 30559 28860
rect 30495 28800 30559 28804
rect 30575 28860 30639 28864
rect 30575 28804 30579 28860
rect 30579 28804 30635 28860
rect 30635 28804 30639 28860
rect 30575 28800 30639 28804
rect 30655 28860 30719 28864
rect 30655 28804 30659 28860
rect 30659 28804 30715 28860
rect 30715 28804 30719 28860
rect 30655 28800 30719 28804
rect 30735 28860 30799 28864
rect 30735 28804 30739 28860
rect 30739 28804 30795 28860
rect 30795 28804 30799 28860
rect 30735 28800 30799 28804
rect 9392 28316 9456 28320
rect 9392 28260 9396 28316
rect 9396 28260 9452 28316
rect 9452 28260 9456 28316
rect 9392 28256 9456 28260
rect 9472 28316 9536 28320
rect 9472 28260 9476 28316
rect 9476 28260 9532 28316
rect 9532 28260 9536 28316
rect 9472 28256 9536 28260
rect 9552 28316 9616 28320
rect 9552 28260 9556 28316
rect 9556 28260 9612 28316
rect 9612 28260 9616 28316
rect 9552 28256 9616 28260
rect 9632 28316 9696 28320
rect 9632 28260 9636 28316
rect 9636 28260 9692 28316
rect 9692 28260 9696 28316
rect 9632 28256 9696 28260
rect 17833 28316 17897 28320
rect 17833 28260 17837 28316
rect 17837 28260 17893 28316
rect 17893 28260 17897 28316
rect 17833 28256 17897 28260
rect 17913 28316 17977 28320
rect 17913 28260 17917 28316
rect 17917 28260 17973 28316
rect 17973 28260 17977 28316
rect 17913 28256 17977 28260
rect 17993 28316 18057 28320
rect 17993 28260 17997 28316
rect 17997 28260 18053 28316
rect 18053 28260 18057 28316
rect 17993 28256 18057 28260
rect 18073 28316 18137 28320
rect 18073 28260 18077 28316
rect 18077 28260 18133 28316
rect 18133 28260 18137 28316
rect 18073 28256 18137 28260
rect 26274 28316 26338 28320
rect 26274 28260 26278 28316
rect 26278 28260 26334 28316
rect 26334 28260 26338 28316
rect 26274 28256 26338 28260
rect 26354 28316 26418 28320
rect 26354 28260 26358 28316
rect 26358 28260 26414 28316
rect 26414 28260 26418 28316
rect 26354 28256 26418 28260
rect 26434 28316 26498 28320
rect 26434 28260 26438 28316
rect 26438 28260 26494 28316
rect 26494 28260 26498 28316
rect 26434 28256 26498 28260
rect 26514 28316 26578 28320
rect 26514 28260 26518 28316
rect 26518 28260 26574 28316
rect 26574 28260 26578 28316
rect 26514 28256 26578 28260
rect 34715 28316 34779 28320
rect 34715 28260 34719 28316
rect 34719 28260 34775 28316
rect 34775 28260 34779 28316
rect 34715 28256 34779 28260
rect 34795 28316 34859 28320
rect 34795 28260 34799 28316
rect 34799 28260 34855 28316
rect 34855 28260 34859 28316
rect 34795 28256 34859 28260
rect 34875 28316 34939 28320
rect 34875 28260 34879 28316
rect 34879 28260 34935 28316
rect 34935 28260 34939 28316
rect 34875 28256 34939 28260
rect 34955 28316 35019 28320
rect 34955 28260 34959 28316
rect 34959 28260 35015 28316
rect 35015 28260 35019 28316
rect 34955 28256 35019 28260
rect 5172 27772 5236 27776
rect 5172 27716 5176 27772
rect 5176 27716 5232 27772
rect 5232 27716 5236 27772
rect 5172 27712 5236 27716
rect 5252 27772 5316 27776
rect 5252 27716 5256 27772
rect 5256 27716 5312 27772
rect 5312 27716 5316 27772
rect 5252 27712 5316 27716
rect 5332 27772 5396 27776
rect 5332 27716 5336 27772
rect 5336 27716 5392 27772
rect 5392 27716 5396 27772
rect 5332 27712 5396 27716
rect 5412 27772 5476 27776
rect 5412 27716 5416 27772
rect 5416 27716 5472 27772
rect 5472 27716 5476 27772
rect 5412 27712 5476 27716
rect 13613 27772 13677 27776
rect 13613 27716 13617 27772
rect 13617 27716 13673 27772
rect 13673 27716 13677 27772
rect 13613 27712 13677 27716
rect 13693 27772 13757 27776
rect 13693 27716 13697 27772
rect 13697 27716 13753 27772
rect 13753 27716 13757 27772
rect 13693 27712 13757 27716
rect 13773 27772 13837 27776
rect 13773 27716 13777 27772
rect 13777 27716 13833 27772
rect 13833 27716 13837 27772
rect 13773 27712 13837 27716
rect 13853 27772 13917 27776
rect 13853 27716 13857 27772
rect 13857 27716 13913 27772
rect 13913 27716 13917 27772
rect 13853 27712 13917 27716
rect 22054 27772 22118 27776
rect 22054 27716 22058 27772
rect 22058 27716 22114 27772
rect 22114 27716 22118 27772
rect 22054 27712 22118 27716
rect 22134 27772 22198 27776
rect 22134 27716 22138 27772
rect 22138 27716 22194 27772
rect 22194 27716 22198 27772
rect 22134 27712 22198 27716
rect 22214 27772 22278 27776
rect 22214 27716 22218 27772
rect 22218 27716 22274 27772
rect 22274 27716 22278 27772
rect 22214 27712 22278 27716
rect 22294 27772 22358 27776
rect 22294 27716 22298 27772
rect 22298 27716 22354 27772
rect 22354 27716 22358 27772
rect 22294 27712 22358 27716
rect 30495 27772 30559 27776
rect 30495 27716 30499 27772
rect 30499 27716 30555 27772
rect 30555 27716 30559 27772
rect 30495 27712 30559 27716
rect 30575 27772 30639 27776
rect 30575 27716 30579 27772
rect 30579 27716 30635 27772
rect 30635 27716 30639 27772
rect 30575 27712 30639 27716
rect 30655 27772 30719 27776
rect 30655 27716 30659 27772
rect 30659 27716 30715 27772
rect 30715 27716 30719 27772
rect 30655 27712 30719 27716
rect 30735 27772 30799 27776
rect 30735 27716 30739 27772
rect 30739 27716 30795 27772
rect 30795 27716 30799 27772
rect 30735 27712 30799 27716
rect 9392 27228 9456 27232
rect 9392 27172 9396 27228
rect 9396 27172 9452 27228
rect 9452 27172 9456 27228
rect 9392 27168 9456 27172
rect 9472 27228 9536 27232
rect 9472 27172 9476 27228
rect 9476 27172 9532 27228
rect 9532 27172 9536 27228
rect 9472 27168 9536 27172
rect 9552 27228 9616 27232
rect 9552 27172 9556 27228
rect 9556 27172 9612 27228
rect 9612 27172 9616 27228
rect 9552 27168 9616 27172
rect 9632 27228 9696 27232
rect 9632 27172 9636 27228
rect 9636 27172 9692 27228
rect 9692 27172 9696 27228
rect 9632 27168 9696 27172
rect 17833 27228 17897 27232
rect 17833 27172 17837 27228
rect 17837 27172 17893 27228
rect 17893 27172 17897 27228
rect 17833 27168 17897 27172
rect 17913 27228 17977 27232
rect 17913 27172 17917 27228
rect 17917 27172 17973 27228
rect 17973 27172 17977 27228
rect 17913 27168 17977 27172
rect 17993 27228 18057 27232
rect 17993 27172 17997 27228
rect 17997 27172 18053 27228
rect 18053 27172 18057 27228
rect 17993 27168 18057 27172
rect 18073 27228 18137 27232
rect 18073 27172 18077 27228
rect 18077 27172 18133 27228
rect 18133 27172 18137 27228
rect 18073 27168 18137 27172
rect 26274 27228 26338 27232
rect 26274 27172 26278 27228
rect 26278 27172 26334 27228
rect 26334 27172 26338 27228
rect 26274 27168 26338 27172
rect 26354 27228 26418 27232
rect 26354 27172 26358 27228
rect 26358 27172 26414 27228
rect 26414 27172 26418 27228
rect 26354 27168 26418 27172
rect 26434 27228 26498 27232
rect 26434 27172 26438 27228
rect 26438 27172 26494 27228
rect 26494 27172 26498 27228
rect 26434 27168 26498 27172
rect 26514 27228 26578 27232
rect 26514 27172 26518 27228
rect 26518 27172 26574 27228
rect 26574 27172 26578 27228
rect 26514 27168 26578 27172
rect 34715 27228 34779 27232
rect 34715 27172 34719 27228
rect 34719 27172 34775 27228
rect 34775 27172 34779 27228
rect 34715 27168 34779 27172
rect 34795 27228 34859 27232
rect 34795 27172 34799 27228
rect 34799 27172 34855 27228
rect 34855 27172 34859 27228
rect 34795 27168 34859 27172
rect 34875 27228 34939 27232
rect 34875 27172 34879 27228
rect 34879 27172 34935 27228
rect 34935 27172 34939 27228
rect 34875 27168 34939 27172
rect 34955 27228 35019 27232
rect 34955 27172 34959 27228
rect 34959 27172 35015 27228
rect 35015 27172 35019 27228
rect 34955 27168 35019 27172
rect 5172 26684 5236 26688
rect 5172 26628 5176 26684
rect 5176 26628 5232 26684
rect 5232 26628 5236 26684
rect 5172 26624 5236 26628
rect 5252 26684 5316 26688
rect 5252 26628 5256 26684
rect 5256 26628 5312 26684
rect 5312 26628 5316 26684
rect 5252 26624 5316 26628
rect 5332 26684 5396 26688
rect 5332 26628 5336 26684
rect 5336 26628 5392 26684
rect 5392 26628 5396 26684
rect 5332 26624 5396 26628
rect 5412 26684 5476 26688
rect 5412 26628 5416 26684
rect 5416 26628 5472 26684
rect 5472 26628 5476 26684
rect 5412 26624 5476 26628
rect 13613 26684 13677 26688
rect 13613 26628 13617 26684
rect 13617 26628 13673 26684
rect 13673 26628 13677 26684
rect 13613 26624 13677 26628
rect 13693 26684 13757 26688
rect 13693 26628 13697 26684
rect 13697 26628 13753 26684
rect 13753 26628 13757 26684
rect 13693 26624 13757 26628
rect 13773 26684 13837 26688
rect 13773 26628 13777 26684
rect 13777 26628 13833 26684
rect 13833 26628 13837 26684
rect 13773 26624 13837 26628
rect 13853 26684 13917 26688
rect 13853 26628 13857 26684
rect 13857 26628 13913 26684
rect 13913 26628 13917 26684
rect 13853 26624 13917 26628
rect 22054 26684 22118 26688
rect 22054 26628 22058 26684
rect 22058 26628 22114 26684
rect 22114 26628 22118 26684
rect 22054 26624 22118 26628
rect 22134 26684 22198 26688
rect 22134 26628 22138 26684
rect 22138 26628 22194 26684
rect 22194 26628 22198 26684
rect 22134 26624 22198 26628
rect 22214 26684 22278 26688
rect 22214 26628 22218 26684
rect 22218 26628 22274 26684
rect 22274 26628 22278 26684
rect 22214 26624 22278 26628
rect 22294 26684 22358 26688
rect 22294 26628 22298 26684
rect 22298 26628 22354 26684
rect 22354 26628 22358 26684
rect 22294 26624 22358 26628
rect 30495 26684 30559 26688
rect 30495 26628 30499 26684
rect 30499 26628 30555 26684
rect 30555 26628 30559 26684
rect 30495 26624 30559 26628
rect 30575 26684 30639 26688
rect 30575 26628 30579 26684
rect 30579 26628 30635 26684
rect 30635 26628 30639 26684
rect 30575 26624 30639 26628
rect 30655 26684 30719 26688
rect 30655 26628 30659 26684
rect 30659 26628 30715 26684
rect 30715 26628 30719 26684
rect 30655 26624 30719 26628
rect 30735 26684 30799 26688
rect 30735 26628 30739 26684
rect 30739 26628 30795 26684
rect 30795 26628 30799 26684
rect 30735 26624 30799 26628
rect 9392 26140 9456 26144
rect 9392 26084 9396 26140
rect 9396 26084 9452 26140
rect 9452 26084 9456 26140
rect 9392 26080 9456 26084
rect 9472 26140 9536 26144
rect 9472 26084 9476 26140
rect 9476 26084 9532 26140
rect 9532 26084 9536 26140
rect 9472 26080 9536 26084
rect 9552 26140 9616 26144
rect 9552 26084 9556 26140
rect 9556 26084 9612 26140
rect 9612 26084 9616 26140
rect 9552 26080 9616 26084
rect 9632 26140 9696 26144
rect 9632 26084 9636 26140
rect 9636 26084 9692 26140
rect 9692 26084 9696 26140
rect 9632 26080 9696 26084
rect 17833 26140 17897 26144
rect 17833 26084 17837 26140
rect 17837 26084 17893 26140
rect 17893 26084 17897 26140
rect 17833 26080 17897 26084
rect 17913 26140 17977 26144
rect 17913 26084 17917 26140
rect 17917 26084 17973 26140
rect 17973 26084 17977 26140
rect 17913 26080 17977 26084
rect 17993 26140 18057 26144
rect 17993 26084 17997 26140
rect 17997 26084 18053 26140
rect 18053 26084 18057 26140
rect 17993 26080 18057 26084
rect 18073 26140 18137 26144
rect 18073 26084 18077 26140
rect 18077 26084 18133 26140
rect 18133 26084 18137 26140
rect 18073 26080 18137 26084
rect 26274 26140 26338 26144
rect 26274 26084 26278 26140
rect 26278 26084 26334 26140
rect 26334 26084 26338 26140
rect 26274 26080 26338 26084
rect 26354 26140 26418 26144
rect 26354 26084 26358 26140
rect 26358 26084 26414 26140
rect 26414 26084 26418 26140
rect 26354 26080 26418 26084
rect 26434 26140 26498 26144
rect 26434 26084 26438 26140
rect 26438 26084 26494 26140
rect 26494 26084 26498 26140
rect 26434 26080 26498 26084
rect 26514 26140 26578 26144
rect 26514 26084 26518 26140
rect 26518 26084 26574 26140
rect 26574 26084 26578 26140
rect 26514 26080 26578 26084
rect 34715 26140 34779 26144
rect 34715 26084 34719 26140
rect 34719 26084 34775 26140
rect 34775 26084 34779 26140
rect 34715 26080 34779 26084
rect 34795 26140 34859 26144
rect 34795 26084 34799 26140
rect 34799 26084 34855 26140
rect 34855 26084 34859 26140
rect 34795 26080 34859 26084
rect 34875 26140 34939 26144
rect 34875 26084 34879 26140
rect 34879 26084 34935 26140
rect 34935 26084 34939 26140
rect 34875 26080 34939 26084
rect 34955 26140 35019 26144
rect 34955 26084 34959 26140
rect 34959 26084 35015 26140
rect 35015 26084 35019 26140
rect 34955 26080 35019 26084
rect 5172 25596 5236 25600
rect 5172 25540 5176 25596
rect 5176 25540 5232 25596
rect 5232 25540 5236 25596
rect 5172 25536 5236 25540
rect 5252 25596 5316 25600
rect 5252 25540 5256 25596
rect 5256 25540 5312 25596
rect 5312 25540 5316 25596
rect 5252 25536 5316 25540
rect 5332 25596 5396 25600
rect 5332 25540 5336 25596
rect 5336 25540 5392 25596
rect 5392 25540 5396 25596
rect 5332 25536 5396 25540
rect 5412 25596 5476 25600
rect 5412 25540 5416 25596
rect 5416 25540 5472 25596
rect 5472 25540 5476 25596
rect 5412 25536 5476 25540
rect 13613 25596 13677 25600
rect 13613 25540 13617 25596
rect 13617 25540 13673 25596
rect 13673 25540 13677 25596
rect 13613 25536 13677 25540
rect 13693 25596 13757 25600
rect 13693 25540 13697 25596
rect 13697 25540 13753 25596
rect 13753 25540 13757 25596
rect 13693 25536 13757 25540
rect 13773 25596 13837 25600
rect 13773 25540 13777 25596
rect 13777 25540 13833 25596
rect 13833 25540 13837 25596
rect 13773 25536 13837 25540
rect 13853 25596 13917 25600
rect 13853 25540 13857 25596
rect 13857 25540 13913 25596
rect 13913 25540 13917 25596
rect 13853 25536 13917 25540
rect 22054 25596 22118 25600
rect 22054 25540 22058 25596
rect 22058 25540 22114 25596
rect 22114 25540 22118 25596
rect 22054 25536 22118 25540
rect 22134 25596 22198 25600
rect 22134 25540 22138 25596
rect 22138 25540 22194 25596
rect 22194 25540 22198 25596
rect 22134 25536 22198 25540
rect 22214 25596 22278 25600
rect 22214 25540 22218 25596
rect 22218 25540 22274 25596
rect 22274 25540 22278 25596
rect 22214 25536 22278 25540
rect 22294 25596 22358 25600
rect 22294 25540 22298 25596
rect 22298 25540 22354 25596
rect 22354 25540 22358 25596
rect 22294 25536 22358 25540
rect 30495 25596 30559 25600
rect 30495 25540 30499 25596
rect 30499 25540 30555 25596
rect 30555 25540 30559 25596
rect 30495 25536 30559 25540
rect 30575 25596 30639 25600
rect 30575 25540 30579 25596
rect 30579 25540 30635 25596
rect 30635 25540 30639 25596
rect 30575 25536 30639 25540
rect 30655 25596 30719 25600
rect 30655 25540 30659 25596
rect 30659 25540 30715 25596
rect 30715 25540 30719 25596
rect 30655 25536 30719 25540
rect 30735 25596 30799 25600
rect 30735 25540 30739 25596
rect 30739 25540 30795 25596
rect 30795 25540 30799 25596
rect 30735 25536 30799 25540
rect 9392 25052 9456 25056
rect 9392 24996 9396 25052
rect 9396 24996 9452 25052
rect 9452 24996 9456 25052
rect 9392 24992 9456 24996
rect 9472 25052 9536 25056
rect 9472 24996 9476 25052
rect 9476 24996 9532 25052
rect 9532 24996 9536 25052
rect 9472 24992 9536 24996
rect 9552 25052 9616 25056
rect 9552 24996 9556 25052
rect 9556 24996 9612 25052
rect 9612 24996 9616 25052
rect 9552 24992 9616 24996
rect 9632 25052 9696 25056
rect 9632 24996 9636 25052
rect 9636 24996 9692 25052
rect 9692 24996 9696 25052
rect 9632 24992 9696 24996
rect 17833 25052 17897 25056
rect 17833 24996 17837 25052
rect 17837 24996 17893 25052
rect 17893 24996 17897 25052
rect 17833 24992 17897 24996
rect 17913 25052 17977 25056
rect 17913 24996 17917 25052
rect 17917 24996 17973 25052
rect 17973 24996 17977 25052
rect 17913 24992 17977 24996
rect 17993 25052 18057 25056
rect 17993 24996 17997 25052
rect 17997 24996 18053 25052
rect 18053 24996 18057 25052
rect 17993 24992 18057 24996
rect 18073 25052 18137 25056
rect 18073 24996 18077 25052
rect 18077 24996 18133 25052
rect 18133 24996 18137 25052
rect 18073 24992 18137 24996
rect 26274 25052 26338 25056
rect 26274 24996 26278 25052
rect 26278 24996 26334 25052
rect 26334 24996 26338 25052
rect 26274 24992 26338 24996
rect 26354 25052 26418 25056
rect 26354 24996 26358 25052
rect 26358 24996 26414 25052
rect 26414 24996 26418 25052
rect 26354 24992 26418 24996
rect 26434 25052 26498 25056
rect 26434 24996 26438 25052
rect 26438 24996 26494 25052
rect 26494 24996 26498 25052
rect 26434 24992 26498 24996
rect 26514 25052 26578 25056
rect 26514 24996 26518 25052
rect 26518 24996 26574 25052
rect 26574 24996 26578 25052
rect 26514 24992 26578 24996
rect 34715 25052 34779 25056
rect 34715 24996 34719 25052
rect 34719 24996 34775 25052
rect 34775 24996 34779 25052
rect 34715 24992 34779 24996
rect 34795 25052 34859 25056
rect 34795 24996 34799 25052
rect 34799 24996 34855 25052
rect 34855 24996 34859 25052
rect 34795 24992 34859 24996
rect 34875 25052 34939 25056
rect 34875 24996 34879 25052
rect 34879 24996 34935 25052
rect 34935 24996 34939 25052
rect 34875 24992 34939 24996
rect 34955 25052 35019 25056
rect 34955 24996 34959 25052
rect 34959 24996 35015 25052
rect 35015 24996 35019 25052
rect 34955 24992 35019 24996
rect 5172 24508 5236 24512
rect 5172 24452 5176 24508
rect 5176 24452 5232 24508
rect 5232 24452 5236 24508
rect 5172 24448 5236 24452
rect 5252 24508 5316 24512
rect 5252 24452 5256 24508
rect 5256 24452 5312 24508
rect 5312 24452 5316 24508
rect 5252 24448 5316 24452
rect 5332 24508 5396 24512
rect 5332 24452 5336 24508
rect 5336 24452 5392 24508
rect 5392 24452 5396 24508
rect 5332 24448 5396 24452
rect 5412 24508 5476 24512
rect 5412 24452 5416 24508
rect 5416 24452 5472 24508
rect 5472 24452 5476 24508
rect 5412 24448 5476 24452
rect 13613 24508 13677 24512
rect 13613 24452 13617 24508
rect 13617 24452 13673 24508
rect 13673 24452 13677 24508
rect 13613 24448 13677 24452
rect 13693 24508 13757 24512
rect 13693 24452 13697 24508
rect 13697 24452 13753 24508
rect 13753 24452 13757 24508
rect 13693 24448 13757 24452
rect 13773 24508 13837 24512
rect 13773 24452 13777 24508
rect 13777 24452 13833 24508
rect 13833 24452 13837 24508
rect 13773 24448 13837 24452
rect 13853 24508 13917 24512
rect 13853 24452 13857 24508
rect 13857 24452 13913 24508
rect 13913 24452 13917 24508
rect 13853 24448 13917 24452
rect 22054 24508 22118 24512
rect 22054 24452 22058 24508
rect 22058 24452 22114 24508
rect 22114 24452 22118 24508
rect 22054 24448 22118 24452
rect 22134 24508 22198 24512
rect 22134 24452 22138 24508
rect 22138 24452 22194 24508
rect 22194 24452 22198 24508
rect 22134 24448 22198 24452
rect 22214 24508 22278 24512
rect 22214 24452 22218 24508
rect 22218 24452 22274 24508
rect 22274 24452 22278 24508
rect 22214 24448 22278 24452
rect 22294 24508 22358 24512
rect 22294 24452 22298 24508
rect 22298 24452 22354 24508
rect 22354 24452 22358 24508
rect 22294 24448 22358 24452
rect 30495 24508 30559 24512
rect 30495 24452 30499 24508
rect 30499 24452 30555 24508
rect 30555 24452 30559 24508
rect 30495 24448 30559 24452
rect 30575 24508 30639 24512
rect 30575 24452 30579 24508
rect 30579 24452 30635 24508
rect 30635 24452 30639 24508
rect 30575 24448 30639 24452
rect 30655 24508 30719 24512
rect 30655 24452 30659 24508
rect 30659 24452 30715 24508
rect 30715 24452 30719 24508
rect 30655 24448 30719 24452
rect 30735 24508 30799 24512
rect 30735 24452 30739 24508
rect 30739 24452 30795 24508
rect 30795 24452 30799 24508
rect 30735 24448 30799 24452
rect 9392 23964 9456 23968
rect 9392 23908 9396 23964
rect 9396 23908 9452 23964
rect 9452 23908 9456 23964
rect 9392 23904 9456 23908
rect 9472 23964 9536 23968
rect 9472 23908 9476 23964
rect 9476 23908 9532 23964
rect 9532 23908 9536 23964
rect 9472 23904 9536 23908
rect 9552 23964 9616 23968
rect 9552 23908 9556 23964
rect 9556 23908 9612 23964
rect 9612 23908 9616 23964
rect 9552 23904 9616 23908
rect 9632 23964 9696 23968
rect 9632 23908 9636 23964
rect 9636 23908 9692 23964
rect 9692 23908 9696 23964
rect 9632 23904 9696 23908
rect 17833 23964 17897 23968
rect 17833 23908 17837 23964
rect 17837 23908 17893 23964
rect 17893 23908 17897 23964
rect 17833 23904 17897 23908
rect 17913 23964 17977 23968
rect 17913 23908 17917 23964
rect 17917 23908 17973 23964
rect 17973 23908 17977 23964
rect 17913 23904 17977 23908
rect 17993 23964 18057 23968
rect 17993 23908 17997 23964
rect 17997 23908 18053 23964
rect 18053 23908 18057 23964
rect 17993 23904 18057 23908
rect 18073 23964 18137 23968
rect 18073 23908 18077 23964
rect 18077 23908 18133 23964
rect 18133 23908 18137 23964
rect 18073 23904 18137 23908
rect 26274 23964 26338 23968
rect 26274 23908 26278 23964
rect 26278 23908 26334 23964
rect 26334 23908 26338 23964
rect 26274 23904 26338 23908
rect 26354 23964 26418 23968
rect 26354 23908 26358 23964
rect 26358 23908 26414 23964
rect 26414 23908 26418 23964
rect 26354 23904 26418 23908
rect 26434 23964 26498 23968
rect 26434 23908 26438 23964
rect 26438 23908 26494 23964
rect 26494 23908 26498 23964
rect 26434 23904 26498 23908
rect 26514 23964 26578 23968
rect 26514 23908 26518 23964
rect 26518 23908 26574 23964
rect 26574 23908 26578 23964
rect 26514 23904 26578 23908
rect 34715 23964 34779 23968
rect 34715 23908 34719 23964
rect 34719 23908 34775 23964
rect 34775 23908 34779 23964
rect 34715 23904 34779 23908
rect 34795 23964 34859 23968
rect 34795 23908 34799 23964
rect 34799 23908 34855 23964
rect 34855 23908 34859 23964
rect 34795 23904 34859 23908
rect 34875 23964 34939 23968
rect 34875 23908 34879 23964
rect 34879 23908 34935 23964
rect 34935 23908 34939 23964
rect 34875 23904 34939 23908
rect 34955 23964 35019 23968
rect 34955 23908 34959 23964
rect 34959 23908 35015 23964
rect 35015 23908 35019 23964
rect 34955 23904 35019 23908
rect 5172 23420 5236 23424
rect 5172 23364 5176 23420
rect 5176 23364 5232 23420
rect 5232 23364 5236 23420
rect 5172 23360 5236 23364
rect 5252 23420 5316 23424
rect 5252 23364 5256 23420
rect 5256 23364 5312 23420
rect 5312 23364 5316 23420
rect 5252 23360 5316 23364
rect 5332 23420 5396 23424
rect 5332 23364 5336 23420
rect 5336 23364 5392 23420
rect 5392 23364 5396 23420
rect 5332 23360 5396 23364
rect 5412 23420 5476 23424
rect 5412 23364 5416 23420
rect 5416 23364 5472 23420
rect 5472 23364 5476 23420
rect 5412 23360 5476 23364
rect 13613 23420 13677 23424
rect 13613 23364 13617 23420
rect 13617 23364 13673 23420
rect 13673 23364 13677 23420
rect 13613 23360 13677 23364
rect 13693 23420 13757 23424
rect 13693 23364 13697 23420
rect 13697 23364 13753 23420
rect 13753 23364 13757 23420
rect 13693 23360 13757 23364
rect 13773 23420 13837 23424
rect 13773 23364 13777 23420
rect 13777 23364 13833 23420
rect 13833 23364 13837 23420
rect 13773 23360 13837 23364
rect 13853 23420 13917 23424
rect 13853 23364 13857 23420
rect 13857 23364 13913 23420
rect 13913 23364 13917 23420
rect 13853 23360 13917 23364
rect 22054 23420 22118 23424
rect 22054 23364 22058 23420
rect 22058 23364 22114 23420
rect 22114 23364 22118 23420
rect 22054 23360 22118 23364
rect 22134 23420 22198 23424
rect 22134 23364 22138 23420
rect 22138 23364 22194 23420
rect 22194 23364 22198 23420
rect 22134 23360 22198 23364
rect 22214 23420 22278 23424
rect 22214 23364 22218 23420
rect 22218 23364 22274 23420
rect 22274 23364 22278 23420
rect 22214 23360 22278 23364
rect 22294 23420 22358 23424
rect 22294 23364 22298 23420
rect 22298 23364 22354 23420
rect 22354 23364 22358 23420
rect 22294 23360 22358 23364
rect 30495 23420 30559 23424
rect 30495 23364 30499 23420
rect 30499 23364 30555 23420
rect 30555 23364 30559 23420
rect 30495 23360 30559 23364
rect 30575 23420 30639 23424
rect 30575 23364 30579 23420
rect 30579 23364 30635 23420
rect 30635 23364 30639 23420
rect 30575 23360 30639 23364
rect 30655 23420 30719 23424
rect 30655 23364 30659 23420
rect 30659 23364 30715 23420
rect 30715 23364 30719 23420
rect 30655 23360 30719 23364
rect 30735 23420 30799 23424
rect 30735 23364 30739 23420
rect 30739 23364 30795 23420
rect 30795 23364 30799 23420
rect 30735 23360 30799 23364
rect 24900 23156 24964 23220
rect 9392 22876 9456 22880
rect 9392 22820 9396 22876
rect 9396 22820 9452 22876
rect 9452 22820 9456 22876
rect 9392 22816 9456 22820
rect 9472 22876 9536 22880
rect 9472 22820 9476 22876
rect 9476 22820 9532 22876
rect 9532 22820 9536 22876
rect 9472 22816 9536 22820
rect 9552 22876 9616 22880
rect 9552 22820 9556 22876
rect 9556 22820 9612 22876
rect 9612 22820 9616 22876
rect 9552 22816 9616 22820
rect 9632 22876 9696 22880
rect 9632 22820 9636 22876
rect 9636 22820 9692 22876
rect 9692 22820 9696 22876
rect 9632 22816 9696 22820
rect 17833 22876 17897 22880
rect 17833 22820 17837 22876
rect 17837 22820 17893 22876
rect 17893 22820 17897 22876
rect 17833 22816 17897 22820
rect 17913 22876 17977 22880
rect 17913 22820 17917 22876
rect 17917 22820 17973 22876
rect 17973 22820 17977 22876
rect 17913 22816 17977 22820
rect 17993 22876 18057 22880
rect 17993 22820 17997 22876
rect 17997 22820 18053 22876
rect 18053 22820 18057 22876
rect 17993 22816 18057 22820
rect 18073 22876 18137 22880
rect 18073 22820 18077 22876
rect 18077 22820 18133 22876
rect 18133 22820 18137 22876
rect 18073 22816 18137 22820
rect 26274 22876 26338 22880
rect 26274 22820 26278 22876
rect 26278 22820 26334 22876
rect 26334 22820 26338 22876
rect 26274 22816 26338 22820
rect 26354 22876 26418 22880
rect 26354 22820 26358 22876
rect 26358 22820 26414 22876
rect 26414 22820 26418 22876
rect 26354 22816 26418 22820
rect 26434 22876 26498 22880
rect 26434 22820 26438 22876
rect 26438 22820 26494 22876
rect 26494 22820 26498 22876
rect 26434 22816 26498 22820
rect 26514 22876 26578 22880
rect 26514 22820 26518 22876
rect 26518 22820 26574 22876
rect 26574 22820 26578 22876
rect 26514 22816 26578 22820
rect 34715 22876 34779 22880
rect 34715 22820 34719 22876
rect 34719 22820 34775 22876
rect 34775 22820 34779 22876
rect 34715 22816 34779 22820
rect 34795 22876 34859 22880
rect 34795 22820 34799 22876
rect 34799 22820 34855 22876
rect 34855 22820 34859 22876
rect 34795 22816 34859 22820
rect 34875 22876 34939 22880
rect 34875 22820 34879 22876
rect 34879 22820 34935 22876
rect 34935 22820 34939 22876
rect 34875 22816 34939 22820
rect 34955 22876 35019 22880
rect 34955 22820 34959 22876
rect 34959 22820 35015 22876
rect 35015 22820 35019 22876
rect 34955 22816 35019 22820
rect 5172 22332 5236 22336
rect 5172 22276 5176 22332
rect 5176 22276 5232 22332
rect 5232 22276 5236 22332
rect 5172 22272 5236 22276
rect 5252 22332 5316 22336
rect 5252 22276 5256 22332
rect 5256 22276 5312 22332
rect 5312 22276 5316 22332
rect 5252 22272 5316 22276
rect 5332 22332 5396 22336
rect 5332 22276 5336 22332
rect 5336 22276 5392 22332
rect 5392 22276 5396 22332
rect 5332 22272 5396 22276
rect 5412 22332 5476 22336
rect 5412 22276 5416 22332
rect 5416 22276 5472 22332
rect 5472 22276 5476 22332
rect 5412 22272 5476 22276
rect 13613 22332 13677 22336
rect 13613 22276 13617 22332
rect 13617 22276 13673 22332
rect 13673 22276 13677 22332
rect 13613 22272 13677 22276
rect 13693 22332 13757 22336
rect 13693 22276 13697 22332
rect 13697 22276 13753 22332
rect 13753 22276 13757 22332
rect 13693 22272 13757 22276
rect 13773 22332 13837 22336
rect 13773 22276 13777 22332
rect 13777 22276 13833 22332
rect 13833 22276 13837 22332
rect 13773 22272 13837 22276
rect 13853 22332 13917 22336
rect 13853 22276 13857 22332
rect 13857 22276 13913 22332
rect 13913 22276 13917 22332
rect 13853 22272 13917 22276
rect 22054 22332 22118 22336
rect 22054 22276 22058 22332
rect 22058 22276 22114 22332
rect 22114 22276 22118 22332
rect 22054 22272 22118 22276
rect 22134 22332 22198 22336
rect 22134 22276 22138 22332
rect 22138 22276 22194 22332
rect 22194 22276 22198 22332
rect 22134 22272 22198 22276
rect 22214 22332 22278 22336
rect 22214 22276 22218 22332
rect 22218 22276 22274 22332
rect 22274 22276 22278 22332
rect 22214 22272 22278 22276
rect 22294 22332 22358 22336
rect 22294 22276 22298 22332
rect 22298 22276 22354 22332
rect 22354 22276 22358 22332
rect 22294 22272 22358 22276
rect 30495 22332 30559 22336
rect 30495 22276 30499 22332
rect 30499 22276 30555 22332
rect 30555 22276 30559 22332
rect 30495 22272 30559 22276
rect 30575 22332 30639 22336
rect 30575 22276 30579 22332
rect 30579 22276 30635 22332
rect 30635 22276 30639 22332
rect 30575 22272 30639 22276
rect 30655 22332 30719 22336
rect 30655 22276 30659 22332
rect 30659 22276 30715 22332
rect 30715 22276 30719 22332
rect 30655 22272 30719 22276
rect 30735 22332 30799 22336
rect 30735 22276 30739 22332
rect 30739 22276 30795 22332
rect 30795 22276 30799 22332
rect 30735 22272 30799 22276
rect 9392 21788 9456 21792
rect 9392 21732 9396 21788
rect 9396 21732 9452 21788
rect 9452 21732 9456 21788
rect 9392 21728 9456 21732
rect 9472 21788 9536 21792
rect 9472 21732 9476 21788
rect 9476 21732 9532 21788
rect 9532 21732 9536 21788
rect 9472 21728 9536 21732
rect 9552 21788 9616 21792
rect 9552 21732 9556 21788
rect 9556 21732 9612 21788
rect 9612 21732 9616 21788
rect 9552 21728 9616 21732
rect 9632 21788 9696 21792
rect 9632 21732 9636 21788
rect 9636 21732 9692 21788
rect 9692 21732 9696 21788
rect 9632 21728 9696 21732
rect 17833 21788 17897 21792
rect 17833 21732 17837 21788
rect 17837 21732 17893 21788
rect 17893 21732 17897 21788
rect 17833 21728 17897 21732
rect 17913 21788 17977 21792
rect 17913 21732 17917 21788
rect 17917 21732 17973 21788
rect 17973 21732 17977 21788
rect 17913 21728 17977 21732
rect 17993 21788 18057 21792
rect 17993 21732 17997 21788
rect 17997 21732 18053 21788
rect 18053 21732 18057 21788
rect 17993 21728 18057 21732
rect 18073 21788 18137 21792
rect 18073 21732 18077 21788
rect 18077 21732 18133 21788
rect 18133 21732 18137 21788
rect 18073 21728 18137 21732
rect 26274 21788 26338 21792
rect 26274 21732 26278 21788
rect 26278 21732 26334 21788
rect 26334 21732 26338 21788
rect 26274 21728 26338 21732
rect 26354 21788 26418 21792
rect 26354 21732 26358 21788
rect 26358 21732 26414 21788
rect 26414 21732 26418 21788
rect 26354 21728 26418 21732
rect 26434 21788 26498 21792
rect 26434 21732 26438 21788
rect 26438 21732 26494 21788
rect 26494 21732 26498 21788
rect 26434 21728 26498 21732
rect 26514 21788 26578 21792
rect 26514 21732 26518 21788
rect 26518 21732 26574 21788
rect 26574 21732 26578 21788
rect 26514 21728 26578 21732
rect 34715 21788 34779 21792
rect 34715 21732 34719 21788
rect 34719 21732 34775 21788
rect 34775 21732 34779 21788
rect 34715 21728 34779 21732
rect 34795 21788 34859 21792
rect 34795 21732 34799 21788
rect 34799 21732 34855 21788
rect 34855 21732 34859 21788
rect 34795 21728 34859 21732
rect 34875 21788 34939 21792
rect 34875 21732 34879 21788
rect 34879 21732 34935 21788
rect 34935 21732 34939 21788
rect 34875 21728 34939 21732
rect 34955 21788 35019 21792
rect 34955 21732 34959 21788
rect 34959 21732 35015 21788
rect 35015 21732 35019 21788
rect 34955 21728 35019 21732
rect 5172 21244 5236 21248
rect 5172 21188 5176 21244
rect 5176 21188 5232 21244
rect 5232 21188 5236 21244
rect 5172 21184 5236 21188
rect 5252 21244 5316 21248
rect 5252 21188 5256 21244
rect 5256 21188 5312 21244
rect 5312 21188 5316 21244
rect 5252 21184 5316 21188
rect 5332 21244 5396 21248
rect 5332 21188 5336 21244
rect 5336 21188 5392 21244
rect 5392 21188 5396 21244
rect 5332 21184 5396 21188
rect 5412 21244 5476 21248
rect 5412 21188 5416 21244
rect 5416 21188 5472 21244
rect 5472 21188 5476 21244
rect 5412 21184 5476 21188
rect 13613 21244 13677 21248
rect 13613 21188 13617 21244
rect 13617 21188 13673 21244
rect 13673 21188 13677 21244
rect 13613 21184 13677 21188
rect 13693 21244 13757 21248
rect 13693 21188 13697 21244
rect 13697 21188 13753 21244
rect 13753 21188 13757 21244
rect 13693 21184 13757 21188
rect 13773 21244 13837 21248
rect 13773 21188 13777 21244
rect 13777 21188 13833 21244
rect 13833 21188 13837 21244
rect 13773 21184 13837 21188
rect 13853 21244 13917 21248
rect 13853 21188 13857 21244
rect 13857 21188 13913 21244
rect 13913 21188 13917 21244
rect 13853 21184 13917 21188
rect 22054 21244 22118 21248
rect 22054 21188 22058 21244
rect 22058 21188 22114 21244
rect 22114 21188 22118 21244
rect 22054 21184 22118 21188
rect 22134 21244 22198 21248
rect 22134 21188 22138 21244
rect 22138 21188 22194 21244
rect 22194 21188 22198 21244
rect 22134 21184 22198 21188
rect 22214 21244 22278 21248
rect 22214 21188 22218 21244
rect 22218 21188 22274 21244
rect 22274 21188 22278 21244
rect 22214 21184 22278 21188
rect 22294 21244 22358 21248
rect 22294 21188 22298 21244
rect 22298 21188 22354 21244
rect 22354 21188 22358 21244
rect 22294 21184 22358 21188
rect 30495 21244 30559 21248
rect 30495 21188 30499 21244
rect 30499 21188 30555 21244
rect 30555 21188 30559 21244
rect 30495 21184 30559 21188
rect 30575 21244 30639 21248
rect 30575 21188 30579 21244
rect 30579 21188 30635 21244
rect 30635 21188 30639 21244
rect 30575 21184 30639 21188
rect 30655 21244 30719 21248
rect 30655 21188 30659 21244
rect 30659 21188 30715 21244
rect 30715 21188 30719 21244
rect 30655 21184 30719 21188
rect 30735 21244 30799 21248
rect 30735 21188 30739 21244
rect 30739 21188 30795 21244
rect 30795 21188 30799 21244
rect 30735 21184 30799 21188
rect 9392 20700 9456 20704
rect 9392 20644 9396 20700
rect 9396 20644 9452 20700
rect 9452 20644 9456 20700
rect 9392 20640 9456 20644
rect 9472 20700 9536 20704
rect 9472 20644 9476 20700
rect 9476 20644 9532 20700
rect 9532 20644 9536 20700
rect 9472 20640 9536 20644
rect 9552 20700 9616 20704
rect 9552 20644 9556 20700
rect 9556 20644 9612 20700
rect 9612 20644 9616 20700
rect 9552 20640 9616 20644
rect 9632 20700 9696 20704
rect 9632 20644 9636 20700
rect 9636 20644 9692 20700
rect 9692 20644 9696 20700
rect 9632 20640 9696 20644
rect 17833 20700 17897 20704
rect 17833 20644 17837 20700
rect 17837 20644 17893 20700
rect 17893 20644 17897 20700
rect 17833 20640 17897 20644
rect 17913 20700 17977 20704
rect 17913 20644 17917 20700
rect 17917 20644 17973 20700
rect 17973 20644 17977 20700
rect 17913 20640 17977 20644
rect 17993 20700 18057 20704
rect 17993 20644 17997 20700
rect 17997 20644 18053 20700
rect 18053 20644 18057 20700
rect 17993 20640 18057 20644
rect 18073 20700 18137 20704
rect 18073 20644 18077 20700
rect 18077 20644 18133 20700
rect 18133 20644 18137 20700
rect 18073 20640 18137 20644
rect 26274 20700 26338 20704
rect 26274 20644 26278 20700
rect 26278 20644 26334 20700
rect 26334 20644 26338 20700
rect 26274 20640 26338 20644
rect 26354 20700 26418 20704
rect 26354 20644 26358 20700
rect 26358 20644 26414 20700
rect 26414 20644 26418 20700
rect 26354 20640 26418 20644
rect 26434 20700 26498 20704
rect 26434 20644 26438 20700
rect 26438 20644 26494 20700
rect 26494 20644 26498 20700
rect 26434 20640 26498 20644
rect 26514 20700 26578 20704
rect 26514 20644 26518 20700
rect 26518 20644 26574 20700
rect 26574 20644 26578 20700
rect 26514 20640 26578 20644
rect 34715 20700 34779 20704
rect 34715 20644 34719 20700
rect 34719 20644 34775 20700
rect 34775 20644 34779 20700
rect 34715 20640 34779 20644
rect 34795 20700 34859 20704
rect 34795 20644 34799 20700
rect 34799 20644 34855 20700
rect 34855 20644 34859 20700
rect 34795 20640 34859 20644
rect 34875 20700 34939 20704
rect 34875 20644 34879 20700
rect 34879 20644 34935 20700
rect 34935 20644 34939 20700
rect 34875 20640 34939 20644
rect 34955 20700 35019 20704
rect 34955 20644 34959 20700
rect 34959 20644 35015 20700
rect 35015 20644 35019 20700
rect 34955 20640 35019 20644
rect 5172 20156 5236 20160
rect 5172 20100 5176 20156
rect 5176 20100 5232 20156
rect 5232 20100 5236 20156
rect 5172 20096 5236 20100
rect 5252 20156 5316 20160
rect 5252 20100 5256 20156
rect 5256 20100 5312 20156
rect 5312 20100 5316 20156
rect 5252 20096 5316 20100
rect 5332 20156 5396 20160
rect 5332 20100 5336 20156
rect 5336 20100 5392 20156
rect 5392 20100 5396 20156
rect 5332 20096 5396 20100
rect 5412 20156 5476 20160
rect 5412 20100 5416 20156
rect 5416 20100 5472 20156
rect 5472 20100 5476 20156
rect 5412 20096 5476 20100
rect 13613 20156 13677 20160
rect 13613 20100 13617 20156
rect 13617 20100 13673 20156
rect 13673 20100 13677 20156
rect 13613 20096 13677 20100
rect 13693 20156 13757 20160
rect 13693 20100 13697 20156
rect 13697 20100 13753 20156
rect 13753 20100 13757 20156
rect 13693 20096 13757 20100
rect 13773 20156 13837 20160
rect 13773 20100 13777 20156
rect 13777 20100 13833 20156
rect 13833 20100 13837 20156
rect 13773 20096 13837 20100
rect 13853 20156 13917 20160
rect 13853 20100 13857 20156
rect 13857 20100 13913 20156
rect 13913 20100 13917 20156
rect 13853 20096 13917 20100
rect 22054 20156 22118 20160
rect 22054 20100 22058 20156
rect 22058 20100 22114 20156
rect 22114 20100 22118 20156
rect 22054 20096 22118 20100
rect 22134 20156 22198 20160
rect 22134 20100 22138 20156
rect 22138 20100 22194 20156
rect 22194 20100 22198 20156
rect 22134 20096 22198 20100
rect 22214 20156 22278 20160
rect 22214 20100 22218 20156
rect 22218 20100 22274 20156
rect 22274 20100 22278 20156
rect 22214 20096 22278 20100
rect 22294 20156 22358 20160
rect 22294 20100 22298 20156
rect 22298 20100 22354 20156
rect 22354 20100 22358 20156
rect 22294 20096 22358 20100
rect 30495 20156 30559 20160
rect 30495 20100 30499 20156
rect 30499 20100 30555 20156
rect 30555 20100 30559 20156
rect 30495 20096 30559 20100
rect 30575 20156 30639 20160
rect 30575 20100 30579 20156
rect 30579 20100 30635 20156
rect 30635 20100 30639 20156
rect 30575 20096 30639 20100
rect 30655 20156 30719 20160
rect 30655 20100 30659 20156
rect 30659 20100 30715 20156
rect 30715 20100 30719 20156
rect 30655 20096 30719 20100
rect 30735 20156 30799 20160
rect 30735 20100 30739 20156
rect 30739 20100 30795 20156
rect 30795 20100 30799 20156
rect 30735 20096 30799 20100
rect 9392 19612 9456 19616
rect 9392 19556 9396 19612
rect 9396 19556 9452 19612
rect 9452 19556 9456 19612
rect 9392 19552 9456 19556
rect 9472 19612 9536 19616
rect 9472 19556 9476 19612
rect 9476 19556 9532 19612
rect 9532 19556 9536 19612
rect 9472 19552 9536 19556
rect 9552 19612 9616 19616
rect 9552 19556 9556 19612
rect 9556 19556 9612 19612
rect 9612 19556 9616 19612
rect 9552 19552 9616 19556
rect 9632 19612 9696 19616
rect 9632 19556 9636 19612
rect 9636 19556 9692 19612
rect 9692 19556 9696 19612
rect 9632 19552 9696 19556
rect 17833 19612 17897 19616
rect 17833 19556 17837 19612
rect 17837 19556 17893 19612
rect 17893 19556 17897 19612
rect 17833 19552 17897 19556
rect 17913 19612 17977 19616
rect 17913 19556 17917 19612
rect 17917 19556 17973 19612
rect 17973 19556 17977 19612
rect 17913 19552 17977 19556
rect 17993 19612 18057 19616
rect 17993 19556 17997 19612
rect 17997 19556 18053 19612
rect 18053 19556 18057 19612
rect 17993 19552 18057 19556
rect 18073 19612 18137 19616
rect 18073 19556 18077 19612
rect 18077 19556 18133 19612
rect 18133 19556 18137 19612
rect 18073 19552 18137 19556
rect 26274 19612 26338 19616
rect 26274 19556 26278 19612
rect 26278 19556 26334 19612
rect 26334 19556 26338 19612
rect 26274 19552 26338 19556
rect 26354 19612 26418 19616
rect 26354 19556 26358 19612
rect 26358 19556 26414 19612
rect 26414 19556 26418 19612
rect 26354 19552 26418 19556
rect 26434 19612 26498 19616
rect 26434 19556 26438 19612
rect 26438 19556 26494 19612
rect 26494 19556 26498 19612
rect 26434 19552 26498 19556
rect 26514 19612 26578 19616
rect 26514 19556 26518 19612
rect 26518 19556 26574 19612
rect 26574 19556 26578 19612
rect 26514 19552 26578 19556
rect 34715 19612 34779 19616
rect 34715 19556 34719 19612
rect 34719 19556 34775 19612
rect 34775 19556 34779 19612
rect 34715 19552 34779 19556
rect 34795 19612 34859 19616
rect 34795 19556 34799 19612
rect 34799 19556 34855 19612
rect 34855 19556 34859 19612
rect 34795 19552 34859 19556
rect 34875 19612 34939 19616
rect 34875 19556 34879 19612
rect 34879 19556 34935 19612
rect 34935 19556 34939 19612
rect 34875 19552 34939 19556
rect 34955 19612 35019 19616
rect 34955 19556 34959 19612
rect 34959 19556 35015 19612
rect 35015 19556 35019 19612
rect 34955 19552 35019 19556
rect 5172 19068 5236 19072
rect 5172 19012 5176 19068
rect 5176 19012 5232 19068
rect 5232 19012 5236 19068
rect 5172 19008 5236 19012
rect 5252 19068 5316 19072
rect 5252 19012 5256 19068
rect 5256 19012 5312 19068
rect 5312 19012 5316 19068
rect 5252 19008 5316 19012
rect 5332 19068 5396 19072
rect 5332 19012 5336 19068
rect 5336 19012 5392 19068
rect 5392 19012 5396 19068
rect 5332 19008 5396 19012
rect 5412 19068 5476 19072
rect 5412 19012 5416 19068
rect 5416 19012 5472 19068
rect 5472 19012 5476 19068
rect 5412 19008 5476 19012
rect 13613 19068 13677 19072
rect 13613 19012 13617 19068
rect 13617 19012 13673 19068
rect 13673 19012 13677 19068
rect 13613 19008 13677 19012
rect 13693 19068 13757 19072
rect 13693 19012 13697 19068
rect 13697 19012 13753 19068
rect 13753 19012 13757 19068
rect 13693 19008 13757 19012
rect 13773 19068 13837 19072
rect 13773 19012 13777 19068
rect 13777 19012 13833 19068
rect 13833 19012 13837 19068
rect 13773 19008 13837 19012
rect 13853 19068 13917 19072
rect 13853 19012 13857 19068
rect 13857 19012 13913 19068
rect 13913 19012 13917 19068
rect 13853 19008 13917 19012
rect 22054 19068 22118 19072
rect 22054 19012 22058 19068
rect 22058 19012 22114 19068
rect 22114 19012 22118 19068
rect 22054 19008 22118 19012
rect 22134 19068 22198 19072
rect 22134 19012 22138 19068
rect 22138 19012 22194 19068
rect 22194 19012 22198 19068
rect 22134 19008 22198 19012
rect 22214 19068 22278 19072
rect 22214 19012 22218 19068
rect 22218 19012 22274 19068
rect 22274 19012 22278 19068
rect 22214 19008 22278 19012
rect 22294 19068 22358 19072
rect 22294 19012 22298 19068
rect 22298 19012 22354 19068
rect 22354 19012 22358 19068
rect 22294 19008 22358 19012
rect 30495 19068 30559 19072
rect 30495 19012 30499 19068
rect 30499 19012 30555 19068
rect 30555 19012 30559 19068
rect 30495 19008 30559 19012
rect 30575 19068 30639 19072
rect 30575 19012 30579 19068
rect 30579 19012 30635 19068
rect 30635 19012 30639 19068
rect 30575 19008 30639 19012
rect 30655 19068 30719 19072
rect 30655 19012 30659 19068
rect 30659 19012 30715 19068
rect 30715 19012 30719 19068
rect 30655 19008 30719 19012
rect 30735 19068 30799 19072
rect 30735 19012 30739 19068
rect 30739 19012 30795 19068
rect 30795 19012 30799 19068
rect 30735 19008 30799 19012
rect 9392 18524 9456 18528
rect 9392 18468 9396 18524
rect 9396 18468 9452 18524
rect 9452 18468 9456 18524
rect 9392 18464 9456 18468
rect 9472 18524 9536 18528
rect 9472 18468 9476 18524
rect 9476 18468 9532 18524
rect 9532 18468 9536 18524
rect 9472 18464 9536 18468
rect 9552 18524 9616 18528
rect 9552 18468 9556 18524
rect 9556 18468 9612 18524
rect 9612 18468 9616 18524
rect 9552 18464 9616 18468
rect 9632 18524 9696 18528
rect 9632 18468 9636 18524
rect 9636 18468 9692 18524
rect 9692 18468 9696 18524
rect 9632 18464 9696 18468
rect 17833 18524 17897 18528
rect 17833 18468 17837 18524
rect 17837 18468 17893 18524
rect 17893 18468 17897 18524
rect 17833 18464 17897 18468
rect 17913 18524 17977 18528
rect 17913 18468 17917 18524
rect 17917 18468 17973 18524
rect 17973 18468 17977 18524
rect 17913 18464 17977 18468
rect 17993 18524 18057 18528
rect 17993 18468 17997 18524
rect 17997 18468 18053 18524
rect 18053 18468 18057 18524
rect 17993 18464 18057 18468
rect 18073 18524 18137 18528
rect 18073 18468 18077 18524
rect 18077 18468 18133 18524
rect 18133 18468 18137 18524
rect 18073 18464 18137 18468
rect 26274 18524 26338 18528
rect 26274 18468 26278 18524
rect 26278 18468 26334 18524
rect 26334 18468 26338 18524
rect 26274 18464 26338 18468
rect 26354 18524 26418 18528
rect 26354 18468 26358 18524
rect 26358 18468 26414 18524
rect 26414 18468 26418 18524
rect 26354 18464 26418 18468
rect 26434 18524 26498 18528
rect 26434 18468 26438 18524
rect 26438 18468 26494 18524
rect 26494 18468 26498 18524
rect 26434 18464 26498 18468
rect 26514 18524 26578 18528
rect 26514 18468 26518 18524
rect 26518 18468 26574 18524
rect 26574 18468 26578 18524
rect 26514 18464 26578 18468
rect 34715 18524 34779 18528
rect 34715 18468 34719 18524
rect 34719 18468 34775 18524
rect 34775 18468 34779 18524
rect 34715 18464 34779 18468
rect 34795 18524 34859 18528
rect 34795 18468 34799 18524
rect 34799 18468 34855 18524
rect 34855 18468 34859 18524
rect 34795 18464 34859 18468
rect 34875 18524 34939 18528
rect 34875 18468 34879 18524
rect 34879 18468 34935 18524
rect 34935 18468 34939 18524
rect 34875 18464 34939 18468
rect 34955 18524 35019 18528
rect 34955 18468 34959 18524
rect 34959 18468 35015 18524
rect 35015 18468 35019 18524
rect 34955 18464 35019 18468
rect 5172 17980 5236 17984
rect 5172 17924 5176 17980
rect 5176 17924 5232 17980
rect 5232 17924 5236 17980
rect 5172 17920 5236 17924
rect 5252 17980 5316 17984
rect 5252 17924 5256 17980
rect 5256 17924 5312 17980
rect 5312 17924 5316 17980
rect 5252 17920 5316 17924
rect 5332 17980 5396 17984
rect 5332 17924 5336 17980
rect 5336 17924 5392 17980
rect 5392 17924 5396 17980
rect 5332 17920 5396 17924
rect 5412 17980 5476 17984
rect 5412 17924 5416 17980
rect 5416 17924 5472 17980
rect 5472 17924 5476 17980
rect 5412 17920 5476 17924
rect 13613 17980 13677 17984
rect 13613 17924 13617 17980
rect 13617 17924 13673 17980
rect 13673 17924 13677 17980
rect 13613 17920 13677 17924
rect 13693 17980 13757 17984
rect 13693 17924 13697 17980
rect 13697 17924 13753 17980
rect 13753 17924 13757 17980
rect 13693 17920 13757 17924
rect 13773 17980 13837 17984
rect 13773 17924 13777 17980
rect 13777 17924 13833 17980
rect 13833 17924 13837 17980
rect 13773 17920 13837 17924
rect 13853 17980 13917 17984
rect 13853 17924 13857 17980
rect 13857 17924 13913 17980
rect 13913 17924 13917 17980
rect 13853 17920 13917 17924
rect 22054 17980 22118 17984
rect 22054 17924 22058 17980
rect 22058 17924 22114 17980
rect 22114 17924 22118 17980
rect 22054 17920 22118 17924
rect 22134 17980 22198 17984
rect 22134 17924 22138 17980
rect 22138 17924 22194 17980
rect 22194 17924 22198 17980
rect 22134 17920 22198 17924
rect 22214 17980 22278 17984
rect 22214 17924 22218 17980
rect 22218 17924 22274 17980
rect 22274 17924 22278 17980
rect 22214 17920 22278 17924
rect 22294 17980 22358 17984
rect 22294 17924 22298 17980
rect 22298 17924 22354 17980
rect 22354 17924 22358 17980
rect 22294 17920 22358 17924
rect 30495 17980 30559 17984
rect 30495 17924 30499 17980
rect 30499 17924 30555 17980
rect 30555 17924 30559 17980
rect 30495 17920 30559 17924
rect 30575 17980 30639 17984
rect 30575 17924 30579 17980
rect 30579 17924 30635 17980
rect 30635 17924 30639 17980
rect 30575 17920 30639 17924
rect 30655 17980 30719 17984
rect 30655 17924 30659 17980
rect 30659 17924 30715 17980
rect 30715 17924 30719 17980
rect 30655 17920 30719 17924
rect 30735 17980 30799 17984
rect 30735 17924 30739 17980
rect 30739 17924 30795 17980
rect 30795 17924 30799 17980
rect 30735 17920 30799 17924
rect 9392 17436 9456 17440
rect 9392 17380 9396 17436
rect 9396 17380 9452 17436
rect 9452 17380 9456 17436
rect 9392 17376 9456 17380
rect 9472 17436 9536 17440
rect 9472 17380 9476 17436
rect 9476 17380 9532 17436
rect 9532 17380 9536 17436
rect 9472 17376 9536 17380
rect 9552 17436 9616 17440
rect 9552 17380 9556 17436
rect 9556 17380 9612 17436
rect 9612 17380 9616 17436
rect 9552 17376 9616 17380
rect 9632 17436 9696 17440
rect 9632 17380 9636 17436
rect 9636 17380 9692 17436
rect 9692 17380 9696 17436
rect 9632 17376 9696 17380
rect 17833 17436 17897 17440
rect 17833 17380 17837 17436
rect 17837 17380 17893 17436
rect 17893 17380 17897 17436
rect 17833 17376 17897 17380
rect 17913 17436 17977 17440
rect 17913 17380 17917 17436
rect 17917 17380 17973 17436
rect 17973 17380 17977 17436
rect 17913 17376 17977 17380
rect 17993 17436 18057 17440
rect 17993 17380 17997 17436
rect 17997 17380 18053 17436
rect 18053 17380 18057 17436
rect 17993 17376 18057 17380
rect 18073 17436 18137 17440
rect 18073 17380 18077 17436
rect 18077 17380 18133 17436
rect 18133 17380 18137 17436
rect 18073 17376 18137 17380
rect 26274 17436 26338 17440
rect 26274 17380 26278 17436
rect 26278 17380 26334 17436
rect 26334 17380 26338 17436
rect 26274 17376 26338 17380
rect 26354 17436 26418 17440
rect 26354 17380 26358 17436
rect 26358 17380 26414 17436
rect 26414 17380 26418 17436
rect 26354 17376 26418 17380
rect 26434 17436 26498 17440
rect 26434 17380 26438 17436
rect 26438 17380 26494 17436
rect 26494 17380 26498 17436
rect 26434 17376 26498 17380
rect 26514 17436 26578 17440
rect 26514 17380 26518 17436
rect 26518 17380 26574 17436
rect 26574 17380 26578 17436
rect 26514 17376 26578 17380
rect 34715 17436 34779 17440
rect 34715 17380 34719 17436
rect 34719 17380 34775 17436
rect 34775 17380 34779 17436
rect 34715 17376 34779 17380
rect 34795 17436 34859 17440
rect 34795 17380 34799 17436
rect 34799 17380 34855 17436
rect 34855 17380 34859 17436
rect 34795 17376 34859 17380
rect 34875 17436 34939 17440
rect 34875 17380 34879 17436
rect 34879 17380 34935 17436
rect 34935 17380 34939 17436
rect 34875 17376 34939 17380
rect 34955 17436 35019 17440
rect 34955 17380 34959 17436
rect 34959 17380 35015 17436
rect 35015 17380 35019 17436
rect 34955 17376 35019 17380
rect 5172 16892 5236 16896
rect 5172 16836 5176 16892
rect 5176 16836 5232 16892
rect 5232 16836 5236 16892
rect 5172 16832 5236 16836
rect 5252 16892 5316 16896
rect 5252 16836 5256 16892
rect 5256 16836 5312 16892
rect 5312 16836 5316 16892
rect 5252 16832 5316 16836
rect 5332 16892 5396 16896
rect 5332 16836 5336 16892
rect 5336 16836 5392 16892
rect 5392 16836 5396 16892
rect 5332 16832 5396 16836
rect 5412 16892 5476 16896
rect 5412 16836 5416 16892
rect 5416 16836 5472 16892
rect 5472 16836 5476 16892
rect 5412 16832 5476 16836
rect 13613 16892 13677 16896
rect 13613 16836 13617 16892
rect 13617 16836 13673 16892
rect 13673 16836 13677 16892
rect 13613 16832 13677 16836
rect 13693 16892 13757 16896
rect 13693 16836 13697 16892
rect 13697 16836 13753 16892
rect 13753 16836 13757 16892
rect 13693 16832 13757 16836
rect 13773 16892 13837 16896
rect 13773 16836 13777 16892
rect 13777 16836 13833 16892
rect 13833 16836 13837 16892
rect 13773 16832 13837 16836
rect 13853 16892 13917 16896
rect 13853 16836 13857 16892
rect 13857 16836 13913 16892
rect 13913 16836 13917 16892
rect 13853 16832 13917 16836
rect 22054 16892 22118 16896
rect 22054 16836 22058 16892
rect 22058 16836 22114 16892
rect 22114 16836 22118 16892
rect 22054 16832 22118 16836
rect 22134 16892 22198 16896
rect 22134 16836 22138 16892
rect 22138 16836 22194 16892
rect 22194 16836 22198 16892
rect 22134 16832 22198 16836
rect 22214 16892 22278 16896
rect 22214 16836 22218 16892
rect 22218 16836 22274 16892
rect 22274 16836 22278 16892
rect 22214 16832 22278 16836
rect 22294 16892 22358 16896
rect 22294 16836 22298 16892
rect 22298 16836 22354 16892
rect 22354 16836 22358 16892
rect 22294 16832 22358 16836
rect 30495 16892 30559 16896
rect 30495 16836 30499 16892
rect 30499 16836 30555 16892
rect 30555 16836 30559 16892
rect 30495 16832 30559 16836
rect 30575 16892 30639 16896
rect 30575 16836 30579 16892
rect 30579 16836 30635 16892
rect 30635 16836 30639 16892
rect 30575 16832 30639 16836
rect 30655 16892 30719 16896
rect 30655 16836 30659 16892
rect 30659 16836 30715 16892
rect 30715 16836 30719 16892
rect 30655 16832 30719 16836
rect 30735 16892 30799 16896
rect 30735 16836 30739 16892
rect 30739 16836 30795 16892
rect 30795 16836 30799 16892
rect 30735 16832 30799 16836
rect 9392 16348 9456 16352
rect 9392 16292 9396 16348
rect 9396 16292 9452 16348
rect 9452 16292 9456 16348
rect 9392 16288 9456 16292
rect 9472 16348 9536 16352
rect 9472 16292 9476 16348
rect 9476 16292 9532 16348
rect 9532 16292 9536 16348
rect 9472 16288 9536 16292
rect 9552 16348 9616 16352
rect 9552 16292 9556 16348
rect 9556 16292 9612 16348
rect 9612 16292 9616 16348
rect 9552 16288 9616 16292
rect 9632 16348 9696 16352
rect 9632 16292 9636 16348
rect 9636 16292 9692 16348
rect 9692 16292 9696 16348
rect 9632 16288 9696 16292
rect 17833 16348 17897 16352
rect 17833 16292 17837 16348
rect 17837 16292 17893 16348
rect 17893 16292 17897 16348
rect 17833 16288 17897 16292
rect 17913 16348 17977 16352
rect 17913 16292 17917 16348
rect 17917 16292 17973 16348
rect 17973 16292 17977 16348
rect 17913 16288 17977 16292
rect 17993 16348 18057 16352
rect 17993 16292 17997 16348
rect 17997 16292 18053 16348
rect 18053 16292 18057 16348
rect 17993 16288 18057 16292
rect 18073 16348 18137 16352
rect 18073 16292 18077 16348
rect 18077 16292 18133 16348
rect 18133 16292 18137 16348
rect 18073 16288 18137 16292
rect 26274 16348 26338 16352
rect 26274 16292 26278 16348
rect 26278 16292 26334 16348
rect 26334 16292 26338 16348
rect 26274 16288 26338 16292
rect 26354 16348 26418 16352
rect 26354 16292 26358 16348
rect 26358 16292 26414 16348
rect 26414 16292 26418 16348
rect 26354 16288 26418 16292
rect 26434 16348 26498 16352
rect 26434 16292 26438 16348
rect 26438 16292 26494 16348
rect 26494 16292 26498 16348
rect 26434 16288 26498 16292
rect 26514 16348 26578 16352
rect 26514 16292 26518 16348
rect 26518 16292 26574 16348
rect 26574 16292 26578 16348
rect 26514 16288 26578 16292
rect 34715 16348 34779 16352
rect 34715 16292 34719 16348
rect 34719 16292 34775 16348
rect 34775 16292 34779 16348
rect 34715 16288 34779 16292
rect 34795 16348 34859 16352
rect 34795 16292 34799 16348
rect 34799 16292 34855 16348
rect 34855 16292 34859 16348
rect 34795 16288 34859 16292
rect 34875 16348 34939 16352
rect 34875 16292 34879 16348
rect 34879 16292 34935 16348
rect 34935 16292 34939 16348
rect 34875 16288 34939 16292
rect 34955 16348 35019 16352
rect 34955 16292 34959 16348
rect 34959 16292 35015 16348
rect 35015 16292 35019 16348
rect 34955 16288 35019 16292
rect 5172 15804 5236 15808
rect 5172 15748 5176 15804
rect 5176 15748 5232 15804
rect 5232 15748 5236 15804
rect 5172 15744 5236 15748
rect 5252 15804 5316 15808
rect 5252 15748 5256 15804
rect 5256 15748 5312 15804
rect 5312 15748 5316 15804
rect 5252 15744 5316 15748
rect 5332 15804 5396 15808
rect 5332 15748 5336 15804
rect 5336 15748 5392 15804
rect 5392 15748 5396 15804
rect 5332 15744 5396 15748
rect 5412 15804 5476 15808
rect 5412 15748 5416 15804
rect 5416 15748 5472 15804
rect 5472 15748 5476 15804
rect 5412 15744 5476 15748
rect 13613 15804 13677 15808
rect 13613 15748 13617 15804
rect 13617 15748 13673 15804
rect 13673 15748 13677 15804
rect 13613 15744 13677 15748
rect 13693 15804 13757 15808
rect 13693 15748 13697 15804
rect 13697 15748 13753 15804
rect 13753 15748 13757 15804
rect 13693 15744 13757 15748
rect 13773 15804 13837 15808
rect 13773 15748 13777 15804
rect 13777 15748 13833 15804
rect 13833 15748 13837 15804
rect 13773 15744 13837 15748
rect 13853 15804 13917 15808
rect 13853 15748 13857 15804
rect 13857 15748 13913 15804
rect 13913 15748 13917 15804
rect 13853 15744 13917 15748
rect 22054 15804 22118 15808
rect 22054 15748 22058 15804
rect 22058 15748 22114 15804
rect 22114 15748 22118 15804
rect 22054 15744 22118 15748
rect 22134 15804 22198 15808
rect 22134 15748 22138 15804
rect 22138 15748 22194 15804
rect 22194 15748 22198 15804
rect 22134 15744 22198 15748
rect 22214 15804 22278 15808
rect 22214 15748 22218 15804
rect 22218 15748 22274 15804
rect 22274 15748 22278 15804
rect 22214 15744 22278 15748
rect 22294 15804 22358 15808
rect 22294 15748 22298 15804
rect 22298 15748 22354 15804
rect 22354 15748 22358 15804
rect 22294 15744 22358 15748
rect 30495 15804 30559 15808
rect 30495 15748 30499 15804
rect 30499 15748 30555 15804
rect 30555 15748 30559 15804
rect 30495 15744 30559 15748
rect 30575 15804 30639 15808
rect 30575 15748 30579 15804
rect 30579 15748 30635 15804
rect 30635 15748 30639 15804
rect 30575 15744 30639 15748
rect 30655 15804 30719 15808
rect 30655 15748 30659 15804
rect 30659 15748 30715 15804
rect 30715 15748 30719 15804
rect 30655 15744 30719 15748
rect 30735 15804 30799 15808
rect 30735 15748 30739 15804
rect 30739 15748 30795 15804
rect 30795 15748 30799 15804
rect 30735 15744 30799 15748
rect 9392 15260 9456 15264
rect 9392 15204 9396 15260
rect 9396 15204 9452 15260
rect 9452 15204 9456 15260
rect 9392 15200 9456 15204
rect 9472 15260 9536 15264
rect 9472 15204 9476 15260
rect 9476 15204 9532 15260
rect 9532 15204 9536 15260
rect 9472 15200 9536 15204
rect 9552 15260 9616 15264
rect 9552 15204 9556 15260
rect 9556 15204 9612 15260
rect 9612 15204 9616 15260
rect 9552 15200 9616 15204
rect 9632 15260 9696 15264
rect 9632 15204 9636 15260
rect 9636 15204 9692 15260
rect 9692 15204 9696 15260
rect 9632 15200 9696 15204
rect 17833 15260 17897 15264
rect 17833 15204 17837 15260
rect 17837 15204 17893 15260
rect 17893 15204 17897 15260
rect 17833 15200 17897 15204
rect 17913 15260 17977 15264
rect 17913 15204 17917 15260
rect 17917 15204 17973 15260
rect 17973 15204 17977 15260
rect 17913 15200 17977 15204
rect 17993 15260 18057 15264
rect 17993 15204 17997 15260
rect 17997 15204 18053 15260
rect 18053 15204 18057 15260
rect 17993 15200 18057 15204
rect 18073 15260 18137 15264
rect 18073 15204 18077 15260
rect 18077 15204 18133 15260
rect 18133 15204 18137 15260
rect 18073 15200 18137 15204
rect 26274 15260 26338 15264
rect 26274 15204 26278 15260
rect 26278 15204 26334 15260
rect 26334 15204 26338 15260
rect 26274 15200 26338 15204
rect 26354 15260 26418 15264
rect 26354 15204 26358 15260
rect 26358 15204 26414 15260
rect 26414 15204 26418 15260
rect 26354 15200 26418 15204
rect 26434 15260 26498 15264
rect 26434 15204 26438 15260
rect 26438 15204 26494 15260
rect 26494 15204 26498 15260
rect 26434 15200 26498 15204
rect 26514 15260 26578 15264
rect 26514 15204 26518 15260
rect 26518 15204 26574 15260
rect 26574 15204 26578 15260
rect 26514 15200 26578 15204
rect 34715 15260 34779 15264
rect 34715 15204 34719 15260
rect 34719 15204 34775 15260
rect 34775 15204 34779 15260
rect 34715 15200 34779 15204
rect 34795 15260 34859 15264
rect 34795 15204 34799 15260
rect 34799 15204 34855 15260
rect 34855 15204 34859 15260
rect 34795 15200 34859 15204
rect 34875 15260 34939 15264
rect 34875 15204 34879 15260
rect 34879 15204 34935 15260
rect 34935 15204 34939 15260
rect 34875 15200 34939 15204
rect 34955 15260 35019 15264
rect 34955 15204 34959 15260
rect 34959 15204 35015 15260
rect 35015 15204 35019 15260
rect 34955 15200 35019 15204
rect 5172 14716 5236 14720
rect 5172 14660 5176 14716
rect 5176 14660 5232 14716
rect 5232 14660 5236 14716
rect 5172 14656 5236 14660
rect 5252 14716 5316 14720
rect 5252 14660 5256 14716
rect 5256 14660 5312 14716
rect 5312 14660 5316 14716
rect 5252 14656 5316 14660
rect 5332 14716 5396 14720
rect 5332 14660 5336 14716
rect 5336 14660 5392 14716
rect 5392 14660 5396 14716
rect 5332 14656 5396 14660
rect 5412 14716 5476 14720
rect 5412 14660 5416 14716
rect 5416 14660 5472 14716
rect 5472 14660 5476 14716
rect 5412 14656 5476 14660
rect 13613 14716 13677 14720
rect 13613 14660 13617 14716
rect 13617 14660 13673 14716
rect 13673 14660 13677 14716
rect 13613 14656 13677 14660
rect 13693 14716 13757 14720
rect 13693 14660 13697 14716
rect 13697 14660 13753 14716
rect 13753 14660 13757 14716
rect 13693 14656 13757 14660
rect 13773 14716 13837 14720
rect 13773 14660 13777 14716
rect 13777 14660 13833 14716
rect 13833 14660 13837 14716
rect 13773 14656 13837 14660
rect 13853 14716 13917 14720
rect 13853 14660 13857 14716
rect 13857 14660 13913 14716
rect 13913 14660 13917 14716
rect 13853 14656 13917 14660
rect 22054 14716 22118 14720
rect 22054 14660 22058 14716
rect 22058 14660 22114 14716
rect 22114 14660 22118 14716
rect 22054 14656 22118 14660
rect 22134 14716 22198 14720
rect 22134 14660 22138 14716
rect 22138 14660 22194 14716
rect 22194 14660 22198 14716
rect 22134 14656 22198 14660
rect 22214 14716 22278 14720
rect 22214 14660 22218 14716
rect 22218 14660 22274 14716
rect 22274 14660 22278 14716
rect 22214 14656 22278 14660
rect 22294 14716 22358 14720
rect 22294 14660 22298 14716
rect 22298 14660 22354 14716
rect 22354 14660 22358 14716
rect 22294 14656 22358 14660
rect 30495 14716 30559 14720
rect 30495 14660 30499 14716
rect 30499 14660 30555 14716
rect 30555 14660 30559 14716
rect 30495 14656 30559 14660
rect 30575 14716 30639 14720
rect 30575 14660 30579 14716
rect 30579 14660 30635 14716
rect 30635 14660 30639 14716
rect 30575 14656 30639 14660
rect 30655 14716 30719 14720
rect 30655 14660 30659 14716
rect 30659 14660 30715 14716
rect 30715 14660 30719 14716
rect 30655 14656 30719 14660
rect 30735 14716 30799 14720
rect 30735 14660 30739 14716
rect 30739 14660 30795 14716
rect 30795 14660 30799 14716
rect 30735 14656 30799 14660
rect 9392 14172 9456 14176
rect 9392 14116 9396 14172
rect 9396 14116 9452 14172
rect 9452 14116 9456 14172
rect 9392 14112 9456 14116
rect 9472 14172 9536 14176
rect 9472 14116 9476 14172
rect 9476 14116 9532 14172
rect 9532 14116 9536 14172
rect 9472 14112 9536 14116
rect 9552 14172 9616 14176
rect 9552 14116 9556 14172
rect 9556 14116 9612 14172
rect 9612 14116 9616 14172
rect 9552 14112 9616 14116
rect 9632 14172 9696 14176
rect 9632 14116 9636 14172
rect 9636 14116 9692 14172
rect 9692 14116 9696 14172
rect 9632 14112 9696 14116
rect 17833 14172 17897 14176
rect 17833 14116 17837 14172
rect 17837 14116 17893 14172
rect 17893 14116 17897 14172
rect 17833 14112 17897 14116
rect 17913 14172 17977 14176
rect 17913 14116 17917 14172
rect 17917 14116 17973 14172
rect 17973 14116 17977 14172
rect 17913 14112 17977 14116
rect 17993 14172 18057 14176
rect 17993 14116 17997 14172
rect 17997 14116 18053 14172
rect 18053 14116 18057 14172
rect 17993 14112 18057 14116
rect 18073 14172 18137 14176
rect 18073 14116 18077 14172
rect 18077 14116 18133 14172
rect 18133 14116 18137 14172
rect 18073 14112 18137 14116
rect 26274 14172 26338 14176
rect 26274 14116 26278 14172
rect 26278 14116 26334 14172
rect 26334 14116 26338 14172
rect 26274 14112 26338 14116
rect 26354 14172 26418 14176
rect 26354 14116 26358 14172
rect 26358 14116 26414 14172
rect 26414 14116 26418 14172
rect 26354 14112 26418 14116
rect 26434 14172 26498 14176
rect 26434 14116 26438 14172
rect 26438 14116 26494 14172
rect 26494 14116 26498 14172
rect 26434 14112 26498 14116
rect 26514 14172 26578 14176
rect 26514 14116 26518 14172
rect 26518 14116 26574 14172
rect 26574 14116 26578 14172
rect 26514 14112 26578 14116
rect 34715 14172 34779 14176
rect 34715 14116 34719 14172
rect 34719 14116 34775 14172
rect 34775 14116 34779 14172
rect 34715 14112 34779 14116
rect 34795 14172 34859 14176
rect 34795 14116 34799 14172
rect 34799 14116 34855 14172
rect 34855 14116 34859 14172
rect 34795 14112 34859 14116
rect 34875 14172 34939 14176
rect 34875 14116 34879 14172
rect 34879 14116 34935 14172
rect 34935 14116 34939 14172
rect 34875 14112 34939 14116
rect 34955 14172 35019 14176
rect 34955 14116 34959 14172
rect 34959 14116 35015 14172
rect 35015 14116 35019 14172
rect 34955 14112 35019 14116
rect 5172 13628 5236 13632
rect 5172 13572 5176 13628
rect 5176 13572 5232 13628
rect 5232 13572 5236 13628
rect 5172 13568 5236 13572
rect 5252 13628 5316 13632
rect 5252 13572 5256 13628
rect 5256 13572 5312 13628
rect 5312 13572 5316 13628
rect 5252 13568 5316 13572
rect 5332 13628 5396 13632
rect 5332 13572 5336 13628
rect 5336 13572 5392 13628
rect 5392 13572 5396 13628
rect 5332 13568 5396 13572
rect 5412 13628 5476 13632
rect 5412 13572 5416 13628
rect 5416 13572 5472 13628
rect 5472 13572 5476 13628
rect 5412 13568 5476 13572
rect 13613 13628 13677 13632
rect 13613 13572 13617 13628
rect 13617 13572 13673 13628
rect 13673 13572 13677 13628
rect 13613 13568 13677 13572
rect 13693 13628 13757 13632
rect 13693 13572 13697 13628
rect 13697 13572 13753 13628
rect 13753 13572 13757 13628
rect 13693 13568 13757 13572
rect 13773 13628 13837 13632
rect 13773 13572 13777 13628
rect 13777 13572 13833 13628
rect 13833 13572 13837 13628
rect 13773 13568 13837 13572
rect 13853 13628 13917 13632
rect 13853 13572 13857 13628
rect 13857 13572 13913 13628
rect 13913 13572 13917 13628
rect 13853 13568 13917 13572
rect 22054 13628 22118 13632
rect 22054 13572 22058 13628
rect 22058 13572 22114 13628
rect 22114 13572 22118 13628
rect 22054 13568 22118 13572
rect 22134 13628 22198 13632
rect 22134 13572 22138 13628
rect 22138 13572 22194 13628
rect 22194 13572 22198 13628
rect 22134 13568 22198 13572
rect 22214 13628 22278 13632
rect 22214 13572 22218 13628
rect 22218 13572 22274 13628
rect 22274 13572 22278 13628
rect 22214 13568 22278 13572
rect 22294 13628 22358 13632
rect 22294 13572 22298 13628
rect 22298 13572 22354 13628
rect 22354 13572 22358 13628
rect 22294 13568 22358 13572
rect 30495 13628 30559 13632
rect 30495 13572 30499 13628
rect 30499 13572 30555 13628
rect 30555 13572 30559 13628
rect 30495 13568 30559 13572
rect 30575 13628 30639 13632
rect 30575 13572 30579 13628
rect 30579 13572 30635 13628
rect 30635 13572 30639 13628
rect 30575 13568 30639 13572
rect 30655 13628 30719 13632
rect 30655 13572 30659 13628
rect 30659 13572 30715 13628
rect 30715 13572 30719 13628
rect 30655 13568 30719 13572
rect 30735 13628 30799 13632
rect 30735 13572 30739 13628
rect 30739 13572 30795 13628
rect 30795 13572 30799 13628
rect 30735 13568 30799 13572
rect 9392 13084 9456 13088
rect 9392 13028 9396 13084
rect 9396 13028 9452 13084
rect 9452 13028 9456 13084
rect 9392 13024 9456 13028
rect 9472 13084 9536 13088
rect 9472 13028 9476 13084
rect 9476 13028 9532 13084
rect 9532 13028 9536 13084
rect 9472 13024 9536 13028
rect 9552 13084 9616 13088
rect 9552 13028 9556 13084
rect 9556 13028 9612 13084
rect 9612 13028 9616 13084
rect 9552 13024 9616 13028
rect 9632 13084 9696 13088
rect 9632 13028 9636 13084
rect 9636 13028 9692 13084
rect 9692 13028 9696 13084
rect 9632 13024 9696 13028
rect 17833 13084 17897 13088
rect 17833 13028 17837 13084
rect 17837 13028 17893 13084
rect 17893 13028 17897 13084
rect 17833 13024 17897 13028
rect 17913 13084 17977 13088
rect 17913 13028 17917 13084
rect 17917 13028 17973 13084
rect 17973 13028 17977 13084
rect 17913 13024 17977 13028
rect 17993 13084 18057 13088
rect 17993 13028 17997 13084
rect 17997 13028 18053 13084
rect 18053 13028 18057 13084
rect 17993 13024 18057 13028
rect 18073 13084 18137 13088
rect 18073 13028 18077 13084
rect 18077 13028 18133 13084
rect 18133 13028 18137 13084
rect 18073 13024 18137 13028
rect 26274 13084 26338 13088
rect 26274 13028 26278 13084
rect 26278 13028 26334 13084
rect 26334 13028 26338 13084
rect 26274 13024 26338 13028
rect 26354 13084 26418 13088
rect 26354 13028 26358 13084
rect 26358 13028 26414 13084
rect 26414 13028 26418 13084
rect 26354 13024 26418 13028
rect 26434 13084 26498 13088
rect 26434 13028 26438 13084
rect 26438 13028 26494 13084
rect 26494 13028 26498 13084
rect 26434 13024 26498 13028
rect 26514 13084 26578 13088
rect 26514 13028 26518 13084
rect 26518 13028 26574 13084
rect 26574 13028 26578 13084
rect 26514 13024 26578 13028
rect 34715 13084 34779 13088
rect 34715 13028 34719 13084
rect 34719 13028 34775 13084
rect 34775 13028 34779 13084
rect 34715 13024 34779 13028
rect 34795 13084 34859 13088
rect 34795 13028 34799 13084
rect 34799 13028 34855 13084
rect 34855 13028 34859 13084
rect 34795 13024 34859 13028
rect 34875 13084 34939 13088
rect 34875 13028 34879 13084
rect 34879 13028 34935 13084
rect 34935 13028 34939 13084
rect 34875 13024 34939 13028
rect 34955 13084 35019 13088
rect 34955 13028 34959 13084
rect 34959 13028 35015 13084
rect 35015 13028 35019 13084
rect 34955 13024 35019 13028
rect 5172 12540 5236 12544
rect 5172 12484 5176 12540
rect 5176 12484 5232 12540
rect 5232 12484 5236 12540
rect 5172 12480 5236 12484
rect 5252 12540 5316 12544
rect 5252 12484 5256 12540
rect 5256 12484 5312 12540
rect 5312 12484 5316 12540
rect 5252 12480 5316 12484
rect 5332 12540 5396 12544
rect 5332 12484 5336 12540
rect 5336 12484 5392 12540
rect 5392 12484 5396 12540
rect 5332 12480 5396 12484
rect 5412 12540 5476 12544
rect 5412 12484 5416 12540
rect 5416 12484 5472 12540
rect 5472 12484 5476 12540
rect 5412 12480 5476 12484
rect 13613 12540 13677 12544
rect 13613 12484 13617 12540
rect 13617 12484 13673 12540
rect 13673 12484 13677 12540
rect 13613 12480 13677 12484
rect 13693 12540 13757 12544
rect 13693 12484 13697 12540
rect 13697 12484 13753 12540
rect 13753 12484 13757 12540
rect 13693 12480 13757 12484
rect 13773 12540 13837 12544
rect 13773 12484 13777 12540
rect 13777 12484 13833 12540
rect 13833 12484 13837 12540
rect 13773 12480 13837 12484
rect 13853 12540 13917 12544
rect 13853 12484 13857 12540
rect 13857 12484 13913 12540
rect 13913 12484 13917 12540
rect 13853 12480 13917 12484
rect 22054 12540 22118 12544
rect 22054 12484 22058 12540
rect 22058 12484 22114 12540
rect 22114 12484 22118 12540
rect 22054 12480 22118 12484
rect 22134 12540 22198 12544
rect 22134 12484 22138 12540
rect 22138 12484 22194 12540
rect 22194 12484 22198 12540
rect 22134 12480 22198 12484
rect 22214 12540 22278 12544
rect 22214 12484 22218 12540
rect 22218 12484 22274 12540
rect 22274 12484 22278 12540
rect 22214 12480 22278 12484
rect 22294 12540 22358 12544
rect 22294 12484 22298 12540
rect 22298 12484 22354 12540
rect 22354 12484 22358 12540
rect 22294 12480 22358 12484
rect 30495 12540 30559 12544
rect 30495 12484 30499 12540
rect 30499 12484 30555 12540
rect 30555 12484 30559 12540
rect 30495 12480 30559 12484
rect 30575 12540 30639 12544
rect 30575 12484 30579 12540
rect 30579 12484 30635 12540
rect 30635 12484 30639 12540
rect 30575 12480 30639 12484
rect 30655 12540 30719 12544
rect 30655 12484 30659 12540
rect 30659 12484 30715 12540
rect 30715 12484 30719 12540
rect 30655 12480 30719 12484
rect 30735 12540 30799 12544
rect 30735 12484 30739 12540
rect 30739 12484 30795 12540
rect 30795 12484 30799 12540
rect 30735 12480 30799 12484
rect 9392 11996 9456 12000
rect 9392 11940 9396 11996
rect 9396 11940 9452 11996
rect 9452 11940 9456 11996
rect 9392 11936 9456 11940
rect 9472 11996 9536 12000
rect 9472 11940 9476 11996
rect 9476 11940 9532 11996
rect 9532 11940 9536 11996
rect 9472 11936 9536 11940
rect 9552 11996 9616 12000
rect 9552 11940 9556 11996
rect 9556 11940 9612 11996
rect 9612 11940 9616 11996
rect 9552 11936 9616 11940
rect 9632 11996 9696 12000
rect 9632 11940 9636 11996
rect 9636 11940 9692 11996
rect 9692 11940 9696 11996
rect 9632 11936 9696 11940
rect 17833 11996 17897 12000
rect 17833 11940 17837 11996
rect 17837 11940 17893 11996
rect 17893 11940 17897 11996
rect 17833 11936 17897 11940
rect 17913 11996 17977 12000
rect 17913 11940 17917 11996
rect 17917 11940 17973 11996
rect 17973 11940 17977 11996
rect 17913 11936 17977 11940
rect 17993 11996 18057 12000
rect 17993 11940 17997 11996
rect 17997 11940 18053 11996
rect 18053 11940 18057 11996
rect 17993 11936 18057 11940
rect 18073 11996 18137 12000
rect 18073 11940 18077 11996
rect 18077 11940 18133 11996
rect 18133 11940 18137 11996
rect 18073 11936 18137 11940
rect 26274 11996 26338 12000
rect 26274 11940 26278 11996
rect 26278 11940 26334 11996
rect 26334 11940 26338 11996
rect 26274 11936 26338 11940
rect 26354 11996 26418 12000
rect 26354 11940 26358 11996
rect 26358 11940 26414 11996
rect 26414 11940 26418 11996
rect 26354 11936 26418 11940
rect 26434 11996 26498 12000
rect 26434 11940 26438 11996
rect 26438 11940 26494 11996
rect 26494 11940 26498 11996
rect 26434 11936 26498 11940
rect 26514 11996 26578 12000
rect 26514 11940 26518 11996
rect 26518 11940 26574 11996
rect 26574 11940 26578 11996
rect 26514 11936 26578 11940
rect 34715 11996 34779 12000
rect 34715 11940 34719 11996
rect 34719 11940 34775 11996
rect 34775 11940 34779 11996
rect 34715 11936 34779 11940
rect 34795 11996 34859 12000
rect 34795 11940 34799 11996
rect 34799 11940 34855 11996
rect 34855 11940 34859 11996
rect 34795 11936 34859 11940
rect 34875 11996 34939 12000
rect 34875 11940 34879 11996
rect 34879 11940 34935 11996
rect 34935 11940 34939 11996
rect 34875 11936 34939 11940
rect 34955 11996 35019 12000
rect 34955 11940 34959 11996
rect 34959 11940 35015 11996
rect 35015 11940 35019 11996
rect 34955 11936 35019 11940
rect 5172 11452 5236 11456
rect 5172 11396 5176 11452
rect 5176 11396 5232 11452
rect 5232 11396 5236 11452
rect 5172 11392 5236 11396
rect 5252 11452 5316 11456
rect 5252 11396 5256 11452
rect 5256 11396 5312 11452
rect 5312 11396 5316 11452
rect 5252 11392 5316 11396
rect 5332 11452 5396 11456
rect 5332 11396 5336 11452
rect 5336 11396 5392 11452
rect 5392 11396 5396 11452
rect 5332 11392 5396 11396
rect 5412 11452 5476 11456
rect 5412 11396 5416 11452
rect 5416 11396 5472 11452
rect 5472 11396 5476 11452
rect 5412 11392 5476 11396
rect 13613 11452 13677 11456
rect 13613 11396 13617 11452
rect 13617 11396 13673 11452
rect 13673 11396 13677 11452
rect 13613 11392 13677 11396
rect 13693 11452 13757 11456
rect 13693 11396 13697 11452
rect 13697 11396 13753 11452
rect 13753 11396 13757 11452
rect 13693 11392 13757 11396
rect 13773 11452 13837 11456
rect 13773 11396 13777 11452
rect 13777 11396 13833 11452
rect 13833 11396 13837 11452
rect 13773 11392 13837 11396
rect 13853 11452 13917 11456
rect 13853 11396 13857 11452
rect 13857 11396 13913 11452
rect 13913 11396 13917 11452
rect 13853 11392 13917 11396
rect 22054 11452 22118 11456
rect 22054 11396 22058 11452
rect 22058 11396 22114 11452
rect 22114 11396 22118 11452
rect 22054 11392 22118 11396
rect 22134 11452 22198 11456
rect 22134 11396 22138 11452
rect 22138 11396 22194 11452
rect 22194 11396 22198 11452
rect 22134 11392 22198 11396
rect 22214 11452 22278 11456
rect 22214 11396 22218 11452
rect 22218 11396 22274 11452
rect 22274 11396 22278 11452
rect 22214 11392 22278 11396
rect 22294 11452 22358 11456
rect 22294 11396 22298 11452
rect 22298 11396 22354 11452
rect 22354 11396 22358 11452
rect 22294 11392 22358 11396
rect 30495 11452 30559 11456
rect 30495 11396 30499 11452
rect 30499 11396 30555 11452
rect 30555 11396 30559 11452
rect 30495 11392 30559 11396
rect 30575 11452 30639 11456
rect 30575 11396 30579 11452
rect 30579 11396 30635 11452
rect 30635 11396 30639 11452
rect 30575 11392 30639 11396
rect 30655 11452 30719 11456
rect 30655 11396 30659 11452
rect 30659 11396 30715 11452
rect 30715 11396 30719 11452
rect 30655 11392 30719 11396
rect 30735 11452 30799 11456
rect 30735 11396 30739 11452
rect 30739 11396 30795 11452
rect 30795 11396 30799 11452
rect 30735 11392 30799 11396
rect 9392 10908 9456 10912
rect 9392 10852 9396 10908
rect 9396 10852 9452 10908
rect 9452 10852 9456 10908
rect 9392 10848 9456 10852
rect 9472 10908 9536 10912
rect 9472 10852 9476 10908
rect 9476 10852 9532 10908
rect 9532 10852 9536 10908
rect 9472 10848 9536 10852
rect 9552 10908 9616 10912
rect 9552 10852 9556 10908
rect 9556 10852 9612 10908
rect 9612 10852 9616 10908
rect 9552 10848 9616 10852
rect 9632 10908 9696 10912
rect 9632 10852 9636 10908
rect 9636 10852 9692 10908
rect 9692 10852 9696 10908
rect 9632 10848 9696 10852
rect 17833 10908 17897 10912
rect 17833 10852 17837 10908
rect 17837 10852 17893 10908
rect 17893 10852 17897 10908
rect 17833 10848 17897 10852
rect 17913 10908 17977 10912
rect 17913 10852 17917 10908
rect 17917 10852 17973 10908
rect 17973 10852 17977 10908
rect 17913 10848 17977 10852
rect 17993 10908 18057 10912
rect 17993 10852 17997 10908
rect 17997 10852 18053 10908
rect 18053 10852 18057 10908
rect 17993 10848 18057 10852
rect 18073 10908 18137 10912
rect 18073 10852 18077 10908
rect 18077 10852 18133 10908
rect 18133 10852 18137 10908
rect 18073 10848 18137 10852
rect 26274 10908 26338 10912
rect 26274 10852 26278 10908
rect 26278 10852 26334 10908
rect 26334 10852 26338 10908
rect 26274 10848 26338 10852
rect 26354 10908 26418 10912
rect 26354 10852 26358 10908
rect 26358 10852 26414 10908
rect 26414 10852 26418 10908
rect 26354 10848 26418 10852
rect 26434 10908 26498 10912
rect 26434 10852 26438 10908
rect 26438 10852 26494 10908
rect 26494 10852 26498 10908
rect 26434 10848 26498 10852
rect 26514 10908 26578 10912
rect 26514 10852 26518 10908
rect 26518 10852 26574 10908
rect 26574 10852 26578 10908
rect 26514 10848 26578 10852
rect 34715 10908 34779 10912
rect 34715 10852 34719 10908
rect 34719 10852 34775 10908
rect 34775 10852 34779 10908
rect 34715 10848 34779 10852
rect 34795 10908 34859 10912
rect 34795 10852 34799 10908
rect 34799 10852 34855 10908
rect 34855 10852 34859 10908
rect 34795 10848 34859 10852
rect 34875 10908 34939 10912
rect 34875 10852 34879 10908
rect 34879 10852 34935 10908
rect 34935 10852 34939 10908
rect 34875 10848 34939 10852
rect 34955 10908 35019 10912
rect 34955 10852 34959 10908
rect 34959 10852 35015 10908
rect 35015 10852 35019 10908
rect 34955 10848 35019 10852
rect 5172 10364 5236 10368
rect 5172 10308 5176 10364
rect 5176 10308 5232 10364
rect 5232 10308 5236 10364
rect 5172 10304 5236 10308
rect 5252 10364 5316 10368
rect 5252 10308 5256 10364
rect 5256 10308 5312 10364
rect 5312 10308 5316 10364
rect 5252 10304 5316 10308
rect 5332 10364 5396 10368
rect 5332 10308 5336 10364
rect 5336 10308 5392 10364
rect 5392 10308 5396 10364
rect 5332 10304 5396 10308
rect 5412 10364 5476 10368
rect 5412 10308 5416 10364
rect 5416 10308 5472 10364
rect 5472 10308 5476 10364
rect 5412 10304 5476 10308
rect 13613 10364 13677 10368
rect 13613 10308 13617 10364
rect 13617 10308 13673 10364
rect 13673 10308 13677 10364
rect 13613 10304 13677 10308
rect 13693 10364 13757 10368
rect 13693 10308 13697 10364
rect 13697 10308 13753 10364
rect 13753 10308 13757 10364
rect 13693 10304 13757 10308
rect 13773 10364 13837 10368
rect 13773 10308 13777 10364
rect 13777 10308 13833 10364
rect 13833 10308 13837 10364
rect 13773 10304 13837 10308
rect 13853 10364 13917 10368
rect 13853 10308 13857 10364
rect 13857 10308 13913 10364
rect 13913 10308 13917 10364
rect 13853 10304 13917 10308
rect 22054 10364 22118 10368
rect 22054 10308 22058 10364
rect 22058 10308 22114 10364
rect 22114 10308 22118 10364
rect 22054 10304 22118 10308
rect 22134 10364 22198 10368
rect 22134 10308 22138 10364
rect 22138 10308 22194 10364
rect 22194 10308 22198 10364
rect 22134 10304 22198 10308
rect 22214 10364 22278 10368
rect 22214 10308 22218 10364
rect 22218 10308 22274 10364
rect 22274 10308 22278 10364
rect 22214 10304 22278 10308
rect 22294 10364 22358 10368
rect 22294 10308 22298 10364
rect 22298 10308 22354 10364
rect 22354 10308 22358 10364
rect 22294 10304 22358 10308
rect 30495 10364 30559 10368
rect 30495 10308 30499 10364
rect 30499 10308 30555 10364
rect 30555 10308 30559 10364
rect 30495 10304 30559 10308
rect 30575 10364 30639 10368
rect 30575 10308 30579 10364
rect 30579 10308 30635 10364
rect 30635 10308 30639 10364
rect 30575 10304 30639 10308
rect 30655 10364 30719 10368
rect 30655 10308 30659 10364
rect 30659 10308 30715 10364
rect 30715 10308 30719 10364
rect 30655 10304 30719 10308
rect 30735 10364 30799 10368
rect 30735 10308 30739 10364
rect 30739 10308 30795 10364
rect 30795 10308 30799 10364
rect 30735 10304 30799 10308
rect 9392 9820 9456 9824
rect 9392 9764 9396 9820
rect 9396 9764 9452 9820
rect 9452 9764 9456 9820
rect 9392 9760 9456 9764
rect 9472 9820 9536 9824
rect 9472 9764 9476 9820
rect 9476 9764 9532 9820
rect 9532 9764 9536 9820
rect 9472 9760 9536 9764
rect 9552 9820 9616 9824
rect 9552 9764 9556 9820
rect 9556 9764 9612 9820
rect 9612 9764 9616 9820
rect 9552 9760 9616 9764
rect 9632 9820 9696 9824
rect 9632 9764 9636 9820
rect 9636 9764 9692 9820
rect 9692 9764 9696 9820
rect 9632 9760 9696 9764
rect 17833 9820 17897 9824
rect 17833 9764 17837 9820
rect 17837 9764 17893 9820
rect 17893 9764 17897 9820
rect 17833 9760 17897 9764
rect 17913 9820 17977 9824
rect 17913 9764 17917 9820
rect 17917 9764 17973 9820
rect 17973 9764 17977 9820
rect 17913 9760 17977 9764
rect 17993 9820 18057 9824
rect 17993 9764 17997 9820
rect 17997 9764 18053 9820
rect 18053 9764 18057 9820
rect 17993 9760 18057 9764
rect 18073 9820 18137 9824
rect 18073 9764 18077 9820
rect 18077 9764 18133 9820
rect 18133 9764 18137 9820
rect 18073 9760 18137 9764
rect 26274 9820 26338 9824
rect 26274 9764 26278 9820
rect 26278 9764 26334 9820
rect 26334 9764 26338 9820
rect 26274 9760 26338 9764
rect 26354 9820 26418 9824
rect 26354 9764 26358 9820
rect 26358 9764 26414 9820
rect 26414 9764 26418 9820
rect 26354 9760 26418 9764
rect 26434 9820 26498 9824
rect 26434 9764 26438 9820
rect 26438 9764 26494 9820
rect 26494 9764 26498 9820
rect 26434 9760 26498 9764
rect 26514 9820 26578 9824
rect 26514 9764 26518 9820
rect 26518 9764 26574 9820
rect 26574 9764 26578 9820
rect 26514 9760 26578 9764
rect 34715 9820 34779 9824
rect 34715 9764 34719 9820
rect 34719 9764 34775 9820
rect 34775 9764 34779 9820
rect 34715 9760 34779 9764
rect 34795 9820 34859 9824
rect 34795 9764 34799 9820
rect 34799 9764 34855 9820
rect 34855 9764 34859 9820
rect 34795 9760 34859 9764
rect 34875 9820 34939 9824
rect 34875 9764 34879 9820
rect 34879 9764 34935 9820
rect 34935 9764 34939 9820
rect 34875 9760 34939 9764
rect 34955 9820 35019 9824
rect 34955 9764 34959 9820
rect 34959 9764 35015 9820
rect 35015 9764 35019 9820
rect 34955 9760 35019 9764
rect 5172 9276 5236 9280
rect 5172 9220 5176 9276
rect 5176 9220 5232 9276
rect 5232 9220 5236 9276
rect 5172 9216 5236 9220
rect 5252 9276 5316 9280
rect 5252 9220 5256 9276
rect 5256 9220 5312 9276
rect 5312 9220 5316 9276
rect 5252 9216 5316 9220
rect 5332 9276 5396 9280
rect 5332 9220 5336 9276
rect 5336 9220 5392 9276
rect 5392 9220 5396 9276
rect 5332 9216 5396 9220
rect 5412 9276 5476 9280
rect 5412 9220 5416 9276
rect 5416 9220 5472 9276
rect 5472 9220 5476 9276
rect 5412 9216 5476 9220
rect 13613 9276 13677 9280
rect 13613 9220 13617 9276
rect 13617 9220 13673 9276
rect 13673 9220 13677 9276
rect 13613 9216 13677 9220
rect 13693 9276 13757 9280
rect 13693 9220 13697 9276
rect 13697 9220 13753 9276
rect 13753 9220 13757 9276
rect 13693 9216 13757 9220
rect 13773 9276 13837 9280
rect 13773 9220 13777 9276
rect 13777 9220 13833 9276
rect 13833 9220 13837 9276
rect 13773 9216 13837 9220
rect 13853 9276 13917 9280
rect 13853 9220 13857 9276
rect 13857 9220 13913 9276
rect 13913 9220 13917 9276
rect 13853 9216 13917 9220
rect 22054 9276 22118 9280
rect 22054 9220 22058 9276
rect 22058 9220 22114 9276
rect 22114 9220 22118 9276
rect 22054 9216 22118 9220
rect 22134 9276 22198 9280
rect 22134 9220 22138 9276
rect 22138 9220 22194 9276
rect 22194 9220 22198 9276
rect 22134 9216 22198 9220
rect 22214 9276 22278 9280
rect 22214 9220 22218 9276
rect 22218 9220 22274 9276
rect 22274 9220 22278 9276
rect 22214 9216 22278 9220
rect 22294 9276 22358 9280
rect 22294 9220 22298 9276
rect 22298 9220 22354 9276
rect 22354 9220 22358 9276
rect 22294 9216 22358 9220
rect 30495 9276 30559 9280
rect 30495 9220 30499 9276
rect 30499 9220 30555 9276
rect 30555 9220 30559 9276
rect 30495 9216 30559 9220
rect 30575 9276 30639 9280
rect 30575 9220 30579 9276
rect 30579 9220 30635 9276
rect 30635 9220 30639 9276
rect 30575 9216 30639 9220
rect 30655 9276 30719 9280
rect 30655 9220 30659 9276
rect 30659 9220 30715 9276
rect 30715 9220 30719 9276
rect 30655 9216 30719 9220
rect 30735 9276 30799 9280
rect 30735 9220 30739 9276
rect 30739 9220 30795 9276
rect 30795 9220 30799 9276
rect 30735 9216 30799 9220
rect 9392 8732 9456 8736
rect 9392 8676 9396 8732
rect 9396 8676 9452 8732
rect 9452 8676 9456 8732
rect 9392 8672 9456 8676
rect 9472 8732 9536 8736
rect 9472 8676 9476 8732
rect 9476 8676 9532 8732
rect 9532 8676 9536 8732
rect 9472 8672 9536 8676
rect 9552 8732 9616 8736
rect 9552 8676 9556 8732
rect 9556 8676 9612 8732
rect 9612 8676 9616 8732
rect 9552 8672 9616 8676
rect 9632 8732 9696 8736
rect 9632 8676 9636 8732
rect 9636 8676 9692 8732
rect 9692 8676 9696 8732
rect 9632 8672 9696 8676
rect 17833 8732 17897 8736
rect 17833 8676 17837 8732
rect 17837 8676 17893 8732
rect 17893 8676 17897 8732
rect 17833 8672 17897 8676
rect 17913 8732 17977 8736
rect 17913 8676 17917 8732
rect 17917 8676 17973 8732
rect 17973 8676 17977 8732
rect 17913 8672 17977 8676
rect 17993 8732 18057 8736
rect 17993 8676 17997 8732
rect 17997 8676 18053 8732
rect 18053 8676 18057 8732
rect 17993 8672 18057 8676
rect 18073 8732 18137 8736
rect 18073 8676 18077 8732
rect 18077 8676 18133 8732
rect 18133 8676 18137 8732
rect 18073 8672 18137 8676
rect 26274 8732 26338 8736
rect 26274 8676 26278 8732
rect 26278 8676 26334 8732
rect 26334 8676 26338 8732
rect 26274 8672 26338 8676
rect 26354 8732 26418 8736
rect 26354 8676 26358 8732
rect 26358 8676 26414 8732
rect 26414 8676 26418 8732
rect 26354 8672 26418 8676
rect 26434 8732 26498 8736
rect 26434 8676 26438 8732
rect 26438 8676 26494 8732
rect 26494 8676 26498 8732
rect 26434 8672 26498 8676
rect 26514 8732 26578 8736
rect 26514 8676 26518 8732
rect 26518 8676 26574 8732
rect 26574 8676 26578 8732
rect 26514 8672 26578 8676
rect 34715 8732 34779 8736
rect 34715 8676 34719 8732
rect 34719 8676 34775 8732
rect 34775 8676 34779 8732
rect 34715 8672 34779 8676
rect 34795 8732 34859 8736
rect 34795 8676 34799 8732
rect 34799 8676 34855 8732
rect 34855 8676 34859 8732
rect 34795 8672 34859 8676
rect 34875 8732 34939 8736
rect 34875 8676 34879 8732
rect 34879 8676 34935 8732
rect 34935 8676 34939 8732
rect 34875 8672 34939 8676
rect 34955 8732 35019 8736
rect 34955 8676 34959 8732
rect 34959 8676 35015 8732
rect 35015 8676 35019 8732
rect 34955 8672 35019 8676
rect 5172 8188 5236 8192
rect 5172 8132 5176 8188
rect 5176 8132 5232 8188
rect 5232 8132 5236 8188
rect 5172 8128 5236 8132
rect 5252 8188 5316 8192
rect 5252 8132 5256 8188
rect 5256 8132 5312 8188
rect 5312 8132 5316 8188
rect 5252 8128 5316 8132
rect 5332 8188 5396 8192
rect 5332 8132 5336 8188
rect 5336 8132 5392 8188
rect 5392 8132 5396 8188
rect 5332 8128 5396 8132
rect 5412 8188 5476 8192
rect 5412 8132 5416 8188
rect 5416 8132 5472 8188
rect 5472 8132 5476 8188
rect 5412 8128 5476 8132
rect 13613 8188 13677 8192
rect 13613 8132 13617 8188
rect 13617 8132 13673 8188
rect 13673 8132 13677 8188
rect 13613 8128 13677 8132
rect 13693 8188 13757 8192
rect 13693 8132 13697 8188
rect 13697 8132 13753 8188
rect 13753 8132 13757 8188
rect 13693 8128 13757 8132
rect 13773 8188 13837 8192
rect 13773 8132 13777 8188
rect 13777 8132 13833 8188
rect 13833 8132 13837 8188
rect 13773 8128 13837 8132
rect 13853 8188 13917 8192
rect 13853 8132 13857 8188
rect 13857 8132 13913 8188
rect 13913 8132 13917 8188
rect 13853 8128 13917 8132
rect 22054 8188 22118 8192
rect 22054 8132 22058 8188
rect 22058 8132 22114 8188
rect 22114 8132 22118 8188
rect 22054 8128 22118 8132
rect 22134 8188 22198 8192
rect 22134 8132 22138 8188
rect 22138 8132 22194 8188
rect 22194 8132 22198 8188
rect 22134 8128 22198 8132
rect 22214 8188 22278 8192
rect 22214 8132 22218 8188
rect 22218 8132 22274 8188
rect 22274 8132 22278 8188
rect 22214 8128 22278 8132
rect 22294 8188 22358 8192
rect 22294 8132 22298 8188
rect 22298 8132 22354 8188
rect 22354 8132 22358 8188
rect 22294 8128 22358 8132
rect 30495 8188 30559 8192
rect 30495 8132 30499 8188
rect 30499 8132 30555 8188
rect 30555 8132 30559 8188
rect 30495 8128 30559 8132
rect 30575 8188 30639 8192
rect 30575 8132 30579 8188
rect 30579 8132 30635 8188
rect 30635 8132 30639 8188
rect 30575 8128 30639 8132
rect 30655 8188 30719 8192
rect 30655 8132 30659 8188
rect 30659 8132 30715 8188
rect 30715 8132 30719 8188
rect 30655 8128 30719 8132
rect 30735 8188 30799 8192
rect 30735 8132 30739 8188
rect 30739 8132 30795 8188
rect 30795 8132 30799 8188
rect 30735 8128 30799 8132
rect 9392 7644 9456 7648
rect 9392 7588 9396 7644
rect 9396 7588 9452 7644
rect 9452 7588 9456 7644
rect 9392 7584 9456 7588
rect 9472 7644 9536 7648
rect 9472 7588 9476 7644
rect 9476 7588 9532 7644
rect 9532 7588 9536 7644
rect 9472 7584 9536 7588
rect 9552 7644 9616 7648
rect 9552 7588 9556 7644
rect 9556 7588 9612 7644
rect 9612 7588 9616 7644
rect 9552 7584 9616 7588
rect 9632 7644 9696 7648
rect 9632 7588 9636 7644
rect 9636 7588 9692 7644
rect 9692 7588 9696 7644
rect 9632 7584 9696 7588
rect 17833 7644 17897 7648
rect 17833 7588 17837 7644
rect 17837 7588 17893 7644
rect 17893 7588 17897 7644
rect 17833 7584 17897 7588
rect 17913 7644 17977 7648
rect 17913 7588 17917 7644
rect 17917 7588 17973 7644
rect 17973 7588 17977 7644
rect 17913 7584 17977 7588
rect 17993 7644 18057 7648
rect 17993 7588 17997 7644
rect 17997 7588 18053 7644
rect 18053 7588 18057 7644
rect 17993 7584 18057 7588
rect 18073 7644 18137 7648
rect 18073 7588 18077 7644
rect 18077 7588 18133 7644
rect 18133 7588 18137 7644
rect 18073 7584 18137 7588
rect 26274 7644 26338 7648
rect 26274 7588 26278 7644
rect 26278 7588 26334 7644
rect 26334 7588 26338 7644
rect 26274 7584 26338 7588
rect 26354 7644 26418 7648
rect 26354 7588 26358 7644
rect 26358 7588 26414 7644
rect 26414 7588 26418 7644
rect 26354 7584 26418 7588
rect 26434 7644 26498 7648
rect 26434 7588 26438 7644
rect 26438 7588 26494 7644
rect 26494 7588 26498 7644
rect 26434 7584 26498 7588
rect 26514 7644 26578 7648
rect 26514 7588 26518 7644
rect 26518 7588 26574 7644
rect 26574 7588 26578 7644
rect 26514 7584 26578 7588
rect 34715 7644 34779 7648
rect 34715 7588 34719 7644
rect 34719 7588 34775 7644
rect 34775 7588 34779 7644
rect 34715 7584 34779 7588
rect 34795 7644 34859 7648
rect 34795 7588 34799 7644
rect 34799 7588 34855 7644
rect 34855 7588 34859 7644
rect 34795 7584 34859 7588
rect 34875 7644 34939 7648
rect 34875 7588 34879 7644
rect 34879 7588 34935 7644
rect 34935 7588 34939 7644
rect 34875 7584 34939 7588
rect 34955 7644 35019 7648
rect 34955 7588 34959 7644
rect 34959 7588 35015 7644
rect 35015 7588 35019 7644
rect 34955 7584 35019 7588
rect 5172 7100 5236 7104
rect 5172 7044 5176 7100
rect 5176 7044 5232 7100
rect 5232 7044 5236 7100
rect 5172 7040 5236 7044
rect 5252 7100 5316 7104
rect 5252 7044 5256 7100
rect 5256 7044 5312 7100
rect 5312 7044 5316 7100
rect 5252 7040 5316 7044
rect 5332 7100 5396 7104
rect 5332 7044 5336 7100
rect 5336 7044 5392 7100
rect 5392 7044 5396 7100
rect 5332 7040 5396 7044
rect 5412 7100 5476 7104
rect 5412 7044 5416 7100
rect 5416 7044 5472 7100
rect 5472 7044 5476 7100
rect 5412 7040 5476 7044
rect 13613 7100 13677 7104
rect 13613 7044 13617 7100
rect 13617 7044 13673 7100
rect 13673 7044 13677 7100
rect 13613 7040 13677 7044
rect 13693 7100 13757 7104
rect 13693 7044 13697 7100
rect 13697 7044 13753 7100
rect 13753 7044 13757 7100
rect 13693 7040 13757 7044
rect 13773 7100 13837 7104
rect 13773 7044 13777 7100
rect 13777 7044 13833 7100
rect 13833 7044 13837 7100
rect 13773 7040 13837 7044
rect 13853 7100 13917 7104
rect 13853 7044 13857 7100
rect 13857 7044 13913 7100
rect 13913 7044 13917 7100
rect 13853 7040 13917 7044
rect 22054 7100 22118 7104
rect 22054 7044 22058 7100
rect 22058 7044 22114 7100
rect 22114 7044 22118 7100
rect 22054 7040 22118 7044
rect 22134 7100 22198 7104
rect 22134 7044 22138 7100
rect 22138 7044 22194 7100
rect 22194 7044 22198 7100
rect 22134 7040 22198 7044
rect 22214 7100 22278 7104
rect 22214 7044 22218 7100
rect 22218 7044 22274 7100
rect 22274 7044 22278 7100
rect 22214 7040 22278 7044
rect 22294 7100 22358 7104
rect 22294 7044 22298 7100
rect 22298 7044 22354 7100
rect 22354 7044 22358 7100
rect 22294 7040 22358 7044
rect 30495 7100 30559 7104
rect 30495 7044 30499 7100
rect 30499 7044 30555 7100
rect 30555 7044 30559 7100
rect 30495 7040 30559 7044
rect 30575 7100 30639 7104
rect 30575 7044 30579 7100
rect 30579 7044 30635 7100
rect 30635 7044 30639 7100
rect 30575 7040 30639 7044
rect 30655 7100 30719 7104
rect 30655 7044 30659 7100
rect 30659 7044 30715 7100
rect 30715 7044 30719 7100
rect 30655 7040 30719 7044
rect 30735 7100 30799 7104
rect 30735 7044 30739 7100
rect 30739 7044 30795 7100
rect 30795 7044 30799 7100
rect 30735 7040 30799 7044
rect 9392 6556 9456 6560
rect 9392 6500 9396 6556
rect 9396 6500 9452 6556
rect 9452 6500 9456 6556
rect 9392 6496 9456 6500
rect 9472 6556 9536 6560
rect 9472 6500 9476 6556
rect 9476 6500 9532 6556
rect 9532 6500 9536 6556
rect 9472 6496 9536 6500
rect 9552 6556 9616 6560
rect 9552 6500 9556 6556
rect 9556 6500 9612 6556
rect 9612 6500 9616 6556
rect 9552 6496 9616 6500
rect 9632 6556 9696 6560
rect 9632 6500 9636 6556
rect 9636 6500 9692 6556
rect 9692 6500 9696 6556
rect 9632 6496 9696 6500
rect 17833 6556 17897 6560
rect 17833 6500 17837 6556
rect 17837 6500 17893 6556
rect 17893 6500 17897 6556
rect 17833 6496 17897 6500
rect 17913 6556 17977 6560
rect 17913 6500 17917 6556
rect 17917 6500 17973 6556
rect 17973 6500 17977 6556
rect 17913 6496 17977 6500
rect 17993 6556 18057 6560
rect 17993 6500 17997 6556
rect 17997 6500 18053 6556
rect 18053 6500 18057 6556
rect 17993 6496 18057 6500
rect 18073 6556 18137 6560
rect 18073 6500 18077 6556
rect 18077 6500 18133 6556
rect 18133 6500 18137 6556
rect 18073 6496 18137 6500
rect 26274 6556 26338 6560
rect 26274 6500 26278 6556
rect 26278 6500 26334 6556
rect 26334 6500 26338 6556
rect 26274 6496 26338 6500
rect 26354 6556 26418 6560
rect 26354 6500 26358 6556
rect 26358 6500 26414 6556
rect 26414 6500 26418 6556
rect 26354 6496 26418 6500
rect 26434 6556 26498 6560
rect 26434 6500 26438 6556
rect 26438 6500 26494 6556
rect 26494 6500 26498 6556
rect 26434 6496 26498 6500
rect 26514 6556 26578 6560
rect 26514 6500 26518 6556
rect 26518 6500 26574 6556
rect 26574 6500 26578 6556
rect 26514 6496 26578 6500
rect 34715 6556 34779 6560
rect 34715 6500 34719 6556
rect 34719 6500 34775 6556
rect 34775 6500 34779 6556
rect 34715 6496 34779 6500
rect 34795 6556 34859 6560
rect 34795 6500 34799 6556
rect 34799 6500 34855 6556
rect 34855 6500 34859 6556
rect 34795 6496 34859 6500
rect 34875 6556 34939 6560
rect 34875 6500 34879 6556
rect 34879 6500 34935 6556
rect 34935 6500 34939 6556
rect 34875 6496 34939 6500
rect 34955 6556 35019 6560
rect 34955 6500 34959 6556
rect 34959 6500 35015 6556
rect 35015 6500 35019 6556
rect 34955 6496 35019 6500
rect 5172 6012 5236 6016
rect 5172 5956 5176 6012
rect 5176 5956 5232 6012
rect 5232 5956 5236 6012
rect 5172 5952 5236 5956
rect 5252 6012 5316 6016
rect 5252 5956 5256 6012
rect 5256 5956 5312 6012
rect 5312 5956 5316 6012
rect 5252 5952 5316 5956
rect 5332 6012 5396 6016
rect 5332 5956 5336 6012
rect 5336 5956 5392 6012
rect 5392 5956 5396 6012
rect 5332 5952 5396 5956
rect 5412 6012 5476 6016
rect 5412 5956 5416 6012
rect 5416 5956 5472 6012
rect 5472 5956 5476 6012
rect 5412 5952 5476 5956
rect 13613 6012 13677 6016
rect 13613 5956 13617 6012
rect 13617 5956 13673 6012
rect 13673 5956 13677 6012
rect 13613 5952 13677 5956
rect 13693 6012 13757 6016
rect 13693 5956 13697 6012
rect 13697 5956 13753 6012
rect 13753 5956 13757 6012
rect 13693 5952 13757 5956
rect 13773 6012 13837 6016
rect 13773 5956 13777 6012
rect 13777 5956 13833 6012
rect 13833 5956 13837 6012
rect 13773 5952 13837 5956
rect 13853 6012 13917 6016
rect 13853 5956 13857 6012
rect 13857 5956 13913 6012
rect 13913 5956 13917 6012
rect 13853 5952 13917 5956
rect 22054 6012 22118 6016
rect 22054 5956 22058 6012
rect 22058 5956 22114 6012
rect 22114 5956 22118 6012
rect 22054 5952 22118 5956
rect 22134 6012 22198 6016
rect 22134 5956 22138 6012
rect 22138 5956 22194 6012
rect 22194 5956 22198 6012
rect 22134 5952 22198 5956
rect 22214 6012 22278 6016
rect 22214 5956 22218 6012
rect 22218 5956 22274 6012
rect 22274 5956 22278 6012
rect 22214 5952 22278 5956
rect 22294 6012 22358 6016
rect 22294 5956 22298 6012
rect 22298 5956 22354 6012
rect 22354 5956 22358 6012
rect 22294 5952 22358 5956
rect 30495 6012 30559 6016
rect 30495 5956 30499 6012
rect 30499 5956 30555 6012
rect 30555 5956 30559 6012
rect 30495 5952 30559 5956
rect 30575 6012 30639 6016
rect 30575 5956 30579 6012
rect 30579 5956 30635 6012
rect 30635 5956 30639 6012
rect 30575 5952 30639 5956
rect 30655 6012 30719 6016
rect 30655 5956 30659 6012
rect 30659 5956 30715 6012
rect 30715 5956 30719 6012
rect 30655 5952 30719 5956
rect 30735 6012 30799 6016
rect 30735 5956 30739 6012
rect 30739 5956 30795 6012
rect 30795 5956 30799 6012
rect 30735 5952 30799 5956
rect 9392 5468 9456 5472
rect 9392 5412 9396 5468
rect 9396 5412 9452 5468
rect 9452 5412 9456 5468
rect 9392 5408 9456 5412
rect 9472 5468 9536 5472
rect 9472 5412 9476 5468
rect 9476 5412 9532 5468
rect 9532 5412 9536 5468
rect 9472 5408 9536 5412
rect 9552 5468 9616 5472
rect 9552 5412 9556 5468
rect 9556 5412 9612 5468
rect 9612 5412 9616 5468
rect 9552 5408 9616 5412
rect 9632 5468 9696 5472
rect 9632 5412 9636 5468
rect 9636 5412 9692 5468
rect 9692 5412 9696 5468
rect 9632 5408 9696 5412
rect 17833 5468 17897 5472
rect 17833 5412 17837 5468
rect 17837 5412 17893 5468
rect 17893 5412 17897 5468
rect 17833 5408 17897 5412
rect 17913 5468 17977 5472
rect 17913 5412 17917 5468
rect 17917 5412 17973 5468
rect 17973 5412 17977 5468
rect 17913 5408 17977 5412
rect 17993 5468 18057 5472
rect 17993 5412 17997 5468
rect 17997 5412 18053 5468
rect 18053 5412 18057 5468
rect 17993 5408 18057 5412
rect 18073 5468 18137 5472
rect 18073 5412 18077 5468
rect 18077 5412 18133 5468
rect 18133 5412 18137 5468
rect 18073 5408 18137 5412
rect 26274 5468 26338 5472
rect 26274 5412 26278 5468
rect 26278 5412 26334 5468
rect 26334 5412 26338 5468
rect 26274 5408 26338 5412
rect 26354 5468 26418 5472
rect 26354 5412 26358 5468
rect 26358 5412 26414 5468
rect 26414 5412 26418 5468
rect 26354 5408 26418 5412
rect 26434 5468 26498 5472
rect 26434 5412 26438 5468
rect 26438 5412 26494 5468
rect 26494 5412 26498 5468
rect 26434 5408 26498 5412
rect 26514 5468 26578 5472
rect 26514 5412 26518 5468
rect 26518 5412 26574 5468
rect 26574 5412 26578 5468
rect 26514 5408 26578 5412
rect 34715 5468 34779 5472
rect 34715 5412 34719 5468
rect 34719 5412 34775 5468
rect 34775 5412 34779 5468
rect 34715 5408 34779 5412
rect 34795 5468 34859 5472
rect 34795 5412 34799 5468
rect 34799 5412 34855 5468
rect 34855 5412 34859 5468
rect 34795 5408 34859 5412
rect 34875 5468 34939 5472
rect 34875 5412 34879 5468
rect 34879 5412 34935 5468
rect 34935 5412 34939 5468
rect 34875 5408 34939 5412
rect 34955 5468 35019 5472
rect 34955 5412 34959 5468
rect 34959 5412 35015 5468
rect 35015 5412 35019 5468
rect 34955 5408 35019 5412
rect 5172 4924 5236 4928
rect 5172 4868 5176 4924
rect 5176 4868 5232 4924
rect 5232 4868 5236 4924
rect 5172 4864 5236 4868
rect 5252 4924 5316 4928
rect 5252 4868 5256 4924
rect 5256 4868 5312 4924
rect 5312 4868 5316 4924
rect 5252 4864 5316 4868
rect 5332 4924 5396 4928
rect 5332 4868 5336 4924
rect 5336 4868 5392 4924
rect 5392 4868 5396 4924
rect 5332 4864 5396 4868
rect 5412 4924 5476 4928
rect 5412 4868 5416 4924
rect 5416 4868 5472 4924
rect 5472 4868 5476 4924
rect 5412 4864 5476 4868
rect 13613 4924 13677 4928
rect 13613 4868 13617 4924
rect 13617 4868 13673 4924
rect 13673 4868 13677 4924
rect 13613 4864 13677 4868
rect 13693 4924 13757 4928
rect 13693 4868 13697 4924
rect 13697 4868 13753 4924
rect 13753 4868 13757 4924
rect 13693 4864 13757 4868
rect 13773 4924 13837 4928
rect 13773 4868 13777 4924
rect 13777 4868 13833 4924
rect 13833 4868 13837 4924
rect 13773 4864 13837 4868
rect 13853 4924 13917 4928
rect 13853 4868 13857 4924
rect 13857 4868 13913 4924
rect 13913 4868 13917 4924
rect 13853 4864 13917 4868
rect 22054 4924 22118 4928
rect 22054 4868 22058 4924
rect 22058 4868 22114 4924
rect 22114 4868 22118 4924
rect 22054 4864 22118 4868
rect 22134 4924 22198 4928
rect 22134 4868 22138 4924
rect 22138 4868 22194 4924
rect 22194 4868 22198 4924
rect 22134 4864 22198 4868
rect 22214 4924 22278 4928
rect 22214 4868 22218 4924
rect 22218 4868 22274 4924
rect 22274 4868 22278 4924
rect 22214 4864 22278 4868
rect 22294 4924 22358 4928
rect 22294 4868 22298 4924
rect 22298 4868 22354 4924
rect 22354 4868 22358 4924
rect 22294 4864 22358 4868
rect 30495 4924 30559 4928
rect 30495 4868 30499 4924
rect 30499 4868 30555 4924
rect 30555 4868 30559 4924
rect 30495 4864 30559 4868
rect 30575 4924 30639 4928
rect 30575 4868 30579 4924
rect 30579 4868 30635 4924
rect 30635 4868 30639 4924
rect 30575 4864 30639 4868
rect 30655 4924 30719 4928
rect 30655 4868 30659 4924
rect 30659 4868 30715 4924
rect 30715 4868 30719 4924
rect 30655 4864 30719 4868
rect 30735 4924 30799 4928
rect 30735 4868 30739 4924
rect 30739 4868 30795 4924
rect 30795 4868 30799 4924
rect 30735 4864 30799 4868
rect 9392 4380 9456 4384
rect 9392 4324 9396 4380
rect 9396 4324 9452 4380
rect 9452 4324 9456 4380
rect 9392 4320 9456 4324
rect 9472 4380 9536 4384
rect 9472 4324 9476 4380
rect 9476 4324 9532 4380
rect 9532 4324 9536 4380
rect 9472 4320 9536 4324
rect 9552 4380 9616 4384
rect 9552 4324 9556 4380
rect 9556 4324 9612 4380
rect 9612 4324 9616 4380
rect 9552 4320 9616 4324
rect 9632 4380 9696 4384
rect 9632 4324 9636 4380
rect 9636 4324 9692 4380
rect 9692 4324 9696 4380
rect 9632 4320 9696 4324
rect 17833 4380 17897 4384
rect 17833 4324 17837 4380
rect 17837 4324 17893 4380
rect 17893 4324 17897 4380
rect 17833 4320 17897 4324
rect 17913 4380 17977 4384
rect 17913 4324 17917 4380
rect 17917 4324 17973 4380
rect 17973 4324 17977 4380
rect 17913 4320 17977 4324
rect 17993 4380 18057 4384
rect 17993 4324 17997 4380
rect 17997 4324 18053 4380
rect 18053 4324 18057 4380
rect 17993 4320 18057 4324
rect 18073 4380 18137 4384
rect 18073 4324 18077 4380
rect 18077 4324 18133 4380
rect 18133 4324 18137 4380
rect 18073 4320 18137 4324
rect 26274 4380 26338 4384
rect 26274 4324 26278 4380
rect 26278 4324 26334 4380
rect 26334 4324 26338 4380
rect 26274 4320 26338 4324
rect 26354 4380 26418 4384
rect 26354 4324 26358 4380
rect 26358 4324 26414 4380
rect 26414 4324 26418 4380
rect 26354 4320 26418 4324
rect 26434 4380 26498 4384
rect 26434 4324 26438 4380
rect 26438 4324 26494 4380
rect 26494 4324 26498 4380
rect 26434 4320 26498 4324
rect 26514 4380 26578 4384
rect 26514 4324 26518 4380
rect 26518 4324 26574 4380
rect 26574 4324 26578 4380
rect 26514 4320 26578 4324
rect 34715 4380 34779 4384
rect 34715 4324 34719 4380
rect 34719 4324 34775 4380
rect 34775 4324 34779 4380
rect 34715 4320 34779 4324
rect 34795 4380 34859 4384
rect 34795 4324 34799 4380
rect 34799 4324 34855 4380
rect 34855 4324 34859 4380
rect 34795 4320 34859 4324
rect 34875 4380 34939 4384
rect 34875 4324 34879 4380
rect 34879 4324 34935 4380
rect 34935 4324 34939 4380
rect 34875 4320 34939 4324
rect 34955 4380 35019 4384
rect 34955 4324 34959 4380
rect 34959 4324 35015 4380
rect 35015 4324 35019 4380
rect 34955 4320 35019 4324
rect 5172 3836 5236 3840
rect 5172 3780 5176 3836
rect 5176 3780 5232 3836
rect 5232 3780 5236 3836
rect 5172 3776 5236 3780
rect 5252 3836 5316 3840
rect 5252 3780 5256 3836
rect 5256 3780 5312 3836
rect 5312 3780 5316 3836
rect 5252 3776 5316 3780
rect 5332 3836 5396 3840
rect 5332 3780 5336 3836
rect 5336 3780 5392 3836
rect 5392 3780 5396 3836
rect 5332 3776 5396 3780
rect 5412 3836 5476 3840
rect 5412 3780 5416 3836
rect 5416 3780 5472 3836
rect 5472 3780 5476 3836
rect 5412 3776 5476 3780
rect 13613 3836 13677 3840
rect 13613 3780 13617 3836
rect 13617 3780 13673 3836
rect 13673 3780 13677 3836
rect 13613 3776 13677 3780
rect 13693 3836 13757 3840
rect 13693 3780 13697 3836
rect 13697 3780 13753 3836
rect 13753 3780 13757 3836
rect 13693 3776 13757 3780
rect 13773 3836 13837 3840
rect 13773 3780 13777 3836
rect 13777 3780 13833 3836
rect 13833 3780 13837 3836
rect 13773 3776 13837 3780
rect 13853 3836 13917 3840
rect 13853 3780 13857 3836
rect 13857 3780 13913 3836
rect 13913 3780 13917 3836
rect 13853 3776 13917 3780
rect 22054 3836 22118 3840
rect 22054 3780 22058 3836
rect 22058 3780 22114 3836
rect 22114 3780 22118 3836
rect 22054 3776 22118 3780
rect 22134 3836 22198 3840
rect 22134 3780 22138 3836
rect 22138 3780 22194 3836
rect 22194 3780 22198 3836
rect 22134 3776 22198 3780
rect 22214 3836 22278 3840
rect 22214 3780 22218 3836
rect 22218 3780 22274 3836
rect 22274 3780 22278 3836
rect 22214 3776 22278 3780
rect 22294 3836 22358 3840
rect 22294 3780 22298 3836
rect 22298 3780 22354 3836
rect 22354 3780 22358 3836
rect 22294 3776 22358 3780
rect 30495 3836 30559 3840
rect 30495 3780 30499 3836
rect 30499 3780 30555 3836
rect 30555 3780 30559 3836
rect 30495 3776 30559 3780
rect 30575 3836 30639 3840
rect 30575 3780 30579 3836
rect 30579 3780 30635 3836
rect 30635 3780 30639 3836
rect 30575 3776 30639 3780
rect 30655 3836 30719 3840
rect 30655 3780 30659 3836
rect 30659 3780 30715 3836
rect 30715 3780 30719 3836
rect 30655 3776 30719 3780
rect 30735 3836 30799 3840
rect 30735 3780 30739 3836
rect 30739 3780 30795 3836
rect 30795 3780 30799 3836
rect 30735 3776 30799 3780
rect 9392 3292 9456 3296
rect 9392 3236 9396 3292
rect 9396 3236 9452 3292
rect 9452 3236 9456 3292
rect 9392 3232 9456 3236
rect 9472 3292 9536 3296
rect 9472 3236 9476 3292
rect 9476 3236 9532 3292
rect 9532 3236 9536 3292
rect 9472 3232 9536 3236
rect 9552 3292 9616 3296
rect 9552 3236 9556 3292
rect 9556 3236 9612 3292
rect 9612 3236 9616 3292
rect 9552 3232 9616 3236
rect 9632 3292 9696 3296
rect 9632 3236 9636 3292
rect 9636 3236 9692 3292
rect 9692 3236 9696 3292
rect 9632 3232 9696 3236
rect 17833 3292 17897 3296
rect 17833 3236 17837 3292
rect 17837 3236 17893 3292
rect 17893 3236 17897 3292
rect 17833 3232 17897 3236
rect 17913 3292 17977 3296
rect 17913 3236 17917 3292
rect 17917 3236 17973 3292
rect 17973 3236 17977 3292
rect 17913 3232 17977 3236
rect 17993 3292 18057 3296
rect 17993 3236 17997 3292
rect 17997 3236 18053 3292
rect 18053 3236 18057 3292
rect 17993 3232 18057 3236
rect 18073 3292 18137 3296
rect 18073 3236 18077 3292
rect 18077 3236 18133 3292
rect 18133 3236 18137 3292
rect 18073 3232 18137 3236
rect 26274 3292 26338 3296
rect 26274 3236 26278 3292
rect 26278 3236 26334 3292
rect 26334 3236 26338 3292
rect 26274 3232 26338 3236
rect 26354 3292 26418 3296
rect 26354 3236 26358 3292
rect 26358 3236 26414 3292
rect 26414 3236 26418 3292
rect 26354 3232 26418 3236
rect 26434 3292 26498 3296
rect 26434 3236 26438 3292
rect 26438 3236 26494 3292
rect 26494 3236 26498 3292
rect 26434 3232 26498 3236
rect 26514 3292 26578 3296
rect 26514 3236 26518 3292
rect 26518 3236 26574 3292
rect 26574 3236 26578 3292
rect 26514 3232 26578 3236
rect 34715 3292 34779 3296
rect 34715 3236 34719 3292
rect 34719 3236 34775 3292
rect 34775 3236 34779 3292
rect 34715 3232 34779 3236
rect 34795 3292 34859 3296
rect 34795 3236 34799 3292
rect 34799 3236 34855 3292
rect 34855 3236 34859 3292
rect 34795 3232 34859 3236
rect 34875 3292 34939 3296
rect 34875 3236 34879 3292
rect 34879 3236 34935 3292
rect 34935 3236 34939 3292
rect 34875 3232 34939 3236
rect 34955 3292 35019 3296
rect 34955 3236 34959 3292
rect 34959 3236 35015 3292
rect 35015 3236 35019 3292
rect 34955 3232 35019 3236
rect 5172 2748 5236 2752
rect 5172 2692 5176 2748
rect 5176 2692 5232 2748
rect 5232 2692 5236 2748
rect 5172 2688 5236 2692
rect 5252 2748 5316 2752
rect 5252 2692 5256 2748
rect 5256 2692 5312 2748
rect 5312 2692 5316 2748
rect 5252 2688 5316 2692
rect 5332 2748 5396 2752
rect 5332 2692 5336 2748
rect 5336 2692 5392 2748
rect 5392 2692 5396 2748
rect 5332 2688 5396 2692
rect 5412 2748 5476 2752
rect 5412 2692 5416 2748
rect 5416 2692 5472 2748
rect 5472 2692 5476 2748
rect 5412 2688 5476 2692
rect 13613 2748 13677 2752
rect 13613 2692 13617 2748
rect 13617 2692 13673 2748
rect 13673 2692 13677 2748
rect 13613 2688 13677 2692
rect 13693 2748 13757 2752
rect 13693 2692 13697 2748
rect 13697 2692 13753 2748
rect 13753 2692 13757 2748
rect 13693 2688 13757 2692
rect 13773 2748 13837 2752
rect 13773 2692 13777 2748
rect 13777 2692 13833 2748
rect 13833 2692 13837 2748
rect 13773 2688 13837 2692
rect 13853 2748 13917 2752
rect 13853 2692 13857 2748
rect 13857 2692 13913 2748
rect 13913 2692 13917 2748
rect 13853 2688 13917 2692
rect 22054 2748 22118 2752
rect 22054 2692 22058 2748
rect 22058 2692 22114 2748
rect 22114 2692 22118 2748
rect 22054 2688 22118 2692
rect 22134 2748 22198 2752
rect 22134 2692 22138 2748
rect 22138 2692 22194 2748
rect 22194 2692 22198 2748
rect 22134 2688 22198 2692
rect 22214 2748 22278 2752
rect 22214 2692 22218 2748
rect 22218 2692 22274 2748
rect 22274 2692 22278 2748
rect 22214 2688 22278 2692
rect 22294 2748 22358 2752
rect 22294 2692 22298 2748
rect 22298 2692 22354 2748
rect 22354 2692 22358 2748
rect 22294 2688 22358 2692
rect 30495 2748 30559 2752
rect 30495 2692 30499 2748
rect 30499 2692 30555 2748
rect 30555 2692 30559 2748
rect 30495 2688 30559 2692
rect 30575 2748 30639 2752
rect 30575 2692 30579 2748
rect 30579 2692 30635 2748
rect 30635 2692 30639 2748
rect 30575 2688 30639 2692
rect 30655 2748 30719 2752
rect 30655 2692 30659 2748
rect 30659 2692 30715 2748
rect 30715 2692 30719 2748
rect 30655 2688 30719 2692
rect 30735 2748 30799 2752
rect 30735 2692 30739 2748
rect 30739 2692 30795 2748
rect 30795 2692 30799 2748
rect 30735 2688 30799 2692
rect 9392 2204 9456 2208
rect 9392 2148 9396 2204
rect 9396 2148 9452 2204
rect 9452 2148 9456 2204
rect 9392 2144 9456 2148
rect 9472 2204 9536 2208
rect 9472 2148 9476 2204
rect 9476 2148 9532 2204
rect 9532 2148 9536 2204
rect 9472 2144 9536 2148
rect 9552 2204 9616 2208
rect 9552 2148 9556 2204
rect 9556 2148 9612 2204
rect 9612 2148 9616 2204
rect 9552 2144 9616 2148
rect 9632 2204 9696 2208
rect 9632 2148 9636 2204
rect 9636 2148 9692 2204
rect 9692 2148 9696 2204
rect 9632 2144 9696 2148
rect 17833 2204 17897 2208
rect 17833 2148 17837 2204
rect 17837 2148 17893 2204
rect 17893 2148 17897 2204
rect 17833 2144 17897 2148
rect 17913 2204 17977 2208
rect 17913 2148 17917 2204
rect 17917 2148 17973 2204
rect 17973 2148 17977 2204
rect 17913 2144 17977 2148
rect 17993 2204 18057 2208
rect 17993 2148 17997 2204
rect 17997 2148 18053 2204
rect 18053 2148 18057 2204
rect 17993 2144 18057 2148
rect 18073 2204 18137 2208
rect 18073 2148 18077 2204
rect 18077 2148 18133 2204
rect 18133 2148 18137 2204
rect 18073 2144 18137 2148
rect 26274 2204 26338 2208
rect 26274 2148 26278 2204
rect 26278 2148 26334 2204
rect 26334 2148 26338 2204
rect 26274 2144 26338 2148
rect 26354 2204 26418 2208
rect 26354 2148 26358 2204
rect 26358 2148 26414 2204
rect 26414 2148 26418 2204
rect 26354 2144 26418 2148
rect 26434 2204 26498 2208
rect 26434 2148 26438 2204
rect 26438 2148 26494 2204
rect 26494 2148 26498 2204
rect 26434 2144 26498 2148
rect 26514 2204 26578 2208
rect 26514 2148 26518 2204
rect 26518 2148 26574 2204
rect 26574 2148 26578 2204
rect 26514 2144 26578 2148
rect 34715 2204 34779 2208
rect 34715 2148 34719 2204
rect 34719 2148 34775 2204
rect 34775 2148 34779 2204
rect 34715 2144 34779 2148
rect 34795 2204 34859 2208
rect 34795 2148 34799 2204
rect 34799 2148 34855 2204
rect 34855 2148 34859 2204
rect 34795 2144 34859 2148
rect 34875 2204 34939 2208
rect 34875 2148 34879 2204
rect 34879 2148 34935 2204
rect 34935 2148 34939 2204
rect 34875 2144 34939 2148
rect 34955 2204 35019 2208
rect 34955 2148 34959 2204
rect 34959 2148 35015 2204
rect 35015 2148 35019 2204
rect 34955 2144 35019 2148
<< metal4 >>
rect 5164 33216 5484 33776
rect 5164 33152 5172 33216
rect 5236 33152 5252 33216
rect 5316 33152 5332 33216
rect 5396 33152 5412 33216
rect 5476 33152 5484 33216
rect 5164 32128 5484 33152
rect 5164 32064 5172 32128
rect 5236 32064 5252 32128
rect 5316 32064 5332 32128
rect 5396 32064 5412 32128
rect 5476 32064 5484 32128
rect 5164 31040 5484 32064
rect 5164 30976 5172 31040
rect 5236 30976 5252 31040
rect 5316 30976 5332 31040
rect 5396 30976 5412 31040
rect 5476 30976 5484 31040
rect 5164 29952 5484 30976
rect 5164 29888 5172 29952
rect 5236 29888 5252 29952
rect 5316 29888 5332 29952
rect 5396 29888 5412 29952
rect 5476 29888 5484 29952
rect 5164 28864 5484 29888
rect 5164 28800 5172 28864
rect 5236 28800 5252 28864
rect 5316 28800 5332 28864
rect 5396 28800 5412 28864
rect 5476 28800 5484 28864
rect 5164 27776 5484 28800
rect 5164 27712 5172 27776
rect 5236 27712 5252 27776
rect 5316 27712 5332 27776
rect 5396 27712 5412 27776
rect 5476 27712 5484 27776
rect 5164 26688 5484 27712
rect 5164 26624 5172 26688
rect 5236 26624 5252 26688
rect 5316 26624 5332 26688
rect 5396 26624 5412 26688
rect 5476 26624 5484 26688
rect 5164 25600 5484 26624
rect 5164 25536 5172 25600
rect 5236 25536 5252 25600
rect 5316 25536 5332 25600
rect 5396 25536 5412 25600
rect 5476 25536 5484 25600
rect 5164 24512 5484 25536
rect 5164 24448 5172 24512
rect 5236 24448 5252 24512
rect 5316 24448 5332 24512
rect 5396 24448 5412 24512
rect 5476 24448 5484 24512
rect 5164 23424 5484 24448
rect 5164 23360 5172 23424
rect 5236 23360 5252 23424
rect 5316 23360 5332 23424
rect 5396 23360 5412 23424
rect 5476 23360 5484 23424
rect 5164 22336 5484 23360
rect 5164 22272 5172 22336
rect 5236 22272 5252 22336
rect 5316 22272 5332 22336
rect 5396 22272 5412 22336
rect 5476 22272 5484 22336
rect 5164 21248 5484 22272
rect 5164 21184 5172 21248
rect 5236 21184 5252 21248
rect 5316 21184 5332 21248
rect 5396 21184 5412 21248
rect 5476 21184 5484 21248
rect 5164 20160 5484 21184
rect 5164 20096 5172 20160
rect 5236 20096 5252 20160
rect 5316 20096 5332 20160
rect 5396 20096 5412 20160
rect 5476 20096 5484 20160
rect 5164 19072 5484 20096
rect 5164 19008 5172 19072
rect 5236 19008 5252 19072
rect 5316 19008 5332 19072
rect 5396 19008 5412 19072
rect 5476 19008 5484 19072
rect 5164 17984 5484 19008
rect 5164 17920 5172 17984
rect 5236 17920 5252 17984
rect 5316 17920 5332 17984
rect 5396 17920 5412 17984
rect 5476 17920 5484 17984
rect 5164 16896 5484 17920
rect 5164 16832 5172 16896
rect 5236 16832 5252 16896
rect 5316 16832 5332 16896
rect 5396 16832 5412 16896
rect 5476 16832 5484 16896
rect 5164 15808 5484 16832
rect 5164 15744 5172 15808
rect 5236 15744 5252 15808
rect 5316 15744 5332 15808
rect 5396 15744 5412 15808
rect 5476 15744 5484 15808
rect 5164 14720 5484 15744
rect 5164 14656 5172 14720
rect 5236 14656 5252 14720
rect 5316 14656 5332 14720
rect 5396 14656 5412 14720
rect 5476 14656 5484 14720
rect 5164 13632 5484 14656
rect 5164 13568 5172 13632
rect 5236 13568 5252 13632
rect 5316 13568 5332 13632
rect 5396 13568 5412 13632
rect 5476 13568 5484 13632
rect 5164 12544 5484 13568
rect 5164 12480 5172 12544
rect 5236 12480 5252 12544
rect 5316 12480 5332 12544
rect 5396 12480 5412 12544
rect 5476 12480 5484 12544
rect 5164 11456 5484 12480
rect 5164 11392 5172 11456
rect 5236 11392 5252 11456
rect 5316 11392 5332 11456
rect 5396 11392 5412 11456
rect 5476 11392 5484 11456
rect 5164 10368 5484 11392
rect 5164 10304 5172 10368
rect 5236 10304 5252 10368
rect 5316 10304 5332 10368
rect 5396 10304 5412 10368
rect 5476 10304 5484 10368
rect 5164 9280 5484 10304
rect 5164 9216 5172 9280
rect 5236 9216 5252 9280
rect 5316 9216 5332 9280
rect 5396 9216 5412 9280
rect 5476 9216 5484 9280
rect 5164 8192 5484 9216
rect 5164 8128 5172 8192
rect 5236 8128 5252 8192
rect 5316 8128 5332 8192
rect 5396 8128 5412 8192
rect 5476 8128 5484 8192
rect 5164 7104 5484 8128
rect 5164 7040 5172 7104
rect 5236 7040 5252 7104
rect 5316 7040 5332 7104
rect 5396 7040 5412 7104
rect 5476 7040 5484 7104
rect 5164 6016 5484 7040
rect 5164 5952 5172 6016
rect 5236 5952 5252 6016
rect 5316 5952 5332 6016
rect 5396 5952 5412 6016
rect 5476 5952 5484 6016
rect 5164 4928 5484 5952
rect 5164 4864 5172 4928
rect 5236 4864 5252 4928
rect 5316 4864 5332 4928
rect 5396 4864 5412 4928
rect 5476 4864 5484 4928
rect 5164 3840 5484 4864
rect 5164 3776 5172 3840
rect 5236 3776 5252 3840
rect 5316 3776 5332 3840
rect 5396 3776 5412 3840
rect 5476 3776 5484 3840
rect 5164 2752 5484 3776
rect 5164 2688 5172 2752
rect 5236 2688 5252 2752
rect 5316 2688 5332 2752
rect 5396 2688 5412 2752
rect 5476 2688 5484 2752
rect 5164 2128 5484 2688
rect 9384 33760 9704 33776
rect 9384 33696 9392 33760
rect 9456 33696 9472 33760
rect 9536 33696 9552 33760
rect 9616 33696 9632 33760
rect 9696 33696 9704 33760
rect 9384 32672 9704 33696
rect 9384 32608 9392 32672
rect 9456 32608 9472 32672
rect 9536 32608 9552 32672
rect 9616 32608 9632 32672
rect 9696 32608 9704 32672
rect 9384 31584 9704 32608
rect 9384 31520 9392 31584
rect 9456 31520 9472 31584
rect 9536 31520 9552 31584
rect 9616 31520 9632 31584
rect 9696 31520 9704 31584
rect 9384 30496 9704 31520
rect 9384 30432 9392 30496
rect 9456 30432 9472 30496
rect 9536 30432 9552 30496
rect 9616 30432 9632 30496
rect 9696 30432 9704 30496
rect 9384 29408 9704 30432
rect 9384 29344 9392 29408
rect 9456 29344 9472 29408
rect 9536 29344 9552 29408
rect 9616 29344 9632 29408
rect 9696 29344 9704 29408
rect 9384 28320 9704 29344
rect 9384 28256 9392 28320
rect 9456 28256 9472 28320
rect 9536 28256 9552 28320
rect 9616 28256 9632 28320
rect 9696 28256 9704 28320
rect 9384 27232 9704 28256
rect 9384 27168 9392 27232
rect 9456 27168 9472 27232
rect 9536 27168 9552 27232
rect 9616 27168 9632 27232
rect 9696 27168 9704 27232
rect 9384 26144 9704 27168
rect 9384 26080 9392 26144
rect 9456 26080 9472 26144
rect 9536 26080 9552 26144
rect 9616 26080 9632 26144
rect 9696 26080 9704 26144
rect 9384 25056 9704 26080
rect 9384 24992 9392 25056
rect 9456 24992 9472 25056
rect 9536 24992 9552 25056
rect 9616 24992 9632 25056
rect 9696 24992 9704 25056
rect 9384 23968 9704 24992
rect 9384 23904 9392 23968
rect 9456 23904 9472 23968
rect 9536 23904 9552 23968
rect 9616 23904 9632 23968
rect 9696 23904 9704 23968
rect 9384 22880 9704 23904
rect 9384 22816 9392 22880
rect 9456 22816 9472 22880
rect 9536 22816 9552 22880
rect 9616 22816 9632 22880
rect 9696 22816 9704 22880
rect 9384 21792 9704 22816
rect 9384 21728 9392 21792
rect 9456 21728 9472 21792
rect 9536 21728 9552 21792
rect 9616 21728 9632 21792
rect 9696 21728 9704 21792
rect 9384 20704 9704 21728
rect 9384 20640 9392 20704
rect 9456 20640 9472 20704
rect 9536 20640 9552 20704
rect 9616 20640 9632 20704
rect 9696 20640 9704 20704
rect 9384 19616 9704 20640
rect 9384 19552 9392 19616
rect 9456 19552 9472 19616
rect 9536 19552 9552 19616
rect 9616 19552 9632 19616
rect 9696 19552 9704 19616
rect 9384 18528 9704 19552
rect 9384 18464 9392 18528
rect 9456 18464 9472 18528
rect 9536 18464 9552 18528
rect 9616 18464 9632 18528
rect 9696 18464 9704 18528
rect 9384 17440 9704 18464
rect 9384 17376 9392 17440
rect 9456 17376 9472 17440
rect 9536 17376 9552 17440
rect 9616 17376 9632 17440
rect 9696 17376 9704 17440
rect 9384 16352 9704 17376
rect 9384 16288 9392 16352
rect 9456 16288 9472 16352
rect 9536 16288 9552 16352
rect 9616 16288 9632 16352
rect 9696 16288 9704 16352
rect 9384 15264 9704 16288
rect 9384 15200 9392 15264
rect 9456 15200 9472 15264
rect 9536 15200 9552 15264
rect 9616 15200 9632 15264
rect 9696 15200 9704 15264
rect 9384 14176 9704 15200
rect 9384 14112 9392 14176
rect 9456 14112 9472 14176
rect 9536 14112 9552 14176
rect 9616 14112 9632 14176
rect 9696 14112 9704 14176
rect 9384 13088 9704 14112
rect 9384 13024 9392 13088
rect 9456 13024 9472 13088
rect 9536 13024 9552 13088
rect 9616 13024 9632 13088
rect 9696 13024 9704 13088
rect 9384 12000 9704 13024
rect 9384 11936 9392 12000
rect 9456 11936 9472 12000
rect 9536 11936 9552 12000
rect 9616 11936 9632 12000
rect 9696 11936 9704 12000
rect 9384 10912 9704 11936
rect 9384 10848 9392 10912
rect 9456 10848 9472 10912
rect 9536 10848 9552 10912
rect 9616 10848 9632 10912
rect 9696 10848 9704 10912
rect 9384 9824 9704 10848
rect 9384 9760 9392 9824
rect 9456 9760 9472 9824
rect 9536 9760 9552 9824
rect 9616 9760 9632 9824
rect 9696 9760 9704 9824
rect 9384 8736 9704 9760
rect 9384 8672 9392 8736
rect 9456 8672 9472 8736
rect 9536 8672 9552 8736
rect 9616 8672 9632 8736
rect 9696 8672 9704 8736
rect 9384 7648 9704 8672
rect 9384 7584 9392 7648
rect 9456 7584 9472 7648
rect 9536 7584 9552 7648
rect 9616 7584 9632 7648
rect 9696 7584 9704 7648
rect 9384 6560 9704 7584
rect 9384 6496 9392 6560
rect 9456 6496 9472 6560
rect 9536 6496 9552 6560
rect 9616 6496 9632 6560
rect 9696 6496 9704 6560
rect 9384 5472 9704 6496
rect 9384 5408 9392 5472
rect 9456 5408 9472 5472
rect 9536 5408 9552 5472
rect 9616 5408 9632 5472
rect 9696 5408 9704 5472
rect 9384 4384 9704 5408
rect 9384 4320 9392 4384
rect 9456 4320 9472 4384
rect 9536 4320 9552 4384
rect 9616 4320 9632 4384
rect 9696 4320 9704 4384
rect 9384 3296 9704 4320
rect 9384 3232 9392 3296
rect 9456 3232 9472 3296
rect 9536 3232 9552 3296
rect 9616 3232 9632 3296
rect 9696 3232 9704 3296
rect 9384 2208 9704 3232
rect 9384 2144 9392 2208
rect 9456 2144 9472 2208
rect 9536 2144 9552 2208
rect 9616 2144 9632 2208
rect 9696 2144 9704 2208
rect 9384 2128 9704 2144
rect 13605 33216 13925 33776
rect 13605 33152 13613 33216
rect 13677 33152 13693 33216
rect 13757 33152 13773 33216
rect 13837 33152 13853 33216
rect 13917 33152 13925 33216
rect 13605 32128 13925 33152
rect 13605 32064 13613 32128
rect 13677 32064 13693 32128
rect 13757 32064 13773 32128
rect 13837 32064 13853 32128
rect 13917 32064 13925 32128
rect 13605 31040 13925 32064
rect 13605 30976 13613 31040
rect 13677 30976 13693 31040
rect 13757 30976 13773 31040
rect 13837 30976 13853 31040
rect 13917 30976 13925 31040
rect 13605 29952 13925 30976
rect 13605 29888 13613 29952
rect 13677 29888 13693 29952
rect 13757 29888 13773 29952
rect 13837 29888 13853 29952
rect 13917 29888 13925 29952
rect 13605 28864 13925 29888
rect 13605 28800 13613 28864
rect 13677 28800 13693 28864
rect 13757 28800 13773 28864
rect 13837 28800 13853 28864
rect 13917 28800 13925 28864
rect 13605 27776 13925 28800
rect 13605 27712 13613 27776
rect 13677 27712 13693 27776
rect 13757 27712 13773 27776
rect 13837 27712 13853 27776
rect 13917 27712 13925 27776
rect 13605 26688 13925 27712
rect 13605 26624 13613 26688
rect 13677 26624 13693 26688
rect 13757 26624 13773 26688
rect 13837 26624 13853 26688
rect 13917 26624 13925 26688
rect 13605 25600 13925 26624
rect 13605 25536 13613 25600
rect 13677 25536 13693 25600
rect 13757 25536 13773 25600
rect 13837 25536 13853 25600
rect 13917 25536 13925 25600
rect 13605 24512 13925 25536
rect 13605 24448 13613 24512
rect 13677 24448 13693 24512
rect 13757 24448 13773 24512
rect 13837 24448 13853 24512
rect 13917 24448 13925 24512
rect 13605 23424 13925 24448
rect 13605 23360 13613 23424
rect 13677 23360 13693 23424
rect 13757 23360 13773 23424
rect 13837 23360 13853 23424
rect 13917 23360 13925 23424
rect 13605 22336 13925 23360
rect 13605 22272 13613 22336
rect 13677 22272 13693 22336
rect 13757 22272 13773 22336
rect 13837 22272 13853 22336
rect 13917 22272 13925 22336
rect 13605 21248 13925 22272
rect 13605 21184 13613 21248
rect 13677 21184 13693 21248
rect 13757 21184 13773 21248
rect 13837 21184 13853 21248
rect 13917 21184 13925 21248
rect 13605 20160 13925 21184
rect 13605 20096 13613 20160
rect 13677 20096 13693 20160
rect 13757 20096 13773 20160
rect 13837 20096 13853 20160
rect 13917 20096 13925 20160
rect 13605 19072 13925 20096
rect 13605 19008 13613 19072
rect 13677 19008 13693 19072
rect 13757 19008 13773 19072
rect 13837 19008 13853 19072
rect 13917 19008 13925 19072
rect 13605 17984 13925 19008
rect 13605 17920 13613 17984
rect 13677 17920 13693 17984
rect 13757 17920 13773 17984
rect 13837 17920 13853 17984
rect 13917 17920 13925 17984
rect 13605 16896 13925 17920
rect 13605 16832 13613 16896
rect 13677 16832 13693 16896
rect 13757 16832 13773 16896
rect 13837 16832 13853 16896
rect 13917 16832 13925 16896
rect 13605 15808 13925 16832
rect 13605 15744 13613 15808
rect 13677 15744 13693 15808
rect 13757 15744 13773 15808
rect 13837 15744 13853 15808
rect 13917 15744 13925 15808
rect 13605 14720 13925 15744
rect 13605 14656 13613 14720
rect 13677 14656 13693 14720
rect 13757 14656 13773 14720
rect 13837 14656 13853 14720
rect 13917 14656 13925 14720
rect 13605 13632 13925 14656
rect 13605 13568 13613 13632
rect 13677 13568 13693 13632
rect 13757 13568 13773 13632
rect 13837 13568 13853 13632
rect 13917 13568 13925 13632
rect 13605 12544 13925 13568
rect 13605 12480 13613 12544
rect 13677 12480 13693 12544
rect 13757 12480 13773 12544
rect 13837 12480 13853 12544
rect 13917 12480 13925 12544
rect 13605 11456 13925 12480
rect 13605 11392 13613 11456
rect 13677 11392 13693 11456
rect 13757 11392 13773 11456
rect 13837 11392 13853 11456
rect 13917 11392 13925 11456
rect 13605 10368 13925 11392
rect 13605 10304 13613 10368
rect 13677 10304 13693 10368
rect 13757 10304 13773 10368
rect 13837 10304 13853 10368
rect 13917 10304 13925 10368
rect 13605 9280 13925 10304
rect 13605 9216 13613 9280
rect 13677 9216 13693 9280
rect 13757 9216 13773 9280
rect 13837 9216 13853 9280
rect 13917 9216 13925 9280
rect 13605 8192 13925 9216
rect 13605 8128 13613 8192
rect 13677 8128 13693 8192
rect 13757 8128 13773 8192
rect 13837 8128 13853 8192
rect 13917 8128 13925 8192
rect 13605 7104 13925 8128
rect 13605 7040 13613 7104
rect 13677 7040 13693 7104
rect 13757 7040 13773 7104
rect 13837 7040 13853 7104
rect 13917 7040 13925 7104
rect 13605 6016 13925 7040
rect 13605 5952 13613 6016
rect 13677 5952 13693 6016
rect 13757 5952 13773 6016
rect 13837 5952 13853 6016
rect 13917 5952 13925 6016
rect 13605 4928 13925 5952
rect 13605 4864 13613 4928
rect 13677 4864 13693 4928
rect 13757 4864 13773 4928
rect 13837 4864 13853 4928
rect 13917 4864 13925 4928
rect 13605 3840 13925 4864
rect 13605 3776 13613 3840
rect 13677 3776 13693 3840
rect 13757 3776 13773 3840
rect 13837 3776 13853 3840
rect 13917 3776 13925 3840
rect 13605 2752 13925 3776
rect 13605 2688 13613 2752
rect 13677 2688 13693 2752
rect 13757 2688 13773 2752
rect 13837 2688 13853 2752
rect 13917 2688 13925 2752
rect 13605 2128 13925 2688
rect 17825 33760 18145 33776
rect 17825 33696 17833 33760
rect 17897 33696 17913 33760
rect 17977 33696 17993 33760
rect 18057 33696 18073 33760
rect 18137 33696 18145 33760
rect 17825 32672 18145 33696
rect 17825 32608 17833 32672
rect 17897 32608 17913 32672
rect 17977 32608 17993 32672
rect 18057 32608 18073 32672
rect 18137 32608 18145 32672
rect 17825 31584 18145 32608
rect 17825 31520 17833 31584
rect 17897 31520 17913 31584
rect 17977 31520 17993 31584
rect 18057 31520 18073 31584
rect 18137 31520 18145 31584
rect 17825 30496 18145 31520
rect 17825 30432 17833 30496
rect 17897 30432 17913 30496
rect 17977 30432 17993 30496
rect 18057 30432 18073 30496
rect 18137 30432 18145 30496
rect 17825 29408 18145 30432
rect 17825 29344 17833 29408
rect 17897 29344 17913 29408
rect 17977 29344 17993 29408
rect 18057 29344 18073 29408
rect 18137 29344 18145 29408
rect 17825 28320 18145 29344
rect 17825 28256 17833 28320
rect 17897 28256 17913 28320
rect 17977 28256 17993 28320
rect 18057 28256 18073 28320
rect 18137 28256 18145 28320
rect 17825 27232 18145 28256
rect 17825 27168 17833 27232
rect 17897 27168 17913 27232
rect 17977 27168 17993 27232
rect 18057 27168 18073 27232
rect 18137 27168 18145 27232
rect 17825 26144 18145 27168
rect 17825 26080 17833 26144
rect 17897 26080 17913 26144
rect 17977 26080 17993 26144
rect 18057 26080 18073 26144
rect 18137 26080 18145 26144
rect 17825 25056 18145 26080
rect 17825 24992 17833 25056
rect 17897 24992 17913 25056
rect 17977 24992 17993 25056
rect 18057 24992 18073 25056
rect 18137 24992 18145 25056
rect 17825 23968 18145 24992
rect 17825 23904 17833 23968
rect 17897 23904 17913 23968
rect 17977 23904 17993 23968
rect 18057 23904 18073 23968
rect 18137 23904 18145 23968
rect 17825 22880 18145 23904
rect 17825 22816 17833 22880
rect 17897 22816 17913 22880
rect 17977 22816 17993 22880
rect 18057 22816 18073 22880
rect 18137 22816 18145 22880
rect 17825 21792 18145 22816
rect 17825 21728 17833 21792
rect 17897 21728 17913 21792
rect 17977 21728 17993 21792
rect 18057 21728 18073 21792
rect 18137 21728 18145 21792
rect 17825 20704 18145 21728
rect 17825 20640 17833 20704
rect 17897 20640 17913 20704
rect 17977 20640 17993 20704
rect 18057 20640 18073 20704
rect 18137 20640 18145 20704
rect 17825 19616 18145 20640
rect 17825 19552 17833 19616
rect 17897 19552 17913 19616
rect 17977 19552 17993 19616
rect 18057 19552 18073 19616
rect 18137 19552 18145 19616
rect 17825 18528 18145 19552
rect 17825 18464 17833 18528
rect 17897 18464 17913 18528
rect 17977 18464 17993 18528
rect 18057 18464 18073 18528
rect 18137 18464 18145 18528
rect 17825 17440 18145 18464
rect 17825 17376 17833 17440
rect 17897 17376 17913 17440
rect 17977 17376 17993 17440
rect 18057 17376 18073 17440
rect 18137 17376 18145 17440
rect 17825 16352 18145 17376
rect 17825 16288 17833 16352
rect 17897 16288 17913 16352
rect 17977 16288 17993 16352
rect 18057 16288 18073 16352
rect 18137 16288 18145 16352
rect 17825 15264 18145 16288
rect 17825 15200 17833 15264
rect 17897 15200 17913 15264
rect 17977 15200 17993 15264
rect 18057 15200 18073 15264
rect 18137 15200 18145 15264
rect 17825 14176 18145 15200
rect 17825 14112 17833 14176
rect 17897 14112 17913 14176
rect 17977 14112 17993 14176
rect 18057 14112 18073 14176
rect 18137 14112 18145 14176
rect 17825 13088 18145 14112
rect 17825 13024 17833 13088
rect 17897 13024 17913 13088
rect 17977 13024 17993 13088
rect 18057 13024 18073 13088
rect 18137 13024 18145 13088
rect 17825 12000 18145 13024
rect 17825 11936 17833 12000
rect 17897 11936 17913 12000
rect 17977 11936 17993 12000
rect 18057 11936 18073 12000
rect 18137 11936 18145 12000
rect 17825 10912 18145 11936
rect 17825 10848 17833 10912
rect 17897 10848 17913 10912
rect 17977 10848 17993 10912
rect 18057 10848 18073 10912
rect 18137 10848 18145 10912
rect 17825 9824 18145 10848
rect 17825 9760 17833 9824
rect 17897 9760 17913 9824
rect 17977 9760 17993 9824
rect 18057 9760 18073 9824
rect 18137 9760 18145 9824
rect 17825 8736 18145 9760
rect 17825 8672 17833 8736
rect 17897 8672 17913 8736
rect 17977 8672 17993 8736
rect 18057 8672 18073 8736
rect 18137 8672 18145 8736
rect 17825 7648 18145 8672
rect 17825 7584 17833 7648
rect 17897 7584 17913 7648
rect 17977 7584 17993 7648
rect 18057 7584 18073 7648
rect 18137 7584 18145 7648
rect 17825 6560 18145 7584
rect 17825 6496 17833 6560
rect 17897 6496 17913 6560
rect 17977 6496 17993 6560
rect 18057 6496 18073 6560
rect 18137 6496 18145 6560
rect 17825 5472 18145 6496
rect 17825 5408 17833 5472
rect 17897 5408 17913 5472
rect 17977 5408 17993 5472
rect 18057 5408 18073 5472
rect 18137 5408 18145 5472
rect 17825 4384 18145 5408
rect 17825 4320 17833 4384
rect 17897 4320 17913 4384
rect 17977 4320 17993 4384
rect 18057 4320 18073 4384
rect 18137 4320 18145 4384
rect 17825 3296 18145 4320
rect 17825 3232 17833 3296
rect 17897 3232 17913 3296
rect 17977 3232 17993 3296
rect 18057 3232 18073 3296
rect 18137 3232 18145 3296
rect 17825 2208 18145 3232
rect 17825 2144 17833 2208
rect 17897 2144 17913 2208
rect 17977 2144 17993 2208
rect 18057 2144 18073 2208
rect 18137 2144 18145 2208
rect 17825 2128 18145 2144
rect 22046 33216 22366 33776
rect 22046 33152 22054 33216
rect 22118 33152 22134 33216
rect 22198 33152 22214 33216
rect 22278 33152 22294 33216
rect 22358 33152 22366 33216
rect 22046 32128 22366 33152
rect 22046 32064 22054 32128
rect 22118 32064 22134 32128
rect 22198 32064 22214 32128
rect 22278 32064 22294 32128
rect 22358 32064 22366 32128
rect 22046 31040 22366 32064
rect 22046 30976 22054 31040
rect 22118 30976 22134 31040
rect 22198 30976 22214 31040
rect 22278 30976 22294 31040
rect 22358 30976 22366 31040
rect 22046 29952 22366 30976
rect 26266 33760 26586 33776
rect 26266 33696 26274 33760
rect 26338 33696 26354 33760
rect 26418 33696 26434 33760
rect 26498 33696 26514 33760
rect 26578 33696 26586 33760
rect 26266 32672 26586 33696
rect 26266 32608 26274 32672
rect 26338 32608 26354 32672
rect 26418 32608 26434 32672
rect 26498 32608 26514 32672
rect 26578 32608 26586 32672
rect 26266 31584 26586 32608
rect 26266 31520 26274 31584
rect 26338 31520 26354 31584
rect 26418 31520 26434 31584
rect 26498 31520 26514 31584
rect 26578 31520 26586 31584
rect 24899 30836 24965 30837
rect 24899 30772 24900 30836
rect 24964 30772 24965 30836
rect 24899 30771 24965 30772
rect 22046 29888 22054 29952
rect 22118 29888 22134 29952
rect 22198 29888 22214 29952
rect 22278 29888 22294 29952
rect 22358 29888 22366 29952
rect 22046 28864 22366 29888
rect 22046 28800 22054 28864
rect 22118 28800 22134 28864
rect 22198 28800 22214 28864
rect 22278 28800 22294 28864
rect 22358 28800 22366 28864
rect 22046 27776 22366 28800
rect 22046 27712 22054 27776
rect 22118 27712 22134 27776
rect 22198 27712 22214 27776
rect 22278 27712 22294 27776
rect 22358 27712 22366 27776
rect 22046 26688 22366 27712
rect 22046 26624 22054 26688
rect 22118 26624 22134 26688
rect 22198 26624 22214 26688
rect 22278 26624 22294 26688
rect 22358 26624 22366 26688
rect 22046 25600 22366 26624
rect 22046 25536 22054 25600
rect 22118 25536 22134 25600
rect 22198 25536 22214 25600
rect 22278 25536 22294 25600
rect 22358 25536 22366 25600
rect 22046 24512 22366 25536
rect 22046 24448 22054 24512
rect 22118 24448 22134 24512
rect 22198 24448 22214 24512
rect 22278 24448 22294 24512
rect 22358 24448 22366 24512
rect 22046 23424 22366 24448
rect 22046 23360 22054 23424
rect 22118 23360 22134 23424
rect 22198 23360 22214 23424
rect 22278 23360 22294 23424
rect 22358 23360 22366 23424
rect 22046 22336 22366 23360
rect 24902 23221 24962 30771
rect 26266 30496 26586 31520
rect 26266 30432 26274 30496
rect 26338 30432 26354 30496
rect 26418 30432 26434 30496
rect 26498 30432 26514 30496
rect 26578 30432 26586 30496
rect 26266 29408 26586 30432
rect 26266 29344 26274 29408
rect 26338 29344 26354 29408
rect 26418 29344 26434 29408
rect 26498 29344 26514 29408
rect 26578 29344 26586 29408
rect 26266 28320 26586 29344
rect 26266 28256 26274 28320
rect 26338 28256 26354 28320
rect 26418 28256 26434 28320
rect 26498 28256 26514 28320
rect 26578 28256 26586 28320
rect 26266 27232 26586 28256
rect 26266 27168 26274 27232
rect 26338 27168 26354 27232
rect 26418 27168 26434 27232
rect 26498 27168 26514 27232
rect 26578 27168 26586 27232
rect 26266 26144 26586 27168
rect 26266 26080 26274 26144
rect 26338 26080 26354 26144
rect 26418 26080 26434 26144
rect 26498 26080 26514 26144
rect 26578 26080 26586 26144
rect 26266 25056 26586 26080
rect 26266 24992 26274 25056
rect 26338 24992 26354 25056
rect 26418 24992 26434 25056
rect 26498 24992 26514 25056
rect 26578 24992 26586 25056
rect 26266 23968 26586 24992
rect 26266 23904 26274 23968
rect 26338 23904 26354 23968
rect 26418 23904 26434 23968
rect 26498 23904 26514 23968
rect 26578 23904 26586 23968
rect 24899 23220 24965 23221
rect 24899 23156 24900 23220
rect 24964 23156 24965 23220
rect 24899 23155 24965 23156
rect 22046 22272 22054 22336
rect 22118 22272 22134 22336
rect 22198 22272 22214 22336
rect 22278 22272 22294 22336
rect 22358 22272 22366 22336
rect 22046 21248 22366 22272
rect 22046 21184 22054 21248
rect 22118 21184 22134 21248
rect 22198 21184 22214 21248
rect 22278 21184 22294 21248
rect 22358 21184 22366 21248
rect 22046 20160 22366 21184
rect 22046 20096 22054 20160
rect 22118 20096 22134 20160
rect 22198 20096 22214 20160
rect 22278 20096 22294 20160
rect 22358 20096 22366 20160
rect 22046 19072 22366 20096
rect 22046 19008 22054 19072
rect 22118 19008 22134 19072
rect 22198 19008 22214 19072
rect 22278 19008 22294 19072
rect 22358 19008 22366 19072
rect 22046 17984 22366 19008
rect 22046 17920 22054 17984
rect 22118 17920 22134 17984
rect 22198 17920 22214 17984
rect 22278 17920 22294 17984
rect 22358 17920 22366 17984
rect 22046 16896 22366 17920
rect 22046 16832 22054 16896
rect 22118 16832 22134 16896
rect 22198 16832 22214 16896
rect 22278 16832 22294 16896
rect 22358 16832 22366 16896
rect 22046 15808 22366 16832
rect 22046 15744 22054 15808
rect 22118 15744 22134 15808
rect 22198 15744 22214 15808
rect 22278 15744 22294 15808
rect 22358 15744 22366 15808
rect 22046 14720 22366 15744
rect 22046 14656 22054 14720
rect 22118 14656 22134 14720
rect 22198 14656 22214 14720
rect 22278 14656 22294 14720
rect 22358 14656 22366 14720
rect 22046 13632 22366 14656
rect 22046 13568 22054 13632
rect 22118 13568 22134 13632
rect 22198 13568 22214 13632
rect 22278 13568 22294 13632
rect 22358 13568 22366 13632
rect 22046 12544 22366 13568
rect 22046 12480 22054 12544
rect 22118 12480 22134 12544
rect 22198 12480 22214 12544
rect 22278 12480 22294 12544
rect 22358 12480 22366 12544
rect 22046 11456 22366 12480
rect 22046 11392 22054 11456
rect 22118 11392 22134 11456
rect 22198 11392 22214 11456
rect 22278 11392 22294 11456
rect 22358 11392 22366 11456
rect 22046 10368 22366 11392
rect 22046 10304 22054 10368
rect 22118 10304 22134 10368
rect 22198 10304 22214 10368
rect 22278 10304 22294 10368
rect 22358 10304 22366 10368
rect 22046 9280 22366 10304
rect 22046 9216 22054 9280
rect 22118 9216 22134 9280
rect 22198 9216 22214 9280
rect 22278 9216 22294 9280
rect 22358 9216 22366 9280
rect 22046 8192 22366 9216
rect 22046 8128 22054 8192
rect 22118 8128 22134 8192
rect 22198 8128 22214 8192
rect 22278 8128 22294 8192
rect 22358 8128 22366 8192
rect 22046 7104 22366 8128
rect 22046 7040 22054 7104
rect 22118 7040 22134 7104
rect 22198 7040 22214 7104
rect 22278 7040 22294 7104
rect 22358 7040 22366 7104
rect 22046 6016 22366 7040
rect 22046 5952 22054 6016
rect 22118 5952 22134 6016
rect 22198 5952 22214 6016
rect 22278 5952 22294 6016
rect 22358 5952 22366 6016
rect 22046 4928 22366 5952
rect 22046 4864 22054 4928
rect 22118 4864 22134 4928
rect 22198 4864 22214 4928
rect 22278 4864 22294 4928
rect 22358 4864 22366 4928
rect 22046 3840 22366 4864
rect 22046 3776 22054 3840
rect 22118 3776 22134 3840
rect 22198 3776 22214 3840
rect 22278 3776 22294 3840
rect 22358 3776 22366 3840
rect 22046 2752 22366 3776
rect 22046 2688 22054 2752
rect 22118 2688 22134 2752
rect 22198 2688 22214 2752
rect 22278 2688 22294 2752
rect 22358 2688 22366 2752
rect 22046 2128 22366 2688
rect 26266 22880 26586 23904
rect 26266 22816 26274 22880
rect 26338 22816 26354 22880
rect 26418 22816 26434 22880
rect 26498 22816 26514 22880
rect 26578 22816 26586 22880
rect 26266 21792 26586 22816
rect 26266 21728 26274 21792
rect 26338 21728 26354 21792
rect 26418 21728 26434 21792
rect 26498 21728 26514 21792
rect 26578 21728 26586 21792
rect 26266 20704 26586 21728
rect 26266 20640 26274 20704
rect 26338 20640 26354 20704
rect 26418 20640 26434 20704
rect 26498 20640 26514 20704
rect 26578 20640 26586 20704
rect 26266 19616 26586 20640
rect 26266 19552 26274 19616
rect 26338 19552 26354 19616
rect 26418 19552 26434 19616
rect 26498 19552 26514 19616
rect 26578 19552 26586 19616
rect 26266 18528 26586 19552
rect 26266 18464 26274 18528
rect 26338 18464 26354 18528
rect 26418 18464 26434 18528
rect 26498 18464 26514 18528
rect 26578 18464 26586 18528
rect 26266 17440 26586 18464
rect 26266 17376 26274 17440
rect 26338 17376 26354 17440
rect 26418 17376 26434 17440
rect 26498 17376 26514 17440
rect 26578 17376 26586 17440
rect 26266 16352 26586 17376
rect 26266 16288 26274 16352
rect 26338 16288 26354 16352
rect 26418 16288 26434 16352
rect 26498 16288 26514 16352
rect 26578 16288 26586 16352
rect 26266 15264 26586 16288
rect 26266 15200 26274 15264
rect 26338 15200 26354 15264
rect 26418 15200 26434 15264
rect 26498 15200 26514 15264
rect 26578 15200 26586 15264
rect 26266 14176 26586 15200
rect 26266 14112 26274 14176
rect 26338 14112 26354 14176
rect 26418 14112 26434 14176
rect 26498 14112 26514 14176
rect 26578 14112 26586 14176
rect 26266 13088 26586 14112
rect 26266 13024 26274 13088
rect 26338 13024 26354 13088
rect 26418 13024 26434 13088
rect 26498 13024 26514 13088
rect 26578 13024 26586 13088
rect 26266 12000 26586 13024
rect 26266 11936 26274 12000
rect 26338 11936 26354 12000
rect 26418 11936 26434 12000
rect 26498 11936 26514 12000
rect 26578 11936 26586 12000
rect 26266 10912 26586 11936
rect 26266 10848 26274 10912
rect 26338 10848 26354 10912
rect 26418 10848 26434 10912
rect 26498 10848 26514 10912
rect 26578 10848 26586 10912
rect 26266 9824 26586 10848
rect 26266 9760 26274 9824
rect 26338 9760 26354 9824
rect 26418 9760 26434 9824
rect 26498 9760 26514 9824
rect 26578 9760 26586 9824
rect 26266 8736 26586 9760
rect 26266 8672 26274 8736
rect 26338 8672 26354 8736
rect 26418 8672 26434 8736
rect 26498 8672 26514 8736
rect 26578 8672 26586 8736
rect 26266 7648 26586 8672
rect 26266 7584 26274 7648
rect 26338 7584 26354 7648
rect 26418 7584 26434 7648
rect 26498 7584 26514 7648
rect 26578 7584 26586 7648
rect 26266 6560 26586 7584
rect 26266 6496 26274 6560
rect 26338 6496 26354 6560
rect 26418 6496 26434 6560
rect 26498 6496 26514 6560
rect 26578 6496 26586 6560
rect 26266 5472 26586 6496
rect 26266 5408 26274 5472
rect 26338 5408 26354 5472
rect 26418 5408 26434 5472
rect 26498 5408 26514 5472
rect 26578 5408 26586 5472
rect 26266 4384 26586 5408
rect 26266 4320 26274 4384
rect 26338 4320 26354 4384
rect 26418 4320 26434 4384
rect 26498 4320 26514 4384
rect 26578 4320 26586 4384
rect 26266 3296 26586 4320
rect 26266 3232 26274 3296
rect 26338 3232 26354 3296
rect 26418 3232 26434 3296
rect 26498 3232 26514 3296
rect 26578 3232 26586 3296
rect 26266 2208 26586 3232
rect 26266 2144 26274 2208
rect 26338 2144 26354 2208
rect 26418 2144 26434 2208
rect 26498 2144 26514 2208
rect 26578 2144 26586 2208
rect 26266 2128 26586 2144
rect 30487 33216 30807 33776
rect 30487 33152 30495 33216
rect 30559 33152 30575 33216
rect 30639 33152 30655 33216
rect 30719 33152 30735 33216
rect 30799 33152 30807 33216
rect 30487 32128 30807 33152
rect 30487 32064 30495 32128
rect 30559 32064 30575 32128
rect 30639 32064 30655 32128
rect 30719 32064 30735 32128
rect 30799 32064 30807 32128
rect 30487 31040 30807 32064
rect 30487 30976 30495 31040
rect 30559 30976 30575 31040
rect 30639 30976 30655 31040
rect 30719 30976 30735 31040
rect 30799 30976 30807 31040
rect 30487 29952 30807 30976
rect 30487 29888 30495 29952
rect 30559 29888 30575 29952
rect 30639 29888 30655 29952
rect 30719 29888 30735 29952
rect 30799 29888 30807 29952
rect 30487 28864 30807 29888
rect 30487 28800 30495 28864
rect 30559 28800 30575 28864
rect 30639 28800 30655 28864
rect 30719 28800 30735 28864
rect 30799 28800 30807 28864
rect 30487 27776 30807 28800
rect 30487 27712 30495 27776
rect 30559 27712 30575 27776
rect 30639 27712 30655 27776
rect 30719 27712 30735 27776
rect 30799 27712 30807 27776
rect 30487 26688 30807 27712
rect 30487 26624 30495 26688
rect 30559 26624 30575 26688
rect 30639 26624 30655 26688
rect 30719 26624 30735 26688
rect 30799 26624 30807 26688
rect 30487 25600 30807 26624
rect 30487 25536 30495 25600
rect 30559 25536 30575 25600
rect 30639 25536 30655 25600
rect 30719 25536 30735 25600
rect 30799 25536 30807 25600
rect 30487 24512 30807 25536
rect 30487 24448 30495 24512
rect 30559 24448 30575 24512
rect 30639 24448 30655 24512
rect 30719 24448 30735 24512
rect 30799 24448 30807 24512
rect 30487 23424 30807 24448
rect 30487 23360 30495 23424
rect 30559 23360 30575 23424
rect 30639 23360 30655 23424
rect 30719 23360 30735 23424
rect 30799 23360 30807 23424
rect 30487 22336 30807 23360
rect 30487 22272 30495 22336
rect 30559 22272 30575 22336
rect 30639 22272 30655 22336
rect 30719 22272 30735 22336
rect 30799 22272 30807 22336
rect 30487 21248 30807 22272
rect 30487 21184 30495 21248
rect 30559 21184 30575 21248
rect 30639 21184 30655 21248
rect 30719 21184 30735 21248
rect 30799 21184 30807 21248
rect 30487 20160 30807 21184
rect 30487 20096 30495 20160
rect 30559 20096 30575 20160
rect 30639 20096 30655 20160
rect 30719 20096 30735 20160
rect 30799 20096 30807 20160
rect 30487 19072 30807 20096
rect 30487 19008 30495 19072
rect 30559 19008 30575 19072
rect 30639 19008 30655 19072
rect 30719 19008 30735 19072
rect 30799 19008 30807 19072
rect 30487 17984 30807 19008
rect 30487 17920 30495 17984
rect 30559 17920 30575 17984
rect 30639 17920 30655 17984
rect 30719 17920 30735 17984
rect 30799 17920 30807 17984
rect 30487 16896 30807 17920
rect 30487 16832 30495 16896
rect 30559 16832 30575 16896
rect 30639 16832 30655 16896
rect 30719 16832 30735 16896
rect 30799 16832 30807 16896
rect 30487 15808 30807 16832
rect 30487 15744 30495 15808
rect 30559 15744 30575 15808
rect 30639 15744 30655 15808
rect 30719 15744 30735 15808
rect 30799 15744 30807 15808
rect 30487 14720 30807 15744
rect 30487 14656 30495 14720
rect 30559 14656 30575 14720
rect 30639 14656 30655 14720
rect 30719 14656 30735 14720
rect 30799 14656 30807 14720
rect 30487 13632 30807 14656
rect 30487 13568 30495 13632
rect 30559 13568 30575 13632
rect 30639 13568 30655 13632
rect 30719 13568 30735 13632
rect 30799 13568 30807 13632
rect 30487 12544 30807 13568
rect 30487 12480 30495 12544
rect 30559 12480 30575 12544
rect 30639 12480 30655 12544
rect 30719 12480 30735 12544
rect 30799 12480 30807 12544
rect 30487 11456 30807 12480
rect 30487 11392 30495 11456
rect 30559 11392 30575 11456
rect 30639 11392 30655 11456
rect 30719 11392 30735 11456
rect 30799 11392 30807 11456
rect 30487 10368 30807 11392
rect 30487 10304 30495 10368
rect 30559 10304 30575 10368
rect 30639 10304 30655 10368
rect 30719 10304 30735 10368
rect 30799 10304 30807 10368
rect 30487 9280 30807 10304
rect 30487 9216 30495 9280
rect 30559 9216 30575 9280
rect 30639 9216 30655 9280
rect 30719 9216 30735 9280
rect 30799 9216 30807 9280
rect 30487 8192 30807 9216
rect 30487 8128 30495 8192
rect 30559 8128 30575 8192
rect 30639 8128 30655 8192
rect 30719 8128 30735 8192
rect 30799 8128 30807 8192
rect 30487 7104 30807 8128
rect 30487 7040 30495 7104
rect 30559 7040 30575 7104
rect 30639 7040 30655 7104
rect 30719 7040 30735 7104
rect 30799 7040 30807 7104
rect 30487 6016 30807 7040
rect 30487 5952 30495 6016
rect 30559 5952 30575 6016
rect 30639 5952 30655 6016
rect 30719 5952 30735 6016
rect 30799 5952 30807 6016
rect 30487 4928 30807 5952
rect 30487 4864 30495 4928
rect 30559 4864 30575 4928
rect 30639 4864 30655 4928
rect 30719 4864 30735 4928
rect 30799 4864 30807 4928
rect 30487 3840 30807 4864
rect 30487 3776 30495 3840
rect 30559 3776 30575 3840
rect 30639 3776 30655 3840
rect 30719 3776 30735 3840
rect 30799 3776 30807 3840
rect 30487 2752 30807 3776
rect 30487 2688 30495 2752
rect 30559 2688 30575 2752
rect 30639 2688 30655 2752
rect 30719 2688 30735 2752
rect 30799 2688 30807 2752
rect 30487 2128 30807 2688
rect 34707 33760 35027 33776
rect 34707 33696 34715 33760
rect 34779 33696 34795 33760
rect 34859 33696 34875 33760
rect 34939 33696 34955 33760
rect 35019 33696 35027 33760
rect 34707 32672 35027 33696
rect 34707 32608 34715 32672
rect 34779 32608 34795 32672
rect 34859 32608 34875 32672
rect 34939 32608 34955 32672
rect 35019 32608 35027 32672
rect 34707 31584 35027 32608
rect 34707 31520 34715 31584
rect 34779 31520 34795 31584
rect 34859 31520 34875 31584
rect 34939 31520 34955 31584
rect 35019 31520 35027 31584
rect 34707 30496 35027 31520
rect 34707 30432 34715 30496
rect 34779 30432 34795 30496
rect 34859 30432 34875 30496
rect 34939 30432 34955 30496
rect 35019 30432 35027 30496
rect 34707 29408 35027 30432
rect 34707 29344 34715 29408
rect 34779 29344 34795 29408
rect 34859 29344 34875 29408
rect 34939 29344 34955 29408
rect 35019 29344 35027 29408
rect 34707 28320 35027 29344
rect 34707 28256 34715 28320
rect 34779 28256 34795 28320
rect 34859 28256 34875 28320
rect 34939 28256 34955 28320
rect 35019 28256 35027 28320
rect 34707 27232 35027 28256
rect 34707 27168 34715 27232
rect 34779 27168 34795 27232
rect 34859 27168 34875 27232
rect 34939 27168 34955 27232
rect 35019 27168 35027 27232
rect 34707 26144 35027 27168
rect 34707 26080 34715 26144
rect 34779 26080 34795 26144
rect 34859 26080 34875 26144
rect 34939 26080 34955 26144
rect 35019 26080 35027 26144
rect 34707 25056 35027 26080
rect 34707 24992 34715 25056
rect 34779 24992 34795 25056
rect 34859 24992 34875 25056
rect 34939 24992 34955 25056
rect 35019 24992 35027 25056
rect 34707 23968 35027 24992
rect 34707 23904 34715 23968
rect 34779 23904 34795 23968
rect 34859 23904 34875 23968
rect 34939 23904 34955 23968
rect 35019 23904 35027 23968
rect 34707 22880 35027 23904
rect 34707 22816 34715 22880
rect 34779 22816 34795 22880
rect 34859 22816 34875 22880
rect 34939 22816 34955 22880
rect 35019 22816 35027 22880
rect 34707 21792 35027 22816
rect 34707 21728 34715 21792
rect 34779 21728 34795 21792
rect 34859 21728 34875 21792
rect 34939 21728 34955 21792
rect 35019 21728 35027 21792
rect 34707 20704 35027 21728
rect 34707 20640 34715 20704
rect 34779 20640 34795 20704
rect 34859 20640 34875 20704
rect 34939 20640 34955 20704
rect 35019 20640 35027 20704
rect 34707 19616 35027 20640
rect 34707 19552 34715 19616
rect 34779 19552 34795 19616
rect 34859 19552 34875 19616
rect 34939 19552 34955 19616
rect 35019 19552 35027 19616
rect 34707 18528 35027 19552
rect 34707 18464 34715 18528
rect 34779 18464 34795 18528
rect 34859 18464 34875 18528
rect 34939 18464 34955 18528
rect 35019 18464 35027 18528
rect 34707 17440 35027 18464
rect 34707 17376 34715 17440
rect 34779 17376 34795 17440
rect 34859 17376 34875 17440
rect 34939 17376 34955 17440
rect 35019 17376 35027 17440
rect 34707 16352 35027 17376
rect 34707 16288 34715 16352
rect 34779 16288 34795 16352
rect 34859 16288 34875 16352
rect 34939 16288 34955 16352
rect 35019 16288 35027 16352
rect 34707 15264 35027 16288
rect 34707 15200 34715 15264
rect 34779 15200 34795 15264
rect 34859 15200 34875 15264
rect 34939 15200 34955 15264
rect 35019 15200 35027 15264
rect 34707 14176 35027 15200
rect 34707 14112 34715 14176
rect 34779 14112 34795 14176
rect 34859 14112 34875 14176
rect 34939 14112 34955 14176
rect 35019 14112 35027 14176
rect 34707 13088 35027 14112
rect 34707 13024 34715 13088
rect 34779 13024 34795 13088
rect 34859 13024 34875 13088
rect 34939 13024 34955 13088
rect 35019 13024 35027 13088
rect 34707 12000 35027 13024
rect 34707 11936 34715 12000
rect 34779 11936 34795 12000
rect 34859 11936 34875 12000
rect 34939 11936 34955 12000
rect 35019 11936 35027 12000
rect 34707 10912 35027 11936
rect 34707 10848 34715 10912
rect 34779 10848 34795 10912
rect 34859 10848 34875 10912
rect 34939 10848 34955 10912
rect 35019 10848 35027 10912
rect 34707 9824 35027 10848
rect 34707 9760 34715 9824
rect 34779 9760 34795 9824
rect 34859 9760 34875 9824
rect 34939 9760 34955 9824
rect 35019 9760 35027 9824
rect 34707 8736 35027 9760
rect 34707 8672 34715 8736
rect 34779 8672 34795 8736
rect 34859 8672 34875 8736
rect 34939 8672 34955 8736
rect 35019 8672 35027 8736
rect 34707 7648 35027 8672
rect 34707 7584 34715 7648
rect 34779 7584 34795 7648
rect 34859 7584 34875 7648
rect 34939 7584 34955 7648
rect 35019 7584 35027 7648
rect 34707 6560 35027 7584
rect 34707 6496 34715 6560
rect 34779 6496 34795 6560
rect 34859 6496 34875 6560
rect 34939 6496 34955 6560
rect 35019 6496 35027 6560
rect 34707 5472 35027 6496
rect 34707 5408 34715 5472
rect 34779 5408 34795 5472
rect 34859 5408 34875 5472
rect 34939 5408 34955 5472
rect 35019 5408 35027 5472
rect 34707 4384 35027 5408
rect 34707 4320 34715 4384
rect 34779 4320 34795 4384
rect 34859 4320 34875 4384
rect 34939 4320 34955 4384
rect 35019 4320 35027 4384
rect 34707 3296 35027 4320
rect 34707 3232 34715 3296
rect 34779 3232 34795 3296
rect 34859 3232 34875 3296
rect 34939 3232 34955 3296
rect 35019 3232 35027 3296
rect 34707 2208 35027 3232
rect 34707 2144 34715 2208
rect 34779 2144 34795 2208
rect 34859 2144 34875 2208
rect 34939 2144 34955 2208
rect 35019 2144 35027 2208
rect 34707 2128 35027 2144
use sky130_fd_sc_hd__fill_2  FILLER_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 1380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 2116 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 2484 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 3128 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29
timestamp 1666464484
transform 1 0 3772 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37
timestamp 1666464484
transform 1 0 4508 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43
timestamp 1666464484
transform 1 0 5060 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50
timestamp 1666464484
transform 1 0 5704 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57
timestamp 1666464484
transform 1 0 6348 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_62 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 6808 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_70
timestamp 1666464484
transform 1 0 7544 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_75
timestamp 1666464484
transform 1 0 8004 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_83
timestamp 1666464484
transform 1 0 8740 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_85
timestamp 1666464484
transform 1 0 8924 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_90
timestamp 1666464484
transform 1 0 9384 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_98
timestamp 1666464484
transform 1 0 10120 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_103
timestamp 1666464484
transform 1 0 10580 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_111
timestamp 1666464484
transform 1 0 11316 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_113
timestamp 1666464484
transform 1 0 11500 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_118
timestamp 1666464484
transform 1 0 11960 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_126
timestamp 1666464484
transform 1 0 12696 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_131
timestamp 1666464484
transform 1 0 13156 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_139
timestamp 1666464484
transform 1 0 13892 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_141
timestamp 1666464484
transform 1 0 14076 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_149
timestamp 1666464484
transform 1 0 14812 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_155
timestamp 1666464484
transform 1 0 15364 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_162
timestamp 1666464484
transform 1 0 16008 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_169
timestamp 1666464484
transform 1 0 16652 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_177
timestamp 1666464484
transform 1 0 17388 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_183
timestamp 1666464484
transform 1 0 17940 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_190
timestamp 1666464484
transform 1 0 18584 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_197
timestamp 1666464484
transform 1 0 19228 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_205
timestamp 1666464484
transform 1 0 19964 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_211
timestamp 1666464484
transform 1 0 20516 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_218
timestamp 1666464484
transform 1 0 21160 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_225
timestamp 1666464484
transform 1 0 21804 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_233
timestamp 1666464484
transform 1 0 22540 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_239
timestamp 1666464484
transform 1 0 23092 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_246
timestamp 1666464484
transform 1 0 23736 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_253
timestamp 1666464484
transform 1 0 24380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_261
timestamp 1666464484
transform 1 0 25116 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_267
timestamp 1666464484
transform 1 0 25668 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_274
timestamp 1666464484
transform 1 0 26312 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_281
timestamp 1666464484
transform 1 0 26956 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_289
timestamp 1666464484
transform 1 0 27692 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_295
timestamp 1666464484
transform 1 0 28244 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_302
timestamp 1666464484
transform 1 0 28888 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_309
timestamp 1666464484
transform 1 0 29532 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_314
timestamp 1666464484
transform 1 0 29992 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_322
timestamp 1666464484
transform 1 0 30728 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_327
timestamp 1666464484
transform 1 0 31188 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_335
timestamp 1666464484
transform 1 0 31924 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_337
timestamp 1666464484
transform 1 0 32108 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_342
timestamp 1666464484
transform 1 0 32568 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_350
timestamp 1666464484
transform 1 0 33304 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_355
timestamp 1666464484
transform 1 0 33764 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_362
timestamp 1666464484
transform 1 0 34408 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_15
timestamp 1666464484
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_27
timestamp 1666464484
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_39
timestamp 1666464484
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_51
timestamp 1666464484
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1666464484
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_57
timestamp 1666464484
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_69
timestamp 1666464484
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_81
timestamp 1666464484
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_93
timestamp 1666464484
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_105
timestamp 1666464484
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 1666464484
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_113
timestamp 1666464484
transform 1 0 11500 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_121
timestamp 1666464484
transform 1 0 12236 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_126
timestamp 1666464484
transform 1 0 12696 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_138
timestamp 1666464484
transform 1 0 13800 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_149
timestamp 1666464484
transform 1 0 14812 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_156
timestamp 1666464484
transform 1 0 15456 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_1_169 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 16652 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_1_181
timestamp 1666464484
transform 1 0 17756 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_193
timestamp 1666464484
transform 1 0 18860 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_1_204
timestamp 1666464484
transform 1 0 19872 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_212
timestamp 1666464484
transform 1 0 20608 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_219
timestamp 1666464484
transform 1 0 21252 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_223
timestamp 1666464484
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_225
timestamp 1666464484
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_237
timestamp 1666464484
transform 1 0 22908 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_249
timestamp 1666464484
transform 1 0 24012 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_272
timestamp 1666464484
transform 1 0 26128 0 -1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_1_281
timestamp 1666464484
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_293
timestamp 1666464484
transform 1 0 28060 0 -1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_1_319
timestamp 1666464484
transform 1 0 30452 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_331
timestamp 1666464484
transform 1 0 31556 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_335
timestamp 1666464484
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_337
timestamp 1666464484
transform 1 0 32108 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_349
timestamp 1666464484
transform 1 0 33212 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_1_361
timestamp 1666464484
transform 1 0 34316 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3
timestamp 1666464484
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_15
timestamp 1666464484
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1666464484
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1666464484
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_41
timestamp 1666464484
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_53
timestamp 1666464484
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_65
timestamp 1666464484
transform 1 0 7084 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_2_78
timestamp 1666464484
transform 1 0 8280 0 1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 1666464484
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_97
timestamp 1666464484
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_109
timestamp 1666464484
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_121
timestamp 1666464484
transform 1 0 12236 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_138
timestamp 1666464484
transform 1 0 13800 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_141
timestamp 1666464484
transform 1 0 14076 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_159
timestamp 1666464484
transform 1 0 15732 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_167
timestamp 1666464484
transform 1 0 16468 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_185
timestamp 1666464484
transform 1 0 18124 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_193
timestamp 1666464484
transform 1 0 18860 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_197
timestamp 1666464484
transform 1 0 19228 0 1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_2_216
timestamp 1666464484
transform 1 0 20976 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_237
timestamp 1666464484
transform 1 0 22908 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_2_249
timestamp 1666464484
transform 1 0 24012 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_253
timestamp 1666464484
transform 1 0 24380 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_271
timestamp 1666464484
transform 1 0 26036 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_286
timestamp 1666464484
transform 1 0 27416 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_296
timestamp 1666464484
transform 1 0 28336 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_309
timestamp 1666464484
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_321
timestamp 1666464484
transform 1 0 30636 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_333
timestamp 1666464484
transform 1 0 31740 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_345
timestamp 1666464484
transform 1 0 32844 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_357
timestamp 1666464484
transform 1 0 33948 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_363
timestamp 1666464484
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 1666464484
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_15
timestamp 1666464484
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_27
timestamp 1666464484
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_39
timestamp 1666464484
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_51
timestamp 1666464484
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1666464484
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_57
timestamp 1666464484
transform 1 0 6348 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_63
timestamp 1666464484
transform 1 0 6900 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_84
timestamp 1666464484
transform 1 0 8832 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_97
timestamp 1666464484
transform 1 0 10028 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_106
timestamp 1666464484
transform 1 0 10856 0 -1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 1666464484
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_125
timestamp 1666464484
transform 1 0 12604 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_3_138
timestamp 1666464484
transform 1 0 13800 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_166
timestamp 1666464484
transform 1 0 16376 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_169
timestamp 1666464484
transform 1 0 16652 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_3_174
timestamp 1666464484
transform 1 0 17112 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_3_196
timestamp 1666464484
transform 1 0 19136 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_204
timestamp 1666464484
transform 1 0 19872 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_222
timestamp 1666464484
transform 1 0 21528 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_225
timestamp 1666464484
transform 1 0 21804 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_243
timestamp 1666464484
transform 1 0 23460 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_251
timestamp 1666464484
transform 1 0 24196 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_268
timestamp 1666464484
transform 1 0 25760 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_278
timestamp 1666464484
transform 1 0 26680 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_281
timestamp 1666464484
transform 1 0 26956 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_299
timestamp 1666464484
transform 1 0 28612 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_311
timestamp 1666464484
transform 1 0 29716 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_323
timestamp 1666464484
transform 1 0 30820 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_335
timestamp 1666464484
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_337
timestamp 1666464484
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_349
timestamp 1666464484
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_3_361
timestamp 1666464484
transform 1 0 34316 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1666464484
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 1666464484
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1666464484
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1666464484
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1666464484
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_53
timestamp 1666464484
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_65
timestamp 1666464484
transform 1 0 7084 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_82
timestamp 1666464484
transform 1 0 8648 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_85
timestamp 1666464484
transform 1 0 8924 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_107
timestamp 1666464484
transform 1 0 10948 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_115
timestamp 1666464484
transform 1 0 11684 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_124
timestamp 1666464484
transform 1 0 12512 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_136
timestamp 1666464484
transform 1 0 13616 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_141
timestamp 1666464484
transform 1 0 14076 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_147
timestamp 1666464484
transform 1 0 14628 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_155
timestamp 1666464484
transform 1 0 15364 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_166
timestamp 1666464484
transform 1 0 16376 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_174
timestamp 1666464484
transform 1 0 17112 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_180
timestamp 1666464484
transform 1 0 17664 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_4_193
timestamp 1666464484
transform 1 0 18860 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_4_197
timestamp 1666464484
transform 1 0 19228 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_4_212
timestamp 1666464484
transform 1 0 20608 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_220
timestamp 1666464484
transform 1 0 21344 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_224
timestamp 1666464484
transform 1 0 21712 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_231
timestamp 1666464484
transform 1 0 22356 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_243
timestamp 1666464484
transform 1 0 23460 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_251
timestamp 1666464484
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_253
timestamp 1666464484
transform 1 0 24380 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_261
timestamp 1666464484
transform 1 0 25116 0 1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_4_285
timestamp 1666464484
transform 1 0 27324 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_297
timestamp 1666464484
transform 1 0 28428 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_305
timestamp 1666464484
transform 1 0 29164 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_309
timestamp 1666464484
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_321
timestamp 1666464484
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_333
timestamp 1666464484
transform 1 0 31740 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_345
timestamp 1666464484
transform 1 0 32844 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_357
timestamp 1666464484
transform 1 0 33948 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_363
timestamp 1666464484
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3
timestamp 1666464484
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_15
timestamp 1666464484
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_27
timestamp 1666464484
transform 1 0 3588 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_36
timestamp 1666464484
transform 1 0 4416 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_44
timestamp 1666464484
transform 1 0 5152 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_51
timestamp 1666464484
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1666464484
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1666464484
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1666464484
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_81
timestamp 1666464484
transform 1 0 8556 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_96
timestamp 1666464484
transform 1 0 9936 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_103
timestamp 1666464484
transform 1 0 10580 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1666464484
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_113
timestamp 1666464484
transform 1 0 11500 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_131
timestamp 1666464484
transform 1 0 13156 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_143
timestamp 1666464484
transform 1 0 14260 0 -1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_5_154
timestamp 1666464484
transform 1 0 15272 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_166
timestamp 1666464484
transform 1 0 16376 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_169
timestamp 1666464484
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_181
timestamp 1666464484
transform 1 0 17756 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_185
timestamp 1666464484
transform 1 0 18124 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_206
timestamp 1666464484
transform 1 0 20056 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_218
timestamp 1666464484
transform 1 0 21160 0 -1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_5_225
timestamp 1666464484
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_237
timestamp 1666464484
transform 1 0 22908 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_241
timestamp 1666464484
transform 1 0 23276 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_262
timestamp 1666464484
transform 1 0 25208 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_271
timestamp 1666464484
transform 1 0 26036 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_279
timestamp 1666464484
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_281
timestamp 1666464484
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_293
timestamp 1666464484
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_305
timestamp 1666464484
transform 1 0 29164 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_317
timestamp 1666464484
transform 1 0 30268 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_329
timestamp 1666464484
transform 1 0 31372 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_335
timestamp 1666464484
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_337
timestamp 1666464484
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_349
timestamp 1666464484
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_5_361
timestamp 1666464484
transform 1 0 34316 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3
timestamp 1666464484
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_15
timestamp 1666464484
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1666464484
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_29
timestamp 1666464484
transform 1 0 3772 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_55
timestamp 1666464484
transform 1 0 6164 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_67
timestamp 1666464484
transform 1 0 7268 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_79
timestamp 1666464484
transform 1 0 8372 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1666464484
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1666464484
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_97
timestamp 1666464484
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_109
timestamp 1666464484
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_121
timestamp 1666464484
transform 1 0 12236 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_129
timestamp 1666464484
transform 1 0 12972 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_6_137
timestamp 1666464484
transform 1 0 13708 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_6_141
timestamp 1666464484
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_153
timestamp 1666464484
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_165
timestamp 1666464484
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_177
timestamp 1666464484
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_189
timestamp 1666464484
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1666464484
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_197
timestamp 1666464484
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_209
timestamp 1666464484
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_221
timestamp 1666464484
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_233
timestamp 1666464484
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_245
timestamp 1666464484
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp 1666464484
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_253
timestamp 1666464484
transform 1 0 24380 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_271
timestamp 1666464484
transform 1 0 26036 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_283
timestamp 1666464484
transform 1 0 27140 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_295
timestamp 1666464484
transform 1 0 28244 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_299
timestamp 1666464484
transform 1 0 28612 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_306
timestamp 1666464484
transform 1 0 29256 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_309
timestamp 1666464484
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_321
timestamp 1666464484
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_333
timestamp 1666464484
transform 1 0 31740 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_345
timestamp 1666464484
transform 1 0 32844 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_357
timestamp 1666464484
transform 1 0 33948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_363
timestamp 1666464484
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 1666464484
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_7_15
timestamp 1666464484
transform 1 0 2484 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_23
timestamp 1666464484
transform 1 0 3220 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_31
timestamp 1666464484
transform 1 0 3956 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_43
timestamp 1666464484
transform 1 0 5060 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1666464484
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_57
timestamp 1666464484
transform 1 0 6348 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_68
timestamp 1666464484
transform 1 0 7360 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_80
timestamp 1666464484
transform 1 0 8464 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_92
timestamp 1666464484
transform 1 0 9568 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_104
timestamp 1666464484
transform 1 0 10672 0 -1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_7_113
timestamp 1666464484
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_134
timestamp 1666464484
transform 1 0 13432 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_146
timestamp 1666464484
transform 1 0 14536 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_158
timestamp 1666464484
transform 1 0 15640 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_166
timestamp 1666464484
transform 1 0 16376 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_169
timestamp 1666464484
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_181
timestamp 1666464484
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_193
timestamp 1666464484
transform 1 0 18860 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_199
timestamp 1666464484
transform 1 0 19412 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_216
timestamp 1666464484
transform 1 0 20976 0 -1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_7_225
timestamp 1666464484
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_237
timestamp 1666464484
transform 1 0 22908 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_243
timestamp 1666464484
transform 1 0 23460 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_260
timestamp 1666464484
transform 1 0 25024 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_272
timestamp 1666464484
transform 1 0 26128 0 -1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_7_281
timestamp 1666464484
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_293
timestamp 1666464484
transform 1 0 28060 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_313
timestamp 1666464484
transform 1 0 29900 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_325
timestamp 1666464484
transform 1 0 31004 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_7_333
timestamp 1666464484
transform 1 0 31740 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_7_337
timestamp 1666464484
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_349
timestamp 1666464484
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_7_361
timestamp 1666464484
transform 1 0 34316 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_3
timestamp 1666464484
transform 1 0 1380 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_26
timestamp 1666464484
transform 1 0 3496 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1666464484
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_41
timestamp 1666464484
transform 1 0 4876 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_8_63
timestamp 1666464484
transform 1 0 6900 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_76
timestamp 1666464484
transform 1 0 8096 0 1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_8_85
timestamp 1666464484
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_109
timestamp 1666464484
transform 1 0 11132 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_8_131
timestamp 1666464484
transform 1 0 13156 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_138
timestamp 1666464484
transform 1 0 13800 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_141
timestamp 1666464484
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_153
timestamp 1666464484
transform 1 0 15180 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_173
timestamp 1666464484
transform 1 0 17020 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_8_183
timestamp 1666464484
transform 1 0 17940 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1666464484
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_197
timestamp 1666464484
transform 1 0 19228 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_215
timestamp 1666464484
transform 1 0 20884 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_235
timestamp 1666464484
transform 1 0 22724 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_243
timestamp 1666464484
transform 1 0 23460 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_250
timestamp 1666464484
transform 1 0 24104 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_253
timestamp 1666464484
transform 1 0 24380 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_271
timestamp 1666464484
transform 1 0 26036 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_283
timestamp 1666464484
transform 1 0 27140 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_289
timestamp 1666464484
transform 1 0 27692 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_306
timestamp 1666464484
transform 1 0 29256 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_8_309
timestamp 1666464484
transform 1 0 29532 0 1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_8_331
timestamp 1666464484
transform 1 0 31556 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_343
timestamp 1666464484
transform 1 0 32660 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_355
timestamp 1666464484
transform 1 0 33764 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_363
timestamp 1666464484
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3
timestamp 1666464484
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_18
timestamp 1666464484
transform 1 0 2760 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_30
timestamp 1666464484
transform 1 0 3864 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_42
timestamp 1666464484
transform 1 0 4968 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_54
timestamp 1666464484
transform 1 0 6072 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_57
timestamp 1666464484
transform 1 0 6348 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_9_79
timestamp 1666464484
transform 1 0 8372 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp 1666464484
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1666464484
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_9_113
timestamp 1666464484
transform 1 0 11500 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_125
timestamp 1666464484
transform 1 0 12604 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_149
timestamp 1666464484
transform 1 0 14812 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_155
timestamp 1666464484
transform 1 0 15364 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_162
timestamp 1666464484
transform 1 0 16008 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_9_169
timestamp 1666464484
transform 1 0 16652 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_175
timestamp 1666464484
transform 1 0 17204 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_182
timestamp 1666464484
transform 1 0 17848 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_206
timestamp 1666464484
transform 1 0 20056 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_216
timestamp 1666464484
transform 1 0 20976 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_225
timestamp 1666464484
transform 1 0 21804 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_233
timestamp 1666464484
transform 1 0 22540 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_241
timestamp 1666464484
transform 1 0 23276 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_262
timestamp 1666464484
transform 1 0 25208 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_272
timestamp 1666464484
transform 1 0 26128 0 -1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_9_281
timestamp 1666464484
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_293
timestamp 1666464484
transform 1 0 28060 0 -1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_9_319
timestamp 1666464484
transform 1 0 30452 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_331
timestamp 1666464484
transform 1 0 31556 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_335
timestamp 1666464484
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_337
timestamp 1666464484
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_349
timestamp 1666464484
transform 1 0 33212 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_361
timestamp 1666464484
transform 1 0 34316 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3
timestamp 1666464484
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_15
timestamp 1666464484
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1666464484
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_29
timestamp 1666464484
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_41
timestamp 1666464484
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_53
timestamp 1666464484
transform 1 0 5980 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_61
timestamp 1666464484
transform 1 0 6716 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_10_69
timestamp 1666464484
transform 1 0 7452 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_10_81
timestamp 1666464484
transform 1 0 8556 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_10_85
timestamp 1666464484
transform 1 0 8924 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_93
timestamp 1666464484
transform 1 0 9660 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_100
timestamp 1666464484
transform 1 0 10304 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_112
timestamp 1666464484
transform 1 0 11408 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_124
timestamp 1666464484
transform 1 0 12512 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_136
timestamp 1666464484
transform 1 0 13616 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_10_141
timestamp 1666464484
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_153
timestamp 1666464484
transform 1 0 15180 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_161
timestamp 1666464484
transform 1 0 15916 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_184
timestamp 1666464484
transform 1 0 18032 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_194
timestamp 1666464484
transform 1 0 18952 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_197
timestamp 1666464484
transform 1 0 19228 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_219
timestamp 1666464484
transform 1 0 21252 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_243
timestamp 1666464484
transform 1 0 23460 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_251
timestamp 1666464484
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_253
timestamp 1666464484
transform 1 0 24380 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_275
timestamp 1666464484
transform 1 0 26404 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_287
timestamp 1666464484
transform 1 0 27508 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_10_299
timestamp 1666464484
transform 1 0 28612 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_307
timestamp 1666464484
transform 1 0 29348 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_309
timestamp 1666464484
transform 1 0 29532 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_331
timestamp 1666464484
transform 1 0 31556 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_355
timestamp 1666464484
transform 1 0 33764 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_363
timestamp 1666464484
transform 1 0 34500 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3
timestamp 1666464484
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_15
timestamp 1666464484
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_27
timestamp 1666464484
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_39
timestamp 1666464484
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_51
timestamp 1666464484
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1666464484
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_57
timestamp 1666464484
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_69
timestamp 1666464484
transform 1 0 7452 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_11_93
timestamp 1666464484
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_105
timestamp 1666464484
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1666464484
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_113
timestamp 1666464484
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_125
timestamp 1666464484
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_137
timestamp 1666464484
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_11_149
timestamp 1666464484
transform 1 0 14812 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_166
timestamp 1666464484
transform 1 0 16376 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_11_169
timestamp 1666464484
transform 1 0 16652 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_175
timestamp 1666464484
transform 1 0 17204 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_182
timestamp 1666464484
transform 1 0 17848 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_206
timestamp 1666464484
transform 1 0 20056 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_217
timestamp 1666464484
transform 1 0 21068 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_223
timestamp 1666464484
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_225
timestamp 1666464484
transform 1 0 21804 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_233
timestamp 1666464484
transform 1 0 22540 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_241
timestamp 1666464484
transform 1 0 23276 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_261
timestamp 1666464484
transform 1 0 25116 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_271
timestamp 1666464484
transform 1 0 26036 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_279
timestamp 1666464484
transform 1 0 26772 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_281
timestamp 1666464484
transform 1 0 26956 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_293
timestamp 1666464484
transform 1 0 28060 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_11_315
timestamp 1666464484
transform 1 0 30084 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_325
timestamp 1666464484
transform 1 0 31004 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_333
timestamp 1666464484
transform 1 0 31740 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_337
timestamp 1666464484
transform 1 0 32108 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_355
timestamp 1666464484
transform 1 0 33764 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_363
timestamp 1666464484
transform 1 0 34500 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3
timestamp 1666464484
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_15
timestamp 1666464484
transform 1 0 2484 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_25
timestamp 1666464484
transform 1 0 3404 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_29
timestamp 1666464484
transform 1 0 3772 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_37
timestamp 1666464484
transform 1 0 4508 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_49
timestamp 1666464484
transform 1 0 5612 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_61
timestamp 1666464484
transform 1 0 6716 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_73
timestamp 1666464484
transform 1 0 7820 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_12_81
timestamp 1666464484
transform 1 0 8556 0 1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_12_85
timestamp 1666464484
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_97
timestamp 1666464484
transform 1 0 10028 0 1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_12_121
timestamp 1666464484
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_133
timestamp 1666464484
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1666464484
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_141
timestamp 1666464484
transform 1 0 14076 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_149
timestamp 1666464484
transform 1 0 14812 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_167
timestamp 1666464484
transform 1 0 16468 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_187
timestamp 1666464484
transform 1 0 18308 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_195
timestamp 1666464484
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_197
timestamp 1666464484
transform 1 0 19228 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_203
timestamp 1666464484
transform 1 0 19780 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_220
timestamp 1666464484
transform 1 0 21344 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_238
timestamp 1666464484
transform 1 0 23000 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_250
timestamp 1666464484
transform 1 0 24104 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_253
timestamp 1666464484
transform 1 0 24380 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_261
timestamp 1666464484
transform 1 0 25116 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_273
timestamp 1666464484
transform 1 0 26220 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_285
timestamp 1666464484
transform 1 0 27324 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_12_297
timestamp 1666464484
transform 1 0 28428 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_306
timestamp 1666464484
transform 1 0 29256 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_309
timestamp 1666464484
transform 1 0 29532 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_317
timestamp 1666464484
transform 1 0 30268 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_329
timestamp 1666464484
transform 1 0 31372 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_337
timestamp 1666464484
transform 1 0 32108 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_355
timestamp 1666464484
transform 1 0 33764 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_363
timestamp 1666464484
transform 1 0 34500 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_3
timestamp 1666464484
transform 1 0 1380 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_13_15
timestamp 1666464484
transform 1 0 2484 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_28
timestamp 1666464484
transform 1 0 3680 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_35
timestamp 1666464484
transform 1 0 4324 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_42
timestamp 1666464484
transform 1 0 4968 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_54
timestamp 1666464484
transform 1 0 6072 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_57
timestamp 1666464484
transform 1 0 6348 0 -1 9792
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_13_81
timestamp 1666464484
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_93
timestamp 1666464484
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_105
timestamp 1666464484
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1666464484
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_113
timestamp 1666464484
transform 1 0 11500 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_131
timestamp 1666464484
transform 1 0 13156 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_143
timestamp 1666464484
transform 1 0 14260 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_155
timestamp 1666464484
transform 1 0 15364 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1666464484
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_169
timestamp 1666464484
transform 1 0 16652 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_177
timestamp 1666464484
transform 1 0 17388 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_185
timestamp 1666464484
transform 1 0 18124 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_193
timestamp 1666464484
transform 1 0 18860 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_13_206
timestamp 1666464484
transform 1 0 20056 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_13_220
timestamp 1666464484
transform 1 0 21344 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_225
timestamp 1666464484
transform 1 0 21804 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_233
timestamp 1666464484
transform 1 0 22540 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_245
timestamp 1666464484
transform 1 0 23644 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_257
timestamp 1666464484
transform 1 0 24748 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_269
timestamp 1666464484
transform 1 0 25852 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_277
timestamp 1666464484
transform 1 0 26588 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_281
timestamp 1666464484
transform 1 0 26956 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_290
timestamp 1666464484
transform 1 0 27784 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_302
timestamp 1666464484
transform 1 0 28888 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_314
timestamp 1666464484
transform 1 0 29992 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_326
timestamp 1666464484
transform 1 0 31096 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_334
timestamp 1666464484
transform 1 0 31832 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_337
timestamp 1666464484
transform 1 0 32108 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_359
timestamp 1666464484
transform 1 0 34132 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_363
timestamp 1666464484
transform 1 0 34500 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_3
timestamp 1666464484
transform 1 0 1380 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_13
timestamp 1666464484
transform 1 0 2300 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_14_25
timestamp 1666464484
transform 1 0 3404 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_29
timestamp 1666464484
transform 1 0 3772 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_37
timestamp 1666464484
transform 1 0 4508 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_45
timestamp 1666464484
transform 1 0 5244 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_62
timestamp 1666464484
transform 1 0 6808 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_82
timestamp 1666464484
transform 1 0 8648 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_85
timestamp 1666464484
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_97
timestamp 1666464484
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_109
timestamp 1666464484
transform 1 0 11132 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_126
timestamp 1666464484
transform 1 0 12696 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_138
timestamp 1666464484
transform 1 0 13800 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_141
timestamp 1666464484
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_153
timestamp 1666464484
transform 1 0 15180 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_165
timestamp 1666464484
transform 1 0 16284 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_177
timestamp 1666464484
transform 1 0 17388 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_189
timestamp 1666464484
transform 1 0 18492 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_195
timestamp 1666464484
transform 1 0 19044 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_197
timestamp 1666464484
transform 1 0 19228 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_209
timestamp 1666464484
transform 1 0 20332 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_213
timestamp 1666464484
transform 1 0 20700 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_234
timestamp 1666464484
transform 1 0 22632 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_246
timestamp 1666464484
transform 1 0 23736 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_14_253
timestamp 1666464484
transform 1 0 24380 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_14_267
timestamp 1666464484
transform 1 0 25668 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_291
timestamp 1666464484
transform 1 0 27876 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_303
timestamp 1666464484
transform 1 0 28980 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_307
timestamp 1666464484
transform 1 0 29348 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_309
timestamp 1666464484
transform 1 0 29532 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_318
timestamp 1666464484
transform 1 0 30360 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_326
timestamp 1666464484
transform 1 0 31096 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_347
timestamp 1666464484
transform 1 0 33028 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_357
timestamp 1666464484
transform 1 0 33948 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_363
timestamp 1666464484
transform 1 0 34500 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_3
timestamp 1666464484
transform 1 0 1380 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_11
timestamp 1666464484
transform 1 0 2116 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_16
timestamp 1666464484
transform 1 0 2576 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_27
timestamp 1666464484
transform 1 0 3588 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_36
timestamp 1666464484
transform 1 0 4416 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_48
timestamp 1666464484
transform 1 0 5520 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_57
timestamp 1666464484
transform 1 0 6348 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_77
timestamp 1666464484
transform 1 0 8188 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_99
timestamp 1666464484
transform 1 0 10212 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1666464484
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_113
timestamp 1666464484
transform 1 0 11500 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_121
timestamp 1666464484
transform 1 0 12236 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_140
timestamp 1666464484
transform 1 0 13984 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_152
timestamp 1666464484
transform 1 0 15088 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_164
timestamp 1666464484
transform 1 0 16192 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_169
timestamp 1666464484
transform 1 0 16652 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_181
timestamp 1666464484
transform 1 0 17756 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_185
timestamp 1666464484
transform 1 0 18124 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_206
timestamp 1666464484
transform 1 0 20056 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_216
timestamp 1666464484
transform 1 0 20976 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_15_225
timestamp 1666464484
transform 1 0 21804 0 -1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_15_238
timestamp 1666464484
transform 1 0 23000 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_250
timestamp 1666464484
transform 1 0 24104 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_254
timestamp 1666464484
transform 1 0 24472 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_271
timestamp 1666464484
transform 1 0 26036 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_279
timestamp 1666464484
transform 1 0 26772 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_281
timestamp 1666464484
transform 1 0 26956 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_301
timestamp 1666464484
transform 1 0 28796 0 -1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_15_313
timestamp 1666464484
transform 1 0 29900 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_325
timestamp 1666464484
transform 1 0 31004 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_333
timestamp 1666464484
transform 1 0 31740 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_337
timestamp 1666464484
transform 1 0 32108 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_355
timestamp 1666464484
transform 1 0 33764 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_363
timestamp 1666464484
transform 1 0 34500 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3
timestamp 1666464484
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_15
timestamp 1666464484
transform 1 0 2484 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_26
timestamp 1666464484
transform 1 0 3496 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_29
timestamp 1666464484
transform 1 0 3772 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_36
timestamp 1666464484
transform 1 0 4416 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_64
timestamp 1666464484
transform 1 0 6992 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_76
timestamp 1666464484
transform 1 0 8096 0 1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_16_85
timestamp 1666464484
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_16_97
timestamp 1666464484
transform 1 0 10028 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_116
timestamp 1666464484
transform 1 0 11776 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_138
timestamp 1666464484
transform 1 0 13800 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_141
timestamp 1666464484
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_153
timestamp 1666464484
transform 1 0 15180 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_165
timestamp 1666464484
transform 1 0 16284 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_169
timestamp 1666464484
transform 1 0 16652 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_175
timestamp 1666464484
transform 1 0 17204 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_188
timestamp 1666464484
transform 1 0 18400 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_16_197
timestamp 1666464484
transform 1 0 19228 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_16_213
timestamp 1666464484
transform 1 0 20700 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_223
timestamp 1666464484
transform 1 0 21620 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_16_237
timestamp 1666464484
transform 1 0 22908 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_243
timestamp 1666464484
transform 1 0 23460 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_250
timestamp 1666464484
transform 1 0 24104 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_253
timestamp 1666464484
transform 1 0 24380 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_265
timestamp 1666464484
transform 1 0 25484 0 1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_16_291
timestamp 1666464484
transform 1 0 27876 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_303
timestamp 1666464484
transform 1 0 28980 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_307
timestamp 1666464484
transform 1 0 29348 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_309
timestamp 1666464484
transform 1 0 29532 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_317
timestamp 1666464484
transform 1 0 30268 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_329
timestamp 1666464484
transform 1 0 31372 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_346
timestamp 1666464484
transform 1 0 32936 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_358
timestamp 1666464484
transform 1 0 34040 0 1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3
timestamp 1666464484
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_15
timestamp 1666464484
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_27
timestamp 1666464484
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_39
timestamp 1666464484
transform 1 0 4692 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_51
timestamp 1666464484
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1666464484
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_57
timestamp 1666464484
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_69
timestamp 1666464484
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_81
timestamp 1666464484
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_93
timestamp 1666464484
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_105
timestamp 1666464484
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1666464484
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_113
timestamp 1666464484
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_125
timestamp 1666464484
transform 1 0 12604 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_137
timestamp 1666464484
transform 1 0 13708 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_149
timestamp 1666464484
transform 1 0 14812 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_157
timestamp 1666464484
transform 1 0 15548 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_166
timestamp 1666464484
transform 1 0 16376 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_169
timestamp 1666464484
transform 1 0 16652 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_177
timestamp 1666464484
transform 1 0 17388 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_190
timestamp 1666464484
transform 1 0 18584 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_218
timestamp 1666464484
transform 1 0 21160 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_17_225
timestamp 1666464484
transform 1 0 21804 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_243
timestamp 1666464484
transform 1 0 23460 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_263
timestamp 1666464484
transform 1 0 25300 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_273
timestamp 1666464484
transform 1 0 26220 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_279
timestamp 1666464484
transform 1 0 26772 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_281
timestamp 1666464484
transform 1 0 26956 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_301
timestamp 1666464484
transform 1 0 28796 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_313
timestamp 1666464484
transform 1 0 29900 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_325
timestamp 1666464484
transform 1 0 31004 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_333
timestamp 1666464484
transform 1 0 31740 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_337
timestamp 1666464484
transform 1 0 32108 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_345
timestamp 1666464484
transform 1 0 32844 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_357
timestamp 1666464484
transform 1 0 33948 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_363
timestamp 1666464484
transform 1 0 34500 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3
timestamp 1666464484
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_15
timestamp 1666464484
transform 1 0 2484 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_18_26
timestamp 1666464484
transform 1 0 3496 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_29
timestamp 1666464484
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_41
timestamp 1666464484
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_53
timestamp 1666464484
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_65
timestamp 1666464484
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_77
timestamp 1666464484
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1666464484
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_85
timestamp 1666464484
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_97
timestamp 1666464484
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_109
timestamp 1666464484
transform 1 0 11132 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_121
timestamp 1666464484
transform 1 0 12236 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_133
timestamp 1666464484
transform 1 0 13340 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_139
timestamp 1666464484
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_141
timestamp 1666464484
transform 1 0 14076 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_145
timestamp 1666464484
transform 1 0 14444 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_157
timestamp 1666464484
transform 1 0 15548 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_172
timestamp 1666464484
transform 1 0 16928 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_18_187
timestamp 1666464484
transform 1 0 18308 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_195
timestamp 1666464484
transform 1 0 19044 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_197
timestamp 1666464484
transform 1 0 19228 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_209
timestamp 1666464484
transform 1 0 20332 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_213
timestamp 1666464484
transform 1 0 20700 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_234
timestamp 1666464484
transform 1 0 22632 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_246
timestamp 1666464484
transform 1 0 23736 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_18_253
timestamp 1666464484
transform 1 0 24380 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_261
timestamp 1666464484
transform 1 0 25116 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_273
timestamp 1666464484
transform 1 0 26220 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_285
timestamp 1666464484
transform 1 0 27324 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_18_299
timestamp 1666464484
transform 1 0 28612 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_307
timestamp 1666464484
transform 1 0 29348 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_309
timestamp 1666464484
transform 1 0 29532 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_321
timestamp 1666464484
transform 1 0 30636 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_333
timestamp 1666464484
transform 1 0 31740 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_345
timestamp 1666464484
transform 1 0 32844 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_357
timestamp 1666464484
transform 1 0 33948 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_363
timestamp 1666464484
transform 1 0 34500 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_3
timestamp 1666464484
transform 1 0 1380 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_19_31
timestamp 1666464484
transform 1 0 3956 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_38
timestamp 1666464484
transform 1 0 4600 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_50
timestamp 1666464484
transform 1 0 5704 0 -1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_19_57
timestamp 1666464484
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_69
timestamp 1666464484
transform 1 0 7452 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_73
timestamp 1666464484
transform 1 0 7820 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_95
timestamp 1666464484
transform 1 0 9844 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_107
timestamp 1666464484
transform 1 0 10948 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1666464484
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_113
timestamp 1666464484
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_125
timestamp 1666464484
transform 1 0 12604 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_149
timestamp 1666464484
transform 1 0 14812 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_19_166
timestamp 1666464484
transform 1 0 16376 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_169
timestamp 1666464484
transform 1 0 16652 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_176
timestamp 1666464484
transform 1 0 17296 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_189
timestamp 1666464484
transform 1 0 18492 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_201
timestamp 1666464484
transform 1 0 19596 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_209
timestamp 1666464484
transform 1 0 20332 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_217
timestamp 1666464484
transform 1 0 21068 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_223
timestamp 1666464484
transform 1 0 21620 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_225
timestamp 1666464484
transform 1 0 21804 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_237
timestamp 1666464484
transform 1 0 22908 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_249
timestamp 1666464484
transform 1 0 24012 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_261
timestamp 1666464484
transform 1 0 25116 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_273
timestamp 1666464484
transform 1 0 26220 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_279
timestamp 1666464484
transform 1 0 26772 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_19_281
timestamp 1666464484
transform 1 0 26956 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_292
timestamp 1666464484
transform 1 0 27968 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_302
timestamp 1666464484
transform 1 0 28888 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_312
timestamp 1666464484
transform 1 0 29808 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_324
timestamp 1666464484
transform 1 0 30912 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_337
timestamp 1666464484
transform 1 0 32108 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_345
timestamp 1666464484
transform 1 0 32844 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_357
timestamp 1666464484
transform 1 0 33948 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_363
timestamp 1666464484
transform 1 0 34500 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_3
timestamp 1666464484
transform 1 0 1380 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_11
timestamp 1666464484
transform 1 0 2116 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_16
timestamp 1666464484
transform 1 0 2576 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_26
timestamp 1666464484
transform 1 0 3496 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_29
timestamp 1666464484
transform 1 0 3772 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_40
timestamp 1666464484
transform 1 0 4784 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_49
timestamp 1666464484
transform 1 0 5612 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_61
timestamp 1666464484
transform 1 0 6716 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_73
timestamp 1666464484
transform 1 0 7820 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_82
timestamp 1666464484
transform 1 0 8648 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_85
timestamp 1666464484
transform 1 0 8924 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_108
timestamp 1666464484
transform 1 0 11040 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_137
timestamp 1666464484
transform 1 0 13708 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_141
timestamp 1666464484
transform 1 0 14076 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_20_152
timestamp 1666464484
transform 1 0 15088 0 1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_20_169
timestamp 1666464484
transform 1 0 16652 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_181
timestamp 1666464484
transform 1 0 17756 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_191
timestamp 1666464484
transform 1 0 18676 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_195
timestamp 1666464484
transform 1 0 19044 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_197
timestamp 1666464484
transform 1 0 19228 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_20_209
timestamp 1666464484
transform 1 0 20332 0 1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_20_232
timestamp 1666464484
transform 1 0 22448 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_244
timestamp 1666464484
transform 1 0 23552 0 1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_20_253
timestamp 1666464484
transform 1 0 24380 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_265
timestamp 1666464484
transform 1 0 25484 0 1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_20_291
timestamp 1666464484
transform 1 0 27876 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_303
timestamp 1666464484
transform 1 0 28980 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_307
timestamp 1666464484
transform 1 0 29348 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_309
timestamp 1666464484
transform 1 0 29532 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_321
timestamp 1666464484
transform 1 0 30636 0 1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_20_347
timestamp 1666464484
transform 1 0 33028 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_359
timestamp 1666464484
transform 1 0 34132 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_363
timestamp 1666464484
transform 1 0 34500 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_3
timestamp 1666464484
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_18
timestamp 1666464484
transform 1 0 2760 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_21_30
timestamp 1666464484
transform 1 0 3864 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_54
timestamp 1666464484
transform 1 0 6072 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_57
timestamp 1666464484
transform 1 0 6348 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_65
timestamp 1666464484
transform 1 0 7084 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_21_93
timestamp 1666464484
transform 1 0 9660 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_102
timestamp 1666464484
transform 1 0 10488 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_110
timestamp 1666464484
transform 1 0 11224 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_113
timestamp 1666464484
transform 1 0 11500 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_137
timestamp 1666464484
transform 1 0 13708 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_148
timestamp 1666464484
transform 1 0 14720 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_161
timestamp 1666464484
transform 1 0 15916 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_167
timestamp 1666464484
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_169
timestamp 1666464484
transform 1 0 16652 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_180
timestamp 1666464484
transform 1 0 17664 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_192
timestamp 1666464484
transform 1 0 18768 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_198
timestamp 1666464484
transform 1 0 19320 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_205
timestamp 1666464484
transform 1 0 19964 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_21_215
timestamp 1666464484
transform 1 0 20884 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_223
timestamp 1666464484
transform 1 0 21620 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_225
timestamp 1666464484
transform 1 0 21804 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_237
timestamp 1666464484
transform 1 0 22908 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_249
timestamp 1666464484
transform 1 0 24012 0 -1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_21_261
timestamp 1666464484
transform 1 0 25116 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_273
timestamp 1666464484
transform 1 0 26220 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_279
timestamp 1666464484
transform 1 0 26772 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_21_281
timestamp 1666464484
transform 1 0 26956 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_21_292
timestamp 1666464484
transform 1 0 27968 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_21_306
timestamp 1666464484
transform 1 0 29256 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_316
timestamp 1666464484
transform 1 0 30176 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_334
timestamp 1666464484
transform 1 0 31832 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_337
timestamp 1666464484
transform 1 0 32108 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_358
timestamp 1666464484
transform 1 0 34040 0 -1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_22_3
timestamp 1666464484
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_15
timestamp 1666464484
transform 1 0 2484 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_21
timestamp 1666464484
transform 1 0 3036 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1666464484
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_29
timestamp 1666464484
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_41
timestamp 1666464484
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_53
timestamp 1666464484
transform 1 0 5980 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_60
timestamp 1666464484
transform 1 0 6624 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_69
timestamp 1666464484
transform 1 0 7452 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_82
timestamp 1666464484
transform 1 0 8648 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_85
timestamp 1666464484
transform 1 0 8924 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_96
timestamp 1666464484
transform 1 0 9936 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_108
timestamp 1666464484
transform 1 0 11040 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_120
timestamp 1666464484
transform 1 0 12144 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_22_131
timestamp 1666464484
transform 1 0 13156 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_139
timestamp 1666464484
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_141
timestamp 1666464484
transform 1 0 14076 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_22_148
timestamp 1666464484
transform 1 0 14720 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_156
timestamp 1666464484
transform 1 0 15456 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_177
timestamp 1666464484
transform 1 0 17388 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_190
timestamp 1666464484
transform 1 0 18584 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_22_197
timestamp 1666464484
transform 1 0 19228 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_217
timestamp 1666464484
transform 1 0 21068 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_228
timestamp 1666464484
transform 1 0 22080 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_240
timestamp 1666464484
transform 1 0 23184 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_250
timestamp 1666464484
transform 1 0 24104 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_253
timestamp 1666464484
transform 1 0 24380 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_271
timestamp 1666464484
transform 1 0 26036 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_291
timestamp 1666464484
transform 1 0 27876 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_301
timestamp 1666464484
transform 1 0 28796 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_307
timestamp 1666464484
transform 1 0 29348 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_309
timestamp 1666464484
transform 1 0 29532 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_330
timestamp 1666464484
transform 1 0 31464 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_353
timestamp 1666464484
transform 1 0 33580 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_361
timestamp 1666464484
transform 1 0 34316 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_23_3
timestamp 1666464484
transform 1 0 1380 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_27
timestamp 1666464484
transform 1 0 3588 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_34
timestamp 1666464484
transform 1 0 4232 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_42
timestamp 1666464484
transform 1 0 4968 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_52
timestamp 1666464484
transform 1 0 5888 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_57
timestamp 1666464484
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_69
timestamp 1666464484
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_81
timestamp 1666464484
transform 1 0 8556 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_94
timestamp 1666464484
transform 1 0 9752 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_110
timestamp 1666464484
transform 1 0 11224 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_113
timestamp 1666464484
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_125
timestamp 1666464484
transform 1 0 12604 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_137
timestamp 1666464484
transform 1 0 13708 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_149
timestamp 1666464484
transform 1 0 14812 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_157
timestamp 1666464484
transform 1 0 15548 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_166
timestamp 1666464484
transform 1 0 16376 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_169
timestamp 1666464484
transform 1 0 16652 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_178
timestamp 1666464484
transform 1 0 17480 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_23_206
timestamp 1666464484
transform 1 0 20056 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_216
timestamp 1666464484
transform 1 0 20976 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_225
timestamp 1666464484
transform 1 0 21804 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_233
timestamp 1666464484
transform 1 0 22540 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_243
timestamp 1666464484
transform 1 0 23460 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_247
timestamp 1666464484
transform 1 0 23828 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_264
timestamp 1666464484
transform 1 0 25392 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_276
timestamp 1666464484
transform 1 0 26496 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_281
timestamp 1666464484
transform 1 0 26956 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_293
timestamp 1666464484
transform 1 0 28060 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_305
timestamp 1666464484
transform 1 0 29164 0 -1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_23_315
timestamp 1666464484
transform 1 0 30084 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_327
timestamp 1666464484
transform 1 0 31188 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_335
timestamp 1666464484
transform 1 0 31924 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_337
timestamp 1666464484
transform 1 0 32108 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_359
timestamp 1666464484
transform 1 0 34132 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_363
timestamp 1666464484
transform 1 0 34500 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_3
timestamp 1666464484
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_15
timestamp 1666464484
transform 1 0 2484 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_24_21
timestamp 1666464484
transform 1 0 3036 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1666464484
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_29
timestamp 1666464484
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_41
timestamp 1666464484
transform 1 0 4876 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_24_48
timestamp 1666464484
transform 1 0 5520 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_24_57
timestamp 1666464484
transform 1 0 6348 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_24_64
timestamp 1666464484
transform 1 0 6992 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_76
timestamp 1666464484
transform 1 0 8096 0 1 15232
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_24_85
timestamp 1666464484
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_97
timestamp 1666464484
transform 1 0 10028 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_109
timestamp 1666464484
transform 1 0 11132 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_24_121
timestamp 1666464484
transform 1 0 12236 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_24_127
timestamp 1666464484
transform 1 0 12788 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_24_138
timestamp 1666464484
transform 1 0 13800 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_141
timestamp 1666464484
transform 1 0 14076 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_149
timestamp 1666464484
transform 1 0 14812 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_170
timestamp 1666464484
transform 1 0 16744 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_24_178
timestamp 1666464484
transform 1 0 17480 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_24_188
timestamp 1666464484
transform 1 0 18400 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_24_197
timestamp 1666464484
transform 1 0 19228 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_24_209
timestamp 1666464484
transform 1 0 20332 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_213
timestamp 1666464484
transform 1 0 20700 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_24_234
timestamp 1666464484
transform 1 0 22632 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_24_246
timestamp 1666464484
transform 1 0 23736 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_24_253
timestamp 1666464484
transform 1 0 24380 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_261
timestamp 1666464484
transform 1 0 25116 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_282
timestamp 1666464484
transform 1 0 27048 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_294
timestamp 1666464484
transform 1 0 28152 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_302
timestamp 1666464484
transform 1 0 28888 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_306
timestamp 1666464484
transform 1 0 29256 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_309
timestamp 1666464484
transform 1 0 29532 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_321
timestamp 1666464484
transform 1 0 30636 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_24_347
timestamp 1666464484
transform 1 0 33028 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_357
timestamp 1666464484
transform 1 0 33948 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_363
timestamp 1666464484
transform 1 0 34500 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_3
timestamp 1666464484
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_15
timestamp 1666464484
transform 1 0 2484 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_27
timestamp 1666464484
transform 1 0 3588 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_39
timestamp 1666464484
transform 1 0 4692 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_45
timestamp 1666464484
transform 1 0 5244 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_52
timestamp 1666464484
transform 1 0 5888 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_57
timestamp 1666464484
transform 1 0 6348 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_25_62
timestamp 1666464484
transform 1 0 6808 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_25_75
timestamp 1666464484
transform 1 0 8004 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_83
timestamp 1666464484
transform 1 0 8740 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_87
timestamp 1666464484
transform 1 0 9108 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_110
timestamp 1666464484
transform 1 0 11224 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_113
timestamp 1666464484
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_125
timestamp 1666464484
transform 1 0 12604 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_25_137
timestamp 1666464484
transform 1 0 13708 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_146
timestamp 1666464484
transform 1 0 14536 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_166
timestamp 1666464484
transform 1 0 16376 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_169
timestamp 1666464484
transform 1 0 16652 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_25_182
timestamp 1666464484
transform 1 0 17848 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_206
timestamp 1666464484
transform 1 0 20056 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_218
timestamp 1666464484
transform 1 0 21160 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_25_225
timestamp 1666464484
transform 1 0 21804 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_25_235
timestamp 1666464484
transform 1 0 22724 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_241
timestamp 1666464484
transform 1 0 23276 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_262
timestamp 1666464484
transform 1 0 25208 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_25_276
timestamp 1666464484
transform 1 0 26496 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_281
timestamp 1666464484
transform 1 0 26956 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_289
timestamp 1666464484
transform 1 0 27692 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_299
timestamp 1666464484
transform 1 0 28612 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_25_310
timestamp 1666464484
transform 1 0 29624 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_322
timestamp 1666464484
transform 1 0 30728 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_334
timestamp 1666464484
transform 1 0 31832 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_337
timestamp 1666464484
transform 1 0 32108 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_356
timestamp 1666464484
transform 1 0 33856 0 -1 16320
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_26_3
timestamp 1666464484
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_15
timestamp 1666464484
transform 1 0 2484 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_26_26
timestamp 1666464484
transform 1 0 3496 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_29
timestamp 1666464484
transform 1 0 3772 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_36
timestamp 1666464484
transform 1 0 4416 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_54
timestamp 1666464484
transform 1 0 6072 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_60
timestamp 1666464484
transform 1 0 6624 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_70
timestamp 1666464484
transform 1 0 7544 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_26_82
timestamp 1666464484
transform 1 0 8648 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_85
timestamp 1666464484
transform 1 0 8924 0 1 16320
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_26_100
timestamp 1666464484
transform 1 0 10304 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_112
timestamp 1666464484
transform 1 0 11408 0 1 16320
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_26_125
timestamp 1666464484
transform 1 0 12604 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_26_137
timestamp 1666464484
transform 1 0 13708 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_26_141
timestamp 1666464484
transform 1 0 14076 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_150
timestamp 1666464484
transform 1 0 14904 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_170
timestamp 1666464484
transform 1 0 16744 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_26_183
timestamp 1666464484
transform 1 0 17940 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_195
timestamp 1666464484
transform 1 0 19044 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_197
timestamp 1666464484
transform 1 0 19228 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_205
timestamp 1666464484
transform 1 0 19964 0 1 16320
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_26_229
timestamp 1666464484
transform 1 0 22172 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_241
timestamp 1666464484
transform 1 0 23276 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_26_249
timestamp 1666464484
transform 1 0 24012 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_253
timestamp 1666464484
transform 1 0 24380 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_271
timestamp 1666464484
transform 1 0 26036 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_26_281
timestamp 1666464484
transform 1 0 26956 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_293
timestamp 1666464484
transform 1 0 28060 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_26_305
timestamp 1666464484
transform 1 0 29164 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_309
timestamp 1666464484
transform 1 0 29532 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_319
timestamp 1666464484
transform 1 0 30452 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_26_333
timestamp 1666464484
transform 1 0 31740 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_337
timestamp 1666464484
transform 1 0 32108 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_343
timestamp 1666464484
transform 1 0 32660 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_355
timestamp 1666464484
transform 1 0 33764 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_363
timestamp 1666464484
transform 1 0 34500 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_3
timestamp 1666464484
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_15
timestamp 1666464484
transform 1 0 2484 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_37
timestamp 1666464484
transform 1 0 4508 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_49
timestamp 1666464484
transform 1 0 5612 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_55
timestamp 1666464484
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_57
timestamp 1666464484
transform 1 0 6348 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_71
timestamp 1666464484
transform 1 0 7636 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_27_78
timestamp 1666464484
transform 1 0 8280 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_90
timestamp 1666464484
transform 1 0 9384 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_98
timestamp 1666464484
transform 1 0 10120 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_110
timestamp 1666464484
transform 1 0 11224 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_113
timestamp 1666464484
transform 1 0 11500 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_136
timestamp 1666464484
transform 1 0 13616 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_148
timestamp 1666464484
transform 1 0 14720 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_156
timestamp 1666464484
transform 1 0 15456 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_166
timestamp 1666464484
transform 1 0 16376 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_169
timestamp 1666464484
transform 1 0 16652 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_181
timestamp 1666464484
transform 1 0 17756 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_209
timestamp 1666464484
transform 1 0 20332 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_219
timestamp 1666464484
transform 1 0 21252 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_223
timestamp 1666464484
transform 1 0 21620 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_225
timestamp 1666464484
transform 1 0 21804 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_237
timestamp 1666464484
transform 1 0 22908 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_256
timestamp 1666464484
transform 1 0 24656 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_27_268
timestamp 1666464484
transform 1 0 25760 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_281
timestamp 1666464484
transform 1 0 26956 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_293
timestamp 1666464484
transform 1 0 28060 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_305
timestamp 1666464484
transform 1 0 29164 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_27_314
timestamp 1666464484
transform 1 0 29992 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_318
timestamp 1666464484
transform 1 0 30360 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_326
timestamp 1666464484
transform 1 0 31096 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_334
timestamp 1666464484
transform 1 0 31832 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_337
timestamp 1666464484
transform 1 0 32108 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_344
timestamp 1666464484
transform 1 0 32752 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_27_351
timestamp 1666464484
transform 1 0 33396 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_363
timestamp 1666464484
transform 1 0 34500 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_3
timestamp 1666464484
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_15
timestamp 1666464484
transform 1 0 2484 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_26
timestamp 1666464484
transform 1 0 3496 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_29
timestamp 1666464484
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_41
timestamp 1666464484
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_53
timestamp 1666464484
transform 1 0 5980 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_28_60
timestamp 1666464484
transform 1 0 6624 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_72
timestamp 1666464484
transform 1 0 7728 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_85
timestamp 1666464484
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_97
timestamp 1666464484
transform 1 0 10028 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_109
timestamp 1666464484
transform 1 0 11132 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_131
timestamp 1666464484
transform 1 0 13156 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_139
timestamp 1666464484
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_141
timestamp 1666464484
transform 1 0 14076 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_173
timestamp 1666464484
transform 1 0 17020 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_185
timestamp 1666464484
transform 1 0 18124 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_28_193
timestamp 1666464484
transform 1 0 18860 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_197
timestamp 1666464484
transform 1 0 19228 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_215
timestamp 1666464484
transform 1 0 20884 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_227
timestamp 1666464484
transform 1 0 21988 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_239
timestamp 1666464484
transform 1 0 23092 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_251
timestamp 1666464484
transform 1 0 24196 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_253
timestamp 1666464484
transform 1 0 24380 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_28_263
timestamp 1666464484
transform 1 0 25300 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_275
timestamp 1666464484
transform 1 0 26404 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_28_283
timestamp 1666464484
transform 1 0 27140 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_293
timestamp 1666464484
transform 1 0 28060 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_297
timestamp 1666464484
transform 1 0 28428 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_28_302
timestamp 1666464484
transform 1 0 28888 0 1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_28_309
timestamp 1666464484
transform 1 0 29532 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_321
timestamp 1666464484
transform 1 0 30636 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_28_327
timestamp 1666464484
transform 1 0 31188 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_28_336
timestamp 1666464484
transform 1 0 32016 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_345
timestamp 1666464484
transform 1 0 32844 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_354
timestamp 1666464484
transform 1 0 33672 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_362
timestamp 1666464484
transform 1 0 34408 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_3
timestamp 1666464484
transform 1 0 1380 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_15
timestamp 1666464484
transform 1 0 2484 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_27
timestamp 1666464484
transform 1 0 3588 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_39
timestamp 1666464484
transform 1 0 4692 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_51
timestamp 1666464484
transform 1 0 5796 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_55
timestamp 1666464484
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_29_57
timestamp 1666464484
transform 1 0 6348 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_29_69
timestamp 1666464484
transform 1 0 7452 0 -1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_29_78
timestamp 1666464484
transform 1 0 8280 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_90
timestamp 1666464484
transform 1 0 9384 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_29_101
timestamp 1666464484
transform 1 0 10396 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_109
timestamp 1666464484
transform 1 0 11132 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_29_113
timestamp 1666464484
transform 1 0 11500 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_119
timestamp 1666464484
transform 1 0 12052 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_125
timestamp 1666464484
transform 1 0 12604 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_149
timestamp 1666464484
transform 1 0 14812 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_157
timestamp 1666464484
transform 1 0 15548 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_166
timestamp 1666464484
transform 1 0 16376 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_169
timestamp 1666464484
transform 1 0 16652 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_177
timestamp 1666464484
transform 1 0 17388 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_189
timestamp 1666464484
transform 1 0 18492 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_207
timestamp 1666464484
transform 1 0 20148 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_29_217
timestamp 1666464484
transform 1 0 21068 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_223
timestamp 1666464484
transform 1 0 21620 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_225
timestamp 1666464484
transform 1 0 21804 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_29_237
timestamp 1666464484
transform 1 0 22908 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_259
timestamp 1666464484
transform 1 0 24932 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_29_268
timestamp 1666464484
transform 1 0 25760 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_281
timestamp 1666464484
transform 1 0 26956 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_289
timestamp 1666464484
transform 1 0 27692 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_297
timestamp 1666464484
transform 1 0 28428 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_29_307
timestamp 1666464484
transform 1 0 29348 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_319
timestamp 1666464484
transform 1 0 30452 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_331
timestamp 1666464484
transform 1 0 31556 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_335
timestamp 1666464484
transform 1 0 31924 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_337
timestamp 1666464484
transform 1 0 32108 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_346
timestamp 1666464484
transform 1 0 32936 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_29_358
timestamp 1666464484
transform 1 0 34040 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_362
timestamp 1666464484
transform 1 0 34408 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_3
timestamp 1666464484
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_15
timestamp 1666464484
transform 1 0 2484 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_21
timestamp 1666464484
transform 1 0 3036 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_26
timestamp 1666464484
transform 1 0 3496 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_29
timestamp 1666464484
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_41
timestamp 1666464484
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_53
timestamp 1666464484
transform 1 0 5980 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_65
timestamp 1666464484
transform 1 0 7084 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_30_79
timestamp 1666464484
transform 1 0 8372 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp 1666464484
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_85
timestamp 1666464484
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_97
timestamp 1666464484
transform 1 0 10028 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_30_104
timestamp 1666464484
transform 1 0 10672 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_30_116
timestamp 1666464484
transform 1 0 11776 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_123
timestamp 1666464484
transform 1 0 12420 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_135
timestamp 1666464484
transform 1 0 13524 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_139
timestamp 1666464484
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_141
timestamp 1666464484
transform 1 0 14076 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_169
timestamp 1666464484
transform 1 0 16652 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_181
timestamp 1666464484
transform 1 0 17756 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_187
timestamp 1666464484
transform 1 0 18308 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_194
timestamp 1666464484
transform 1 0 18952 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_197
timestamp 1666464484
transform 1 0 19228 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_219
timestamp 1666464484
transform 1 0 21252 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_231
timestamp 1666464484
transform 1 0 22356 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_243
timestamp 1666464484
transform 1 0 23460 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_250
timestamp 1666464484
transform 1 0 24104 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_253
timestamp 1666464484
transform 1 0 24380 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_30_261
timestamp 1666464484
transform 1 0 25116 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_30_276
timestamp 1666464484
transform 1 0 26496 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_280
timestamp 1666464484
transform 1 0 26864 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_288
timestamp 1666464484
transform 1 0 27600 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_306
timestamp 1666464484
transform 1 0 29256 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_309
timestamp 1666464484
transform 1 0 29532 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_316
timestamp 1666464484
transform 1 0 30176 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_328
timestamp 1666464484
transform 1 0 31280 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_30_339
timestamp 1666464484
transform 1 0 32292 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_30_349
timestamp 1666464484
transform 1 0 33212 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_30_361
timestamp 1666464484
transform 1 0 34316 0 1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_31_3
timestamp 1666464484
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_34
timestamp 1666464484
transform 1 0 4232 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_31_42
timestamp 1666464484
transform 1 0 4968 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_54
timestamp 1666464484
transform 1 0 6072 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_31_57
timestamp 1666464484
transform 1 0 6348 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_31_82
timestamp 1666464484
transform 1 0 8648 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_89
timestamp 1666464484
transform 1 0 9292 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_97
timestamp 1666464484
transform 1 0 10028 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_31_106
timestamp 1666464484
transform 1 0 10856 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_31_113
timestamp 1666464484
transform 1 0 11500 0 -1 19584
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_31_127
timestamp 1666464484
transform 1 0 12788 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_139
timestamp 1666464484
transform 1 0 13892 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_147
timestamp 1666464484
transform 1 0 14628 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_166
timestamp 1666464484
transform 1 0 16376 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_169
timestamp 1666464484
transform 1 0 16652 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_177
timestamp 1666464484
transform 1 0 17388 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_189
timestamp 1666464484
transform 1 0 18492 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_197
timestamp 1666464484
transform 1 0 19228 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_31_215
timestamp 1666464484
transform 1 0 20884 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_223
timestamp 1666464484
transform 1 0 21620 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_225
timestamp 1666464484
transform 1 0 21804 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_31_233
timestamp 1666464484
transform 1 0 22540 0 -1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_31_258
timestamp 1666464484
transform 1 0 24840 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_270
timestamp 1666464484
transform 1 0 25944 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_278
timestamp 1666464484
transform 1 0 26680 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_281
timestamp 1666464484
transform 1 0 26956 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_31_287
timestamp 1666464484
transform 1 0 27508 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_295
timestamp 1666464484
transform 1 0 28244 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_31_315
timestamp 1666464484
transform 1 0 30084 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_323
timestamp 1666464484
transform 1 0 30820 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_331
timestamp 1666464484
transform 1 0 31556 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_335
timestamp 1666464484
transform 1 0 31924 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_337
timestamp 1666464484
transform 1 0 32108 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_346
timestamp 1666464484
transform 1 0 32936 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_358
timestamp 1666464484
transform 1 0 34040 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_32_3
timestamp 1666464484
transform 1 0 1380 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_9
timestamp 1666464484
transform 1 0 1932 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_26
timestamp 1666464484
transform 1 0 3496 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_29
timestamp 1666464484
transform 1 0 3772 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_39
timestamp 1666464484
transform 1 0 4692 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_48
timestamp 1666464484
transform 1 0 5520 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_60
timestamp 1666464484
transform 1 0 6624 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_66
timestamp 1666464484
transform 1 0 7176 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_76
timestamp 1666464484
transform 1 0 8096 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_85
timestamp 1666464484
transform 1 0 8924 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_91
timestamp 1666464484
transform 1 0 9476 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_99
timestamp 1666464484
transform 1 0 10212 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_109
timestamp 1666464484
transform 1 0 11132 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_118
timestamp 1666464484
transform 1 0 11960 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_32_130
timestamp 1666464484
transform 1 0 13064 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_138
timestamp 1666464484
transform 1 0 13800 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_141
timestamp 1666464484
transform 1 0 14076 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_148
timestamp 1666464484
transform 1 0 14720 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_152
timestamp 1666464484
transform 1 0 15088 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_159
timestamp 1666464484
transform 1 0 15732 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_172
timestamp 1666464484
transform 1 0 16928 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_185
timestamp 1666464484
transform 1 0 18124 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_32_193
timestamp 1666464484
transform 1 0 18860 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_197
timestamp 1666464484
transform 1 0 19228 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_32_207
timestamp 1666464484
transform 1 0 20148 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_213
timestamp 1666464484
transform 1 0 20700 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_234
timestamp 1666464484
transform 1 0 22632 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_246
timestamp 1666464484
transform 1 0 23736 0 1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_32_253
timestamp 1666464484
transform 1 0 24380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_265
timestamp 1666464484
transform 1 0 25484 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_277
timestamp 1666464484
transform 1 0 26588 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_289
timestamp 1666464484
transform 1 0 27692 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_295
timestamp 1666464484
transform 1 0 28244 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_304
timestamp 1666464484
transform 1 0 29072 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_309
timestamp 1666464484
transform 1 0 29532 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_321
timestamp 1666464484
transform 1 0 30636 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_333
timestamp 1666464484
transform 1 0 31740 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_345
timestamp 1666464484
transform 1 0 32844 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_357
timestamp 1666464484
transform 1 0 33948 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_363
timestamp 1666464484
transform 1 0 34500 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_3
timestamp 1666464484
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_15
timestamp 1666464484
transform 1 0 2484 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_19
timestamp 1666464484
transform 1 0 2852 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_28
timestamp 1666464484
transform 1 0 3680 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_39
timestamp 1666464484
transform 1 0 4692 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_51
timestamp 1666464484
transform 1 0 5796 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_55
timestamp 1666464484
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_57
timestamp 1666464484
transform 1 0 6348 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_33_65
timestamp 1666464484
transform 1 0 7084 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_33_74
timestamp 1666464484
transform 1 0 7912 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_82
timestamp 1666464484
transform 1 0 8648 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_94
timestamp 1666464484
transform 1 0 9752 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_110
timestamp 1666464484
transform 1 0 11224 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_113
timestamp 1666464484
transform 1 0 11500 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_125
timestamp 1666464484
transform 1 0 12604 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_141
timestamp 1666464484
transform 1 0 14076 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_154
timestamp 1666464484
transform 1 0 15272 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_163
timestamp 1666464484
transform 1 0 16100 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_167
timestamp 1666464484
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_169
timestamp 1666464484
transform 1 0 16652 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_181
timestamp 1666464484
transform 1 0 17756 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_185
timestamp 1666464484
transform 1 0 18124 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_206
timestamp 1666464484
transform 1 0 20056 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_217
timestamp 1666464484
transform 1 0 21068 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_223
timestamp 1666464484
transform 1 0 21620 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_225
timestamp 1666464484
transform 1 0 21804 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_33_233
timestamp 1666464484
transform 1 0 22540 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_239
timestamp 1666464484
transform 1 0 23092 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_260
timestamp 1666464484
transform 1 0 25024 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_272
timestamp 1666464484
transform 1 0 26128 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_33_281
timestamp 1666464484
transform 1 0 26956 0 -1 20672
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_33_293
timestamp 1666464484
transform 1 0 28060 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_305
timestamp 1666464484
transform 1 0 29164 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_317
timestamp 1666464484
transform 1 0 30268 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_329
timestamp 1666464484
transform 1 0 31372 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_334
timestamp 1666464484
transform 1 0 31832 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_337
timestamp 1666464484
transform 1 0 32108 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_348
timestamp 1666464484
transform 1 0 33120 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_360
timestamp 1666464484
transform 1 0 34224 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_34_3
timestamp 1666464484
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_15
timestamp 1666464484
transform 1 0 2484 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_26
timestamp 1666464484
transform 1 0 3496 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_29
timestamp 1666464484
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_41
timestamp 1666464484
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_53
timestamp 1666464484
transform 1 0 5980 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_34_65
timestamp 1666464484
transform 1 0 7084 0 1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_34_72
timestamp 1666464484
transform 1 0 7728 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_85
timestamp 1666464484
transform 1 0 8924 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_34_97
timestamp 1666464484
transform 1 0 10028 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_105
timestamp 1666464484
transform 1 0 10764 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_117
timestamp 1666464484
transform 1 0 11868 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_129
timestamp 1666464484
transform 1 0 12972 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_136
timestamp 1666464484
transform 1 0 13616 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_141
timestamp 1666464484
transform 1 0 14076 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_34_148
timestamp 1666464484
transform 1 0 14720 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_156
timestamp 1666464484
transform 1 0 15456 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_34_178
timestamp 1666464484
transform 1 0 17480 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_186
timestamp 1666464484
transform 1 0 18216 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_194
timestamp 1666464484
transform 1 0 18952 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_197
timestamp 1666464484
transform 1 0 19228 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_209
timestamp 1666464484
transform 1 0 20332 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_213
timestamp 1666464484
transform 1 0 20700 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_34_234
timestamp 1666464484
transform 1 0 22632 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_242
timestamp 1666464484
transform 1 0 23368 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_250
timestamp 1666464484
transform 1 0 24104 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_253
timestamp 1666464484
transform 1 0 24380 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_261
timestamp 1666464484
transform 1 0 25116 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_273
timestamp 1666464484
transform 1 0 26220 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_285
timestamp 1666464484
transform 1 0 27324 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_297
timestamp 1666464484
transform 1 0 28428 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_34_305
timestamp 1666464484
transform 1 0 29164 0 1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_34_309
timestamp 1666464484
transform 1 0 29532 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_321
timestamp 1666464484
transform 1 0 30636 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_327
timestamp 1666464484
transform 1 0 31188 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_333
timestamp 1666464484
transform 1 0 31740 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_342
timestamp 1666464484
transform 1 0 32568 0 1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_34_349
timestamp 1666464484
transform 1 0 33212 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_34_361
timestamp 1666464484
transform 1 0 34316 0 1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_35_3
timestamp 1666464484
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_15
timestamp 1666464484
transform 1 0 2484 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_23
timestamp 1666464484
transform 1 0 3220 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_35_34
timestamp 1666464484
transform 1 0 4232 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_46
timestamp 1666464484
transform 1 0 5336 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_54
timestamp 1666464484
transform 1 0 6072 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_57
timestamp 1666464484
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_69
timestamp 1666464484
transform 1 0 7452 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_81
timestamp 1666464484
transform 1 0 8556 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_93
timestamp 1666464484
transform 1 0 9660 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_105
timestamp 1666464484
transform 1 0 10764 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_111
timestamp 1666464484
transform 1 0 11316 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_113
timestamp 1666464484
transform 1 0 11500 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_120
timestamp 1666464484
transform 1 0 12144 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_132
timestamp 1666464484
transform 1 0 13248 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_35_144
timestamp 1666464484
transform 1 0 14352 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_148
timestamp 1666464484
transform 1 0 14720 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_35_157
timestamp 1666464484
transform 1 0 15548 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_35_165
timestamp 1666464484
transform 1 0 16284 0 -1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_35_169
timestamp 1666464484
transform 1 0 16652 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_181
timestamp 1666464484
transform 1 0 17756 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_193
timestamp 1666464484
transform 1 0 18860 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_35_216
timestamp 1666464484
transform 1 0 20976 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_225
timestamp 1666464484
transform 1 0 21804 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_35_232
timestamp 1666464484
transform 1 0 22448 0 -1 21760
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_35_259
timestamp 1666464484
transform 1 0 24932 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_271
timestamp 1666464484
transform 1 0 26036 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_279
timestamp 1666464484
transform 1 0 26772 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_281
timestamp 1666464484
transform 1 0 26956 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_290
timestamp 1666464484
transform 1 0 27784 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_35_297
timestamp 1666464484
transform 1 0 28428 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_309
timestamp 1666464484
transform 1 0 29532 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_35_321
timestamp 1666464484
transform 1 0 30636 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_329
timestamp 1666464484
transform 1 0 31372 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_35_333
timestamp 1666464484
transform 1 0 31740 0 -1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_35_337
timestamp 1666464484
transform 1 0 32108 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_349
timestamp 1666464484
transform 1 0 33212 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_35_361
timestamp 1666464484
transform 1 0 34316 0 -1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_36_3
timestamp 1666464484
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_15
timestamp 1666464484
transform 1 0 2484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 1666464484
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_29
timestamp 1666464484
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_41
timestamp 1666464484
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_53
timestamp 1666464484
transform 1 0 5980 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_36_61
timestamp 1666464484
transform 1 0 6716 0 1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_36_68
timestamp 1666464484
transform 1 0 7360 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_80
timestamp 1666464484
transform 1 0 8464 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_85
timestamp 1666464484
transform 1 0 8924 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_36_90
timestamp 1666464484
transform 1 0 9384 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_98
timestamp 1666464484
transform 1 0 10120 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_120
timestamp 1666464484
transform 1 0 12144 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_132
timestamp 1666464484
transform 1 0 13248 0 1 21760
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_36_141
timestamp 1666464484
transform 1 0 14076 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_153
timestamp 1666464484
transform 1 0 15180 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_165
timestamp 1666464484
transform 1 0 16284 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_177
timestamp 1666464484
transform 1 0 17388 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_188
timestamp 1666464484
transform 1 0 18400 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_197
timestamp 1666464484
transform 1 0 19228 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_36_205
timestamp 1666464484
transform 1 0 19964 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_213
timestamp 1666464484
transform 1 0 20700 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_234
timestamp 1666464484
transform 1 0 22632 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_243
timestamp 1666464484
transform 1 0 23460 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_251
timestamp 1666464484
transform 1 0 24196 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_36_253
timestamp 1666464484
transform 1 0 24380 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_36_263
timestamp 1666464484
transform 1 0 25300 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_36_274
timestamp 1666464484
transform 1 0 26312 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_291
timestamp 1666464484
transform 1 0 27876 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_300
timestamp 1666464484
transform 1 0 28704 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_309
timestamp 1666464484
transform 1 0 29532 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_36_318
timestamp 1666464484
transform 1 0 30360 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_324
timestamp 1666464484
transform 1 0 30912 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_332
timestamp 1666464484
transform 1 0 31648 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_343
timestamp 1666464484
transform 1 0 32660 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_347
timestamp 1666464484
transform 1 0 33028 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_353
timestamp 1666464484
transform 1 0 33580 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_36_361
timestamp 1666464484
transform 1 0 34316 0 1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_37_3
timestamp 1666464484
transform 1 0 1380 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_15
timestamp 1666464484
transform 1 0 2484 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_32
timestamp 1666464484
transform 1 0 4048 0 -1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_37_43
timestamp 1666464484
transform 1 0 5060 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_37_55
timestamp 1666464484
transform 1 0 6164 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_57
timestamp 1666464484
transform 1 0 6348 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_65
timestamp 1666464484
transform 1 0 7084 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_72
timestamp 1666464484
transform 1 0 7728 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_81
timestamp 1666464484
transform 1 0 8556 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_37_94
timestamp 1666464484
transform 1 0 9752 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_110
timestamp 1666464484
transform 1 0 11224 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_113
timestamp 1666464484
transform 1 0 11500 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_118
timestamp 1666464484
transform 1 0 11960 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_122
timestamp 1666464484
transform 1 0 12328 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_140
timestamp 1666464484
transform 1 0 13984 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_144
timestamp 1666464484
transform 1 0 14352 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_149
timestamp 1666464484
transform 1 0 14812 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_159
timestamp 1666464484
transform 1 0 15732 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_167
timestamp 1666464484
transform 1 0 16468 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_169
timestamp 1666464484
transform 1 0 16652 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_37_180
timestamp 1666464484
transform 1 0 17664 0 -1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_37_192
timestamp 1666464484
transform 1 0 18768 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_211
timestamp 1666464484
transform 1 0 20516 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_37_223
timestamp 1666464484
transform 1 0 21620 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_225
timestamp 1666464484
transform 1 0 21804 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_230
timestamp 1666464484
transform 1 0 22264 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_37_242
timestamp 1666464484
transform 1 0 23368 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_37_247
timestamp 1666464484
transform 1 0 23828 0 -1 22848
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_37_263
timestamp 1666464484
transform 1 0 25300 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_275
timestamp 1666464484
transform 1 0 26404 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_279
timestamp 1666464484
transform 1 0 26772 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_281
timestamp 1666464484
transform 1 0 26956 0 -1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_37_307
timestamp 1666464484
transform 1 0 29348 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_319
timestamp 1666464484
transform 1 0 30452 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_37_330
timestamp 1666464484
transform 1 0 31464 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_37_337
timestamp 1666464484
transform 1 0 32108 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_348
timestamp 1666464484
transform 1 0 33120 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_359
timestamp 1666464484
transform 1 0 34132 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_363
timestamp 1666464484
transform 1 0 34500 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_3
timestamp 1666464484
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_15
timestamp 1666464484
transform 1 0 2484 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_26
timestamp 1666464484
transform 1 0 3496 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_29
timestamp 1666464484
transform 1 0 3772 0 1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_38_40
timestamp 1666464484
transform 1 0 4784 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_52
timestamp 1666464484
transform 1 0 5888 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_38_60
timestamp 1666464484
transform 1 0 6624 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_38_71
timestamp 1666464484
transform 1 0 7636 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_82
timestamp 1666464484
transform 1 0 8648 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_85
timestamp 1666464484
transform 1 0 8924 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_38_91
timestamp 1666464484
transform 1 0 9476 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_38_120
timestamp 1666464484
transform 1 0 12144 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_135
timestamp 1666464484
transform 1 0 13524 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_139
timestamp 1666464484
transform 1 0 13892 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_141
timestamp 1666464484
transform 1 0 14076 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_38_149
timestamp 1666464484
transform 1 0 14812 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_38_159
timestamp 1666464484
transform 1 0 15732 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_169
timestamp 1666464484
transform 1 0 16652 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_175
timestamp 1666464484
transform 1 0 17204 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_192
timestamp 1666464484
transform 1 0 18768 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_197
timestamp 1666464484
transform 1 0 19228 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_38_204
timestamp 1666464484
transform 1 0 19872 0 1 22848
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_38_232
timestamp 1666464484
transform 1 0 22448 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_244
timestamp 1666464484
transform 1 0 23552 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_253
timestamp 1666464484
transform 1 0 24380 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_263
timestamp 1666464484
transform 1 0 25300 0 1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_38_270
timestamp 1666464484
transform 1 0 25944 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_282
timestamp 1666464484
transform 1 0 27048 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_286
timestamp 1666464484
transform 1 0 27416 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_296
timestamp 1666464484
transform 1 0 28336 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_38_305
timestamp 1666464484
transform 1 0 29164 0 1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_38_309
timestamp 1666464484
transform 1 0 29532 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_321
timestamp 1666464484
transform 1 0 30636 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_338
timestamp 1666464484
transform 1 0 32200 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_349
timestamp 1666464484
transform 1 0 33212 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_356
timestamp 1666464484
transform 1 0 33856 0 1 22848
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_39_3
timestamp 1666464484
transform 1 0 1380 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_39_15
timestamp 1666464484
transform 1 0 2484 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_39
timestamp 1666464484
transform 1 0 4692 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_50
timestamp 1666464484
transform 1 0 5704 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_39_57
timestamp 1666464484
transform 1 0 6348 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_61
timestamp 1666464484
transform 1 0 6716 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_81
timestamp 1666464484
transform 1 0 8556 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_91
timestamp 1666464484
transform 1 0 9476 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_39_100
timestamp 1666464484
transform 1 0 10304 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_113
timestamp 1666464484
transform 1 0 11500 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_39_135
timestamp 1666464484
transform 1 0 13524 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_141
timestamp 1666464484
transform 1 0 14076 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_145
timestamp 1666464484
transform 1 0 14444 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_157
timestamp 1666464484
transform 1 0 15548 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_166
timestamp 1666464484
transform 1 0 16376 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_39_169
timestamp 1666464484
transform 1 0 16652 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_181
timestamp 1666464484
transform 1 0 17756 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_185
timestamp 1666464484
transform 1 0 18124 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_206
timestamp 1666464484
transform 1 0 20056 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_215
timestamp 1666464484
transform 1 0 20884 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_223
timestamp 1666464484
transform 1 0 21620 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_225
timestamp 1666464484
transform 1 0 21804 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_39_236
timestamp 1666464484
transform 1 0 22816 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_248
timestamp 1666464484
transform 1 0 23920 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_260
timestamp 1666464484
transform 1 0 25024 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_272
timestamp 1666464484
transform 1 0 26128 0 -1 23936
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_39_281
timestamp 1666464484
transform 1 0 26956 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_293
timestamp 1666464484
transform 1 0 28060 0 -1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_39_319
timestamp 1666464484
transform 1 0 30452 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_331
timestamp 1666464484
transform 1 0 31556 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_335
timestamp 1666464484
transform 1 0 31924 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_337
timestamp 1666464484
transform 1 0 32108 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_349
timestamp 1666464484
transform 1 0 33212 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_39_361
timestamp 1666464484
transform 1 0 34316 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_40_3
timestamp 1666464484
transform 1 0 1380 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_11
timestamp 1666464484
transform 1 0 2116 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_17
timestamp 1666464484
transform 1 0 2668 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_26
timestamp 1666464484
transform 1 0 3496 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_29
timestamp 1666464484
transform 1 0 3772 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_39
timestamp 1666464484
transform 1 0 4692 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_50
timestamp 1666464484
transform 1 0 5704 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_58
timestamp 1666464484
transform 1 0 6440 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_82
timestamp 1666464484
transform 1 0 8648 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_85
timestamp 1666464484
transform 1 0 8924 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_97
timestamp 1666464484
transform 1 0 10028 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_109
timestamp 1666464484
transform 1 0 11132 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_117
timestamp 1666464484
transform 1 0 11868 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_121
timestamp 1666464484
transform 1 0 12236 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_133
timestamp 1666464484
transform 1 0 13340 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_139
timestamp 1666464484
transform 1 0 13892 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_141
timestamp 1666464484
transform 1 0 14076 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_40_150
timestamp 1666464484
transform 1 0 14904 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_156
timestamp 1666464484
transform 1 0 15456 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_40_162
timestamp 1666464484
transform 1 0 16008 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_40_170
timestamp 1666464484
transform 1 0 16744 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_40_176
timestamp 1666464484
transform 1 0 17296 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_186
timestamp 1666464484
transform 1 0 18216 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_194
timestamp 1666464484
transform 1 0 18952 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_197
timestamp 1666464484
transform 1 0 19228 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_40_209
timestamp 1666464484
transform 1 0 20332 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_216
timestamp 1666464484
transform 1 0 20976 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_236
timestamp 1666464484
transform 1 0 22816 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_246
timestamp 1666464484
transform 1 0 23736 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_40_253
timestamp 1666464484
transform 1 0 24380 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_261
timestamp 1666464484
transform 1 0 25116 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_265
timestamp 1666464484
transform 1 0 25484 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_277
timestamp 1666464484
transform 1 0 26588 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_289
timestamp 1666464484
transform 1 0 27692 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_301
timestamp 1666464484
transform 1 0 28796 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_307
timestamp 1666464484
transform 1 0 29348 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_40_309
timestamp 1666464484
transform 1 0 29532 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_317
timestamp 1666464484
transform 1 0 30268 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_325
timestamp 1666464484
transform 1 0 31004 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_337
timestamp 1666464484
transform 1 0 32108 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_349
timestamp 1666464484
transform 1 0 33212 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_40_361
timestamp 1666464484
transform 1 0 34316 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_41_3
timestamp 1666464484
transform 1 0 1380 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_11
timestamp 1666464484
transform 1 0 2116 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_32
timestamp 1666464484
transform 1 0 4048 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_41_49
timestamp 1666464484
transform 1 0 5612 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_55
timestamp 1666464484
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_57
timestamp 1666464484
transform 1 0 6348 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_61
timestamp 1666464484
transform 1 0 6716 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_75
timestamp 1666464484
transform 1 0 8004 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_87
timestamp 1666464484
transform 1 0 9108 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_99
timestamp 1666464484
transform 1 0 10212 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_41_111
timestamp 1666464484
transform 1 0 11316 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_113
timestamp 1666464484
transform 1 0 11500 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_125
timestamp 1666464484
transform 1 0 12604 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_137
timestamp 1666464484
transform 1 0 13708 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_157
timestamp 1666464484
transform 1 0 15548 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_164
timestamp 1666464484
transform 1 0 16192 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_41_169
timestamp 1666464484
transform 1 0 16652 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_41_181
timestamp 1666464484
transform 1 0 17756 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_201
timestamp 1666464484
transform 1 0 19596 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_41_213
timestamp 1666464484
transform 1 0 20700 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_41_222
timestamp 1666464484
transform 1 0 21528 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_225
timestamp 1666464484
transform 1 0 21804 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_41_246
timestamp 1666464484
transform 1 0 23736 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_41_258
timestamp 1666464484
transform 1 0 24840 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_265
timestamp 1666464484
transform 1 0 25484 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_269
timestamp 1666464484
transform 1 0 25852 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_276
timestamp 1666464484
transform 1 0 26496 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_41_281
timestamp 1666464484
transform 1 0 26956 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_293
timestamp 1666464484
transform 1 0 28060 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_41_305
timestamp 1666464484
transform 1 0 29164 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_313
timestamp 1666464484
transform 1 0 29900 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_331
timestamp 1666464484
transform 1 0 31556 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_335
timestamp 1666464484
transform 1 0 31924 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_337
timestamp 1666464484
transform 1 0 32108 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_349
timestamp 1666464484
transform 1 0 33212 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_41_361
timestamp 1666464484
transform 1 0 34316 0 -1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_42_3
timestamp 1666464484
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_15
timestamp 1666464484
transform 1 0 2484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_27
timestamp 1666464484
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_42_29
timestamp 1666464484
transform 1 0 3772 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_35
timestamp 1666464484
transform 1 0 4324 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_47
timestamp 1666464484
transform 1 0 5428 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_42_59
timestamp 1666464484
transform 1 0 6532 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_64
timestamp 1666464484
transform 1 0 6992 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_76
timestamp 1666464484
transform 1 0 8096 0 1 25024
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_42_85
timestamp 1666464484
transform 1 0 8924 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_97
timestamp 1666464484
transform 1 0 10028 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_109
timestamp 1666464484
transform 1 0 11132 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_117
timestamp 1666464484
transform 1 0 11868 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_127
timestamp 1666464484
transform 1 0 12788 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_139
timestamp 1666464484
transform 1 0 13892 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_141
timestamp 1666464484
transform 1 0 14076 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_158
timestamp 1666464484
transform 1 0 15640 0 1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_42_166
timestamp 1666464484
transform 1 0 16376 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_178
timestamp 1666464484
transform 1 0 17480 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_190
timestamp 1666464484
transform 1 0 18584 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_42_197
timestamp 1666464484
transform 1 0 19228 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_42_219
timestamp 1666464484
transform 1 0 21252 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_243
timestamp 1666464484
transform 1 0 23460 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_251
timestamp 1666464484
transform 1 0 24196 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_42_253
timestamp 1666464484
transform 1 0 24380 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_42_261
timestamp 1666464484
transform 1 0 25116 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_269
timestamp 1666464484
transform 1 0 25852 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_278
timestamp 1666464484
transform 1 0 26680 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_42_287
timestamp 1666464484
transform 1 0 27508 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_293
timestamp 1666464484
transform 1 0 28060 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_297
timestamp 1666464484
transform 1 0 28428 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_42_305
timestamp 1666464484
transform 1 0 29164 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_42_309
timestamp 1666464484
transform 1 0 29532 0 1 25024
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_42_332
timestamp 1666464484
transform 1 0 31648 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_344
timestamp 1666464484
transform 1 0 32752 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_356
timestamp 1666464484
transform 1 0 33856 0 1 25024
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_43_3
timestamp 1666464484
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_15
timestamp 1666464484
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_27
timestamp 1666464484
transform 1 0 3588 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_39
timestamp 1666464484
transform 1 0 4692 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_51
timestamp 1666464484
transform 1 0 5796 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_55
timestamp 1666464484
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_57
timestamp 1666464484
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_69
timestamp 1666464484
transform 1 0 7452 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_81
timestamp 1666464484
transform 1 0 8556 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_89
timestamp 1666464484
transform 1 0 9292 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_97
timestamp 1666464484
transform 1 0 10028 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_43_105
timestamp 1666464484
transform 1 0 10764 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_111
timestamp 1666464484
transform 1 0 11316 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_43_113
timestamp 1666464484
transform 1 0 11500 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_43_126
timestamp 1666464484
transform 1 0 12696 0 -1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_43_136
timestamp 1666464484
transform 1 0 13616 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_148
timestamp 1666464484
transform 1 0 14720 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_160
timestamp 1666464484
transform 1 0 15824 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_169
timestamp 1666464484
transform 1 0 16652 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_177
timestamp 1666464484
transform 1 0 17388 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_181
timestamp 1666464484
transform 1 0 17756 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_202
timestamp 1666464484
transform 1 0 19688 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_43_214
timestamp 1666464484
transform 1 0 20792 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_222
timestamp 1666464484
transform 1 0 21528 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_225
timestamp 1666464484
transform 1 0 21804 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_43_246
timestamp 1666464484
transform 1 0 23736 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_43_257
timestamp 1666464484
transform 1 0 24748 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_267
timestamp 1666464484
transform 1 0 25668 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_43_278
timestamp 1666464484
transform 1 0 26680 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_281
timestamp 1666464484
transform 1 0 26956 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_43_290
timestamp 1666464484
transform 1 0 27784 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_298
timestamp 1666464484
transform 1 0 28520 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_319
timestamp 1666464484
transform 1 0 30452 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_331
timestamp 1666464484
transform 1 0 31556 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_335
timestamp 1666464484
transform 1 0 31924 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_43_337
timestamp 1666464484
transform 1 0 32108 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_43_345
timestamp 1666464484
transform 1 0 32844 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_357
timestamp 1666464484
transform 1 0 33948 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_363
timestamp 1666464484
transform 1 0 34500 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_3
timestamp 1666464484
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_15
timestamp 1666464484
transform 1 0 2484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp 1666464484
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_29
timestamp 1666464484
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_41
timestamp 1666464484
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_53
timestamp 1666464484
transform 1 0 5980 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_65
timestamp 1666464484
transform 1 0 7084 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_77
timestamp 1666464484
transform 1 0 8188 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_83
timestamp 1666464484
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_85
timestamp 1666464484
transform 1 0 8924 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_93
timestamp 1666464484
transform 1 0 9660 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_105
timestamp 1666464484
transform 1 0 10764 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_116
timestamp 1666464484
transform 1 0 11776 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_120
timestamp 1666464484
transform 1 0 12144 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_128
timestamp 1666464484
transform 1 0 12880 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_44_137
timestamp 1666464484
transform 1 0 13708 0 1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_44_141
timestamp 1666464484
transform 1 0 14076 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_153
timestamp 1666464484
transform 1 0 15180 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_157
timestamp 1666464484
transform 1 0 15548 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_164
timestamp 1666464484
transform 1 0 16192 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_184
timestamp 1666464484
transform 1 0 18032 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_44_194
timestamp 1666464484
transform 1 0 18952 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_197
timestamp 1666464484
transform 1 0 19228 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_209
timestamp 1666464484
transform 1 0 20332 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_213
timestamp 1666464484
transform 1 0 20700 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_234
timestamp 1666464484
transform 1 0 22632 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_246
timestamp 1666464484
transform 1 0 23736 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_44_253
timestamp 1666464484
transform 1 0 24380 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_44_270
timestamp 1666464484
transform 1 0 25944 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_44_283
timestamp 1666464484
transform 1 0 27140 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_44_293
timestamp 1666464484
transform 1 0 28060 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_299
timestamp 1666464484
transform 1 0 28612 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_306
timestamp 1666464484
transform 1 0 29256 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_309
timestamp 1666464484
transform 1 0 29532 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_313
timestamp 1666464484
transform 1 0 29900 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_334
timestamp 1666464484
transform 1 0 31832 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_346
timestamp 1666464484
transform 1 0 32936 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_358
timestamp 1666464484
transform 1 0 34040 0 1 26112
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_45_3
timestamp 1666464484
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_15
timestamp 1666464484
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_27
timestamp 1666464484
transform 1 0 3588 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_39
timestamp 1666464484
transform 1 0 4692 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_51
timestamp 1666464484
transform 1 0 5796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_55
timestamp 1666464484
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_57
timestamp 1666464484
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_69
timestamp 1666464484
transform 1 0 7452 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_45_81
timestamp 1666464484
transform 1 0 8556 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_45_92
timestamp 1666464484
transform 1 0 9568 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_104
timestamp 1666464484
transform 1 0 10672 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_113
timestamp 1666464484
transform 1 0 11500 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_121
timestamp 1666464484
transform 1 0 12236 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_45_133
timestamp 1666464484
transform 1 0 13340 0 -1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_45_139
timestamp 1666464484
transform 1 0 13892 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_151
timestamp 1666464484
transform 1 0 14996 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_155
timestamp 1666464484
transform 1 0 15364 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_45_161
timestamp 1666464484
transform 1 0 15916 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_167
timestamp 1666464484
transform 1 0 16468 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_169
timestamp 1666464484
transform 1 0 16652 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_181
timestamp 1666464484
transform 1 0 17756 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_185
timestamp 1666464484
transform 1 0 18124 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_45_206
timestamp 1666464484
transform 1 0 20056 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_212
timestamp 1666464484
transform 1 0 20608 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_219
timestamp 1666464484
transform 1 0 21252 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_223
timestamp 1666464484
transform 1 0 21620 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_45_225
timestamp 1666464484
transform 1 0 21804 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_236
timestamp 1666464484
transform 1 0 22816 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_248
timestamp 1666464484
transform 1 0 23920 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_45_256
timestamp 1666464484
transform 1 0 24656 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_45_276
timestamp 1666464484
transform 1 0 26496 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_45_281
timestamp 1666464484
transform 1 0 26956 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_288
timestamp 1666464484
transform 1 0 27600 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_300
timestamp 1666464484
transform 1 0 28704 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_45_308
timestamp 1666464484
transform 1 0 29440 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_45_330
timestamp 1666464484
transform 1 0 31464 0 -1 27200
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_45_337
timestamp 1666464484
transform 1 0 32108 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_349
timestamp 1666464484
transform 1 0 33212 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_45_361
timestamp 1666464484
transform 1 0 34316 0 -1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_46_3
timestamp 1666464484
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_15
timestamp 1666464484
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_27
timestamp 1666464484
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_29
timestamp 1666464484
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_41
timestamp 1666464484
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_53
timestamp 1666464484
transform 1 0 5980 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_65
timestamp 1666464484
transform 1 0 7084 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_77
timestamp 1666464484
transform 1 0 8188 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_83
timestamp 1666464484
transform 1 0 8740 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_46_85
timestamp 1666464484
transform 1 0 8924 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_46_99
timestamp 1666464484
transform 1 0 10212 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_111
timestamp 1666464484
transform 1 0 11316 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_123
timestamp 1666464484
transform 1 0 12420 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_134
timestamp 1666464484
transform 1 0 13432 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_46_141
timestamp 1666464484
transform 1 0 14076 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_46_152
timestamp 1666464484
transform 1 0 15088 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_160
timestamp 1666464484
transform 1 0 15824 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_167
timestamp 1666464484
transform 1 0 16468 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_187
timestamp 1666464484
transform 1 0 18308 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_195
timestamp 1666464484
transform 1 0 19044 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_197
timestamp 1666464484
transform 1 0 19228 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_209
timestamp 1666464484
transform 1 0 20332 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_221
timestamp 1666464484
transform 1 0 21436 0 1 27200
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_46_236
timestamp 1666464484
transform 1 0 22816 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_248
timestamp 1666464484
transform 1 0 23920 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_253
timestamp 1666464484
transform 1 0 24380 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_46_282
timestamp 1666464484
transform 1 0 27048 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_292
timestamp 1666464484
transform 1 0 27968 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_299
timestamp 1666464484
transform 1 0 28612 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_307
timestamp 1666464484
transform 1 0 29348 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_46_309
timestamp 1666464484
transform 1 0 29532 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_46_327
timestamp 1666464484
transform 1 0 31188 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_339
timestamp 1666464484
transform 1 0 32292 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_351
timestamp 1666464484
transform 1 0 33396 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_363
timestamp 1666464484
transform 1 0 34500 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_3
timestamp 1666464484
transform 1 0 1380 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_15
timestamp 1666464484
transform 1 0 2484 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_27
timestamp 1666464484
transform 1 0 3588 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_39
timestamp 1666464484
transform 1 0 4692 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_51
timestamp 1666464484
transform 1 0 5796 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_55
timestamp 1666464484
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_57
timestamp 1666464484
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_47_69
timestamp 1666464484
transform 1 0 7452 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_47_78
timestamp 1666464484
transform 1 0 8280 0 -1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_47_89
timestamp 1666464484
transform 1 0 9292 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_101
timestamp 1666464484
transform 1 0 10396 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_47_109
timestamp 1666464484
transform 1 0 11132 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_47_113
timestamp 1666464484
transform 1 0 11500 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_134
timestamp 1666464484
transform 1 0 13432 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_47_143
timestamp 1666464484
transform 1 0 14260 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_47_151
timestamp 1666464484
transform 1 0 14996 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_47_162
timestamp 1666464484
transform 1 0 16008 0 -1 28288
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_47_169
timestamp 1666464484
transform 1 0 16652 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_181
timestamp 1666464484
transform 1 0 17756 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_193
timestamp 1666464484
transform 1 0 18860 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_47_200
timestamp 1666464484
transform 1 0 19504 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_47_213
timestamp 1666464484
transform 1 0 20700 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_47_221
timestamp 1666464484
transform 1 0 21436 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_47_225
timestamp 1666464484
transform 1 0 21804 0 -1 28288
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_47_237
timestamp 1666464484
transform 1 0 22908 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_249
timestamp 1666464484
transform 1 0 24012 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_257
timestamp 1666464484
transform 1 0 24748 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_47_274
timestamp 1666464484
transform 1 0 26312 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_47_281
timestamp 1666464484
transform 1 0 26956 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_47_288
timestamp 1666464484
transform 1 0 27600 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_300
timestamp 1666464484
transform 1 0 28704 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_47_312
timestamp 1666464484
transform 1 0 29808 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_319
timestamp 1666464484
transform 1 0 30452 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_331
timestamp 1666464484
transform 1 0 31556 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_335
timestamp 1666464484
transform 1 0 31924 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_337
timestamp 1666464484
transform 1 0 32108 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_349
timestamp 1666464484
transform 1 0 33212 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_47_361
timestamp 1666464484
transform 1 0 34316 0 -1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_48_3
timestamp 1666464484
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_15
timestamp 1666464484
transform 1 0 2484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 1666464484
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_29
timestamp 1666464484
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_41
timestamp 1666464484
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_53
timestamp 1666464484
transform 1 0 5980 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_65
timestamp 1666464484
transform 1 0 7084 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_77
timestamp 1666464484
transform 1 0 8188 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_83
timestamp 1666464484
transform 1 0 8740 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_48_85
timestamp 1666464484
transform 1 0 8924 0 1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_48_90
timestamp 1666464484
transform 1 0 9384 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_102
timestamp 1666464484
transform 1 0 10488 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_106
timestamp 1666464484
transform 1 0 10856 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_124
timestamp 1666464484
transform 1 0 12512 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_135
timestamp 1666464484
transform 1 0 13524 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_139
timestamp 1666464484
transform 1 0 13892 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_48_141
timestamp 1666464484
transform 1 0 14076 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_48_157
timestamp 1666464484
transform 1 0 15548 0 1 28288
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_48_170
timestamp 1666464484
transform 1 0 16744 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_182
timestamp 1666464484
transform 1 0 17848 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_48_194
timestamp 1666464484
transform 1 0 18952 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_197
timestamp 1666464484
transform 1 0 19228 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_201
timestamp 1666464484
transform 1 0 19596 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_207
timestamp 1666464484
transform 1 0 20148 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_48_218
timestamp 1666464484
transform 1 0 21160 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_48_226
timestamp 1666464484
transform 1 0 21896 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_250
timestamp 1666464484
transform 1 0 24104 0 1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_48_253
timestamp 1666464484
transform 1 0 24380 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_265
timestamp 1666464484
transform 1 0 25484 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_271
timestamp 1666464484
transform 1 0 26036 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_48_293
timestamp 1666464484
transform 1 0 28060 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_48_304
timestamp 1666464484
transform 1 0 29072 0 1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_48_309
timestamp 1666464484
transform 1 0 29532 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_321
timestamp 1666464484
transform 1 0 30636 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_333
timestamp 1666464484
transform 1 0 31740 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_345
timestamp 1666464484
transform 1 0 32844 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_357
timestamp 1666464484
transform 1 0 33948 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_363
timestamp 1666464484
transform 1 0 34500 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_3
timestamp 1666464484
transform 1 0 1380 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_15
timestamp 1666464484
transform 1 0 2484 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_27
timestamp 1666464484
transform 1 0 3588 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_39
timestamp 1666464484
transform 1 0 4692 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_51
timestamp 1666464484
transform 1 0 5796 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_55
timestamp 1666464484
transform 1 0 6164 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_57
timestamp 1666464484
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_69
timestamp 1666464484
transform 1 0 7452 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_73
timestamp 1666464484
transform 1 0 7820 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_80
timestamp 1666464484
transform 1 0 8464 0 -1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_49_92
timestamp 1666464484
transform 1 0 9568 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_104
timestamp 1666464484
transform 1 0 10672 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_49_113
timestamp 1666464484
transform 1 0 11500 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_49_136
timestamp 1666464484
transform 1 0 13616 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_144
timestamp 1666464484
transform 1 0 14352 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_151
timestamp 1666464484
transform 1 0 14996 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_49_160
timestamp 1666464484
transform 1 0 15824 0 -1 29376
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_49_169
timestamp 1666464484
transform 1 0 16652 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_203
timestamp 1666464484
transform 1 0 19780 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_215
timestamp 1666464484
transform 1 0 20884 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_49_222
timestamp 1666464484
transform 1 0 21528 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_225
timestamp 1666464484
transform 1 0 21804 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_236
timestamp 1666464484
transform 1 0 22816 0 -1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_49_246
timestamp 1666464484
transform 1 0 23736 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_258
timestamp 1666464484
transform 1 0 24840 0 -1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_49_267
timestamp 1666464484
transform 1 0 25668 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_49_279
timestamp 1666464484
transform 1 0 26772 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_281
timestamp 1666464484
transform 1 0 26956 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_285
timestamp 1666464484
transform 1 0 27324 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_289
timestamp 1666464484
transform 1 0 27692 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_298
timestamp 1666464484
transform 1 0 28520 0 -1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_49_307
timestamp 1666464484
transform 1 0 29348 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_319
timestamp 1666464484
transform 1 0 30452 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_331
timestamp 1666464484
transform 1 0 31556 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_335
timestamp 1666464484
transform 1 0 31924 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_337
timestamp 1666464484
transform 1 0 32108 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_349
timestamp 1666464484
transform 1 0 33212 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_49_361
timestamp 1666464484
transform 1 0 34316 0 -1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_50_3
timestamp 1666464484
transform 1 0 1380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_15
timestamp 1666464484
transform 1 0 2484 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_27
timestamp 1666464484
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_29
timestamp 1666464484
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_41
timestamp 1666464484
transform 1 0 4876 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_53
timestamp 1666464484
transform 1 0 5980 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_65
timestamp 1666464484
transform 1 0 7084 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_77
timestamp 1666464484
transform 1 0 8188 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_83
timestamp 1666464484
transform 1 0 8740 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_85
timestamp 1666464484
transform 1 0 8924 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_89
timestamp 1666464484
transform 1 0 9292 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_96
timestamp 1666464484
transform 1 0 9936 0 1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_50_104
timestamp 1666464484
transform 1 0 10672 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_116
timestamp 1666464484
transform 1 0 11776 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_124
timestamp 1666464484
transform 1 0 12512 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_50_132
timestamp 1666464484
transform 1 0 13248 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_50_141
timestamp 1666464484
transform 1 0 14076 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_145
timestamp 1666464484
transform 1 0 14444 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_153
timestamp 1666464484
transform 1 0 15180 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_165
timestamp 1666464484
transform 1 0 16284 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_177
timestamp 1666464484
transform 1 0 17388 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_189
timestamp 1666464484
transform 1 0 18492 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_195
timestamp 1666464484
transform 1 0 19044 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_50_197
timestamp 1666464484
transform 1 0 19228 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_212
timestamp 1666464484
transform 1 0 20608 0 1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_50_223
timestamp 1666464484
transform 1 0 21620 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_235
timestamp 1666464484
transform 1 0 22724 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_247
timestamp 1666464484
transform 1 0 23828 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_251
timestamp 1666464484
transform 1 0 24196 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_253
timestamp 1666464484
transform 1 0 24380 0 1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_50_263
timestamp 1666464484
transform 1 0 25300 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_275
timestamp 1666464484
transform 1 0 26404 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_283
timestamp 1666464484
transform 1 0 27140 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_292
timestamp 1666464484
transform 1 0 27968 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_303
timestamp 1666464484
transform 1 0 28980 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_307
timestamp 1666464484
transform 1 0 29348 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_309
timestamp 1666464484
transform 1 0 29532 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_321
timestamp 1666464484
transform 1 0 30636 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_333
timestamp 1666464484
transform 1 0 31740 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_345
timestamp 1666464484
transform 1 0 32844 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_357
timestamp 1666464484
transform 1 0 33948 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_363
timestamp 1666464484
transform 1 0 34500 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_3
timestamp 1666464484
transform 1 0 1380 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_15
timestamp 1666464484
transform 1 0 2484 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_27
timestamp 1666464484
transform 1 0 3588 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_39
timestamp 1666464484
transform 1 0 4692 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_51
timestamp 1666464484
transform 1 0 5796 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_55
timestamp 1666464484
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_57
timestamp 1666464484
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_69
timestamp 1666464484
transform 1 0 7452 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_81
timestamp 1666464484
transform 1 0 8556 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_93
timestamp 1666464484
transform 1 0 9660 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_105
timestamp 1666464484
transform 1 0 10764 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_111
timestamp 1666464484
transform 1 0 11316 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_113
timestamp 1666464484
transform 1 0 11500 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_125
timestamp 1666464484
transform 1 0 12604 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_133
timestamp 1666464484
transform 1 0 13340 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_156
timestamp 1666464484
transform 1 0 15456 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_169
timestamp 1666464484
transform 1 0 16652 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_181
timestamp 1666464484
transform 1 0 17756 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_187
timestamp 1666464484
transform 1 0 18308 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_210
timestamp 1666464484
transform 1 0 20424 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_51_217
timestamp 1666464484
transform 1 0 21068 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_223
timestamp 1666464484
transform 1 0 21620 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_225
timestamp 1666464484
transform 1 0 21804 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_237
timestamp 1666464484
transform 1 0 22908 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_249
timestamp 1666464484
transform 1 0 24012 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_255
timestamp 1666464484
transform 1 0 24564 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_51_273
timestamp 1666464484
transform 1 0 26220 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_279
timestamp 1666464484
transform 1 0 26772 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_51_281
timestamp 1666464484
transform 1 0 26956 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_292
timestamp 1666464484
transform 1 0 27968 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_304
timestamp 1666464484
transform 1 0 29072 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_314
timestamp 1666464484
transform 1 0 29992 0 -1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_51_323
timestamp 1666464484
transform 1 0 30820 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_51_335
timestamp 1666464484
transform 1 0 31924 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_337
timestamp 1666464484
transform 1 0 32108 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_349
timestamp 1666464484
transform 1 0 33212 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_51_361
timestamp 1666464484
transform 1 0 34316 0 -1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_52_3
timestamp 1666464484
transform 1 0 1380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_15
timestamp 1666464484
transform 1 0 2484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_27
timestamp 1666464484
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_29
timestamp 1666464484
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_41
timestamp 1666464484
transform 1 0 4876 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_53
timestamp 1666464484
transform 1 0 5980 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_65
timestamp 1666464484
transform 1 0 7084 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_77
timestamp 1666464484
transform 1 0 8188 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_83
timestamp 1666464484
transform 1 0 8740 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_85
timestamp 1666464484
transform 1 0 8924 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_92
timestamp 1666464484
transform 1 0 9568 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_99
timestamp 1666464484
transform 1 0 10212 0 1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_52_106
timestamp 1666464484
transform 1 0 10856 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_118
timestamp 1666464484
transform 1 0 11960 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_130
timestamp 1666464484
transform 1 0 13064 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_52_138
timestamp 1666464484
transform 1 0 13800 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_141
timestamp 1666464484
transform 1 0 14076 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_145
timestamp 1666464484
transform 1 0 14444 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_167
timestamp 1666464484
transform 1 0 16468 0 1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_52_174
timestamp 1666464484
transform 1 0 17112 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_186
timestamp 1666464484
transform 1 0 18216 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_52_194
timestamp 1666464484
transform 1 0 18952 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_52_197
timestamp 1666464484
transform 1 0 19228 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_52_209
timestamp 1666464484
transform 1 0 20332 0 1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_52_217
timestamp 1666464484
transform 1 0 21068 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_229
timestamp 1666464484
transform 1 0 22172 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_235
timestamp 1666464484
transform 1 0 22724 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_52_242
timestamp 1666464484
transform 1 0 23368 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_52_250
timestamp 1666464484
transform 1 0 24104 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_52_253
timestamp 1666464484
transform 1 0 24380 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_52_276
timestamp 1666464484
transform 1 0 26496 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_52_284
timestamp 1666464484
transform 1 0 27232 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_303
timestamp 1666464484
transform 1 0 28980 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_307
timestamp 1666464484
transform 1 0 29348 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_309
timestamp 1666464484
transform 1 0 29532 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_321
timestamp 1666464484
transform 1 0 30636 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_333
timestamp 1666464484
transform 1 0 31740 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_345
timestamp 1666464484
transform 1 0 32844 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_357
timestamp 1666464484
transform 1 0 33948 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_363
timestamp 1666464484
transform 1 0 34500 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_3
timestamp 1666464484
transform 1 0 1380 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_15
timestamp 1666464484
transform 1 0 2484 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_27
timestamp 1666464484
transform 1 0 3588 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_39
timestamp 1666464484
transform 1 0 4692 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_51
timestamp 1666464484
transform 1 0 5796 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_55
timestamp 1666464484
transform 1 0 6164 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_57
timestamp 1666464484
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_69
timestamp 1666464484
transform 1 0 7452 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_81
timestamp 1666464484
transform 1 0 8556 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_92
timestamp 1666464484
transform 1 0 9568 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_53_110
timestamp 1666464484
transform 1 0 11224 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_53_113
timestamp 1666464484
transform 1 0 11500 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_125
timestamp 1666464484
transform 1 0 12604 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_136
timestamp 1666464484
transform 1 0 13616 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_53_156
timestamp 1666464484
transform 1 0 15456 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_162
timestamp 1666464484
transform 1 0 16008 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_53_166
timestamp 1666464484
transform 1 0 16376 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_169
timestamp 1666464484
transform 1 0 16652 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_175
timestamp 1666464484
transform 1 0 17204 0 -1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_53_182
timestamp 1666464484
transform 1 0 17848 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_194
timestamp 1666464484
transform 1 0 18952 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_53_222
timestamp 1666464484
transform 1 0 21528 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_225
timestamp 1666464484
transform 1 0 21804 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_246
timestamp 1666464484
transform 1 0 23736 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_250
timestamp 1666464484
transform 1 0 24104 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_258
timestamp 1666464484
transform 1 0 24840 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_53_271
timestamp 1666464484
transform 1 0 26036 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_53_279
timestamp 1666464484
transform 1 0 26772 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_53_281
timestamp 1666464484
transform 1 0 26956 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_292
timestamp 1666464484
transform 1 0 27968 0 -1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_53_305
timestamp 1666464484
transform 1 0 29164 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_317
timestamp 1666464484
transform 1 0 30268 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_329
timestamp 1666464484
transform 1 0 31372 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_335
timestamp 1666464484
transform 1 0 31924 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_337
timestamp 1666464484
transform 1 0 32108 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_349
timestamp 1666464484
transform 1 0 33212 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_53_361
timestamp 1666464484
transform 1 0 34316 0 -1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_54_3
timestamp 1666464484
transform 1 0 1380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_15
timestamp 1666464484
transform 1 0 2484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_27
timestamp 1666464484
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_29
timestamp 1666464484
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_41
timestamp 1666464484
transform 1 0 4876 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_53
timestamp 1666464484
transform 1 0 5980 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_65
timestamp 1666464484
transform 1 0 7084 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_54_77
timestamp 1666464484
transform 1 0 8188 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_82
timestamp 1666464484
transform 1 0 8648 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_85
timestamp 1666464484
transform 1 0 8924 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_54_98
timestamp 1666464484
transform 1 0 10120 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_54_106
timestamp 1666464484
transform 1 0 10856 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_54_117
timestamp 1666464484
transform 1 0 11868 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_54_138
timestamp 1666464484
transform 1 0 13800 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_141
timestamp 1666464484
transform 1 0 14076 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_54_146
timestamp 1666464484
transform 1 0 14536 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_54_154
timestamp 1666464484
transform 1 0 15272 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_54_162
timestamp 1666464484
transform 1 0 16008 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_180
timestamp 1666464484
transform 1 0 17664 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_54_190
timestamp 1666464484
transform 1 0 18584 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_54_197
timestamp 1666464484
transform 1 0 19228 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_212
timestamp 1666464484
transform 1 0 20608 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_54_220
timestamp 1666464484
transform 1 0 21344 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_54_240
timestamp 1666464484
transform 1 0 23184 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_54_249
timestamp 1666464484
transform 1 0 24012 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_54_253
timestamp 1666464484
transform 1 0 24380 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_54_264
timestamp 1666464484
transform 1 0 25392 0 1 31552
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_54_292
timestamp 1666464484
transform 1 0 27968 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_54_304
timestamp 1666464484
transform 1 0 29072 0 1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_54_309
timestamp 1666464484
transform 1 0 29532 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_321
timestamp 1666464484
transform 1 0 30636 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_333
timestamp 1666464484
transform 1 0 31740 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_345
timestamp 1666464484
transform 1 0 32844 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_357
timestamp 1666464484
transform 1 0 33948 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_363
timestamp 1666464484
transform 1 0 34500 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_3
timestamp 1666464484
transform 1 0 1380 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_15
timestamp 1666464484
transform 1 0 2484 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_27
timestamp 1666464484
transform 1 0 3588 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_39
timestamp 1666464484
transform 1 0 4692 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_51
timestamp 1666464484
transform 1 0 5796 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_55
timestamp 1666464484
transform 1 0 6164 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_57
timestamp 1666464484
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_69
timestamp 1666464484
transform 1 0 7452 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_81
timestamp 1666464484
transform 1 0 8556 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_55_89
timestamp 1666464484
transform 1 0 9292 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_55_97
timestamp 1666464484
transform 1 0 10028 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_55_105
timestamp 1666464484
transform 1 0 10764 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_111
timestamp 1666464484
transform 1 0 11316 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_55_113
timestamp 1666464484
transform 1 0 11500 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_124
timestamp 1666464484
transform 1 0 12512 0 -1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_55_137
timestamp 1666464484
transform 1 0 13708 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_149
timestamp 1666464484
transform 1 0 14812 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_161
timestamp 1666464484
transform 1 0 15916 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_167
timestamp 1666464484
transform 1 0 16468 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_55_169
timestamp 1666464484
transform 1 0 16652 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_180
timestamp 1666464484
transform 1 0 17664 0 -1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_55_187
timestamp 1666464484
transform 1 0 18308 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_199
timestamp 1666464484
transform 1 0 19412 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_55_211
timestamp 1666464484
transform 1 0 20516 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_222
timestamp 1666464484
transform 1 0 21528 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_225
timestamp 1666464484
transform 1 0 21804 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_55_230
timestamp 1666464484
transform 1 0 22264 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_236
timestamp 1666464484
transform 1 0 22816 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_242
timestamp 1666464484
transform 1 0 23368 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_257
timestamp 1666464484
transform 1 0 24748 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_269
timestamp 1666464484
transform 1 0 25852 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_55_277
timestamp 1666464484
transform 1 0 26588 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_55_281
timestamp 1666464484
transform 1 0 26956 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_55_305
timestamp 1666464484
transform 1 0 29164 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_55_313
timestamp 1666464484
transform 1 0 29900 0 -1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_55_320
timestamp 1666464484
transform 1 0 30544 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_332
timestamp 1666464484
transform 1 0 31648 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_55_337
timestamp 1666464484
transform 1 0 32108 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_55_345
timestamp 1666464484
transform 1 0 32844 0 -1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_55_352
timestamp 1666464484
transform 1 0 33488 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_3
timestamp 1666464484
transform 1 0 1380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_15
timestamp 1666464484
transform 1 0 2484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_27
timestamp 1666464484
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_29
timestamp 1666464484
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_41
timestamp 1666464484
transform 1 0 4876 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_53
timestamp 1666464484
transform 1 0 5980 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_65
timestamp 1666464484
transform 1 0 7084 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_77
timestamp 1666464484
transform 1 0 8188 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_83
timestamp 1666464484
transform 1 0 8740 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_85
timestamp 1666464484
transform 1 0 8924 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_100
timestamp 1666464484
transform 1 0 10304 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_112
timestamp 1666464484
transform 1 0 11408 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_124
timestamp 1666464484
transform 1 0 12512 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_136
timestamp 1666464484
transform 1 0 13616 0 1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_56_141
timestamp 1666464484
transform 1 0 14076 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_153
timestamp 1666464484
transform 1 0 15180 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_159
timestamp 1666464484
transform 1 0 15732 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_172
timestamp 1666464484
transform 1 0 16928 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_184
timestamp 1666464484
transform 1 0 18032 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_197
timestamp 1666464484
transform 1 0 19228 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_216
timestamp 1666464484
transform 1 0 20976 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_56_228
timestamp 1666464484
transform 1 0 22080 0 1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_56_233
timestamp 1666464484
transform 1 0 22540 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_245
timestamp 1666464484
transform 1 0 23644 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_251
timestamp 1666464484
transform 1 0 24196 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_253
timestamp 1666464484
transform 1 0 24380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_265
timestamp 1666464484
transform 1 0 25484 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_277
timestamp 1666464484
transform 1 0 26588 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_289
timestamp 1666464484
transform 1 0 27692 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_301
timestamp 1666464484
transform 1 0 28796 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_307
timestamp 1666464484
transform 1 0 29348 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_309
timestamp 1666464484
transform 1 0 29532 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_321
timestamp 1666464484
transform 1 0 30636 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_333
timestamp 1666464484
transform 1 0 31740 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_345
timestamp 1666464484
transform 1 0 32844 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_357
timestamp 1666464484
transform 1 0 33948 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_363
timestamp 1666464484
transform 1 0 34500 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_3
timestamp 1666464484
transform 1 0 1380 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_15
timestamp 1666464484
transform 1 0 2484 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_57_27
timestamp 1666464484
transform 1 0 3588 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_57_29
timestamp 1666464484
transform 1 0 3772 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_57_37
timestamp 1666464484
transform 1 0 4508 0 -1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_57_44
timestamp 1666464484
transform 1 0 5152 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_57
timestamp 1666464484
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_57_69
timestamp 1666464484
transform 1 0 7452 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_57_76
timestamp 1666464484
transform 1 0 8096 0 -1 33728
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_57_85
timestamp 1666464484
transform 1 0 8924 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_97
timestamp 1666464484
transform 1 0 10028 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_103
timestamp 1666464484
transform 1 0 10580 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_108
timestamp 1666464484
transform 1 0 11040 0 -1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_57_113
timestamp 1666464484
transform 1 0 11500 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_125
timestamp 1666464484
transform 1 0 12604 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_57_137
timestamp 1666464484
transform 1 0 13708 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_57_141
timestamp 1666464484
transform 1 0 14076 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_57_147
timestamp 1666464484
transform 1 0 14628 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_159
timestamp 1666464484
transform 1 0 15732 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_57_167
timestamp 1666464484
transform 1 0 16468 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_57_169
timestamp 1666464484
transform 1 0 16652 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_57_175
timestamp 1666464484
transform 1 0 17204 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_187
timestamp 1666464484
transform 1 0 18308 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_57_195
timestamp 1666464484
transform 1 0 19044 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_57_197
timestamp 1666464484
transform 1 0 19228 0 -1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_57_204
timestamp 1666464484
transform 1 0 19872 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_216
timestamp 1666464484
transform 1 0 20976 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_57_225
timestamp 1666464484
transform 1 0 21804 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_231
timestamp 1666464484
transform 1 0 22356 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_236
timestamp 1666464484
transform 1 0 22816 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_248
timestamp 1666464484
transform 1 0 23920 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_57_253
timestamp 1666464484
transform 1 0 24380 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_57_261
timestamp 1666464484
transform 1 0 25116 0 -1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_57_268
timestamp 1666464484
transform 1 0 25760 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_281
timestamp 1666464484
transform 1 0 26956 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_57_293
timestamp 1666464484
transform 1 0 28060 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_57_300
timestamp 1666464484
transform 1 0 28704 0 -1 33728
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_57_309
timestamp 1666464484
transform 1 0 29532 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_321
timestamp 1666464484
transform 1 0 30636 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_327
timestamp 1666464484
transform 1 0 31188 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_332
timestamp 1666464484
transform 1 0 31648 0 -1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_57_337
timestamp 1666464484
transform 1 0 32108 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_349
timestamp 1666464484
transform 1 0 33212 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_57_357
timestamp 1666464484
transform 1 0 33948 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_57_362
timestamp 1666464484
transform 1 0 34408 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1666464484
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1666464484
transform -1 0 34868 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1666464484
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1666464484
transform -1 0 34868 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1666464484
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1666464484
transform -1 0 34868 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1666464484
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1666464484
transform -1 0 34868 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1666464484
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1666464484
transform -1 0 34868 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1666464484
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1666464484
transform -1 0 34868 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1666464484
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1666464484
transform -1 0 34868 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1666464484
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1666464484
transform -1 0 34868 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1666464484
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1666464484
transform -1 0 34868 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1666464484
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1666464484
transform -1 0 34868 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1666464484
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1666464484
transform -1 0 34868 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1666464484
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1666464484
transform -1 0 34868 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1666464484
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1666464484
transform -1 0 34868 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1666464484
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1666464484
transform -1 0 34868 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1666464484
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1666464484
transform -1 0 34868 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1666464484
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1666464484
transform -1 0 34868 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1666464484
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1666464484
transform -1 0 34868 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1666464484
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1666464484
transform -1 0 34868 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1666464484
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1666464484
transform -1 0 34868 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1666464484
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1666464484
transform -1 0 34868 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1666464484
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1666464484
transform -1 0 34868 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1666464484
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1666464484
transform -1 0 34868 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1666464484
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1666464484
transform -1 0 34868 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1666464484
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1666464484
transform -1 0 34868 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1666464484
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1666464484
transform -1 0 34868 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1666464484
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1666464484
transform -1 0 34868 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1666464484
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1666464484
transform -1 0 34868 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1666464484
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1666464484
transform -1 0 34868 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1666464484
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1666464484
transform -1 0 34868 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1666464484
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1666464484
transform -1 0 34868 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1666464484
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1666464484
transform -1 0 34868 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1666464484
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1666464484
transform -1 0 34868 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1666464484
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1666464484
transform -1 0 34868 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1666464484
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1666464484
transform -1 0 34868 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1666464484
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1666464484
transform -1 0 34868 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1666464484
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1666464484
transform -1 0 34868 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1666464484
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1666464484
transform -1 0 34868 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1666464484
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1666464484
transform -1 0 34868 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1666464484
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1666464484
transform -1 0 34868 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1666464484
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1666464484
transform -1 0 34868 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1666464484
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1666464484
transform -1 0 34868 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1666464484
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1666464484
transform -1 0 34868 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1666464484
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1666464484
transform -1 0 34868 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1666464484
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1666464484
transform -1 0 34868 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1666464484
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1666464484
transform -1 0 34868 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1666464484
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1666464484
transform -1 0 34868 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1666464484
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1666464484
transform -1 0 34868 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1666464484
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1666464484
transform -1 0 34868 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1666464484
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1666464484
transform -1 0 34868 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1666464484
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1666464484
transform -1 0 34868 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1666464484
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1666464484
transform -1 0 34868 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1666464484
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1666464484
transform -1 0 34868 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1666464484
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1666464484
transform -1 0 34868 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1666464484
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1666464484
transform -1 0 34868 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1666464484
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1666464484
transform -1 0 34868 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1666464484
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1666464484
transform -1 0 34868 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1666464484
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1666464484
transform -1 0 34868 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1666464484
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1666464484
transform -1 0 34868 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1666464484
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1666464484
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1666464484
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1666464484
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1666464484
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1666464484
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1666464484
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1666464484
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1666464484
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1666464484
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1666464484
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1666464484
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1666464484
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1666464484
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1666464484
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1666464484
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1666464484
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1666464484
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1666464484
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1666464484
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1666464484
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1666464484
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1666464484
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1666464484
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1666464484
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1666464484
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1666464484
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1666464484
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1666464484
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1666464484
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1666464484
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1666464484
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1666464484
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1666464484
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1666464484
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1666464484
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1666464484
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1666464484
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1666464484
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1666464484
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1666464484
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1666464484
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1666464484
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1666464484
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1666464484
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1666464484
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1666464484
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1666464484
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1666464484
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1666464484
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1666464484
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1666464484
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1666464484
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1666464484
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1666464484
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1666464484
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1666464484
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1666464484
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1666464484
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1666464484
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1666464484
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1666464484
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1666464484
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1666464484
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1666464484
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1666464484
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1666464484
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1666464484
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1666464484
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1666464484
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1666464484
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1666464484
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1666464484
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1666464484
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1666464484
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1666464484
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1666464484
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1666464484
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1666464484
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1666464484
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1666464484
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1666464484
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1666464484
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1666464484
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1666464484
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1666464484
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1666464484
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1666464484
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1666464484
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1666464484
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1666464484
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1666464484
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1666464484
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1666464484
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1666464484
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1666464484
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1666464484
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1666464484
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1666464484
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1666464484
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1666464484
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1666464484
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1666464484
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1666464484
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1666464484
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1666464484
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1666464484
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1666464484
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1666464484
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1666464484
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1666464484
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1666464484
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1666464484
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1666464484
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1666464484
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1666464484
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1666464484
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1666464484
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1666464484
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1666464484
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1666464484
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1666464484
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1666464484
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1666464484
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1666464484
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1666464484
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1666464484
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1666464484
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1666464484
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1666464484
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1666464484
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1666464484
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1666464484
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1666464484
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1666464484
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1666464484
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1666464484
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1666464484
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1666464484
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1666464484
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1666464484
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1666464484
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1666464484
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1666464484
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1666464484
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1666464484
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1666464484
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1666464484
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1666464484
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1666464484
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1666464484
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1666464484
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1666464484
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1666464484
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1666464484
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1666464484
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1666464484
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1666464484
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1666464484
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1666464484
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1666464484
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1666464484
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1666464484
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1666464484
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1666464484
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1666464484
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1666464484
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1666464484
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1666464484
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1666464484
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1666464484
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1666464484
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1666464484
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1666464484
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1666464484
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1666464484
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1666464484
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1666464484
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1666464484
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1666464484
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1666464484
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1666464484
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1666464484
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1666464484
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1666464484
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1666464484
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1666464484
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1666464484
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1666464484
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1666464484
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1666464484
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1666464484
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1666464484
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1666464484
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1666464484
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1666464484
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1666464484
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1666464484
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1666464484
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1666464484
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1666464484
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1666464484
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1666464484
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1666464484
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1666464484
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1666464484
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1666464484
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1666464484
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1666464484
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1666464484
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1666464484
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1666464484
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1666464484
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1666464484
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1666464484
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1666464484
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1666464484
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1666464484
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1666464484
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1666464484
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1666464484
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1666464484
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1666464484
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1666464484
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1666464484
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1666464484
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1666464484
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1666464484
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1666464484
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1666464484
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1666464484
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1666464484
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1666464484
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1666464484
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1666464484
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1666464484
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1666464484
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1666464484
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1666464484
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1666464484
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1666464484
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1666464484
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1666464484
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1666464484
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1666464484
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1666464484
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1666464484
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1666464484
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1666464484
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1666464484
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1666464484
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1666464484
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1666464484
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1666464484
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1666464484
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1666464484
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1666464484
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1666464484
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1666464484
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1666464484
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1666464484
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1666464484
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1666464484
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1666464484
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1666464484
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1666464484
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1666464484
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1666464484
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1666464484
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1666464484
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1666464484
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1666464484
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1666464484
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1666464484
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1666464484
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1666464484
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1666464484
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1666464484
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1666464484
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1666464484
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1666464484
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1666464484
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1666464484
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1666464484
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1666464484
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1666464484
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1666464484
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1666464484
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1666464484
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1666464484
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1666464484
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1666464484
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1666464484
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1666464484
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1666464484
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1666464484
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1666464484
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1666464484
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1666464484
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1666464484
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1666464484
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1666464484
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1666464484
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1666464484
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1666464484
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1666464484
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1666464484
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1666464484
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1666464484
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1666464484
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1666464484
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1666464484
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1666464484
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1666464484
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1666464484
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1666464484
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1666464484
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1666464484
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1666464484
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1666464484
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1666464484
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1666464484
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1666464484
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1666464484
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1666464484
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1666464484
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1666464484
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1666464484
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1666464484
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1666464484
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1666464484
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1666464484
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1666464484
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1666464484
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1666464484
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1666464484
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1666464484
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1666464484
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1666464484
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1666464484
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1666464484
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1666464484
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1666464484
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1666464484
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1666464484
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1666464484
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1666464484
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1666464484
transform 1 0 3680 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1666464484
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1666464484
transform 1 0 8832 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1666464484
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1666464484
transform 1 0 13984 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1666464484
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1666464484
transform 1 0 19136 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1666464484
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1666464484
transform 1 0 24288 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1666464484
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1666464484
transform 1 0 29440 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1666464484
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0465_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 2484 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0466_
timestamp 1666464484
transform -1 0 4232 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_6  _0467_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 4416 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__inv_4  _0468_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 5796 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0469_
timestamp 1666464484
transform 1 0 14444 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0470_
timestamp 1666464484
transform 1 0 10396 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0471_
timestamp 1666464484
transform 1 0 12512 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0472_
timestamp 1666464484
transform 1 0 14444 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_4  _0473_
timestamp 1666464484
transform 1 0 16284 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__inv_4  _0474_
timestamp 1666464484
transform 1 0 9568 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0475_
timestamp 1666464484
transform 1 0 13616 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_4  _0476_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 26036 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0477_
timestamp 1666464484
transform -1 0 25944 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0478_
timestamp 1666464484
transform -1 0 28428 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0479_
timestamp 1666464484
transform -1 0 29072 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0480_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 33488 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _0481_
timestamp 1666464484
transform -1 0 30544 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0482__1
timestamp 1666464484
transform -1 0 12696 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0483_
timestamp 1666464484
transform 1 0 4692 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0484_
timestamp 1666464484
transform 1 0 4048 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0485_
timestamp 1666464484
transform -1 0 2576 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__or4b_4  _0486_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 26128 0 -1 3264
box -38 -48 1050 592
use sky130_fd_sc_hd__nor2_1  _0487_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 8280 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__and2_2  _0488_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 5336 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0489_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 9568 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _0490_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 10304 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__nor3b_4  _0491_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 11224 0 -1 16320
box -38 -48 1418 592
use sky130_fd_sc_hd__mux2_1  _0492_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 9200 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0493_
timestamp 1666464484
transform -1 0 9936 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0494_
timestamp 1666464484
transform 1 0 22080 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__or3b_1  _0495_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 11868 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _0496_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 12604 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0497_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 14628 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _0498_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 20700 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _0499_
timestamp 1666464484
transform -1 0 12604 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _0500_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 10580 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or4bb_4  _0501_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__nand2_4  _0502_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 15916 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_4  _0503_
timestamp 1666464484
transform 1 0 14260 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_2  _0504_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 14536 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0505_
timestamp 1666464484
transform -1 0 13616 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _0506_
timestamp 1666464484
transform 1 0 13340 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0507_
timestamp 1666464484
transform 1 0 6072 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _0508_
timestamp 1666464484
transform 1 0 7360 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0509_
timestamp 1666464484
transform 1 0 13524 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0510_
timestamp 1666464484
transform -1 0 13432 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0511_
timestamp 1666464484
transform 1 0 19780 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0512_
timestamp 1666464484
transform 1 0 7268 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _0513_
timestamp 1666464484
transform 1 0 6532 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0514_
timestamp 1666464484
transform 1 0 6716 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _0515_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 6624 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _0516_
timestamp 1666464484
transform -1 0 7360 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0517_
timestamp 1666464484
transform 1 0 18032 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux4_2  _0518_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 8556 0 -1 10880
box -38 -48 1694 592
use sky130_fd_sc_hd__mux2_1  _0519_
timestamp 1666464484
transform 1 0 16928 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux4_2  _0520_
timestamp 1666464484
transform 1 0 12144 0 1 10880
box -38 -48 1694 592
use sky130_fd_sc_hd__mux2_1  _0521_
timestamp 1666464484
transform 1 0 15548 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux4_2  _0522_
timestamp 1666464484
transform 1 0 12328 0 -1 10880
box -38 -48 1694 592
use sky130_fd_sc_hd__mux2_1  _0523_
timestamp 1666464484
transform -1 0 14812 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux4_2  _0524_
timestamp 1666464484
transform 1 0 6532 0 -1 10880
box -38 -48 1694 592
use sky130_fd_sc_hd__mux2_1  _0525_
timestamp 1666464484
transform 1 0 12972 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_2  _0526_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 2576 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__or4b_4  _0527_
timestamp 1666464484
transform 1 0 26404 0 1 3264
box -38 -48 1050 592
use sky130_fd_sc_hd__mux2_2  _0528_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 11040 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_2  _0529_
timestamp 1666464484
transform 1 0 11684 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_2  _0530_
timestamp 1666464484
transform 1 0 12880 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_4  _0531_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 16928 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__nand2_2  _0532_
timestamp 1666464484
transform 1 0 2576 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0533_
timestamp 1666464484
transform 1 0 8832 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_2  _0534_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 5888 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0535_
timestamp 1666464484
transform -1 0 3496 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _0536_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 2944 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0537_
timestamp 1666464484
transform 1 0 1932 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0538_
timestamp 1666464484
transform -1 0 2300 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _0539_
timestamp 1666464484
transform 1 0 2852 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__and3b_2  _0540_
timestamp 1666464484
transform -1 0 3404 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__a41o_1  _0541_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 2668 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0542_
timestamp 1666464484
transform -1 0 4600 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0543_
timestamp 1666464484
transform 1 0 2300 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__or4_4  _0544_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 7544 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0545_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 5520 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _0546_
timestamp 1666464484
transform -1 0 15916 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__and2_2  _0547_
timestamp 1666464484
transform -1 0 13248 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_2  _0548_
timestamp 1666464484
transform -1 0 14260 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _0549_
timestamp 1666464484
transform -1 0 25484 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _0550_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 27508 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _0551_
timestamp 1666464484
transform 1 0 25944 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0552_
timestamp 1666464484
transform 1 0 27140 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _0553_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 27140 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0554_
timestamp 1666464484
transform -1 0 28612 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _0555_
timestamp 1666464484
transform -1 0 27600 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0556_
timestamp 1666464484
transform -1 0 24748 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _0557_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 25116 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _0558_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 26680 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_2  _0559_
timestamp 1666464484
transform 1 0 27140 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__o311a_2  _0560_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 25116 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__a211oi_4  _0561_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 26312 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__a32o_4  _0562_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 26496 0 -1 27200
box -38 -48 1602 592
use sky130_fd_sc_hd__and3_1  _0563_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 28060 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_2  _0564_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 28336 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_2  _0565_
timestamp 1666464484
transform 1 0 28888 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__a311oi_4  _0566_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 27048 0 1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__and2_2  _0567_
timestamp 1666464484
transform 1 0 24748 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0568_
timestamp 1666464484
transform 1 0 24472 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _0569_
timestamp 1666464484
transform -1 0 25668 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0570_
timestamp 1666464484
transform -1 0 27968 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_8  _0571_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 26128 0 1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__nor2_4  _0572_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 27968 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _0573_
timestamp 1666464484
transform -1 0 27692 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _0574_
timestamp 1666464484
transform 1 0 30360 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__and2_2  _0575_
timestamp 1666464484
transform -1 0 29992 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _0576_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 28336 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__o2bb2a_2  _0577_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 27140 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__o31ai_4  _0578_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 26496 0 1 30464
box -38 -48 1602 592
use sky130_fd_sc_hd__o31a_2  _0579_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 27232 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__nor4_4  _0580_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 28980 0 1 30464
box -38 -48 1602 592
use sky130_fd_sc_hd__o311a_4  _0581_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 24656 0 -1 30464
box -38 -48 1602 592
use sky130_fd_sc_hd__and2b_1  _0582_
timestamp 1666464484
transform -1 0 22908 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_2  _0583_
timestamp 1666464484
transform -1 0 23368 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__or3_4  _0584_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 28336 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__o311a_2  _0585_
timestamp 1666464484
transform -1 0 26036 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__xor2_4  _0586_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 25944 0 1 31552
box -38 -48 2062 592
use sky130_fd_sc_hd__xnor2_4  _0587_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 29164 0 -1 32640
box -38 -48 2062 592
use sky130_fd_sc_hd__inv_2  _0588_
timestamp 1666464484
transform -1 0 22540 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0589_
timestamp 1666464484
transform -1 0 19504 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _0590_
timestamp 1666464484
transform 1 0 20240 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0591_
timestamp 1666464484
transform -1 0 21068 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _0592_
timestamp 1666464484
transform 1 0 19688 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _0593_
timestamp 1666464484
transform -1 0 23736 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_4  _0594_
timestamp 1666464484
transform -1 0 24104 0 1 28288
box -38 -48 2062 592
use sky130_fd_sc_hd__a21oi_2  _0595_
timestamp 1666464484
transform -1 0 21620 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__o311a_2  _0596_
timestamp 1666464484
transform 1 0 21988 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0597_
timestamp 1666464484
transform 1 0 20608 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _0598_
timestamp 1666464484
transform -1 0 21160 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0599_
timestamp 1666464484
transform -1 0 21344 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _0600_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 24012 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _0601_
timestamp 1666464484
transform 1 0 22816 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_4  _0602_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 22172 0 -1 31552
box -38 -48 1602 592
use sky130_fd_sc_hd__or3b_1  _0603_
timestamp 1666464484
transform 1 0 24196 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0604_
timestamp 1666464484
transform 1 0 24564 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_4  _0605_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 22080 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__nand2_1  _0606_
timestamp 1666464484
transform -1 0 21528 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__a211oi_4  _0607_
timestamp 1666464484
transform 1 0 20056 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__xnor2_2  _0608_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 20608 0 1 31552
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_1  _0609_
timestamp 1666464484
transform -1 0 17848 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _0610_
timestamp 1666464484
transform -1 0 15824 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__and2_2  _0611_
timestamp 1666464484
transform -1 0 14996 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__or2_4  _0612_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 15180 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_4  _0613_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 19412 0 1 29376
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_4  _0614_
timestamp 1666464484
transform -1 0 19780 0 -1 29376
box -38 -48 2062 592
use sky130_fd_sc_hd__o21ai_1  _0615_
timestamp 1666464484
transform -1 0 13800 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_2  _0616_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 20148 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_4  _0617_
timestamp 1666464484
transform -1 0 20424 0 -1 30464
box -38 -48 2062 592
use sky130_fd_sc_hd__nand2_1  _0618_
timestamp 1666464484
transform -1 0 16376 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__o221ai_4  _0619_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 16468 0 1 30464
box -38 -48 1970 592
use sky130_fd_sc_hd__xnor2_1  _0620_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 20332 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0621_
timestamp 1666464484
transform -1 0 22264 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0622_
timestamp 1666464484
transform 1 0 20700 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__o21bai_1  _0623_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 18032 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_4  _0624_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 17664 0 1 31552
box -38 -48 1326 592
use sky130_fd_sc_hd__a21boi_2  _0625_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 16008 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_4  _0626_
timestamp 1666464484
transform -1 0 15548 0 1 28288
box -38 -48 1234 592
use sky130_fd_sc_hd__or2_4  _0627_
timestamp 1666464484
transform -1 0 13432 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0628_
timestamp 1666464484
transform 1 0 12972 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0629_
timestamp 1666464484
transform 1 0 14260 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_2  _0630_
timestamp 1666464484
transform -1 0 13800 0 1 31552
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_2  _0631_
timestamp 1666464484
transform -1 0 10304 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0632_
timestamp 1666464484
transform -1 0 10856 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__nand3b_4  _0633_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 13984 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__xnor2_4  _0634_
timestamp 1666464484
transform -1 0 15456 0 -1 30464
box -38 -48 2062 592
use sky130_fd_sc_hd__nand2_1  _0635_
timestamp 1666464484
transform -1 0 10212 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__o221ai_4  _0636_
timestamp 1666464484
transform 1 0 11684 0 -1 29376
box -38 -48 1970 592
use sky130_fd_sc_hd__nand2_1  _0637_
timestamp 1666464484
transform -1 0 9568 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0638_
timestamp 1666464484
transform 1 0 15548 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0639_
timestamp 1666464484
transform 1 0 16836 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0640_
timestamp 1666464484
transform -1 0 17112 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0641_
timestamp 1666464484
transform -1 0 18308 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0642_
timestamp 1666464484
transform 1 0 16836 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_1  _0643_
timestamp 1666464484
transform 1 0 10396 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_4  _0644_
timestamp 1666464484
transform 1 0 9936 0 -1 31552
box -38 -48 1326 592
use sky130_fd_sc_hd__o211ai_4  _0645_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 12512 0 1 28288
box -38 -48 1602 592
use sky130_fd_sc_hd__a21o_1  _0646_
timestamp 1666464484
transform 1 0 9384 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _0647_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 10672 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_2  _0648_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 9568 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _0649_
timestamp 1666464484
transform 1 0 7912 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0650_
timestamp 1666464484
transform 1 0 9108 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0651_
timestamp 1666464484
transform -1 0 8280 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0652_
timestamp 1666464484
transform 1 0 12880 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__nand4_4  _0653_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 11868 0 -1 28288
box -38 -48 1602 592
use sky130_fd_sc_hd__and3_1  _0654_
timestamp 1666464484
transform -1 0 13708 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0655_
timestamp 1666464484
transform -1 0 17296 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0656_
timestamp 1666464484
transform -1 0 16008 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0657_
timestamp 1666464484
transform -1 0 14444 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0658_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 16376 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0659_
timestamp 1666464484
transform -1 0 15640 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0660_
timestamp 1666464484
transform -1 0 16376 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0661_
timestamp 1666464484
transform -1 0 16192 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_2  _0662_
timestamp 1666464484
transform 1 0 14812 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _0663_
timestamp 1666464484
transform 1 0 11684 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_2  _0664_
timestamp 1666464484
transform 1 0 11132 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0665_
timestamp 1666464484
transform -1 0 8648 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0666_
timestamp 1666464484
transform 1 0 8924 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0667_
timestamp 1666464484
transform 1 0 9292 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__a31o_1  _0668_
timestamp 1666464484
transform -1 0 9292 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_4  _0669_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 10212 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__and2b_1  _0670_
timestamp 1666464484
transform 1 0 9108 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _0671_
timestamp 1666464484
transform -1 0 8556 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _0672_
timestamp 1666464484
transform -1 0 9568 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__or2_4  _0673_
timestamp 1666464484
transform 1 0 14076 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__or2_4  _0674_
timestamp 1666464484
transform -1 0 16376 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0675_
timestamp 1666464484
transform -1 0 10764 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0676_
timestamp 1666464484
transform -1 0 10028 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__nand2b_4  _0677_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 15364 0 -1 13056
box -38 -48 1050 592
use sky130_fd_sc_hd__nor2_4  _0678_
timestamp 1666464484
transform -1 0 16744 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__nand2b_4  _0679_
timestamp 1666464484
transform -1 0 16652 0 1 13056
box -38 -48 1050 592
use sky130_fd_sc_hd__or2_4  _0680_
timestamp 1666464484
transform 1 0 17756 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_2  _0681_
timestamp 1666464484
transform -1 0 32568 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0682_
timestamp 1666464484
transform 1 0 31832 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0683_
timestamp 1666464484
transform -1 0 32660 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0684_
timestamp 1666464484
transform 1 0 32292 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__and4_2  _0685_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 29716 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0686_
timestamp 1666464484
transform -1 0 29256 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_2  _0687_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 31096 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_2  _0688_
timestamp 1666464484
transform 1 0 32292 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a22oi_2  _0689_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 31924 0 1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__and4_1  _0690_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 32292 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0691_
timestamp 1666464484
transform -1 0 33212 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__or3_4  _0692_
timestamp 1666464484
transform -1 0 33120 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _0693_
timestamp 1666464484
transform -1 0 31832 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_2  _0694_
timestamp 1666464484
transform -1 0 32660 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_2  _0695_
timestamp 1666464484
transform -1 0 31648 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__nand2b_1  _0696_
timestamp 1666464484
transform -1 0 31740 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0697_
timestamp 1666464484
transform 1 0 31464 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _0698_
timestamp 1666464484
transform 1 0 31096 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _0699_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 32568 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0700_
timestamp 1666464484
transform 1 0 31464 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0701_
timestamp 1666464484
transform -1 0 33396 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0702_
timestamp 1666464484
transform -1 0 33672 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _0703_
timestamp 1666464484
transform -1 0 33212 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _0704_
timestamp 1666464484
transform 1 0 33120 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__a2bb2o_2  _0705_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 32292 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_2  _0706_
timestamp 1666464484
transform -1 0 32200 0 1 22848
box -38 -48 1234 592
use sky130_fd_sc_hd__nor2_1  _0707_
timestamp 1666464484
transform 1 0 33580 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__or2_4  _0708_
timestamp 1666464484
transform 1 0 33488 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_2  _0709_
timestamp 1666464484
transform -1 0 30176 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__a22oi_4  _0710_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 28520 0 -1 19584
box -38 -48 1602 592
use sky130_fd_sc_hd__o21ba_1  _0711_
timestamp 1666464484
transform 1 0 28336 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _0712_
timestamp 1666464484
transform -1 0 32016 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _0713_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 32384 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__o22a_4  _0714_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 27968 0 1 18496
box -38 -48 1326 592
use sky130_fd_sc_hd__xor2_1  _0715_
timestamp 1666464484
transform -1 0 28428 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a22oi_1  _0716_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 31188 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0717_
timestamp 1666464484
transform 1 0 29716 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0718_
timestamp 1666464484
transform -1 0 31188 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0719_
timestamp 1666464484
transform 1 0 28796 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__or2_4  _0720_
timestamp 1666464484
transform -1 0 27600 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_4  _0721_
timestamp 1666464484
transform -1 0 29348 0 -1 22848
box -38 -48 2062 592
use sky130_fd_sc_hd__nor2_1  _0722_
timestamp 1666464484
transform -1 0 26312 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__o21bai_2  _0723_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 27508 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0724_
timestamp 1666464484
transform 1 0 28704 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _0725_
timestamp 1666464484
transform 1 0 30820 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0726_
timestamp 1666464484
transform -1 0 30636 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0727_
timestamp 1666464484
transform -1 0 27508 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__nand2b_4  _0728_
timestamp 1666464484
transform 1 0 14536 0 1 11968
box -38 -48 1050 592
use sky130_fd_sc_hd__nor2_4  _0729_
timestamp 1666464484
transform 1 0 17756 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__nand2b_4  _0730_
timestamp 1666464484
transform 1 0 15916 0 1 11968
box -38 -48 1050 592
use sky130_fd_sc_hd__nor2_4  _0731_
timestamp 1666464484
transform 1 0 17664 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__or2_4  _0732_
timestamp 1666464484
transform 1 0 15732 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_4  _0733_
timestamp 1666464484
transform 1 0 17756 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _0734_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 30360 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_4  _0735_
timestamp 1666464484
transform 1 0 17572 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_2  _0736_
timestamp 1666464484
transform 1 0 16928 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _0737_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 25668 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_4  _0738_
timestamp 1666464484
transform 1 0 17480 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_2  _0739_
timestamp 1666464484
transform -1 0 17204 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_4  _0740_
timestamp 1666464484
transform 1 0 17848 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_2  _0741_
timestamp 1666464484
transform 1 0 16836 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0742_
timestamp 1666464484
transform -1 0 22080 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0743_
timestamp 1666464484
transform 1 0 20608 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_2  _0744_
timestamp 1666464484
transform 1 0 17388 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_4  _0745_
timestamp 1666464484
transform 1 0 16836 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _0746_
timestamp 1666464484
transform 1 0 20424 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__or2_4  _0747_
timestamp 1666464484
transform 1 0 16836 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0748_
timestamp 1666464484
transform 1 0 23552 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0749_
timestamp 1666464484
transform -1 0 25484 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__a41o_1  _0750_
timestamp 1666464484
transform 1 0 24564 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _0751_
timestamp 1666464484
transform 1 0 25300 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _0752_
timestamp 1666464484
transform 1 0 25852 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_1  _0753_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 19596 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _0754_
timestamp 1666464484
transform -1 0 14720 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_4  _0755_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 12788 0 -1 20672
box -38 -48 1326 592
use sky130_fd_sc_hd__nor2_1  _0756_
timestamp 1666464484
transform 1 0 3220 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_2  _0757_
timestamp 1666464484
transform -1 0 3496 0 1 19584
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_1  _0758_
timestamp 1666464484
transform 1 0 1656 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0759_
timestamp 1666464484
transform -1 0 12880 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _0760_
timestamp 1666464484
transform 1 0 12052 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__a22oi_1  _0761_
timestamp 1666464484
transform 1 0 13064 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _0762_
timestamp 1666464484
transform 1 0 12052 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _0763_
timestamp 1666464484
transform -1 0 30360 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0764_
timestamp 1666464484
transform -1 0 28428 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _0765_
timestamp 1666464484
transform -1 0 28888 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0766_
timestamp 1666464484
transform 1 0 27140 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0767_
timestamp 1666464484
transform -1 0 28980 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0768_
timestamp 1666464484
transform 1 0 18216 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0769_
timestamp 1666464484
transform 1 0 19412 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _0770_
timestamp 1666464484
transform -1 0 25300 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0771_
timestamp 1666464484
transform 1 0 25024 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _0772_
timestamp 1666464484
transform -1 0 28060 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__or3_2  _0773_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 28060 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _0774_
timestamp 1666464484
transform 1 0 14260 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_4  _0775_
timestamp 1666464484
transform 1 0 12236 0 -1 23936
box -38 -48 1326 592
use sky130_fd_sc_hd__inv_2  _0776_
timestamp 1666464484
transform -1 0 3496 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_4  _0777_
timestamp 1666464484
transform 1 0 2668 0 -1 23936
box -38 -48 2062 592
use sky130_fd_sc_hd__nand2_2  _0778_
timestamp 1666464484
transform -1 0 3496 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0779_
timestamp 1666464484
transform -1 0 4048 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _0780_
timestamp 1666464484
transform -1 0 15732 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a41o_1  _0781_
timestamp 1666464484
transform -1 0 15548 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0782_
timestamp 1666464484
transform -1 0 17664 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _0783_
timestamp 1666464484
transform -1 0 16652 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _0784_
timestamp 1666464484
transform -1 0 27784 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0785_
timestamp 1666464484
transform -1 0 29624 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0786_
timestamp 1666464484
transform 1 0 20424 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0787_
timestamp 1666464484
transform -1 0 23000 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0788_
timestamp 1666464484
transform 1 0 27232 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _0789_
timestamp 1666464484
transform 1 0 22172 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _0790_
timestamp 1666464484
transform 1 0 27968 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0791_
timestamp 1666464484
transform 1 0 21988 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_1  _0792_
timestamp 1666464484
transform 1 0 24564 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _0793_
timestamp 1666464484
transform -1 0 23460 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0794_
timestamp 1666464484
transform 1 0 15180 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _0795_
timestamp 1666464484
transform -1 0 14812 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0796_
timestamp 1666464484
transform 1 0 11960 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__o311a_4  _0797_
timestamp 1666464484
transform 1 0 12420 0 -1 22848
box -38 -48 1602 592
use sky130_fd_sc_hd__inv_2  _0798_
timestamp 1666464484
transform -1 0 9384 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_4  _0799_
timestamp 1666464484
transform -1 0 8648 0 1 23936
box -38 -48 2062 592
use sky130_fd_sc_hd__and2_2  _0800_
timestamp 1666464484
transform -1 0 9476 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0801_
timestamp 1666464484
transform -1 0 6992 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _0802_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 18768 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_2  _0803_
timestamp 1666464484
transform 1 0 17756 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0804_
timestamp 1666464484
transform 1 0 21988 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _0805_
timestamp 1666464484
transform 1 0 28244 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_4  _0806_
timestamp 1666464484
transform -1 0 27876 0 1 21760
box -38 -48 1234 592
use sky130_fd_sc_hd__a32o_1  _0807_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 27968 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _0808_
timestamp 1666464484
transform -1 0 28612 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0809_
timestamp 1666464484
transform 1 0 19412 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0810_
timestamp 1666464484
transform 1 0 19964 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _0811_
timestamp 1666464484
transform 1 0 20424 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0812_
timestamp 1666464484
transform 1 0 20424 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _0813_
timestamp 1666464484
transform 1 0 19872 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__o31ai_4  _0814_
timestamp 1666464484
transform -1 0 20976 0 -1 21760
box -38 -48 1602 592
use sky130_fd_sc_hd__nand2_1  _0815_
timestamp 1666464484
transform 1 0 11684 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_2  _0816_
timestamp 1666464484
transform 1 0 12512 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0817_
timestamp 1666464484
transform -1 0 11960 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0818_
timestamp 1666464484
transform -1 0 10396 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0819_
timestamp 1666464484
transform 1 0 10212 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_2  _0820_
timestamp 1666464484
transform 1 0 10396 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0821_
timestamp 1666464484
transform 1 0 8004 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0822_
timestamp 1666464484
transform 1 0 9108 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_1  _0823_
timestamp 1666464484
transform 1 0 8280 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _0824_
timestamp 1666464484
transform -1 0 8096 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _0825_
timestamp 1666464484
transform 1 0 5520 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0826_
timestamp 1666464484
transform 1 0 6348 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _0827_
timestamp 1666464484
transform -1 0 7452 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _0828_
timestamp 1666464484
transform -1 0 7912 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_2  _0829_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 6808 0 -1 25024
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_2  _0830_
timestamp 1666464484
transform 1 0 9844 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_2  _0831_
timestamp 1666464484
transform 1 0 4416 0 -1 25024
box -38 -48 1234 592
use sky130_fd_sc_hd__a21oi_2  _0832_
timestamp 1666464484
transform 1 0 4140 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _0833_
timestamp 1666464484
transform -1 0 4692 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _0834_
timestamp 1666464484
transform 1 0 2852 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_4  _0835_
timestamp 1666464484
transform -1 0 7636 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__clkinv_2  _0836_
timestamp 1666464484
transform 1 0 6992 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0837_
timestamp 1666464484
transform 1 0 3128 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _0838_
timestamp 1666464484
transform -1 0 7728 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0839_
timestamp 1666464484
transform -1 0 7176 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0840_
timestamp 1666464484
transform 1 0 9016 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _0841_
timestamp 1666464484
transform -1 0 10856 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a41o_1  _0842_
timestamp 1666464484
transform 1 0 7636 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _0843_
timestamp 1666464484
transform 1 0 7176 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0844_
timestamp 1666464484
transform -1 0 8648 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0845_
timestamp 1666464484
transform 1 0 9108 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0846_
timestamp 1666464484
transform -1 0 8556 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _0847_
timestamp 1666464484
transform 1 0 6900 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _0848_
timestamp 1666464484
transform 1 0 5060 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _0849_
timestamp 1666464484
transform -1 0 4324 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _0850_
timestamp 1666464484
transform 1 0 5060 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0851_
timestamp 1666464484
transform -1 0 2668 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__a2bb2o_1  _0852_
timestamp 1666464484
transform -1 0 4692 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _0853_
timestamp 1666464484
transform 1 0 4600 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__a311o_1  _0854_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 3956 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__o31a_1  _0855_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 3588 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_1  _0856_
timestamp 1666464484
transform 1 0 2944 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _0857_
timestamp 1666464484
transform -1 0 5520 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _0858_
timestamp 1666464484
transform -1 0 3496 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _0859_
timestamp 1666464484
transform 1 0 3956 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0860_
timestamp 1666464484
transform 1 0 3956 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__and3_2  _0861_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 6532 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__and2_2  _0862_
timestamp 1666464484
transform 1 0 3956 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__and3_2  _0863_
timestamp 1666464484
transform 1 0 3956 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _0864_
timestamp 1666464484
transform 1 0 6992 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_2  _0865_
timestamp 1666464484
transform -1 0 8648 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_4  _0866_
timestamp 1666464484
transform 1 0 10120 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_4  _0867_
timestamp 1666464484
transform 1 0 8648 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_2  _0868_
timestamp 1666464484
transform 1 0 9108 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _0869_
timestamp 1666464484
transform -1 0 3496 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_2  _0870_
timestamp 1666464484
transform -1 0 3496 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_2  _0871_
timestamp 1666464484
transform 1 0 20424 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__and3_2  _0872_
timestamp 1666464484
transform 1 0 29348 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__and3_2  _0873_
timestamp 1666464484
transform 1 0 19412 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__and3_2  _0874_
timestamp 1666464484
transform 1 0 23552 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__and3_2  _0875_
timestamp 1666464484
transform 1 0 28704 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_2  _0876_
timestamp 1666464484
transform 1 0 21988 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _0877_
timestamp 1666464484
transform 1 0 19412 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__and3_2  _0878_
timestamp 1666464484
transform 1 0 28612 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_2  _0879_
timestamp 1666464484
transform 1 0 20516 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__and3_2  _0880_
timestamp 1666464484
transform 1 0 22724 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__and3_2  _0881_
timestamp 1666464484
transform 1 0 25668 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__and3_2  _0882_
timestamp 1666464484
transform -1 0 16008 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__and3_2  _0883_
timestamp 1666464484
transform 1 0 28060 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__and3_2  _0884_
timestamp 1666464484
transform 1 0 18400 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__and3_2  _0885_
timestamp 1666464484
transform -1 0 17388 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__and3_2  _0886_
timestamp 1666464484
transform 1 0 18400 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0887_
timestamp 1666464484
transform -1 0 15548 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0888_
timestamp 1666464484
transform 1 0 25576 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_2  _0889_
timestamp 1666464484
transform 1 0 13340 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0890_
timestamp 1666464484
transform 1 0 25484 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_2  _0891_
timestamp 1666464484
transform 1 0 11960 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0892_
timestamp 1666464484
transform 1 0 28336 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_2  _0893_
timestamp 1666464484
transform 1 0 15640 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0894_
timestamp 1666464484
transform 1 0 24564 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0895_
timestamp 1666464484
transform 1 0 29716 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0896_
timestamp 1666464484
transform -1 0 24104 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0897_
timestamp 1666464484
transform 1 0 17296 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0898_
timestamp 1666464484
transform 1 0 17296 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0899_
timestamp 1666464484
transform 1 0 17388 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0900_
timestamp 1666464484
transform 1 0 16836 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0901_
timestamp 1666464484
transform -1 0 29256 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0902_
timestamp 1666464484
transform 1 0 30452 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0903_
timestamp 1666464484
transform -1 0 29256 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0904_
timestamp 1666464484
transform 1 0 29716 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0905_
timestamp 1666464484
transform 1 0 22448 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0906_
timestamp 1666464484
transform 1 0 21988 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0907_
timestamp 1666464484
transform 1 0 20424 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0908_
timestamp 1666464484
transform 1 0 21988 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0909_
timestamp 1666464484
transform -1 0 31740 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0910_
timestamp 1666464484
transform 1 0 32292 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0911_
timestamp 1666464484
transform -1 0 31832 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0912_
timestamp 1666464484
transform -1 0 33948 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0913_
timestamp 1666464484
transform -1 0 14904 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0914_
timestamp 1666464484
transform 1 0 15824 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0915_
timestamp 1666464484
transform 1 0 16836 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0916_
timestamp 1666464484
transform 1 0 15180 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0917_
timestamp 1666464484
transform 1 0 19412 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0918_
timestamp 1666464484
transform 1 0 20516 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0919_
timestamp 1666464484
transform 1 0 19412 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0920_
timestamp 1666464484
transform -1 0 22540 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0921_
timestamp 1666464484
transform -1 0 26036 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _0922_
timestamp 1666464484
transform 1 0 24564 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _0923_
timestamp 1666464484
transform -1 0 26680 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _0924_
timestamp 1666464484
transform -1 0 28336 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0925_
timestamp 1666464484
transform 1 0 20424 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0926_
timestamp 1666464484
transform -1 0 21620 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0927_
timestamp 1666464484
transform 1 0 22908 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0928_
timestamp 1666464484
transform 1 0 21988 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0929_
timestamp 1666464484
transform 1 0 25944 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0930_
timestamp 1666464484
transform -1 0 28796 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0931_
timestamp 1666464484
transform 1 0 23184 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0932_
timestamp 1666464484
transform -1 0 25116 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0933_
timestamp 1666464484
transform -1 0 30176 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0934_
timestamp 1666464484
transform 1 0 32292 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0935_
timestamp 1666464484
transform -1 0 33948 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0936_
timestamp 1666464484
transform -1 0 31832 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0937_
timestamp 1666464484
transform 1 0 23552 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0938_
timestamp 1666464484
transform 1 0 24564 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0939_
timestamp 1666464484
transform 1 0 23552 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0940_
timestamp 1666464484
transform 1 0 24564 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0941_
timestamp 1666464484
transform 1 0 17664 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0942_
timestamp 1666464484
transform -1 0 16192 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0943_
timestamp 1666464484
transform -1 0 16468 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0944_
timestamp 1666464484
transform 1 0 18400 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0945_
timestamp 1666464484
transform 1 0 29900 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0946_
timestamp 1666464484
transform -1 0 29256 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0947_
timestamp 1666464484
transform 1 0 30452 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0948_
timestamp 1666464484
transform -1 0 32844 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0949_
timestamp 1666464484
transform -1 0 21528 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0950_
timestamp 1666464484
transform 1 0 23184 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0951_
timestamp 1666464484
transform 1 0 20976 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0952_
timestamp 1666464484
transform -1 0 21252 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0953_
timestamp 1666464484
transform -1 0 25116 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0954_
timestamp 1666464484
transform 1 0 23552 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _0955_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 3588 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_2  _0956_
timestamp 1666464484
transform 1 0 3956 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _0957_
timestamp 1666464484
transform -1 0 3220 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0958_
timestamp 1666464484
transform -1 0 2760 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _0959_
timestamp 1666464484
transform -1 0 12144 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _0960_
timestamp 1666464484
transform 1 0 9292 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _0961_
timestamp 1666464484
transform 1 0 12144 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _0962_
timestamp 1666464484
transform -1 0 12604 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _0963_
timestamp 1666464484
transform 1 0 3036 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _0964_
timestamp 1666464484
transform 1 0 7820 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _0965_
timestamp 1666464484
transform -1 0 10856 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _0966_
timestamp 1666464484
transform 1 0 9844 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _0967_
timestamp 1666464484
transform 1 0 6992 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _0968_
timestamp 1666464484
transform 1 0 10028 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _0969_
timestamp 1666464484
transform 1 0 14260 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _0970_
timestamp 1666464484
transform 1 0 12696 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _0971_
timestamp 1666464484
transform 1 0 8188 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _0972_
timestamp 1666464484
transform -1 0 4416 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _0973_
timestamp 1666464484
transform -1 0 5612 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0974__2
timestamp 1666464484
transform 1 0 15180 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0975__3
timestamp 1666464484
transform -1 0 15272 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0976__4
timestamp 1666464484
transform -1 0 17112 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0977__5
timestamp 1666464484
transform 1 0 17388 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0978__6
timestamp 1666464484
transform -1 0 19872 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0979__7
timestamp 1666464484
transform -1 0 21712 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0980__8
timestamp 1666464484
transform -1 0 22356 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0981_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 24564 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0982_
timestamp 1666464484
transform 1 0 24564 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0983_
timestamp 1666464484
transform 1 0 27324 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0984_
timestamp 1666464484
transform 1 0 23828 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0985_
timestamp 1666464484
transform 1 0 27324 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0986_
timestamp 1666464484
transform 1 0 24564 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0987_
timestamp 1666464484
transform 1 0 15548 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0988_
timestamp 1666464484
transform 1 0 16836 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0989_
timestamp 1666464484
transform -1 0 16376 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0990_
timestamp 1666464484
transform 1 0 14996 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0991_
timestamp 1666464484
transform -1 0 29900 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0992_
timestamp 1666464484
transform -1 0 29256 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0993_
timestamp 1666464484
transform 1 0 30084 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0994_
timestamp 1666464484
transform 1 0 28612 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0995_
timestamp 1666464484
transform 1 0 21252 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0996_
timestamp 1666464484
transform 1 0 19504 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0997_
timestamp 1666464484
transform 1 0 19412 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0998_
timestamp 1666464484
transform 1 0 19872 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0999_
timestamp 1666464484
transform -1 0 32936 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1000_
timestamp 1666464484
transform 1 0 32292 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1001_
timestamp 1666464484
transform 1 0 32292 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1002_
timestamp 1666464484
transform -1 0 33764 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1003_
timestamp 1666464484
transform 1 0 14904 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1004_
timestamp 1666464484
transform 1 0 15272 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1005_
timestamp 1666464484
transform 1 0 14904 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1006_
timestamp 1666464484
transform 1 0 15180 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfstp_4  _1007_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 3956 0 1 5440
box -38 -48 2246 592
use sky130_fd_sc_hd__dfrtp_2  _1008_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 3496 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1009_
timestamp 1666464484
transform 1 0 1656 0 -1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1010_
timestamp 1666464484
transform -1 0 12144 0 1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1011_
timestamp 1666464484
transform -1 0 12144 0 1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1012_
timestamp 1666464484
transform -1 0 13616 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1013_
timestamp 1666464484
transform -1 0 13156 0 1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1014_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 2116 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfxtp_1  _1015_
timestamp 1666464484
transform 1 0 7084 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1016_
timestamp 1666464484
transform 1 0 11684 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1017_
timestamp 1666464484
transform 1 0 10764 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1018_
timestamp 1666464484
transform 1 0 5336 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1019_
timestamp 1666464484
transform 1 0 7176 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1020_
timestamp 1666464484
transform 1 0 11684 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1021_
timestamp 1666464484
transform 1 0 11684 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1022_
timestamp 1666464484
transform 1 0 5428 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1023_
timestamp 1666464484
transform 1 0 7176 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1024_
timestamp 1666464484
transform 1 0 11224 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1025_
timestamp 1666464484
transform 1 0 10304 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1026_
timestamp 1666464484
transform 1 0 5520 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfrtp_1  _1027_
timestamp 1666464484
transform 1 0 6992 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1028_
timestamp 1666464484
transform 1 0 9108 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1029_
timestamp 1666464484
transform 1 0 8924 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1030_
timestamp 1666464484
transform 1 0 6532 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1031_
timestamp 1666464484
transform 1 0 9108 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1032_
timestamp 1666464484
transform 1 0 11776 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1033_
timestamp 1666464484
transform 1 0 11776 0 -1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1034_
timestamp 1666464484
transform -1 0 9844 0 -1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dfxtp_4  _1035_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 4048 0 -1 25024
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _1036_
timestamp 1666464484
transform 1 0 6808 0 -1 23936
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_2  _1037_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 7084 0 -1 19584
box -38 -48 1602 592
use sky130_fd_sc_hd__dfrtp_1  _1038_
timestamp 1666464484
transform 1 0 2668 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfxtp_4  _1039_
timestamp 1666464484
transform 1 0 2484 0 -1 19584
box -38 -48 1786 592
use sky130_fd_sc_hd__dfrtp_2  _1040_
timestamp 1666464484
transform 1 0 4140 0 -1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__dfxtp_1  _1041_
timestamp 1666464484
transform 1 0 12328 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1042_
timestamp 1666464484
transform -1 0 15732 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1043_
timestamp 1666464484
transform 1 0 14904 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1044_
timestamp 1666464484
transform 1 0 16652 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1045_
timestamp 1666464484
transform 1 0 17664 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1046_
timestamp 1666464484
transform 1 0 19504 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1047_
timestamp 1666464484
transform -1 0 21528 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1048_
timestamp 1666464484
transform 1 0 21988 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1049_
timestamp 1666464484
transform 1 0 18860 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1050_
timestamp 1666464484
transform 1 0 19412 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1051_
timestamp 1666464484
transform 1 0 18676 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1052_
timestamp 1666464484
transform 1 0 19412 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1053_
timestamp 1666464484
transform -1 0 25760 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1054_
timestamp 1666464484
transform 1 0 24564 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1055_
timestamp 1666464484
transform 1 0 25852 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1056_
timestamp 1666464484
transform -1 0 28612 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1057_
timestamp 1666464484
transform 1 0 19688 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1058_
timestamp 1666464484
transform 1 0 21988 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1059_
timestamp 1666464484
transform 1 0 20700 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1060_
timestamp 1666464484
transform 1 0 19596 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1061_
timestamp 1666464484
transform 1 0 24564 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1062_
timestamp 1666464484
transform 1 0 26404 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1063_
timestamp 1666464484
transform 1 0 24564 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1064_
timestamp 1666464484
transform -1 0 25392 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_4  _1065_
timestamp 1666464484
transform -1 0 31464 0 1 14144
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _1066_
timestamp 1666464484
transform 1 0 31832 0 1 14144
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_2  _1067_
timestamp 1666464484
transform 1 0 32292 0 -1 16320
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_4  _1068_
timestamp 1666464484
transform 1 0 32292 0 -1 14144
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _1069_
timestamp 1666464484
transform 1 0 23184 0 -1 18496
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_2  _1070_
timestamp 1666464484
transform 1 0 23092 0 -1 17408
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_4  _1071_
timestamp 1666464484
transform 1 0 23184 0 -1 21760
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _1072_
timestamp 1666464484
transform 1 0 23092 0 -1 19584
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_1  _1073_
timestamp 1666464484
transform 1 0 17296 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1074_
timestamp 1666464484
transform -1 0 18032 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1075_
timestamp 1666464484
transform -1 0 18308 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_4  _1076_
timestamp 1666464484
transform 1 0 17848 0 -1 25024
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _1077_
timestamp 1666464484
transform 1 0 29716 0 -1 27200
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_1  _1078_
timestamp 1666464484
transform 1 0 29716 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1079_
timestamp 1666464484
transform 1 0 30084 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1080_
timestamp 1666464484
transform 1 0 30084 0 1 25024
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_4  _1081_
timestamp 1666464484
transform 1 0 21988 0 -1 25024
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_1  _1082_
timestamp 1666464484
transform 1 0 21344 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1083_
timestamp 1666464484
transform -1 0 21252 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_4  _1084_
timestamp 1666464484
transform 1 0 21988 0 -1 26112
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_1  _1085_
timestamp 1666464484
transform -1 0 25116 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1086_
timestamp 1666464484
transform -1 0 25024 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_CIRCUIT_1957.int_memory_1.GATES_21.result $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 32292 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_CIRCUIT_1957.int_memory_1.GATES_22.result
timestamp 1666464484
transform 1 0 20608 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_CIRCUIT_1957.int_memory_1.GATES_23.result
timestamp 1666464484
transform 1 0 25208 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_CIRCUIT_1957.int_memory_1.GATES_24.result
timestamp 1666464484
transform 1 0 32292 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_CIRCUIT_1957.int_memory_1.GATES_25.result
timestamp 1666464484
transform 1 0 23184 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_CIRCUIT_1957.int_memory_1.GATES_26.result
timestamp 1666464484
transform -1 0 19688 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_CIRCUIT_1957.int_memory_1.GATES_27.result
timestamp 1666464484
transform 1 0 29992 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_CIRCUIT_1957.int_memory_1.GATES_28.result
timestamp 1666464484
transform 1 0 21620 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_CIRCUIT_1957.int_memory_1.GATES_29.result
timestamp 1666464484
transform 1 0 24564 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_CIRCUIT_1957.int_memory_1.GATES_30.result
timestamp 1666464484
transform 1 0 26036 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_CIRCUIT_1957.int_memory_1.GATES_31.result
timestamp 1666464484
transform 1 0 16192 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_CIRCUIT_1957.int_memory_1.GATES_32.result
timestamp 1666464484
transform 1 0 29716 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_CIRCUIT_1957.int_memory_1.GATES_33.result
timestamp 1666464484
transform 1 0 21620 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_CIRCUIT_1957.int_memory_1.GATES_50.result
timestamp 1666464484
transform -1 0 17020 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_CIRCUIT_1957.int_memory_1.GATES_53.result
timestamp 1666464484
transform 1 0 19412 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0__0460_
timestamp 1666464484
transform 1 0 20608 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk
timestamp 1666464484
transform 1 0 15548 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_CIRCUIT_1957.int_memory_1.GATES_21.result
timestamp 1666464484
transform -1 0 33764 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_CIRCUIT_1957.int_memory_1.GATES_22.result
timestamp 1666464484
transform 1 0 18216 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_CIRCUIT_1957.int_memory_1.GATES_23.result
timestamp 1666464484
transform 1 0 26036 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_CIRCUIT_1957.int_memory_1.GATES_24.result
timestamp 1666464484
transform -1 0 33028 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_CIRCUIT_1957.int_memory_1.GATES_25.result
timestamp 1666464484
transform 1 0 20792 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_CIRCUIT_1957.int_memory_1.GATES_26.result
timestamp 1666464484
transform -1 0 17480 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_CIRCUIT_1957.int_memory_1.GATES_27.result
timestamp 1666464484
transform 1 0 28612 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_CIRCUIT_1957.int_memory_1.GATES_28.result
timestamp 1666464484
transform -1 0 22632 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_CIRCUIT_1957.int_memory_1.GATES_29.result
timestamp 1666464484
transform 1 0 23368 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_CIRCUIT_1957.int_memory_1.GATES_30.result
timestamp 1666464484
transform -1 0 22632 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_CIRCUIT_1957.int_memory_1.GATES_31.result
timestamp 1666464484
transform -1 0 14812 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_CIRCUIT_1957.int_memory_1.GATES_32.result
timestamp 1666464484
transform -1 0 30452 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_CIRCUIT_1957.int_memory_1.GATES_33.result
timestamp 1666464484
transform 1 0 18216 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_CIRCUIT_1957.int_memory_1.GATES_50.result
timestamp 1666464484
transform 1 0 12972 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_CIRCUIT_1957.int_memory_1.GATES_53.result
timestamp 1666464484
transform -1 0 20056 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f__0460_
timestamp 1666464484
transform -1 0 20056 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_CIRCUIT_1957.int_memory_1.GATES_21.result
timestamp 1666464484
transform -1 0 33028 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_CIRCUIT_1957.int_memory_1.GATES_22.result
timestamp 1666464484
transform 1 0 18216 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_CIRCUIT_1957.int_memory_1.GATES_23.result
timestamp 1666464484
transform -1 0 25208 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_CIRCUIT_1957.int_memory_1.GATES_24.result
timestamp 1666464484
transform -1 0 33028 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_CIRCUIT_1957.int_memory_1.GATES_25.result
timestamp 1666464484
transform 1 0 20792 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_CIRCUIT_1957.int_memory_1.GATES_26.result
timestamp 1666464484
transform 1 0 18216 0 -1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_CIRCUIT_1957.int_memory_1.GATES_27.result
timestamp 1666464484
transform 1 0 28612 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_CIRCUIT_1957.int_memory_1.GATES_28.result
timestamp 1666464484
transform -1 0 22632 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_CIRCUIT_1957.int_memory_1.GATES_29.result
timestamp 1666464484
transform 1 0 23368 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_CIRCUIT_1957.int_memory_1.GATES_30.result
timestamp 1666464484
transform 1 0 26036 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_CIRCUIT_1957.int_memory_1.GATES_31.result
timestamp 1666464484
transform 1 0 18216 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_CIRCUIT_1957.int_memory_1.GATES_32.result
timestamp 1666464484
transform -1 0 30452 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_CIRCUIT_1957.int_memory_1.GATES_33.result
timestamp 1666464484
transform 1 0 18216 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_CIRCUIT_1957.int_memory_1.GATES_50.result
timestamp 1666464484
transform 1 0 12972 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_CIRCUIT_1957.int_memory_1.GATES_53.result
timestamp 1666464484
transform -1 0 20056 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f__0460_
timestamp 1666464484
transform 1 0 20792 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_0__f_clk
timestamp 1666464484
transform -1 0 9660 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_1__f_clk
timestamp 1666464484
transform -1 0 9660 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_2__f_clk
timestamp 1666464484
transform 1 0 19412 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_3__f_clk
timestamp 1666464484
transform 1 0 20792 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__buf_6  fanout28 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 21988 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  fanout29
timestamp 1666464484
transform -1 0 15088 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  fanout30
timestamp 1666464484
transform 1 0 21988 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  fanout31 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 27508 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout32
timestamp 1666464484
transform 1 0 24564 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  fanout33
timestamp 1666464484
transform -1 0 22816 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  fanout34
timestamp 1666464484
transform 1 0 17112 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  fanout35 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 16836 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  fanout36
timestamp 1666464484
transform -1 0 16376 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  fanout37
timestamp 1666464484
transform 1 0 20700 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  fanout38
timestamp 1666464484
transform -1 0 18124 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  fanout39
timestamp 1666464484
transform 1 0 21988 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  fanout40
timestamp 1666464484
transform 1 0 16100 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  fanout41
timestamp 1666464484
transform 1 0 18400 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout42
timestamp 1666464484
transform 1 0 20424 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  fanout43
timestamp 1666464484
transform -1 0 15272 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  fanout44
timestamp 1666464484
transform 1 0 14260 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout45 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 20516 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  fanout46
timestamp 1666464484
transform -1 0 12788 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout47
timestamp 1666464484
transform -1 0 20332 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout48
timestamp 1666464484
transform -1 0 29808 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout49
timestamp 1666464484
transform -1 0 25300 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout50
timestamp 1666464484
transform -1 0 30084 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  fanout51
timestamp 1666464484
transform 1 0 26404 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout52
timestamp 1666464484
transform 1 0 13340 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_8  fanout53 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 11224 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_6  fanout54
timestamp 1666464484
transform -1 0 4784 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__buf_8  fanout55
timestamp 1666464484
transform 1 0 10120 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_8  fanout56 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 12512 0 1 22848
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_2  input1
timestamp 1666464484
transform 1 0 7728 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input2
timestamp 1666464484
transform 1 0 10672 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input3
timestamp 1666464484
transform -1 0 14628 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input4
timestamp 1666464484
transform -1 0 17204 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input5
timestamp 1666464484
transform -1 0 19872 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input6
timestamp 1666464484
transform -1 0 22816 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input7
timestamp 1666464484
transform -1 0 25760 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input8
timestamp 1666464484
transform -1 0 28704 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input9
timestamp 1666464484
transform -1 0 31648 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input10
timestamp 1666464484
transform -1 0 34408 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input11
timestamp 1666464484
transform 1 0 4784 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  output12
timestamp 1666464484
transform -1 0 2116 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output13
timestamp 1666464484
transform 1 0 14260 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output14
timestamp 1666464484
transform 1 0 15456 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output15
timestamp 1666464484
transform 1 0 16836 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output16
timestamp 1666464484
transform 1 0 18032 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output17
timestamp 1666464484
transform 1 0 19412 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output18
timestamp 1666464484
transform 1 0 20608 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output19
timestamp 1666464484
transform 1 0 21988 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output20
timestamp 1666464484
transform 1 0 23184 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output21
timestamp 1666464484
transform -1 0 25116 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output22
timestamp 1666464484
transform -1 0 26312 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output23
timestamp 1666464484
transform -1 0 3128 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output24
timestamp 1666464484
transform -1 0 27692 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output25
timestamp 1666464484
transform 1 0 28336 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output26
timestamp 1666464484
transform -1 0 4508 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output27
timestamp 1666464484
transform -1 0 5704 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  tholin_avalonsemi_5401_57 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 6808 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tholin_avalonsemi_5401_58
timestamp 1666464484
transform -1 0 8004 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tholin_avalonsemi_5401_59
timestamp 1666464484
transform -1 0 9384 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tholin_avalonsemi_5401_60
timestamp 1666464484
transform -1 0 10580 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tholin_avalonsemi_5401_61
timestamp 1666464484
transform -1 0 11960 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tholin_avalonsemi_5401_62
timestamp 1666464484
transform -1 0 13156 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tholin_avalonsemi_5401_63
timestamp 1666464484
transform -1 0 29992 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tholin_avalonsemi_5401_64
timestamp 1666464484
transform -1 0 31188 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tholin_avalonsemi_5401_65
timestamp 1666464484
transform -1 0 32568 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tholin_avalonsemi_5401_66
timestamp 1666464484
transform -1 0 33764 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tholin_avalonsemi_5401_67
timestamp 1666464484
transform -1 0 34408 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tholin_avalonsemi_5401_68
timestamp 1666464484
transform -1 0 34408 0 1 2176
box -38 -48 314 592
<< labels >>
flabel metal2 s 1766 35200 1822 36000 0 FreeSans 224 90 0 0 clk
port 0 nsew signal input
flabel metal2 s 7654 35200 7710 36000 0 FreeSans 224 90 0 0 io_in[0]
port 1 nsew signal input
flabel metal2 s 10598 35200 10654 36000 0 FreeSans 224 90 0 0 io_in[1]
port 2 nsew signal input
flabel metal2 s 13542 35200 13598 36000 0 FreeSans 224 90 0 0 io_in[2]
port 3 nsew signal input
flabel metal2 s 16486 35200 16542 36000 0 FreeSans 224 90 0 0 io_in[3]
port 4 nsew signal input
flabel metal2 s 19430 35200 19486 36000 0 FreeSans 224 90 0 0 io_in[4]
port 5 nsew signal input
flabel metal2 s 22374 35200 22430 36000 0 FreeSans 224 90 0 0 io_in[5]
port 6 nsew signal input
flabel metal2 s 25318 35200 25374 36000 0 FreeSans 224 90 0 0 io_in[6]
port 7 nsew signal input
flabel metal2 s 28262 35200 28318 36000 0 FreeSans 224 90 0 0 io_in[7]
port 8 nsew signal input
flabel metal2 s 31206 35200 31262 36000 0 FreeSans 224 90 0 0 io_in[8]
port 9 nsew signal input
flabel metal2 s 34150 35200 34206 36000 0 FreeSans 224 90 0 0 io_in[9]
port 10 nsew signal input
flabel metal3 s 35200 17824 36000 17944 0 FreeSans 480 0 0 0 io_oeb
port 11 nsew signal tristate
flabel metal2 s 1214 0 1270 800 0 FreeSans 224 90 0 0 io_out[0]
port 12 nsew signal tristate
flabel metal2 s 14094 0 14150 800 0 FreeSans 224 90 0 0 io_out[10]
port 13 nsew signal tristate
flabel metal2 s 15382 0 15438 800 0 FreeSans 224 90 0 0 io_out[11]
port 14 nsew signal tristate
flabel metal2 s 16670 0 16726 800 0 FreeSans 224 90 0 0 io_out[12]
port 15 nsew signal tristate
flabel metal2 s 17958 0 18014 800 0 FreeSans 224 90 0 0 io_out[13]
port 16 nsew signal tristate
flabel metal2 s 19246 0 19302 800 0 FreeSans 224 90 0 0 io_out[14]
port 17 nsew signal tristate
flabel metal2 s 20534 0 20590 800 0 FreeSans 224 90 0 0 io_out[15]
port 18 nsew signal tristate
flabel metal2 s 21822 0 21878 800 0 FreeSans 224 90 0 0 io_out[16]
port 19 nsew signal tristate
flabel metal2 s 23110 0 23166 800 0 FreeSans 224 90 0 0 io_out[17]
port 20 nsew signal tristate
flabel metal2 s 24398 0 24454 800 0 FreeSans 224 90 0 0 io_out[18]
port 21 nsew signal tristate
flabel metal2 s 25686 0 25742 800 0 FreeSans 224 90 0 0 io_out[19]
port 22 nsew signal tristate
flabel metal2 s 2502 0 2558 800 0 FreeSans 224 90 0 0 io_out[1]
port 23 nsew signal tristate
flabel metal2 s 26974 0 27030 800 0 FreeSans 224 90 0 0 io_out[20]
port 24 nsew signal tristate
flabel metal2 s 28262 0 28318 800 0 FreeSans 224 90 0 0 io_out[21]
port 25 nsew signal tristate
flabel metal2 s 29550 0 29606 800 0 FreeSans 224 90 0 0 io_out[22]
port 26 nsew signal tristate
flabel metal2 s 30838 0 30894 800 0 FreeSans 224 90 0 0 io_out[23]
port 27 nsew signal tristate
flabel metal2 s 32126 0 32182 800 0 FreeSans 224 90 0 0 io_out[24]
port 28 nsew signal tristate
flabel metal2 s 33414 0 33470 800 0 FreeSans 224 90 0 0 io_out[25]
port 29 nsew signal tristate
flabel metal2 s 34702 0 34758 800 0 FreeSans 224 90 0 0 io_out[26]
port 30 nsew signal tristate
flabel metal2 s 3790 0 3846 800 0 FreeSans 224 90 0 0 io_out[2]
port 31 nsew signal tristate
flabel metal2 s 5078 0 5134 800 0 FreeSans 224 90 0 0 io_out[3]
port 32 nsew signal tristate
flabel metal2 s 6366 0 6422 800 0 FreeSans 224 90 0 0 io_out[4]
port 33 nsew signal tristate
flabel metal2 s 7654 0 7710 800 0 FreeSans 224 90 0 0 io_out[5]
port 34 nsew signal tristate
flabel metal2 s 8942 0 8998 800 0 FreeSans 224 90 0 0 io_out[6]
port 35 nsew signal tristate
flabel metal2 s 10230 0 10286 800 0 FreeSans 224 90 0 0 io_out[7]
port 36 nsew signal tristate
flabel metal2 s 11518 0 11574 800 0 FreeSans 224 90 0 0 io_out[8]
port 37 nsew signal tristate
flabel metal2 s 12806 0 12862 800 0 FreeSans 224 90 0 0 io_out[9]
port 38 nsew signal tristate
flabel metal2 s 4710 35200 4766 36000 0 FreeSans 224 90 0 0 rst
port 39 nsew signal input
flabel metal4 s 5164 2128 5484 33776 0 FreeSans 1920 90 0 0 vccd1
port 40 nsew power bidirectional
flabel metal4 s 13605 2128 13925 33776 0 FreeSans 1920 90 0 0 vccd1
port 40 nsew power bidirectional
flabel metal4 s 22046 2128 22366 33776 0 FreeSans 1920 90 0 0 vccd1
port 40 nsew power bidirectional
flabel metal4 s 30487 2128 30807 33776 0 FreeSans 1920 90 0 0 vccd1
port 40 nsew power bidirectional
flabel metal4 s 9384 2128 9704 33776 0 FreeSans 1920 90 0 0 vssd1
port 41 nsew ground bidirectional
flabel metal4 s 17825 2128 18145 33776 0 FreeSans 1920 90 0 0 vssd1
port 41 nsew ground bidirectional
flabel metal4 s 26266 2128 26586 33776 0 FreeSans 1920 90 0 0 vssd1
port 41 nsew ground bidirectional
flabel metal4 s 34707 2128 35027 33776 0 FreeSans 1920 90 0 0 vssd1
port 41 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 36000 36000
<< end >>
