// This is the unpowered netlist.
module tholin_avalonsemi_tbb1143 (clk,
    rst,
    io_in,
    io_out);
 input clk;
 input rst;
 input [5:0] io_in;
 output [7:0] io_out;

 wire \CIRCUIT_2223.CLK ;
 wire \CIRCUIT_2223.GATES_1.input1[0] ;
 wire \CIRCUIT_2223.GATES_1.input1[1] ;
 wire \CIRCUIT_2223.GATES_1.input1[2] ;
 wire \CIRCUIT_2223.GATES_1.input1[3] ;
 wire \CIRCUIT_2223.GATES_11.input2 ;
 wire \CIRCUIT_2223.GATES_2.input2 ;
 wire \CIRCUIT_2223.GATES_3.input2 ;
 wire \CIRCUIT_2223.GATES_4.input1[0] ;
 wire \CIRCUIT_2223.GATES_4.input1[1] ;
 wire \CIRCUIT_2223.GATES_4.input1[2] ;
 wire \CIRCUIT_2223.GATES_4.input1[3] ;
 wire \CIRCUIT_2223.GATES_5.input2 ;
 wire \CIRCUIT_2223.MEMORY_18.clock ;
 wire \CIRCUIT_2223.MEMORY_18.d ;
 wire \CIRCUIT_2223.MEMORY_18.s_currentState ;
 wire \CIRCUIT_2223.MEMORY_19.d ;
 wire \CIRCUIT_2223.MEMORY_19.s_currentState ;
 wire \CIRCUIT_2223.MEMORY_20.d ;
 wire \CIRCUIT_2223.MEMORY_20.s_currentState ;
 wire \CIRCUIT_2223.MEMORY_21.d ;
 wire \CIRCUIT_2223.MEMORY_21.s_currentState ;
 wire \CIRCUIT_2223.MEMORY_22.d ;
 wire \CIRCUIT_2223.MEMORY_22.s_currentState ;
 wire \CIRCUIT_2223.MEMORY_23.s_currentState ;
 wire \CIRCUIT_2223.MEMORY_24.d ;
 wire \CIRCUIT_2223.MEMORY_24.s_currentState ;
 wire \CIRCUIT_2223.MEMORY_25.d ;
 wire \CIRCUIT_2223.MEMORY_25.s_currentState ;
 wire \CIRCUIT_2223.MEMORY_26.s_currentState ;
 wire \CIRCUIT_2223.s_logisimNet48 ;
 wire \CIRCUIT_2223.tone_generator_1.GATES_1.result ;
 wire \CIRCUIT_2223.tone_generator_1.GATES_2.result ;
 wire \CIRCUIT_2223.tone_generator_1.GATES_3.result ;
 wire \CIRCUIT_2223.tone_generator_1.MEMORY_10.s_currentState ;
 wire \CIRCUIT_2223.tone_generator_1.MEMORY_11.s_currentState ;
 wire \CIRCUIT_2223.tone_generator_1.MEMORY_12.s_currentState ;
 wire \CIRCUIT_2223.tone_generator_1.MEMORY_13.s_currentState ;
 wire \CIRCUIT_2223.tone_generator_1.MEMORY_14.s_currentState ;
 wire \CIRCUIT_2223.tone_generator_1.MEMORY_15.s_currentState ;
 wire \CIRCUIT_2223.tone_generator_1.MEMORY_16.s_currentState ;
 wire \CIRCUIT_2223.tone_generator_1.MEMORY_17.s_currentState ;
 wire \CIRCUIT_2223.tone_generator_1.MEMORY_18.s_currentState ;
 wire \CIRCUIT_2223.tone_generator_1.MEMORY_19.s_currentState ;
 wire \CIRCUIT_2223.tone_generator_1.MEMORY_20.s_currentState ;
 wire \CIRCUIT_2223.tone_generator_1.MEMORY_4.s_currentState ;
 wire \CIRCUIT_2223.tone_generator_1.MEMORY_6.s_currentState ;
 wire \CIRCUIT_2223.tone_generator_1.MEMORY_7.s_currentState ;
 wire \CIRCUIT_2223.tone_generator_1.MEMORY_8.s_currentState ;
 wire \CIRCUIT_2223.tone_generator_1.MEMORY_9.s_currentState ;
 wire \CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_10.input2 ;
 wire \CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_11.input2 ;
 wire \CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_12.input2 ;
 wire \CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_13.input2 ;
 wire \CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_14.input2 ;
 wire \CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_15.input2 ;
 wire \CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_16.input2 ;
 wire \CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_17.input2 ;
 wire \CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_27.result ;
 wire \CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_7.input2 ;
 wire \CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_8.input2 ;
 wire \CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_9.input2 ;
 wire \CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_28.clock ;
 wire \CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_28.d ;
 wire \CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_28.s_currentState ;
 wire \CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_29.d ;
 wire \CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_29.s_currentState ;
 wire \CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_30.d ;
 wire \CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_30.s_currentState ;
 wire \CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_31.d ;
 wire \CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_31.s_currentState ;
 wire \CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_32.d ;
 wire \CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_32.s_currentState ;
 wire \CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_33.d ;
 wire \CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_33.s_currentState ;
 wire \CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_34.d ;
 wire \CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_34.s_currentState ;
 wire \CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_35.d ;
 wire \CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_35.s_currentState ;
 wire \CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_36.d ;
 wire \CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_36.s_currentState ;
 wire \CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_37.d ;
 wire \CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_37.s_currentState ;
 wire \CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_38.s_currentState ;
 wire \CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_39.d ;
 wire \CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_39.s_currentState ;
 wire \CIRCUIT_2223.tone_generator_2_1.GATES_10.input2 ;
 wire \CIRCUIT_2223.tone_generator_2_1.GATES_11.input2 ;
 wire \CIRCUIT_2223.tone_generator_2_1.GATES_12.input2 ;
 wire \CIRCUIT_2223.tone_generator_2_1.GATES_13.input2 ;
 wire \CIRCUIT_2223.tone_generator_2_1.GATES_14.input2 ;
 wire \CIRCUIT_2223.tone_generator_2_1.GATES_15.input2 ;
 wire \CIRCUIT_2223.tone_generator_2_1.GATES_16.input2 ;
 wire \CIRCUIT_2223.tone_generator_2_1.GATES_17.input2 ;
 wire \CIRCUIT_2223.tone_generator_2_1.GATES_27.result ;
 wire \CIRCUIT_2223.tone_generator_2_1.GATES_7.input2 ;
 wire \CIRCUIT_2223.tone_generator_2_1.GATES_8.input2 ;
 wire \CIRCUIT_2223.tone_generator_2_1.GATES_9.input2 ;
 wire \CIRCUIT_2223.tone_generator_2_1.MEMORY_28.clock ;
 wire \CIRCUIT_2223.tone_generator_2_1.MEMORY_28.d ;
 wire \CIRCUIT_2223.tone_generator_2_1.MEMORY_28.s_currentState ;
 wire \CIRCUIT_2223.tone_generator_2_1.MEMORY_29.d ;
 wire \CIRCUIT_2223.tone_generator_2_1.MEMORY_29.s_currentState ;
 wire \CIRCUIT_2223.tone_generator_2_1.MEMORY_30.d ;
 wire \CIRCUIT_2223.tone_generator_2_1.MEMORY_30.s_currentState ;
 wire \CIRCUIT_2223.tone_generator_2_1.MEMORY_31.d ;
 wire \CIRCUIT_2223.tone_generator_2_1.MEMORY_31.s_currentState ;
 wire \CIRCUIT_2223.tone_generator_2_1.MEMORY_32.d ;
 wire \CIRCUIT_2223.tone_generator_2_1.MEMORY_32.s_currentState ;
 wire \CIRCUIT_2223.tone_generator_2_1.MEMORY_33.d ;
 wire \CIRCUIT_2223.tone_generator_2_1.MEMORY_33.s_currentState ;
 wire \CIRCUIT_2223.tone_generator_2_1.MEMORY_34.d ;
 wire \CIRCUIT_2223.tone_generator_2_1.MEMORY_34.s_currentState ;
 wire \CIRCUIT_2223.tone_generator_2_1.MEMORY_35.d ;
 wire \CIRCUIT_2223.tone_generator_2_1.MEMORY_35.s_currentState ;
 wire \CIRCUIT_2223.tone_generator_2_1.MEMORY_36.d ;
 wire \CIRCUIT_2223.tone_generator_2_1.MEMORY_36.s_currentState ;
 wire \CIRCUIT_2223.tone_generator_2_1.MEMORY_37.d ;
 wire \CIRCUIT_2223.tone_generator_2_1.MEMORY_37.s_currentState ;
 wire \CIRCUIT_2223.tone_generator_2_1.MEMORY_38.s_currentState ;
 wire \CIRCUIT_2223.tone_generator_2_1.MEMORY_39.d ;
 wire \CIRCUIT_2223.tone_generator_2_1.MEMORY_39.s_currentState ;
 wire \CIRCUIT_2223.tone_generator_2_2.GATES_10.input2 ;
 wire \CIRCUIT_2223.tone_generator_2_2.GATES_11.input2 ;
 wire \CIRCUIT_2223.tone_generator_2_2.GATES_12.input2 ;
 wire \CIRCUIT_2223.tone_generator_2_2.GATES_13.input2 ;
 wire \CIRCUIT_2223.tone_generator_2_2.GATES_14.input2 ;
 wire \CIRCUIT_2223.tone_generator_2_2.GATES_15.input2 ;
 wire \CIRCUIT_2223.tone_generator_2_2.GATES_16.input2 ;
 wire \CIRCUIT_2223.tone_generator_2_2.GATES_17.input2 ;
 wire \CIRCUIT_2223.tone_generator_2_2.GATES_27.result ;
 wire \CIRCUIT_2223.tone_generator_2_2.GATES_7.input2 ;
 wire \CIRCUIT_2223.tone_generator_2_2.GATES_8.input2 ;
 wire \CIRCUIT_2223.tone_generator_2_2.GATES_9.input2 ;
 wire \CIRCUIT_2223.tone_generator_2_2.MEMORY_28.clock ;
 wire \CIRCUIT_2223.tone_generator_2_2.MEMORY_28.d ;
 wire \CIRCUIT_2223.tone_generator_2_2.MEMORY_28.s_currentState ;
 wire \CIRCUIT_2223.tone_generator_2_2.MEMORY_29.d ;
 wire \CIRCUIT_2223.tone_generator_2_2.MEMORY_29.s_currentState ;
 wire \CIRCUIT_2223.tone_generator_2_2.MEMORY_30.d ;
 wire \CIRCUIT_2223.tone_generator_2_2.MEMORY_30.s_currentState ;
 wire \CIRCUIT_2223.tone_generator_2_2.MEMORY_31.d ;
 wire \CIRCUIT_2223.tone_generator_2_2.MEMORY_31.s_currentState ;
 wire \CIRCUIT_2223.tone_generator_2_2.MEMORY_32.d ;
 wire \CIRCUIT_2223.tone_generator_2_2.MEMORY_32.s_currentState ;
 wire \CIRCUIT_2223.tone_generator_2_2.MEMORY_33.d ;
 wire \CIRCUIT_2223.tone_generator_2_2.MEMORY_33.s_currentState ;
 wire \CIRCUIT_2223.tone_generator_2_2.MEMORY_34.d ;
 wire \CIRCUIT_2223.tone_generator_2_2.MEMORY_34.s_currentState ;
 wire \CIRCUIT_2223.tone_generator_2_2.MEMORY_35.d ;
 wire \CIRCUIT_2223.tone_generator_2_2.MEMORY_35.s_currentState ;
 wire \CIRCUIT_2223.tone_generator_2_2.MEMORY_36.d ;
 wire \CIRCUIT_2223.tone_generator_2_2.MEMORY_36.s_currentState ;
 wire \CIRCUIT_2223.tone_generator_2_2.MEMORY_37.d ;
 wire \CIRCUIT_2223.tone_generator_2_2.MEMORY_37.s_currentState ;
 wire \CIRCUIT_2223.tone_generator_2_2.MEMORY_38.s_currentState ;
 wire \CIRCUIT_2223.tone_generator_2_2.MEMORY_39.d ;
 wire \CIRCUIT_2223.tone_generator_2_2.MEMORY_39.s_currentState ;
 wire \CIRCUIT_2223.triangle_wave_generator_1.GATES_10.input2 ;
 wire \CIRCUIT_2223.triangle_wave_generator_1.GATES_11.input2 ;
 wire \CIRCUIT_2223.triangle_wave_generator_1.GATES_12.input2 ;
 wire \CIRCUIT_2223.triangle_wave_generator_1.GATES_13.input2 ;
 wire \CIRCUIT_2223.triangle_wave_generator_1.GATES_14.input2 ;
 wire \CIRCUIT_2223.triangle_wave_generator_1.GATES_15.input2 ;
 wire \CIRCUIT_2223.triangle_wave_generator_1.GATES_16.input2 ;
 wire \CIRCUIT_2223.triangle_wave_generator_1.GATES_17.input2 ;
 wire \CIRCUIT_2223.triangle_wave_generator_1.GATES_27.result ;
 wire \CIRCUIT_2223.triangle_wave_generator_1.GATES_7.input2 ;
 wire \CIRCUIT_2223.triangle_wave_generator_1.GATES_8.input2 ;
 wire \CIRCUIT_2223.triangle_wave_generator_1.GATES_9.input2 ;
 wire \CIRCUIT_2223.triangle_wave_generator_1.MEMORY_28.clock ;
 wire \CIRCUIT_2223.triangle_wave_generator_1.MEMORY_28.d ;
 wire \CIRCUIT_2223.triangle_wave_generator_1.MEMORY_28.s_currentState ;
 wire \CIRCUIT_2223.triangle_wave_generator_1.MEMORY_29.d ;
 wire \CIRCUIT_2223.triangle_wave_generator_1.MEMORY_29.s_currentState ;
 wire \CIRCUIT_2223.triangle_wave_generator_1.MEMORY_30.d ;
 wire \CIRCUIT_2223.triangle_wave_generator_1.MEMORY_30.s_currentState ;
 wire \CIRCUIT_2223.triangle_wave_generator_1.MEMORY_31.d ;
 wire \CIRCUIT_2223.triangle_wave_generator_1.MEMORY_31.s_currentState ;
 wire \CIRCUIT_2223.triangle_wave_generator_1.MEMORY_32.d ;
 wire \CIRCUIT_2223.triangle_wave_generator_1.MEMORY_32.s_currentState ;
 wire \CIRCUIT_2223.triangle_wave_generator_1.MEMORY_33.d ;
 wire \CIRCUIT_2223.triangle_wave_generator_1.MEMORY_33.s_currentState ;
 wire \CIRCUIT_2223.triangle_wave_generator_1.MEMORY_34.d ;
 wire \CIRCUIT_2223.triangle_wave_generator_1.MEMORY_34.s_currentState ;
 wire \CIRCUIT_2223.triangle_wave_generator_1.MEMORY_35.d ;
 wire \CIRCUIT_2223.triangle_wave_generator_1.MEMORY_35.s_currentState ;
 wire \CIRCUIT_2223.triangle_wave_generator_1.MEMORY_36.d ;
 wire \CIRCUIT_2223.triangle_wave_generator_1.MEMORY_36.s_currentState ;
 wire \CIRCUIT_2223.triangle_wave_generator_1.MEMORY_37.d ;
 wire \CIRCUIT_2223.triangle_wave_generator_1.MEMORY_37.s_currentState ;
 wire \CIRCUIT_2223.triangle_wave_generator_1.MEMORY_38.s_currentState ;
 wire \CIRCUIT_2223.triangle_wave_generator_1.MEMORY_39.d ;
 wire \CIRCUIT_2223.triangle_wave_generator_1.MEMORY_39.s_currentState ;
 wire \CIRCUIT_2223.triangle_wave_generator_1.MEMORY_40.clock ;
 wire \CIRCUIT_2223.triangle_wave_generator_1.MEMORY_40.d ;
 wire \CIRCUIT_2223.triangle_wave_generator_1.MEMORY_40.s_currentState ;
 wire \CIRCUIT_2223.triangle_wave_generator_1.MEMORY_41.clock ;
 wire \CIRCUIT_2223.triangle_wave_generator_1.MEMORY_41.s_currentState ;
 wire \CIRCUIT_2223.triangle_wave_generator_1.MEMORY_42.s_currentState ;
 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire _236_;
 wire _237_;
 wire _238_;
 wire _239_;
 wire _240_;
 wire _241_;
 wire _242_;
 wire _243_;
 wire _244_;
 wire _245_;
 wire _246_;
 wire _247_;
 wire _248_;
 wire _249_;
 wire _250_;
 wire _251_;
 wire _252_;
 wire _253_;
 wire _254_;
 wire _255_;
 wire _256_;
 wire _257_;
 wire _258_;
 wire _259_;
 wire _260_;
 wire _261_;
 wire _262_;
 wire _263_;
 wire _264_;
 wire _265_;
 wire _266_;
 wire _267_;
 wire _268_;
 wire _269_;
 wire _270_;
 wire _271_;
 wire _272_;
 wire _273_;
 wire _274_;
 wire _275_;
 wire _276_;
 wire _277_;
 wire _278_;
 wire _279_;
 wire _280_;
 wire _281_;
 wire _282_;
 wire _283_;
 wire _284_;
 wire _285_;
 wire _286_;
 wire _287_;
 wire _288_;
 wire _289_;
 wire _290_;
 wire _291_;
 wire _292_;
 wire _293_;
 wire _294_;
 wire _295_;
 wire _296_;
 wire _297_;
 wire _298_;
 wire _299_;
 wire _300_;
 wire _301_;
 wire _302_;
 wire _303_;
 wire _304_;
 wire _305_;
 wire _306_;
 wire _307_;
 wire clknet_0__183_;
 wire clknet_0__203_;
 wire clknet_0__222_;
 wire clknet_0__245_;
 wire clknet_0__264_;
 wire clknet_0_clk;
 wire clknet_1_0__leaf__183_;
 wire clknet_1_0__leaf__203_;
 wire clknet_1_0__leaf__222_;
 wire clknet_1_0__leaf__245_;
 wire clknet_1_0__leaf__264_;
 wire clknet_1_0__leaf_clk;
 wire clknet_1_1__leaf__183_;
 wire clknet_1_1__leaf__203_;
 wire clknet_1_1__leaf__222_;
 wire clknet_1_1__leaf__245_;
 wire clknet_1_1__leaf__264_;
 wire clknet_1_1__leaf_clk;
 wire net1;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net2;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net3;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net4;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire \slow_clock[0] ;
 wire \slow_clock[1] ;
 wire \slow_clock[2] ;
 wire \slow_clock[3] ;
 wire \slow_clock[4] ;
 wire \slow_clock[5] ;
 wire \slow_clock[6] ;

 sky130_fd_sc_hd__decap_3 FILLER_0_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_258 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_280 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_216 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_298 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_160 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_212 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_80 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_191 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_50 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_16 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_180 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_23 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_48 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_243 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_25 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_296 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_104 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_152 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_219 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_192 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_68 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_268 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_207 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_219 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_129 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_164 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_188 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_252 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_296 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_43 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_296 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_144 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_191 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_298 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_32 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_72 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_84 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_10 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_122 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_213 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_238 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_128 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_84 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_96 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_152 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_16 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_263 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_31 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_114 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_21 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_271 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_36 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_62 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_215 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_236 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_246 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_124 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_176 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_200 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_254 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_32 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_40 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_96 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_201 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_297 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_187 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_199 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_298 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_49 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_98 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_43 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_296 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_74 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_156 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_298 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_36 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_212 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_254 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_298 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_48 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_213 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_296 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_255 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_36 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_25 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_256 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_171 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_214 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_46 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_124 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_252 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_90 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_156 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_168 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_38 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_94 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_100 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_123 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_162 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_210 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_298 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_127 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_220 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_291 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_36 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_44 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_243 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_32 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_76 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_24 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_114 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_76 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_286 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_36 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_188 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_291 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_206 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_214 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_298 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_50 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_63 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_78 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_295 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_32 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_52 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_95 ();
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_94 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_95 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_96 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_97 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_98 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_99 ();
 sky130_fd_sc_hd__inv_2 _308_ (.A(net24),
    .Y(_117_));
 sky130_fd_sc_hd__inv_2 _309_ (.A(\CIRCUIT_2223.GATES_1.input1[1] ),
    .Y(_179_));
 sky130_fd_sc_hd__inv_2 _310_ (.A(\CIRCUIT_2223.MEMORY_23.s_currentState ),
    .Y(\CIRCUIT_2223.GATES_11.input2 ));
 sky130_fd_sc_hd__inv_2 _311_ (.A(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_38.s_currentState ),
    .Y(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_28.clock ));
 sky130_fd_sc_hd__inv_2 _312_ (.A(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_37.s_currentState ),
    .Y(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_37.d ));
 sky130_fd_sc_hd__inv_2 _313_ (.A(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_36.s_currentState ),
    .Y(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_36.d ));
 sky130_fd_sc_hd__inv_2 _314_ (.A(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_35.s_currentState ),
    .Y(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_35.d ));
 sky130_fd_sc_hd__inv_2 _315_ (.A(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_34.s_currentState ),
    .Y(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_34.d ));
 sky130_fd_sc_hd__inv_2 _316_ (.A(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_33.s_currentState ),
    .Y(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_33.d ));
 sky130_fd_sc_hd__inv_2 _317_ (.A(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_32.s_currentState ),
    .Y(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_32.d ));
 sky130_fd_sc_hd__inv_2 _318_ (.A(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_31.s_currentState ),
    .Y(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_31.d ));
 sky130_fd_sc_hd__inv_2 _319_ (.A(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_30.s_currentState ),
    .Y(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_30.d ));
 sky130_fd_sc_hd__inv_2 _320_ (.A(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_29.s_currentState ),
    .Y(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_29.d ));
 sky130_fd_sc_hd__inv_2 _321_ (.A(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_28.s_currentState ),
    .Y(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_28.d ));
 sky130_fd_sc_hd__inv_2 _322_ (.A(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_39.s_currentState ),
    .Y(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_39.d ));
 sky130_fd_sc_hd__inv_2 _323_ (.A(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_39.s_currentState ),
    .Y(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_39.d ));
 sky130_fd_sc_hd__inv_2 _324_ (.A(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_40.s_currentState ),
    .Y(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_40.d ));
 sky130_fd_sc_hd__inv_2 _325_ (.A(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_41.s_currentState ),
    .Y(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_40.clock ));
 sky130_fd_sc_hd__inv_2 _326_ (.A(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_42.s_currentState ),
    .Y(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_41.clock ));
 sky130_fd_sc_hd__inv_2 _327_ (.A(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_28.s_currentState ),
    .Y(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_28.d ));
 sky130_fd_sc_hd__inv_2 _328_ (.A(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_29.s_currentState ),
    .Y(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_29.d ));
 sky130_fd_sc_hd__inv_2 _329_ (.A(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_30.s_currentState ),
    .Y(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_30.d ));
 sky130_fd_sc_hd__inv_2 _330_ (.A(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_31.s_currentState ),
    .Y(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_31.d ));
 sky130_fd_sc_hd__inv_2 _331_ (.A(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_32.s_currentState ),
    .Y(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_32.d ));
 sky130_fd_sc_hd__inv_2 _332_ (.A(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_33.s_currentState ),
    .Y(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_33.d ));
 sky130_fd_sc_hd__inv_2 _333_ (.A(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_34.s_currentState ),
    .Y(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_34.d ));
 sky130_fd_sc_hd__inv_2 _334_ (.A(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_35.s_currentState ),
    .Y(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_35.d ));
 sky130_fd_sc_hd__inv_2 _335_ (.A(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_36.s_currentState ),
    .Y(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_36.d ));
 sky130_fd_sc_hd__inv_2 _336_ (.A(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_37.s_currentState ),
    .Y(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_37.d ));
 sky130_fd_sc_hd__inv_2 _337_ (.A(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_38.s_currentState ),
    .Y(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_28.clock ));
 sky130_fd_sc_hd__inv_2 _338_ (.A(\CIRCUIT_2223.tone_generator_2_1.MEMORY_39.s_currentState ),
    .Y(\CIRCUIT_2223.tone_generator_2_1.MEMORY_39.d ));
 sky130_fd_sc_hd__inv_2 _339_ (.A(\CIRCUIT_2223.tone_generator_2_1.MEMORY_28.s_currentState ),
    .Y(\CIRCUIT_2223.tone_generator_2_1.MEMORY_28.d ));
 sky130_fd_sc_hd__inv_2 _340_ (.A(\CIRCUIT_2223.tone_generator_2_1.MEMORY_29.s_currentState ),
    .Y(\CIRCUIT_2223.tone_generator_2_1.MEMORY_29.d ));
 sky130_fd_sc_hd__inv_2 _341_ (.A(\CIRCUIT_2223.tone_generator_2_1.MEMORY_30.s_currentState ),
    .Y(\CIRCUIT_2223.tone_generator_2_1.MEMORY_30.d ));
 sky130_fd_sc_hd__inv_2 _342_ (.A(\CIRCUIT_2223.tone_generator_2_1.MEMORY_31.s_currentState ),
    .Y(\CIRCUIT_2223.tone_generator_2_1.MEMORY_31.d ));
 sky130_fd_sc_hd__inv_2 _343_ (.A(\CIRCUIT_2223.tone_generator_2_1.MEMORY_32.s_currentState ),
    .Y(\CIRCUIT_2223.tone_generator_2_1.MEMORY_32.d ));
 sky130_fd_sc_hd__inv_2 _344_ (.A(\CIRCUIT_2223.tone_generator_2_1.MEMORY_33.s_currentState ),
    .Y(\CIRCUIT_2223.tone_generator_2_1.MEMORY_33.d ));
 sky130_fd_sc_hd__inv_2 _345_ (.A(\CIRCUIT_2223.tone_generator_2_1.MEMORY_34.s_currentState ),
    .Y(\CIRCUIT_2223.tone_generator_2_1.MEMORY_34.d ));
 sky130_fd_sc_hd__inv_2 _346_ (.A(\CIRCUIT_2223.tone_generator_2_1.MEMORY_35.s_currentState ),
    .Y(\CIRCUIT_2223.tone_generator_2_1.MEMORY_35.d ));
 sky130_fd_sc_hd__inv_2 _347_ (.A(\CIRCUIT_2223.tone_generator_2_1.MEMORY_36.s_currentState ),
    .Y(\CIRCUIT_2223.tone_generator_2_1.MEMORY_36.d ));
 sky130_fd_sc_hd__inv_2 _348_ (.A(\CIRCUIT_2223.tone_generator_2_1.MEMORY_37.s_currentState ),
    .Y(\CIRCUIT_2223.tone_generator_2_1.MEMORY_37.d ));
 sky130_fd_sc_hd__inv_2 _349_ (.A(\CIRCUIT_2223.tone_generator_2_1.MEMORY_38.s_currentState ),
    .Y(\CIRCUIT_2223.tone_generator_2_1.MEMORY_28.clock ));
 sky130_fd_sc_hd__inv_2 _350_ (.A(\CIRCUIT_2223.tone_generator_2_2.MEMORY_39.s_currentState ),
    .Y(\CIRCUIT_2223.tone_generator_2_2.MEMORY_39.d ));
 sky130_fd_sc_hd__inv_2 _351_ (.A(\CIRCUIT_2223.tone_generator_2_2.MEMORY_28.s_currentState ),
    .Y(\CIRCUIT_2223.tone_generator_2_2.MEMORY_28.d ));
 sky130_fd_sc_hd__inv_2 _352_ (.A(\CIRCUIT_2223.tone_generator_2_2.MEMORY_29.s_currentState ),
    .Y(\CIRCUIT_2223.tone_generator_2_2.MEMORY_29.d ));
 sky130_fd_sc_hd__inv_2 _353_ (.A(\CIRCUIT_2223.tone_generator_2_2.MEMORY_30.s_currentState ),
    .Y(\CIRCUIT_2223.tone_generator_2_2.MEMORY_30.d ));
 sky130_fd_sc_hd__inv_2 _354_ (.A(\CIRCUIT_2223.tone_generator_2_2.MEMORY_31.s_currentState ),
    .Y(\CIRCUIT_2223.tone_generator_2_2.MEMORY_31.d ));
 sky130_fd_sc_hd__inv_2 _355_ (.A(\CIRCUIT_2223.tone_generator_2_2.MEMORY_32.s_currentState ),
    .Y(\CIRCUIT_2223.tone_generator_2_2.MEMORY_32.d ));
 sky130_fd_sc_hd__inv_2 _356_ (.A(\CIRCUIT_2223.tone_generator_2_2.MEMORY_33.s_currentState ),
    .Y(\CIRCUIT_2223.tone_generator_2_2.MEMORY_33.d ));
 sky130_fd_sc_hd__inv_2 _357_ (.A(\CIRCUIT_2223.tone_generator_2_2.MEMORY_34.s_currentState ),
    .Y(\CIRCUIT_2223.tone_generator_2_2.MEMORY_34.d ));
 sky130_fd_sc_hd__inv_2 _358_ (.A(\CIRCUIT_2223.tone_generator_2_2.MEMORY_35.s_currentState ),
    .Y(\CIRCUIT_2223.tone_generator_2_2.MEMORY_35.d ));
 sky130_fd_sc_hd__inv_2 _359_ (.A(\CIRCUIT_2223.tone_generator_2_2.MEMORY_36.s_currentState ),
    .Y(\CIRCUIT_2223.tone_generator_2_2.MEMORY_36.d ));
 sky130_fd_sc_hd__inv_2 _360_ (.A(\CIRCUIT_2223.tone_generator_2_2.MEMORY_37.s_currentState ),
    .Y(\CIRCUIT_2223.tone_generator_2_2.MEMORY_37.d ));
 sky130_fd_sc_hd__inv_2 _361_ (.A(\CIRCUIT_2223.tone_generator_2_2.MEMORY_38.s_currentState ),
    .Y(\CIRCUIT_2223.tone_generator_2_2.MEMORY_28.clock ));
 sky130_fd_sc_hd__inv_2 _362_ (.A(\CIRCUIT_2223.MEMORY_26.s_currentState ),
    .Y(\CIRCUIT_2223.MEMORY_18.clock ));
 sky130_fd_sc_hd__inv_2 _363_ (.A(\CIRCUIT_2223.MEMORY_25.s_currentState ),
    .Y(\CIRCUIT_2223.MEMORY_25.d ));
 sky130_fd_sc_hd__inv_2 _364_ (.A(net17),
    .Y(\CIRCUIT_2223.MEMORY_24.d ));
 sky130_fd_sc_hd__inv_2 _365_ (.A(\CIRCUIT_2223.MEMORY_22.s_currentState ),
    .Y(\CIRCUIT_2223.MEMORY_22.d ));
 sky130_fd_sc_hd__inv_2 _366_ (.A(\CIRCUIT_2223.MEMORY_21.s_currentState ),
    .Y(\CIRCUIT_2223.MEMORY_21.d ));
 sky130_fd_sc_hd__inv_2 _367_ (.A(\CIRCUIT_2223.MEMORY_20.s_currentState ),
    .Y(\CIRCUIT_2223.MEMORY_20.d ));
 sky130_fd_sc_hd__inv_2 _368_ (.A(\CIRCUIT_2223.MEMORY_19.s_currentState ),
    .Y(\CIRCUIT_2223.MEMORY_19.d ));
 sky130_fd_sc_hd__inv_2 _369_ (.A(\CIRCUIT_2223.MEMORY_18.s_currentState ),
    .Y(\CIRCUIT_2223.MEMORY_18.d ));
 sky130_fd_sc_hd__and4_4 _370_ (.A(net2),
    .B(net1),
    .C(\CIRCUIT_2223.GATES_1.input1[0] ),
    .D(\CIRCUIT_2223.GATES_1.input1[1] ),
    .X(_180_));
 sky130_fd_sc_hd__and4_4 _371_ (.A(net2),
    .B(net1),
    .C(\CIRCUIT_2223.GATES_1.input1[2] ),
    .D(\CIRCUIT_2223.GATES_1.input1[3] ),
    .X(_181_));
 sky130_fd_sc_hd__nand2_4 _372_ (.A(_180_),
    .B(_181_),
    .Y(_182_));
 sky130_fd_sc_hd__mux2_1 _373_ (.A0(net6),
    .A1(\CIRCUIT_2223.s_logisimNet48 ),
    .S(_182_),
    .X(_178_));
 sky130_fd_sc_hd__mux2_1 _374_ (.A0(net35),
    .A1(\CIRCUIT_2223.GATES_5.input2 ),
    .S(_182_),
    .X(_177_));
 sky130_fd_sc_hd__mux2_1 _375_ (.A0(net36),
    .A1(\CIRCUIT_2223.GATES_3.input2 ),
    .S(_182_),
    .X(_176_));
 sky130_fd_sc_hd__mux2_1 _376_ (.A0(net37),
    .A1(\CIRCUIT_2223.GATES_2.input2 ),
    .S(_182_),
    .X(_175_));
 sky130_fd_sc_hd__nand2_8 _377_ (.A(net23),
    .B(net33),
    .Y(_000_));
 sky130_fd_sc_hd__nand2_2 _378_ (.A(clknet_1_0__leaf_clk),
    .B(\CIRCUIT_2223.GATES_11.input2 ),
    .Y(_183_));
 sky130_fd_sc_hd__inv_2 _379__1 (.A(clknet_1_0__leaf__183_),
    .Y(net39));
 sky130_fd_sc_hd__inv_2 _379__2 (.A(clknet_1_0__leaf__183_),
    .Y(net40));
 sky130_fd_sc_hd__xor2_1 _380_ (.A(\CIRCUIT_2223.tone_generator_2_2.MEMORY_28.s_currentState ),
    .B(\CIRCUIT_2223.tone_generator_2_2.GATES_7.input2 ),
    .X(_184_));
 sky130_fd_sc_hd__xor2_1 _381_ (.A(\CIRCUIT_2223.tone_generator_2_2.MEMORY_30.s_currentState ),
    .B(\CIRCUIT_2223.tone_generator_2_2.GATES_9.input2 ),
    .X(_185_));
 sky130_fd_sc_hd__or2_1 _382_ (.A(\CIRCUIT_2223.tone_generator_2_2.MEMORY_38.s_currentState ),
    .B(\CIRCUIT_2223.tone_generator_2_2.GATES_17.input2 ),
    .X(_186_));
 sky130_fd_sc_hd__nand2_1 _383_ (.A(\CIRCUIT_2223.tone_generator_2_2.MEMORY_38.s_currentState ),
    .B(\CIRCUIT_2223.tone_generator_2_2.GATES_17.input2 ),
    .Y(_187_));
 sky130_fd_sc_hd__xor2_1 _384_ (.A(\CIRCUIT_2223.tone_generator_2_2.MEMORY_33.s_currentState ),
    .B(\CIRCUIT_2223.tone_generator_2_2.GATES_12.input2 ),
    .X(_188_));
 sky130_fd_sc_hd__xor2_1 _385_ (.A(\CIRCUIT_2223.tone_generator_2_2.MEMORY_34.s_currentState ),
    .B(\CIRCUIT_2223.tone_generator_2_2.GATES_13.input2 ),
    .X(_189_));
 sky130_fd_sc_hd__xor2_1 _386_ (.A(\CIRCUIT_2223.tone_generator_2_2.MEMORY_36.s_currentState ),
    .B(\CIRCUIT_2223.tone_generator_2_2.GATES_15.input2 ),
    .X(_190_));
 sky130_fd_sc_hd__or2_1 _387_ (.A(\CIRCUIT_2223.tone_generator_2_2.MEMORY_29.s_currentState ),
    .B(\CIRCUIT_2223.tone_generator_2_2.GATES_8.input2 ),
    .X(_191_));
 sky130_fd_sc_hd__nand2_1 _388_ (.A(\CIRCUIT_2223.tone_generator_2_2.MEMORY_29.s_currentState ),
    .B(\CIRCUIT_2223.tone_generator_2_2.GATES_8.input2 ),
    .Y(_192_));
 sky130_fd_sc_hd__xor2_1 _389_ (.A(\CIRCUIT_2223.tone_generator_2_2.MEMORY_32.s_currentState ),
    .B(\CIRCUIT_2223.tone_generator_2_2.GATES_11.input2 ),
    .X(_193_));
 sky130_fd_sc_hd__xor2_1 _390_ (.A(\CIRCUIT_2223.tone_generator_2_2.MEMORY_31.s_currentState ),
    .B(\CIRCUIT_2223.tone_generator_2_2.GATES_10.input2 ),
    .X(_194_));
 sky130_fd_sc_hd__or4_1 _391_ (.A(_188_),
    .B(_189_),
    .C(_190_),
    .D(_194_),
    .X(_195_));
 sky130_fd_sc_hd__a221o_1 _392_ (.A1(_186_),
    .A2(_187_),
    .B1(_191_),
    .B2(_192_),
    .C1(_193_),
    .X(_196_));
 sky130_fd_sc_hd__xor2_1 _393_ (.A(\CIRCUIT_2223.tone_generator_2_2.MEMORY_35.s_currentState ),
    .B(\CIRCUIT_2223.tone_generator_2_2.GATES_14.input2 ),
    .X(_197_));
 sky130_fd_sc_hd__xor2_1 _394_ (.A(\CIRCUIT_2223.tone_generator_2_2.MEMORY_37.s_currentState ),
    .B(\CIRCUIT_2223.tone_generator_2_2.GATES_16.input2 ),
    .X(_198_));
 sky130_fd_sc_hd__or4_1 _395_ (.A(_184_),
    .B(_185_),
    .C(_197_),
    .D(_198_),
    .X(_199_));
 sky130_fd_sc_hd__nor3_2 _396_ (.A(_195_),
    .B(_196_),
    .C(_199_),
    .Y(\CIRCUIT_2223.tone_generator_2_2.GATES_27.result ));
 sky130_fd_sc_hd__o211ai_4 _397_ (.A1(\CIRCUIT_2223.GATES_1.input1[2] ),
    .A2(\CIRCUIT_2223.GATES_1.input1[3] ),
    .B1(net2),
    .C1(net1),
    .Y(_200_));
 sky130_fd_sc_hd__o211ai_4 _398_ (.A1(\CIRCUIT_2223.GATES_1.input1[0] ),
    .A2(\CIRCUIT_2223.GATES_1.input1[1] ),
    .B1(net2),
    .C1(net1),
    .Y(_201_));
 sky130_fd_sc_hd__inv_2 _399_ (.A(_201_),
    .Y(_202_));
 sky130_fd_sc_hd__a32o_2 _400_ (.A1(net30),
    .A2(_200_),
    .A3(_202_),
    .B1(clknet_1_1__leaf__183_),
    .B2(\CIRCUIT_2223.tone_generator_2_2.GATES_27.result ),
    .X(_203_));
 sky130_fd_sc_hd__xor2_2 _401_ (.A(net19),
    .B(clknet_1_1__leaf__203_),
    .X(_094_));
 sky130_fd_sc_hd__xor2_1 _402_ (.A(\CIRCUIT_2223.tone_generator_2_1.MEMORY_29.s_currentState ),
    .B(\CIRCUIT_2223.tone_generator_2_1.GATES_8.input2 ),
    .X(_204_));
 sky130_fd_sc_hd__xor2_1 _403_ (.A(\CIRCUIT_2223.tone_generator_2_1.MEMORY_33.s_currentState ),
    .B(\CIRCUIT_2223.tone_generator_2_1.GATES_12.input2 ),
    .X(_205_));
 sky130_fd_sc_hd__xor2_1 _404_ (.A(\CIRCUIT_2223.tone_generator_2_1.MEMORY_30.s_currentState ),
    .B(\CIRCUIT_2223.tone_generator_2_1.GATES_9.input2 ),
    .X(_206_));
 sky130_fd_sc_hd__or2_1 _405_ (.A(\CIRCUIT_2223.tone_generator_2_1.MEMORY_38.s_currentState ),
    .B(\CIRCUIT_2223.tone_generator_2_1.GATES_17.input2 ),
    .X(_207_));
 sky130_fd_sc_hd__nand2_1 _406_ (.A(\CIRCUIT_2223.tone_generator_2_1.MEMORY_38.s_currentState ),
    .B(\CIRCUIT_2223.tone_generator_2_1.GATES_17.input2 ),
    .Y(_208_));
 sky130_fd_sc_hd__xor2_1 _407_ (.A(\CIRCUIT_2223.tone_generator_2_1.MEMORY_37.s_currentState ),
    .B(\CIRCUIT_2223.tone_generator_2_1.GATES_16.input2 ),
    .X(_209_));
 sky130_fd_sc_hd__xor2_1 _408_ (.A(\CIRCUIT_2223.tone_generator_2_1.MEMORY_28.s_currentState ),
    .B(\CIRCUIT_2223.tone_generator_2_1.GATES_7.input2 ),
    .X(_210_));
 sky130_fd_sc_hd__xor2_1 _409_ (.A(\CIRCUIT_2223.tone_generator_2_1.MEMORY_31.s_currentState ),
    .B(\CIRCUIT_2223.tone_generator_2_1.GATES_10.input2 ),
    .X(_211_));
 sky130_fd_sc_hd__xor2_1 _410_ (.A(\CIRCUIT_2223.tone_generator_2_1.MEMORY_36.s_currentState ),
    .B(\CIRCUIT_2223.tone_generator_2_1.GATES_15.input2 ),
    .X(_212_));
 sky130_fd_sc_hd__xor2_1 _411_ (.A(\CIRCUIT_2223.tone_generator_2_1.MEMORY_34.s_currentState ),
    .B(\CIRCUIT_2223.tone_generator_2_1.GATES_13.input2 ),
    .X(_213_));
 sky130_fd_sc_hd__or4_1 _412_ (.A(_205_),
    .B(_211_),
    .C(_212_),
    .D(_213_),
    .X(_214_));
 sky130_fd_sc_hd__nand2_1 _413_ (.A(\CIRCUIT_2223.tone_generator_2_1.MEMORY_32.s_currentState ),
    .B(\CIRCUIT_2223.tone_generator_2_1.GATES_11.input2 ),
    .Y(_215_));
 sky130_fd_sc_hd__or2_1 _414_ (.A(\CIRCUIT_2223.tone_generator_2_1.MEMORY_32.s_currentState ),
    .B(\CIRCUIT_2223.tone_generator_2_1.GATES_11.input2 ),
    .X(_216_));
 sky130_fd_sc_hd__a221o_1 _415_ (.A1(_207_),
    .A2(_208_),
    .B1(_215_),
    .B2(_216_),
    .C1(_204_),
    .X(_217_));
 sky130_fd_sc_hd__xor2_1 _416_ (.A(\CIRCUIT_2223.tone_generator_2_1.MEMORY_35.s_currentState ),
    .B(\CIRCUIT_2223.tone_generator_2_1.GATES_14.input2 ),
    .X(_218_));
 sky130_fd_sc_hd__or4_1 _417_ (.A(_206_),
    .B(_209_),
    .C(_210_),
    .D(_218_),
    .X(_219_));
 sky130_fd_sc_hd__nor3_2 _418_ (.A(_214_),
    .B(_217_),
    .C(_219_),
    .Y(\CIRCUIT_2223.tone_generator_2_1.GATES_27.result ));
 sky130_fd_sc_hd__and4b_4 _419_ (.A_N(\CIRCUIT_2223.GATES_1.input1[3] ),
    .B(\CIRCUIT_2223.GATES_1.input1[2] ),
    .C(net1),
    .D(net2),
    .X(_220_));
 sky130_fd_sc_hd__and3b_1 _420_ (.A_N(_180_),
    .B(_220_),
    .C(net30),
    .X(_221_));
 sky130_fd_sc_hd__a21oi_2 _421_ (.A1(clknet_1_1__leaf__183_),
    .A2(\CIRCUIT_2223.tone_generator_2_1.GATES_27.result ),
    .B1(_221_),
    .Y(_222_));
 sky130_fd_sc_hd__xnor2_2 _422_ (.A(net21),
    .B(clknet_1_1__leaf__222_),
    .Y(_073_));
 sky130_fd_sc_hd__nand2_1 _423_ (.A(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_36.s_currentState ),
    .B(\CIRCUIT_2223.triangle_wave_generator_1.GATES_15.input2 ),
    .Y(_223_));
 sky130_fd_sc_hd__or2_1 _424_ (.A(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_36.s_currentState ),
    .B(\CIRCUIT_2223.triangle_wave_generator_1.GATES_15.input2 ),
    .X(_224_));
 sky130_fd_sc_hd__nand2_1 _425_ (.A(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_33.s_currentState ),
    .B(\CIRCUIT_2223.triangle_wave_generator_1.GATES_12.input2 ),
    .Y(_225_));
 sky130_fd_sc_hd__or2_1 _426_ (.A(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_33.s_currentState ),
    .B(\CIRCUIT_2223.triangle_wave_generator_1.GATES_12.input2 ),
    .X(_226_));
 sky130_fd_sc_hd__a22o_1 _427_ (.A1(_223_),
    .A2(_224_),
    .B1(_225_),
    .B2(_226_),
    .X(_227_));
 sky130_fd_sc_hd__xor2_1 _428_ (.A(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_30.s_currentState ),
    .B(\CIRCUIT_2223.triangle_wave_generator_1.GATES_9.input2 ),
    .X(_228_));
 sky130_fd_sc_hd__xor2_1 _429_ (.A(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_38.s_currentState ),
    .B(\CIRCUIT_2223.triangle_wave_generator_1.GATES_17.input2 ),
    .X(_229_));
 sky130_fd_sc_hd__xor2_1 _430_ (.A(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_37.s_currentState ),
    .B(\CIRCUIT_2223.triangle_wave_generator_1.GATES_16.input2 ),
    .X(_230_));
 sky130_fd_sc_hd__nand2_1 _431_ (.A(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_35.s_currentState ),
    .B(\CIRCUIT_2223.triangle_wave_generator_1.GATES_14.input2 ),
    .Y(_231_));
 sky130_fd_sc_hd__or2_1 _432_ (.A(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_35.s_currentState ),
    .B(\CIRCUIT_2223.triangle_wave_generator_1.GATES_14.input2 ),
    .X(_232_));
 sky130_fd_sc_hd__xor2_1 _433_ (.A(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_29.s_currentState ),
    .B(\CIRCUIT_2223.triangle_wave_generator_1.GATES_8.input2 ),
    .X(_233_));
 sky130_fd_sc_hd__xor2_1 _434_ (.A(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_32.s_currentState ),
    .B(\CIRCUIT_2223.triangle_wave_generator_1.GATES_11.input2 ),
    .X(_234_));
 sky130_fd_sc_hd__or2_1 _435_ (.A(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_28.s_currentState ),
    .B(\CIRCUIT_2223.triangle_wave_generator_1.GATES_7.input2 ),
    .X(_235_));
 sky130_fd_sc_hd__nand2_1 _436_ (.A(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_28.s_currentState ),
    .B(\CIRCUIT_2223.triangle_wave_generator_1.GATES_7.input2 ),
    .Y(_236_));
 sky130_fd_sc_hd__xor2_1 _437_ (.A(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_31.s_currentState ),
    .B(\CIRCUIT_2223.triangle_wave_generator_1.GATES_10.input2 ),
    .X(_237_));
 sky130_fd_sc_hd__xor2_1 _438_ (.A(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_34.s_currentState ),
    .B(\CIRCUIT_2223.triangle_wave_generator_1.GATES_13.input2 ),
    .X(_238_));
 sky130_fd_sc_hd__a221o_1 _439_ (.A1(_231_),
    .A2(_232_),
    .B1(_235_),
    .B2(_236_),
    .C1(_237_),
    .X(_239_));
 sky130_fd_sc_hd__or4_1 _440_ (.A(_228_),
    .B(_233_),
    .C(_234_),
    .D(_238_),
    .X(_240_));
 sky130_fd_sc_hd__or4_2 _441_ (.A(_227_),
    .B(_229_),
    .C(_230_),
    .D(_240_),
    .X(_241_));
 sky130_fd_sc_hd__nor2_1 _442_ (.A(_239_),
    .B(_241_),
    .Y(\CIRCUIT_2223.triangle_wave_generator_1.GATES_27.result ));
 sky130_fd_sc_hd__nand2_4 _443_ (.A(_180_),
    .B(_220_),
    .Y(_242_));
 sky130_fd_sc_hd__and4b_4 _444_ (.A_N(\CIRCUIT_2223.GATES_1.input1[2] ),
    .B(\CIRCUIT_2223.GATES_1.input1[3] ),
    .C(net2),
    .D(net1),
    .X(_243_));
 sky130_fd_sc_hd__a21boi_1 _445_ (.A1(_179_),
    .A2(_243_),
    .B1_N(_242_),
    .Y(_244_));
 sky130_fd_sc_hd__o32a_2 _446_ (.A1(net40),
    .A2(_239_),
    .A3(_241_),
    .B1(_244_),
    .B2(_117_),
    .X(_245_));
 sky130_fd_sc_hd__xnor2_2 _447_ (.A(net18),
    .B(clknet_1_1__leaf__245_),
    .Y(_049_));
 sky130_fd_sc_hd__or2_1 _448_ (.A(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_29.s_currentState ),
    .B(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_8.input2 ),
    .X(_246_));
 sky130_fd_sc_hd__nand2_1 _449_ (.A(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_29.s_currentState ),
    .B(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_8.input2 ),
    .Y(_247_));
 sky130_fd_sc_hd__xor2_1 _450_ (.A(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_28.s_currentState ),
    .B(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_7.input2 ),
    .X(_248_));
 sky130_fd_sc_hd__xor2_1 _451_ (.A(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_33.s_currentState ),
    .B(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_12.input2 ),
    .X(_249_));
 sky130_fd_sc_hd__xor2_1 _452_ (.A(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_30.s_currentState ),
    .B(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_9.input2 ),
    .X(_250_));
 sky130_fd_sc_hd__xor2_1 _453_ (.A(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_38.s_currentState ),
    .B(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_17.input2 ),
    .X(_251_));
 sky130_fd_sc_hd__xor2_1 _454_ (.A(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_35.s_currentState ),
    .B(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_14.input2 ),
    .X(_252_));
 sky130_fd_sc_hd__xor2_1 _455_ (.A(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_31.s_currentState ),
    .B(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_10.input2 ),
    .X(_253_));
 sky130_fd_sc_hd__xor2_1 _456_ (.A(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_36.s_currentState ),
    .B(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_15.input2 ),
    .X(_254_));
 sky130_fd_sc_hd__xor2_1 _457_ (.A(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_34.s_currentState ),
    .B(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_13.input2 ),
    .X(_255_));
 sky130_fd_sc_hd__or4_1 _458_ (.A(_249_),
    .B(_253_),
    .C(_254_),
    .D(_255_),
    .X(_256_));
 sky130_fd_sc_hd__nand2_1 _459_ (.A(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_32.s_currentState ),
    .B(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_11.input2 ),
    .Y(_257_));
 sky130_fd_sc_hd__or2_1 _460_ (.A(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_32.s_currentState ),
    .B(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_11.input2 ),
    .X(_258_));
 sky130_fd_sc_hd__a221o_1 _461_ (.A1(_246_),
    .A2(_247_),
    .B1(_257_),
    .B2(_258_),
    .C1(_251_),
    .X(_259_));
 sky130_fd_sc_hd__xor2_1 _462_ (.A(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_37.s_currentState ),
    .B(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_16.input2 ),
    .X(_260_));
 sky130_fd_sc_hd__or4_1 _463_ (.A(_248_),
    .B(_250_),
    .C(_252_),
    .D(_260_),
    .X(_261_));
 sky130_fd_sc_hd__nor3_2 _464_ (.A(_256_),
    .B(_259_),
    .C(_261_),
    .Y(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_27.result ));
 sky130_fd_sc_hd__nand2_2 _465_ (.A(_181_),
    .B(_201_),
    .Y(_262_));
 sky130_fd_sc_hd__a22o_1 _466_ (.A1(_181_),
    .A2(_201_),
    .B1(_243_),
    .B2(\CIRCUIT_2223.GATES_1.input1[1] ),
    .X(_263_));
 sky130_fd_sc_hd__a22o_2 _467_ (.A1(clknet_1_0__leaf__183_),
    .A2(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_27.result ),
    .B1(_263_),
    .B2(net28),
    .X(_264_));
 sky130_fd_sc_hd__xor2_2 _468_ (.A(net22),
    .B(clknet_1_1__leaf__264_),
    .X(_028_));
 sky130_fd_sc_hd__and4_2 _469_ (.A(\CIRCUIT_2223.s_logisimNet48 ),
    .B(\CIRCUIT_2223.GATES_5.input2 ),
    .C(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_39.s_currentState ),
    .D(\CIRCUIT_2223.GATES_4.input1[0] ),
    .X(_265_));
 sky130_fd_sc_hd__a22o_1 _470_ (.A1(\CIRCUIT_2223.GATES_5.input2 ),
    .A2(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_42.s_currentState ),
    .B1(\CIRCUIT_2223.GATES_4.input1[1] ),
    .B2(\CIRCUIT_2223.s_logisimNet48 ),
    .X(_266_));
 sky130_fd_sc_hd__nand4_1 _471_ (.A(\CIRCUIT_2223.s_logisimNet48 ),
    .B(\CIRCUIT_2223.GATES_5.input2 ),
    .C(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_42.s_currentState ),
    .D(\CIRCUIT_2223.GATES_4.input1[1] ),
    .Y(_267_));
 sky130_fd_sc_hd__nand2_1 _472_ (.A(_266_),
    .B(_267_),
    .Y(_268_));
 sky130_fd_sc_hd__xnor2_1 _473_ (.A(_265_),
    .B(_268_),
    .Y(net9));
 sky130_fd_sc_hd__and4_1 _474_ (.A(\CIRCUIT_2223.s_logisimNet48 ),
    .B(\CIRCUIT_2223.GATES_5.input2 ),
    .C(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_41.s_currentState ),
    .D(\CIRCUIT_2223.GATES_4.input1[2] ),
    .X(_269_));
 sky130_fd_sc_hd__a22oi_1 _475_ (.A1(\CIRCUIT_2223.GATES_5.input2 ),
    .A2(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_41.s_currentState ),
    .B1(\CIRCUIT_2223.GATES_4.input1[2] ),
    .B2(\CIRCUIT_2223.s_logisimNet48 ),
    .Y(_270_));
 sky130_fd_sc_hd__or2_1 _476_ (.A(_269_),
    .B(_270_),
    .X(_271_));
 sky130_fd_sc_hd__a21bo_1 _477_ (.A1(_265_),
    .A2(_266_),
    .B1_N(_267_),
    .X(_272_));
 sky130_fd_sc_hd__and2b_1 _478_ (.A_N(_271_),
    .B(_272_),
    .X(_273_));
 sky130_fd_sc_hd__xnor2_1 _479_ (.A(_271_),
    .B(_272_),
    .Y(net10));
 sky130_fd_sc_hd__and4_1 _480_ (.A(\CIRCUIT_2223.s_logisimNet48 ),
    .B(\CIRCUIT_2223.GATES_5.input2 ),
    .C(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_40.s_currentState ),
    .D(\CIRCUIT_2223.GATES_4.input1[3] ),
    .X(_274_));
 sky130_fd_sc_hd__a22o_1 _481_ (.A1(\CIRCUIT_2223.GATES_5.input2 ),
    .A2(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_40.s_currentState ),
    .B1(\CIRCUIT_2223.GATES_4.input1[3] ),
    .B2(\CIRCUIT_2223.s_logisimNet48 ),
    .X(_275_));
 sky130_fd_sc_hd__and2b_1 _482_ (.A_N(_274_),
    .B(_275_),
    .X(_276_));
 sky130_fd_sc_hd__nor2_1 _483_ (.A(_269_),
    .B(_273_),
    .Y(_277_));
 sky130_fd_sc_hd__xnor2_1 _484_ (.A(_276_),
    .B(_277_),
    .Y(net11));
 sky130_fd_sc_hd__a22oi_2 _485_ (.A1(\CIRCUIT_2223.GATES_3.input2 ),
    .A2(\CIRCUIT_2223.tone_generator_2_1.MEMORY_39.s_currentState ),
    .B1(\CIRCUIT_2223.tone_generator_2_2.MEMORY_39.s_currentState ),
    .B2(\CIRCUIT_2223.GATES_2.input2 ),
    .Y(_278_));
 sky130_fd_sc_hd__and4_1 _486_ (.A(\CIRCUIT_2223.GATES_3.input2 ),
    .B(\CIRCUIT_2223.GATES_2.input2 ),
    .C(\CIRCUIT_2223.tone_generator_2_1.MEMORY_39.s_currentState ),
    .D(\CIRCUIT_2223.tone_generator_2_2.MEMORY_39.s_currentState ),
    .X(_279_));
 sky130_fd_sc_hd__nor2_1 _487_ (.A(_278_),
    .B(_279_),
    .Y(_280_));
 sky130_fd_sc_hd__o31a_2 _488_ (.A1(_269_),
    .A2(_273_),
    .A3(_274_),
    .B1(_275_),
    .X(_281_));
 sky130_fd_sc_hd__xor2_1 _489_ (.A(_280_),
    .B(_281_),
    .X(net12));
 sky130_fd_sc_hd__a21o_1 _490_ (.A1(_280_),
    .A2(_281_),
    .B1(_279_),
    .X(net13));
 sky130_fd_sc_hd__a22oi_2 _491_ (.A1(\CIRCUIT_2223.GATES_5.input2 ),
    .A2(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_39.s_currentState ),
    .B1(\CIRCUIT_2223.GATES_4.input1[0] ),
    .B2(\CIRCUIT_2223.s_logisimNet48 ),
    .Y(_282_));
 sky130_fd_sc_hd__nor2_1 _492_ (.A(_265_),
    .B(_282_),
    .Y(net8));
 sky130_fd_sc_hd__xor2_1 _493_ (.A(\CIRCUIT_2223.tone_generator_1.MEMORY_20.s_currentState ),
    .B(\CIRCUIT_2223.tone_generator_1.MEMORY_6.s_currentState ),
    .X(\CIRCUIT_2223.tone_generator_1.GATES_1.result ));
 sky130_fd_sc_hd__xor2_1 _494_ (.A(\CIRCUIT_2223.tone_generator_1.MEMORY_20.s_currentState ),
    .B(\CIRCUIT_2223.tone_generator_1.MEMORY_7.s_currentState ),
    .X(\CIRCUIT_2223.tone_generator_1.GATES_2.result ));
 sky130_fd_sc_hd__xor2_1 _495_ (.A(\CIRCUIT_2223.tone_generator_1.MEMORY_20.s_currentState ),
    .B(\CIRCUIT_2223.tone_generator_1.MEMORY_9.s_currentState ),
    .X(\CIRCUIT_2223.tone_generator_1.GATES_3.result ));
 sky130_fd_sc_hd__and4_4 _496_ (.A(net2),
    .B(net1),
    .C(\CIRCUIT_2223.GATES_1.input1[0] ),
    .D(_179_),
    .X(_283_));
 sky130_fd_sc_hd__nand2_2 _497_ (.A(_243_),
    .B(_283_),
    .Y(_284_));
 sky130_fd_sc_hd__mux2_1 _498_ (.A0(net37),
    .A1(\CIRCUIT_2223.triangle_wave_generator_1.GATES_8.input2 ),
    .S(_284_),
    .X(_119_));
 sky130_fd_sc_hd__mux2_1 _499_ (.A0(net36),
    .A1(\CIRCUIT_2223.triangle_wave_generator_1.GATES_9.input2 ),
    .S(_284_),
    .X(_120_));
 sky130_fd_sc_hd__mux2_1 _500_ (.A0(net35),
    .A1(\CIRCUIT_2223.triangle_wave_generator_1.GATES_10.input2 ),
    .S(_284_),
    .X(_121_));
 sky130_fd_sc_hd__nor2_1 _501_ (.A(\slow_clock[0] ),
    .B(net34),
    .Y(_122_));
 sky130_fd_sc_hd__a21oi_1 _502_ (.A1(\slow_clock[0] ),
    .A2(\slow_clock[1] ),
    .B1(net34),
    .Y(_285_));
 sky130_fd_sc_hd__o21a_1 _503_ (.A1(\slow_clock[0] ),
    .A2(\slow_clock[1] ),
    .B1(_285_),
    .X(_123_));
 sky130_fd_sc_hd__a21oi_1 _504_ (.A1(\slow_clock[0] ),
    .A2(\slow_clock[1] ),
    .B1(\slow_clock[2] ),
    .Y(_286_));
 sky130_fd_sc_hd__and3_1 _505_ (.A(\slow_clock[0] ),
    .B(\slow_clock[1] ),
    .C(\slow_clock[2] ),
    .X(_287_));
 sky130_fd_sc_hd__nor3_1 _506_ (.A(net34),
    .B(_286_),
    .C(_287_),
    .Y(_124_));
 sky130_fd_sc_hd__and4_1 _507_ (.A(\slow_clock[0] ),
    .B(\slow_clock[1] ),
    .C(\slow_clock[2] ),
    .D(\slow_clock[3] ),
    .X(_288_));
 sky130_fd_sc_hd__nor2_1 _508_ (.A(net34),
    .B(_288_),
    .Y(_289_));
 sky130_fd_sc_hd__o21a_1 _509_ (.A1(\slow_clock[3] ),
    .A2(_287_),
    .B1(_289_),
    .X(_125_));
 sky130_fd_sc_hd__and2_1 _510_ (.A(\slow_clock[4] ),
    .B(_288_),
    .X(_290_));
 sky130_fd_sc_hd__nor2_1 _511_ (.A(net34),
    .B(_290_),
    .Y(_291_));
 sky130_fd_sc_hd__o21a_1 _512_ (.A1(\slow_clock[4] ),
    .A2(_288_),
    .B1(_291_),
    .X(_126_));
 sky130_fd_sc_hd__and3_1 _513_ (.A(\slow_clock[4] ),
    .B(\slow_clock[5] ),
    .C(_288_),
    .X(_292_));
 sky130_fd_sc_hd__nor2_1 _514_ (.A(net34),
    .B(_292_),
    .Y(_293_));
 sky130_fd_sc_hd__o21a_1 _515_ (.A1(\slow_clock[5] ),
    .A2(_290_),
    .B1(_293_),
    .X(_127_));
 sky130_fd_sc_hd__and2_1 _516_ (.A(\slow_clock[6] ),
    .B(_292_),
    .X(_294_));
 sky130_fd_sc_hd__nor2_1 _517_ (.A(net34),
    .B(_294_),
    .Y(_295_));
 sky130_fd_sc_hd__o21a_1 _518_ (.A1(\slow_clock[6] ),
    .A2(_292_),
    .B1(_295_),
    .X(_128_));
 sky130_fd_sc_hd__a21oi_1 _519_ (.A1(net25),
    .A2(_294_),
    .B1(net34),
    .Y(_296_));
 sky130_fd_sc_hd__o21a_1 _520_ (.A1(net25),
    .A2(_294_),
    .B1(_296_),
    .X(_129_));
 sky130_fd_sc_hd__nand2_2 _521_ (.A(_180_),
    .B(_243_),
    .Y(_297_));
 sky130_fd_sc_hd__mux2_1 _522_ (.A0(net37),
    .A1(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_15.input2 ),
    .S(_297_),
    .X(_130_));
 sky130_fd_sc_hd__mux2_1 _523_ (.A0(net36),
    .A1(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_16.input2 ),
    .S(_297_),
    .X(_131_));
 sky130_fd_sc_hd__mux2_1 _524_ (.A0(net35),
    .A1(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_17.input2 ),
    .S(_297_),
    .X(_132_));
 sky130_fd_sc_hd__mux2_1 _525_ (.A0(net6),
    .A1(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_7.input2 ),
    .S(_297_),
    .X(_133_));
 sky130_fd_sc_hd__and4b_4 _526_ (.A_N(\CIRCUIT_2223.GATES_1.input1[0] ),
    .B(\CIRCUIT_2223.GATES_1.input1[1] ),
    .C(net2),
    .D(net1),
    .X(_298_));
 sky130_fd_sc_hd__nand2_2 _527_ (.A(_243_),
    .B(_298_),
    .Y(_299_));
 sky130_fd_sc_hd__mux2_1 _528_ (.A0(net37),
    .A1(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_11.input2 ),
    .S(_299_),
    .X(_134_));
 sky130_fd_sc_hd__mux2_1 _529_ (.A0(net36),
    .A1(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_12.input2 ),
    .S(_299_),
    .X(_135_));
 sky130_fd_sc_hd__mux2_1 _530_ (.A0(net35),
    .A1(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_13.input2 ),
    .S(_299_),
    .X(_136_));
 sky130_fd_sc_hd__mux2_1 _531_ (.A0(net6),
    .A1(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_14.input2 ),
    .S(_299_),
    .X(_137_));
 sky130_fd_sc_hd__nand2b_2 _532_ (.A_N(net1),
    .B(net2),
    .Y(_300_));
 sky130_fd_sc_hd__mux2_1 _533_ (.A0(net37),
    .A1(\CIRCUIT_2223.GATES_1.input1[0] ),
    .S(_300_),
    .X(_138_));
 sky130_fd_sc_hd__mux2_1 _534_ (.A0(net36),
    .A1(\CIRCUIT_2223.GATES_1.input1[1] ),
    .S(_300_),
    .X(_139_));
 sky130_fd_sc_hd__mux2_1 _535_ (.A0(net35),
    .A1(\CIRCUIT_2223.GATES_1.input1[2] ),
    .S(_300_),
    .X(_140_));
 sky130_fd_sc_hd__mux2_1 _536_ (.A0(net6),
    .A1(\CIRCUIT_2223.GATES_1.input1[3] ),
    .S(_300_),
    .X(_141_));
 sky130_fd_sc_hd__nand2_2 _537_ (.A(_180_),
    .B(_200_),
    .Y(_301_));
 sky130_fd_sc_hd__mux2_1 _538_ (.A0(net37),
    .A1(\CIRCUIT_2223.tone_generator_2_2.GATES_8.input2 ),
    .S(_301_),
    .X(_142_));
 sky130_fd_sc_hd__mux2_1 _539_ (.A0(net36),
    .A1(\CIRCUIT_2223.tone_generator_2_2.GATES_9.input2 ),
    .S(_301_),
    .X(_143_));
 sky130_fd_sc_hd__mux2_1 _540_ (.A0(net35),
    .A1(\CIRCUIT_2223.tone_generator_2_2.GATES_10.input2 ),
    .S(_301_),
    .X(_144_));
 sky130_fd_sc_hd__mux2_1 _541_ (.A0(net37),
    .A1(\CIRCUIT_2223.triangle_wave_generator_1.GATES_11.input2 ),
    .S(_242_),
    .X(_145_));
 sky130_fd_sc_hd__mux2_1 _542_ (.A0(net36),
    .A1(\CIRCUIT_2223.triangle_wave_generator_1.GATES_12.input2 ),
    .S(_242_),
    .X(_146_));
 sky130_fd_sc_hd__mux2_1 _543_ (.A0(net35),
    .A1(\CIRCUIT_2223.triangle_wave_generator_1.GATES_13.input2 ),
    .S(_242_),
    .X(_147_));
 sky130_fd_sc_hd__mux2_1 _544_ (.A0(net6),
    .A1(\CIRCUIT_2223.triangle_wave_generator_1.GATES_14.input2 ),
    .S(_242_),
    .X(_148_));
 sky130_fd_sc_hd__nand2_4 _545_ (.A(_201_),
    .B(_243_),
    .Y(_302_));
 sky130_fd_sc_hd__mux2_1 _546_ (.A0(net37),
    .A1(\CIRCUIT_2223.triangle_wave_generator_1.GATES_15.input2 ),
    .S(_302_),
    .X(_149_));
 sky130_fd_sc_hd__mux2_1 _547_ (.A0(net36),
    .A1(\CIRCUIT_2223.triangle_wave_generator_1.GATES_16.input2 ),
    .S(_302_),
    .X(_150_));
 sky130_fd_sc_hd__mux2_1 _548_ (.A0(net35),
    .A1(\CIRCUIT_2223.triangle_wave_generator_1.GATES_17.input2 ),
    .S(_302_),
    .X(_151_));
 sky130_fd_sc_hd__mux2_1 _549_ (.A0(net6),
    .A1(\CIRCUIT_2223.triangle_wave_generator_1.GATES_7.input2 ),
    .S(_302_),
    .X(_152_));
 sky130_fd_sc_hd__mux2_1 _550_ (.A0(net37),
    .A1(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_8.input2 ),
    .S(_262_),
    .X(_153_));
 sky130_fd_sc_hd__mux2_1 _551_ (.A0(net36),
    .A1(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_9.input2 ),
    .S(_262_),
    .X(_154_));
 sky130_fd_sc_hd__mux2_1 _552_ (.A0(net5),
    .A1(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_10.input2 ),
    .S(_262_),
    .X(_155_));
 sky130_fd_sc_hd__nand2_2 _553_ (.A(_201_),
    .B(_220_),
    .Y(_303_));
 sky130_fd_sc_hd__mux2_1 _554_ (.A0(net37),
    .A1(\CIRCUIT_2223.tone_generator_2_1.GATES_11.input2 ),
    .S(_303_),
    .X(_156_));
 sky130_fd_sc_hd__mux2_1 _555_ (.A0(net36),
    .A1(\CIRCUIT_2223.tone_generator_2_1.GATES_12.input2 ),
    .S(_303_),
    .X(_157_));
 sky130_fd_sc_hd__mux2_1 _556_ (.A0(net5),
    .A1(\CIRCUIT_2223.tone_generator_2_1.GATES_13.input2 ),
    .S(_303_),
    .X(_158_));
 sky130_fd_sc_hd__mux2_1 _557_ (.A0(net6),
    .A1(\CIRCUIT_2223.tone_generator_2_1.GATES_14.input2 ),
    .S(_303_),
    .X(_159_));
 sky130_fd_sc_hd__nand2_4 _558_ (.A(_220_),
    .B(_283_),
    .Y(_304_));
 sky130_fd_sc_hd__mux2_1 _559_ (.A0(net38),
    .A1(\CIRCUIT_2223.tone_generator_2_1.GATES_15.input2 ),
    .S(_304_),
    .X(_160_));
 sky130_fd_sc_hd__mux2_1 _560_ (.A0(net4),
    .A1(\CIRCUIT_2223.tone_generator_2_1.GATES_16.input2 ),
    .S(_304_),
    .X(_161_));
 sky130_fd_sc_hd__mux2_1 _561_ (.A0(net5),
    .A1(\CIRCUIT_2223.tone_generator_2_1.GATES_17.input2 ),
    .S(_304_),
    .X(_162_));
 sky130_fd_sc_hd__mux2_1 _562_ (.A0(net6),
    .A1(\CIRCUIT_2223.tone_generator_2_1.GATES_7.input2 ),
    .S(_304_),
    .X(_163_));
 sky130_fd_sc_hd__nand2_2 _563_ (.A(_220_),
    .B(_298_),
    .Y(_305_));
 sky130_fd_sc_hd__mux2_1 _564_ (.A0(net38),
    .A1(\CIRCUIT_2223.tone_generator_2_1.GATES_8.input2 ),
    .S(_305_),
    .X(_164_));
 sky130_fd_sc_hd__mux2_1 _565_ (.A0(net4),
    .A1(\CIRCUIT_2223.tone_generator_2_1.GATES_9.input2 ),
    .S(_305_),
    .X(_165_));
 sky130_fd_sc_hd__mux2_1 _566_ (.A0(net5),
    .A1(\CIRCUIT_2223.tone_generator_2_1.GATES_10.input2 ),
    .S(_305_),
    .X(_166_));
 sky130_fd_sc_hd__nand2_2 _567_ (.A(_200_),
    .B(_283_),
    .Y(_306_));
 sky130_fd_sc_hd__mux2_1 _568_ (.A0(net38),
    .A1(\CIRCUIT_2223.tone_generator_2_2.GATES_11.input2 ),
    .S(_306_),
    .X(_167_));
 sky130_fd_sc_hd__mux2_1 _569_ (.A0(net4),
    .A1(\CIRCUIT_2223.tone_generator_2_2.GATES_12.input2 ),
    .S(_306_),
    .X(_168_));
 sky130_fd_sc_hd__mux2_1 _570_ (.A0(net35),
    .A1(\CIRCUIT_2223.tone_generator_2_2.GATES_13.input2 ),
    .S(_306_),
    .X(_169_));
 sky130_fd_sc_hd__mux2_1 _571_ (.A0(net6),
    .A1(\CIRCUIT_2223.tone_generator_2_2.GATES_14.input2 ),
    .S(_306_),
    .X(_170_));
 sky130_fd_sc_hd__nand2_4 _572_ (.A(_200_),
    .B(_298_),
    .Y(_307_));
 sky130_fd_sc_hd__mux2_1 _573_ (.A0(net38),
    .A1(\CIRCUIT_2223.tone_generator_2_2.GATES_15.input2 ),
    .S(_307_),
    .X(_171_));
 sky130_fd_sc_hd__mux2_1 _574_ (.A0(net4),
    .A1(\CIRCUIT_2223.tone_generator_2_2.GATES_16.input2 ),
    .S(_307_),
    .X(_172_));
 sky130_fd_sc_hd__mux2_1 _575_ (.A0(net35),
    .A1(\CIRCUIT_2223.tone_generator_2_2.GATES_17.input2 ),
    .S(_307_),
    .X(_173_));
 sky130_fd_sc_hd__mux2_1 _576_ (.A0(net6),
    .A1(\CIRCUIT_2223.tone_generator_2_2.GATES_7.input2 ),
    .S(_307_),
    .X(_174_));
 sky130_fd_sc_hd__and2_1 _577_ (.A(_181_),
    .B(_298_),
    .X(_096_));
 sky130_fd_sc_hd__and2_1 _578_ (.A(_181_),
    .B(_283_),
    .X(_097_));
 sky130_fd_sc_hd__inv_2 _579_ (.A(net23),
    .Y(_115_));
 sky130_fd_sc_hd__inv_2 _580_ (.A(net23),
    .Y(_113_));
 sky130_fd_sc_hd__inv_2 _581_ (.A(net25),
    .Y(_111_));
 sky130_fd_sc_hd__inv_2 _582_ (.A(net25),
    .Y(_109_));
 sky130_fd_sc_hd__inv_2 _583_ (.A(net25),
    .Y(_107_));
 sky130_fd_sc_hd__inv_2 _584_ (.A(net23),
    .Y(_104_));
 sky130_fd_sc_hd__inv_2 _585_ (.A(net23),
    .Y(_102_));
 sky130_fd_sc_hd__xor2_2 _586_ (.A(net19),
    .B(clknet_1_1__leaf__203_),
    .X(_092_));
 sky130_fd_sc_hd__xor2_2 _587_ (.A(net19),
    .B(clknet_1_0__leaf__203_),
    .X(_090_));
 sky130_fd_sc_hd__xor2_2 _588_ (.A(net19),
    .B(clknet_1_0__leaf__203_),
    .X(_088_));
 sky130_fd_sc_hd__xor2_2 _589_ (.A(net19),
    .B(clknet_1_0__leaf__203_),
    .X(_086_));
 sky130_fd_sc_hd__xor2_2 _590_ (.A(net19),
    .B(clknet_1_0__leaf__203_),
    .X(_084_));
 sky130_fd_sc_hd__xor2_2 _591_ (.A(net19),
    .B(clknet_1_1__leaf__203_),
    .X(_081_));
 sky130_fd_sc_hd__xor2_2 _592_ (.A(net19),
    .B(clknet_1_1__leaf__203_),
    .X(_079_));
 sky130_fd_sc_hd__xor2_2 _593_ (.A(net19),
    .B(clknet_1_1__leaf__203_),
    .X(_077_));
 sky130_fd_sc_hd__xor2_2 _594_ (.A(net20),
    .B(clknet_1_1__leaf__203_),
    .X(_075_));
 sky130_fd_sc_hd__xnor2_2 _595_ (.A(net21),
    .B(clknet_1_1__leaf__222_),
    .Y(_071_));
 sky130_fd_sc_hd__xnor2_2 _596_ (.A(net21),
    .B(clknet_1_1__leaf__222_),
    .Y(_069_));
 sky130_fd_sc_hd__xnor2_2 _597_ (.A(net21),
    .B(clknet_1_1__leaf__222_),
    .Y(_067_));
 sky130_fd_sc_hd__xnor2_2 _598_ (.A(net21),
    .B(clknet_1_1__leaf__222_),
    .Y(_065_));
 sky130_fd_sc_hd__xnor2_2 _599_ (.A(_000_),
    .B(clknet_1_1__leaf__222_),
    .Y(_063_));
 sky130_fd_sc_hd__xnor2_2 _600_ (.A(net21),
    .B(clknet_1_0__leaf__222_),
    .Y(_060_));
 sky130_fd_sc_hd__xnor2_2 _601_ (.A(net21),
    .B(clknet_1_0__leaf__222_),
    .Y(_058_));
 sky130_fd_sc_hd__xnor2_2 _602_ (.A(net21),
    .B(clknet_1_0__leaf__222_),
    .Y(_056_));
 sky130_fd_sc_hd__xnor2_2 _603_ (.A(net21),
    .B(clknet_1_0__leaf__222_),
    .Y(_054_));
 sky130_fd_sc_hd__xnor2_2 _604_ (.A(net18),
    .B(clknet_1_0__leaf__245_),
    .Y(_047_));
 sky130_fd_sc_hd__xnor2_2 _605_ (.A(net18),
    .B(clknet_1_0__leaf__245_),
    .Y(_045_));
 sky130_fd_sc_hd__xnor2_2 _606_ (.A(net18),
    .B(clknet_1_0__leaf__245_),
    .Y(_043_));
 sky130_fd_sc_hd__xnor2_2 _607_ (.A(net18),
    .B(clknet_1_0__leaf__245_),
    .Y(_041_));
 sky130_fd_sc_hd__xnor2_2 _608_ (.A(net20),
    .B(clknet_1_0__leaf__245_),
    .Y(_039_));
 sky130_fd_sc_hd__xnor2_2 _609_ (.A(net18),
    .B(clknet_1_1__leaf__245_),
    .Y(_036_));
 sky130_fd_sc_hd__xnor2_2 _610_ (.A(net18),
    .B(clknet_1_1__leaf__245_),
    .Y(_034_));
 sky130_fd_sc_hd__xnor2_2 _611_ (.A(net18),
    .B(clknet_1_1__leaf__245_),
    .Y(_032_));
 sky130_fd_sc_hd__xnor2_2 _612_ (.A(net18),
    .B(clknet_1_1__leaf__245_),
    .Y(_030_));
 sky130_fd_sc_hd__xor2_2 _613_ (.A(net22),
    .B(clknet_1_1__leaf__264_),
    .X(_026_));
 sky130_fd_sc_hd__xor2_2 _614_ (.A(net22),
    .B(clknet_1_1__leaf__264_),
    .X(_024_));
 sky130_fd_sc_hd__xor2_2 _615_ (.A(net22),
    .B(clknet_1_1__leaf__264_),
    .X(_022_));
 sky130_fd_sc_hd__xor2_2 _616_ (.A(net20),
    .B(clknet_1_0__leaf__264_),
    .X(_019_));
 sky130_fd_sc_hd__xor2_2 _617_ (.A(net22),
    .B(clknet_1_0__leaf__264_),
    .X(_017_));
 sky130_fd_sc_hd__xor2_2 _618_ (.A(net22),
    .B(clknet_1_0__leaf__264_),
    .X(_015_));
 sky130_fd_sc_hd__xor2_2 _619_ (.A(net22),
    .B(clknet_1_0__leaf__264_),
    .X(_013_));
 sky130_fd_sc_hd__xor2_2 _620_ (.A(net22),
    .B(clknet_1_1__leaf__264_),
    .X(_011_));
 sky130_fd_sc_hd__xor2_2 _621_ (.A(net22),
    .B(clknet_1_1__leaf__264_),
    .X(_009_));
 sky130_fd_sc_hd__nand2_1 _622_ (.A(net28),
    .B(net33),
    .Y(_001_));
 sky130_fd_sc_hd__nand2_1 _623_ (.A(net28),
    .B(net33),
    .Y(_002_));
 sky130_fd_sc_hd__nand2_1 _624_ (.A(net28),
    .B(net33),
    .Y(_003_));
 sky130_fd_sc_hd__nand2_1 _625_ (.A(net27),
    .B(net33),
    .Y(_004_));
 sky130_fd_sc_hd__nand2_1 _626_ (.A(net27),
    .B(net33),
    .Y(_005_));
 sky130_fd_sc_hd__nand2_1 _627_ (.A(net27),
    .B(net33),
    .Y(_006_));
 sky130_fd_sc_hd__nand2_1 _628_ (.A(net27),
    .B(net33),
    .Y(_007_));
 sky130_fd_sc_hd__nand2_1 _629_ (.A(net27),
    .B(net33),
    .Y(_008_));
 sky130_fd_sc_hd__inv_2 _630_ (.A(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_37.s_currentState ),
    .Y(_010_));
 sky130_fd_sc_hd__inv_2 _631_ (.A(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_36.s_currentState ),
    .Y(_012_));
 sky130_fd_sc_hd__inv_2 _632_ (.A(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_35.s_currentState ),
    .Y(_014_));
 sky130_fd_sc_hd__inv_2 _633_ (.A(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_34.s_currentState ),
    .Y(_016_));
 sky130_fd_sc_hd__inv_2 _634_ (.A(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_33.s_currentState ),
    .Y(_018_));
 sky130_fd_sc_hd__inv_2 _635_ (.A(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_32.s_currentState ),
    .Y(_020_));
 sky130_fd_sc_hd__xor2_2 _636_ (.A(net20),
    .B(clknet_1_0__leaf__264_),
    .X(_021_));
 sky130_fd_sc_hd__inv_2 _637_ (.A(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_30.s_currentState ),
    .Y(_023_));
 sky130_fd_sc_hd__inv_2 _638_ (.A(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_29.s_currentState ),
    .Y(_025_));
 sky130_fd_sc_hd__inv_2 _639_ (.A(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_28.s_currentState ),
    .Y(_027_));
 sky130_fd_sc_hd__inv_2 _640_ (.A(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_38.s_currentState ),
    .Y(_029_));
 sky130_fd_sc_hd__inv_2 _641_ (.A(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_38.s_currentState ),
    .Y(_031_));
 sky130_fd_sc_hd__inv_2 _642_ (.A(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_28.s_currentState ),
    .Y(_033_));
 sky130_fd_sc_hd__inv_2 _643_ (.A(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_29.s_currentState ),
    .Y(_035_));
 sky130_fd_sc_hd__inv_2 _644_ (.A(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_30.s_currentState ),
    .Y(_037_));
 sky130_fd_sc_hd__xnor2_2 _645_ (.A(net20),
    .B(clknet_1_0__leaf__245_),
    .Y(_038_));
 sky130_fd_sc_hd__inv_2 _646_ (.A(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_32.s_currentState ),
    .Y(_040_));
 sky130_fd_sc_hd__inv_2 _647_ (.A(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_33.s_currentState ),
    .Y(_042_));
 sky130_fd_sc_hd__inv_2 _648_ (.A(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_34.s_currentState ),
    .Y(_044_));
 sky130_fd_sc_hd__inv_2 _649_ (.A(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_35.s_currentState ),
    .Y(_046_));
 sky130_fd_sc_hd__inv_2 _650_ (.A(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_36.s_currentState ),
    .Y(_048_));
 sky130_fd_sc_hd__inv_2 _651_ (.A(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_37.s_currentState ),
    .Y(_050_));
 sky130_fd_sc_hd__inv_2 _652_ (.A(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_41.s_currentState ),
    .Y(_051_));
 sky130_fd_sc_hd__inv_2 _653_ (.A(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_42.s_currentState ),
    .Y(_052_));
 sky130_fd_sc_hd__inv_2 _654_ (.A(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_39.s_currentState ),
    .Y(_053_));
 sky130_fd_sc_hd__inv_2 _655_ (.A(\CIRCUIT_2223.tone_generator_2_1.MEMORY_38.s_currentState ),
    .Y(_055_));
 sky130_fd_sc_hd__inv_2 _656_ (.A(\CIRCUIT_2223.tone_generator_2_1.MEMORY_28.s_currentState ),
    .Y(_057_));
 sky130_fd_sc_hd__inv_2 _657_ (.A(\CIRCUIT_2223.tone_generator_2_1.MEMORY_29.s_currentState ),
    .Y(_059_));
 sky130_fd_sc_hd__inv_2 _658_ (.A(\CIRCUIT_2223.tone_generator_2_1.MEMORY_30.s_currentState ),
    .Y(_061_));
 sky130_fd_sc_hd__xnor2_2 _659_ (.A(net21),
    .B(clknet_1_0__leaf__222_),
    .Y(_062_));
 sky130_fd_sc_hd__inv_2 _660_ (.A(\CIRCUIT_2223.tone_generator_2_1.MEMORY_32.s_currentState ),
    .Y(_064_));
 sky130_fd_sc_hd__inv_2 _661_ (.A(\CIRCUIT_2223.tone_generator_2_1.MEMORY_33.s_currentState ),
    .Y(_066_));
 sky130_fd_sc_hd__inv_2 _662_ (.A(\CIRCUIT_2223.tone_generator_2_1.MEMORY_34.s_currentState ),
    .Y(_068_));
 sky130_fd_sc_hd__inv_2 _663_ (.A(\CIRCUIT_2223.tone_generator_2_1.MEMORY_35.s_currentState ),
    .Y(_070_));
 sky130_fd_sc_hd__inv_2 _664_ (.A(\CIRCUIT_2223.tone_generator_2_1.MEMORY_36.s_currentState ),
    .Y(_072_));
 sky130_fd_sc_hd__inv_2 _665_ (.A(\CIRCUIT_2223.tone_generator_2_1.MEMORY_37.s_currentState ),
    .Y(_074_));
 sky130_fd_sc_hd__inv_2 _666_ (.A(\CIRCUIT_2223.tone_generator_2_2.MEMORY_38.s_currentState ),
    .Y(_076_));
 sky130_fd_sc_hd__inv_2 _667_ (.A(\CIRCUIT_2223.tone_generator_2_2.MEMORY_28.s_currentState ),
    .Y(_078_));
 sky130_fd_sc_hd__inv_2 _668_ (.A(\CIRCUIT_2223.tone_generator_2_2.MEMORY_29.s_currentState ),
    .Y(_080_));
 sky130_fd_sc_hd__inv_2 _669_ (.A(\CIRCUIT_2223.tone_generator_2_2.MEMORY_30.s_currentState ),
    .Y(_082_));
 sky130_fd_sc_hd__xor2_2 _670_ (.A(net19),
    .B(clknet_1_0__leaf__203_),
    .X(_083_));
 sky130_fd_sc_hd__inv_2 _671_ (.A(\CIRCUIT_2223.tone_generator_2_2.MEMORY_32.s_currentState ),
    .Y(_085_));
 sky130_fd_sc_hd__inv_2 _672_ (.A(\CIRCUIT_2223.tone_generator_2_2.MEMORY_33.s_currentState ),
    .Y(_087_));
 sky130_fd_sc_hd__inv_2 _673_ (.A(\CIRCUIT_2223.tone_generator_2_2.MEMORY_34.s_currentState ),
    .Y(_089_));
 sky130_fd_sc_hd__inv_2 _674_ (.A(\CIRCUIT_2223.tone_generator_2_2.MEMORY_35.s_currentState ),
    .Y(_091_));
 sky130_fd_sc_hd__inv_2 _675_ (.A(\CIRCUIT_2223.tone_generator_2_2.MEMORY_36.s_currentState ),
    .Y(_093_));
 sky130_fd_sc_hd__inv_2 _676_ (.A(\CIRCUIT_2223.tone_generator_2_2.MEMORY_37.s_currentState ),
    .Y(_095_));
 sky130_fd_sc_hd__nand2_1 _677_ (.A(net29),
    .B(net7),
    .Y(_098_));
 sky130_fd_sc_hd__nand2_1 _678_ (.A(net29),
    .B(net7),
    .Y(_099_));
 sky130_fd_sc_hd__nand2_1 _679_ (.A(net27),
    .B(net33),
    .Y(_100_));
 sky130_fd_sc_hd__nand2_1 _680_ (.A(net27),
    .B(net34),
    .Y(_101_));
 sky130_fd_sc_hd__inv_2 _681_ (.A(\CIRCUIT_2223.MEMORY_25.s_currentState ),
    .Y(_103_));
 sky130_fd_sc_hd__inv_2 _682_ (.A(net16),
    .Y(_105_));
 sky130_fd_sc_hd__inv_2 _683_ (.A(net43),
    .Y(_106_));
 sky130_fd_sc_hd__inv_2 _684_ (.A(\CIRCUIT_2223.MEMORY_22.s_currentState ),
    .Y(_108_));
 sky130_fd_sc_hd__inv_2 _685_ (.A(\CIRCUIT_2223.MEMORY_21.s_currentState ),
    .Y(_110_));
 sky130_fd_sc_hd__inv_2 _686_ (.A(\CIRCUIT_2223.MEMORY_20.s_currentState ),
    .Y(_112_));
 sky130_fd_sc_hd__inv_2 _687_ (.A(\CIRCUIT_2223.MEMORY_19.s_currentState ),
    .Y(_114_));
 sky130_fd_sc_hd__inv_2 _688_ (.A(\CIRCUIT_2223.MEMORY_18.s_currentState ),
    .Y(_116_));
 sky130_fd_sc_hd__inv_2 _689_ (.A(\CIRCUIT_2223.MEMORY_26.s_currentState ),
    .Y(_118_));
 sky130_fd_sc_hd__dfxtp_1 _690_ (.CLK(net23),
    .D(_119_),
    .Q(\CIRCUIT_2223.triangle_wave_generator_1.GATES_8.input2 ));
 sky130_fd_sc_hd__dfxtp_1 _691_ (.CLK(net23),
    .D(_120_),
    .Q(\CIRCUIT_2223.triangle_wave_generator_1.GATES_9.input2 ));
 sky130_fd_sc_hd__dfxtp_1 _692_ (.CLK(net24),
    .D(_121_),
    .Q(\CIRCUIT_2223.triangle_wave_generator_1.GATES_10.input2 ));
 sky130_fd_sc_hd__dfxtp_1 _693_ (.CLK(clknet_1_1__leaf_clk),
    .D(_122_),
    .Q(\slow_clock[0] ));
 sky130_fd_sc_hd__dfxtp_1 _694_ (.CLK(clknet_1_1__leaf_clk),
    .D(_123_),
    .Q(\slow_clock[1] ));
 sky130_fd_sc_hd__dfxtp_1 _695_ (.CLK(clknet_1_1__leaf_clk),
    .D(_124_),
    .Q(\slow_clock[2] ));
 sky130_fd_sc_hd__dfxtp_1 _696_ (.CLK(clknet_1_1__leaf_clk),
    .D(_125_),
    .Q(\slow_clock[3] ));
 sky130_fd_sc_hd__dfxtp_1 _697_ (.CLK(clknet_1_0__leaf_clk),
    .D(_126_),
    .Q(\slow_clock[4] ));
 sky130_fd_sc_hd__dfxtp_1 _698_ (.CLK(clknet_1_0__leaf_clk),
    .D(_127_),
    .Q(\slow_clock[5] ));
 sky130_fd_sc_hd__dfxtp_1 _699_ (.CLK(clknet_1_0__leaf_clk),
    .D(_128_),
    .Q(\slow_clock[6] ));
 sky130_fd_sc_hd__dfxtp_1 _700_ (.CLK(clknet_1_0__leaf_clk),
    .D(_129_),
    .Q(\CIRCUIT_2223.CLK ));
 sky130_fd_sc_hd__dfxtp_1 _701_ (.CLK(\CIRCUIT_2223.MEMORY_24.s_currentState ),
    .D(\CIRCUIT_2223.tone_generator_1.MEMORY_20.s_currentState ),
    .Q(\CIRCUIT_2223.tone_generator_1.MEMORY_4.s_currentState ));
 sky130_fd_sc_hd__dfxtp_1 _702_ (.CLK(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_39.s_currentState ),
    .D(\CIRCUIT_2223.tone_generator_1.MEMORY_20.s_currentState ),
    .Q(\CIRCUIT_2223.GATES_4.input1[0] ));
 sky130_fd_sc_hd__dfxtp_1 _703_ (.CLK(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_39.s_currentState ),
    .D(\CIRCUIT_2223.tone_generator_1.MEMORY_19.s_currentState ),
    .Q(\CIRCUIT_2223.GATES_4.input1[1] ));
 sky130_fd_sc_hd__dfxtp_1 _704_ (.CLK(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_39.s_currentState ),
    .D(\CIRCUIT_2223.tone_generator_1.MEMORY_17.s_currentState ),
    .Q(\CIRCUIT_2223.GATES_4.input1[2] ));
 sky130_fd_sc_hd__dfxtp_1 _705_ (.CLK(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_39.s_currentState ),
    .D(\CIRCUIT_2223.tone_generator_1.MEMORY_14.s_currentState ),
    .Q(\CIRCUIT_2223.GATES_4.input1[3] ));
 sky130_fd_sc_hd__dfxtp_1 _706_ (.CLK(net17),
    .D(\CIRCUIT_2223.tone_generator_1.MEMORY_4.s_currentState ),
    .Q(\CIRCUIT_2223.tone_generator_1.MEMORY_6.s_currentState ));
 sky130_fd_sc_hd__dfxtp_1 _707_ (.CLK(net17),
    .D(\CIRCUIT_2223.tone_generator_1.GATES_1.result ),
    .Q(\CIRCUIT_2223.tone_generator_1.MEMORY_7.s_currentState ));
 sky130_fd_sc_hd__dfxtp_1 _708_ (.CLK(net16),
    .D(\CIRCUIT_2223.tone_generator_1.GATES_2.result ),
    .Q(\CIRCUIT_2223.tone_generator_1.MEMORY_8.s_currentState ));
 sky130_fd_sc_hd__dfxtp_1 _709_ (.CLK(net16),
    .D(\CIRCUIT_2223.tone_generator_1.MEMORY_8.s_currentState ),
    .Q(\CIRCUIT_2223.tone_generator_1.MEMORY_9.s_currentState ));
 sky130_fd_sc_hd__dfxtp_1 _710_ (.CLK(net16),
    .D(\CIRCUIT_2223.tone_generator_1.GATES_3.result ),
    .Q(\CIRCUIT_2223.tone_generator_1.MEMORY_10.s_currentState ));
 sky130_fd_sc_hd__dfxtp_1 _711_ (.CLK(net16),
    .D(\CIRCUIT_2223.tone_generator_1.MEMORY_10.s_currentState ),
    .Q(\CIRCUIT_2223.tone_generator_1.MEMORY_11.s_currentState ));
 sky130_fd_sc_hd__dfstp_1 _712_ (.CLK(net16),
    .D(\CIRCUIT_2223.tone_generator_1.MEMORY_11.s_currentState ),
    .SET_B(net18),
    .Q(\CIRCUIT_2223.tone_generator_1.MEMORY_12.s_currentState ));
 sky130_fd_sc_hd__dfrtp_1 _713_ (.CLK(net16),
    .D(\CIRCUIT_2223.tone_generator_1.MEMORY_12.s_currentState ),
    .RESET_B(_001_),
    .Q(\CIRCUIT_2223.tone_generator_1.MEMORY_13.s_currentState ));
 sky130_fd_sc_hd__dfstp_1 _714_ (.CLK(net16),
    .D(\CIRCUIT_2223.tone_generator_1.MEMORY_13.s_currentState ),
    .SET_B(_002_),
    .Q(\CIRCUIT_2223.tone_generator_1.MEMORY_14.s_currentState ));
 sky130_fd_sc_hd__dfrtp_1 _715_ (.CLK(net17),
    .D(\CIRCUIT_2223.tone_generator_1.MEMORY_14.s_currentState ),
    .RESET_B(_003_),
    .Q(\CIRCUIT_2223.tone_generator_1.MEMORY_15.s_currentState ));
 sky130_fd_sc_hd__dfstp_1 _716_ (.CLK(net17),
    .D(\CIRCUIT_2223.tone_generator_1.MEMORY_15.s_currentState ),
    .SET_B(_004_),
    .Q(\CIRCUIT_2223.tone_generator_1.MEMORY_16.s_currentState ));
 sky130_fd_sc_hd__dfrtp_1 _717_ (.CLK(net17),
    .D(\CIRCUIT_2223.tone_generator_1.MEMORY_16.s_currentState ),
    .RESET_B(_005_),
    .Q(\CIRCUIT_2223.tone_generator_1.MEMORY_17.s_currentState ));
 sky130_fd_sc_hd__dfstp_1 _718_ (.CLK(net17),
    .D(\CIRCUIT_2223.tone_generator_1.MEMORY_17.s_currentState ),
    .SET_B(_006_),
    .Q(\CIRCUIT_2223.tone_generator_1.MEMORY_18.s_currentState ));
 sky130_fd_sc_hd__dfstp_1 _719_ (.CLK(net17),
    .D(\CIRCUIT_2223.tone_generator_1.MEMORY_18.s_currentState ),
    .SET_B(_007_),
    .Q(\CIRCUIT_2223.tone_generator_1.MEMORY_19.s_currentState ));
 sky130_fd_sc_hd__dfrtp_2 _720_ (.CLK(net17),
    .D(\CIRCUIT_2223.tone_generator_1.MEMORY_19.s_currentState ),
    .RESET_B(_008_),
    .Q(\CIRCUIT_2223.tone_generator_1.MEMORY_20.s_currentState ));
 sky130_fd_sc_hd__dfxtp_1 _721_ (.CLK(net31),
    .D(_130_),
    .Q(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_15.input2 ));
 sky130_fd_sc_hd__dfxtp_1 _722_ (.CLK(net27),
    .D(_131_),
    .Q(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_16.input2 ));
 sky130_fd_sc_hd__dfxtp_1 _723_ (.CLK(net28),
    .D(_132_),
    .Q(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_17.input2 ));
 sky130_fd_sc_hd__dfxtp_1 _724_ (.CLK(net31),
    .D(_133_),
    .Q(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_7.input2 ));
 sky130_fd_sc_hd__dfxtp_1 _725_ (.CLK(net28),
    .D(_134_),
    .Q(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_11.input2 ));
 sky130_fd_sc_hd__dfxtp_1 _726_ (.CLK(net28),
    .D(_135_),
    .Q(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_12.input2 ));
 sky130_fd_sc_hd__dfxtp_1 _727_ (.CLK(net28),
    .D(_136_),
    .Q(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_13.input2 ));
 sky130_fd_sc_hd__dfxtp_1 _728_ (.CLK(net28),
    .D(_137_),
    .Q(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_14.input2 ));
 sky130_fd_sc_hd__dfxtp_2 _729_ (.CLK(net24),
    .D(_138_),
    .Q(\CIRCUIT_2223.GATES_1.input1[0] ));
 sky130_fd_sc_hd__dfxtp_4 _730_ (.CLK(net24),
    .D(_139_),
    .Q(\CIRCUIT_2223.GATES_1.input1[1] ));
 sky130_fd_sc_hd__dfxtp_2 _731_ (.CLK(net26),
    .D(_140_),
    .Q(\CIRCUIT_2223.GATES_1.input1[2] ));
 sky130_fd_sc_hd__dfxtp_2 _732_ (.CLK(net26),
    .D(_141_),
    .Q(\CIRCUIT_2223.GATES_1.input1[3] ));
 sky130_fd_sc_hd__dfxtp_2 _733_ (.CLK(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_27.result ),
    .D(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_39.d ),
    .Q(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_39.s_currentState ));
 sky130_fd_sc_hd__dfrtp_2 _734_ (.CLK(_010_),
    .D(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_28.clock ),
    .RESET_B(_009_),
    .Q(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_38.s_currentState ));
 sky130_fd_sc_hd__dfrtp_2 _735_ (.CLK(_012_),
    .D(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_37.d ),
    .RESET_B(_011_),
    .Q(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_37.s_currentState ));
 sky130_fd_sc_hd__dfrtp_2 _736_ (.CLK(_014_),
    .D(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_36.d ),
    .RESET_B(_013_),
    .Q(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_36.s_currentState ));
 sky130_fd_sc_hd__dfrtp_2 _737_ (.CLK(_016_),
    .D(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_35.d ),
    .RESET_B(_015_),
    .Q(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_35.s_currentState ));
 sky130_fd_sc_hd__dfrtp_2 _738_ (.CLK(_018_),
    .D(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_34.d ),
    .RESET_B(_017_),
    .Q(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_34.s_currentState ));
 sky130_fd_sc_hd__dfrtp_2 _739_ (.CLK(_020_),
    .D(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_33.d ),
    .RESET_B(_019_),
    .Q(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_33.s_currentState ));
 sky130_fd_sc_hd__dfrtp_2 _740_ (.CLK(net16),
    .D(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_32.d ),
    .RESET_B(_021_),
    .Q(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_32.s_currentState ));
 sky130_fd_sc_hd__dfrtp_4 _741_ (.CLK(_023_),
    .D(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_31.d ),
    .RESET_B(_022_),
    .Q(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_31.s_currentState ));
 sky130_fd_sc_hd__dfrtp_2 _742_ (.CLK(_025_),
    .D(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_30.d ),
    .RESET_B(_024_),
    .Q(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_30.s_currentState ));
 sky130_fd_sc_hd__dfrtp_2 _743_ (.CLK(_027_),
    .D(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_29.d ),
    .RESET_B(_026_),
    .Q(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_29.s_currentState ));
 sky130_fd_sc_hd__dfrtp_2 _744_ (.CLK(_029_),
    .D(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_28.d ),
    .RESET_B(_028_),
    .Q(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_28.s_currentState ));
 sky130_fd_sc_hd__dfrtp_2 _745_ (.CLK(_031_),
    .D(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_28.d ),
    .RESET_B(_030_),
    .Q(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_28.s_currentState ));
 sky130_fd_sc_hd__dfrtp_2 _746_ (.CLK(_033_),
    .D(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_29.d ),
    .RESET_B(_032_),
    .Q(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_29.s_currentState ));
 sky130_fd_sc_hd__dfrtp_2 _747_ (.CLK(_035_),
    .D(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_30.d ),
    .RESET_B(_034_),
    .Q(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_30.s_currentState ));
 sky130_fd_sc_hd__dfrtp_4 _748_ (.CLK(_037_),
    .D(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_31.d ),
    .RESET_B(_036_),
    .Q(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_31.s_currentState ));
 sky130_fd_sc_hd__dfrtp_2 _749_ (.CLK(net16),
    .D(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_32.d ),
    .RESET_B(_038_),
    .Q(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_32.s_currentState ));
 sky130_fd_sc_hd__dfrtp_2 _750_ (.CLK(_040_),
    .D(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_33.d ),
    .RESET_B(_039_),
    .Q(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_33.s_currentState ));
 sky130_fd_sc_hd__dfrtp_2 _751_ (.CLK(_042_),
    .D(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_34.d ),
    .RESET_B(_041_),
    .Q(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_34.s_currentState ));
 sky130_fd_sc_hd__dfrtp_2 _752_ (.CLK(_044_),
    .D(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_35.d ),
    .RESET_B(_043_),
    .Q(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_35.s_currentState ));
 sky130_fd_sc_hd__dfrtp_2 _753_ (.CLK(_046_),
    .D(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_36.d ),
    .RESET_B(_045_),
    .Q(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_36.s_currentState ));
 sky130_fd_sc_hd__dfrtp_2 _754_ (.CLK(_048_),
    .D(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_37.d ),
    .RESET_B(_047_),
    .Q(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_37.s_currentState ));
 sky130_fd_sc_hd__dfrtp_2 _755_ (.CLK(_050_),
    .D(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_28.clock ),
    .RESET_B(_049_),
    .Q(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_38.s_currentState ));
 sky130_fd_sc_hd__dfxtp_2 _756_ (.CLK(\CIRCUIT_2223.triangle_wave_generator_1.GATES_27.result ),
    .D(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_39.d ),
    .Q(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_39.s_currentState ));
 sky130_fd_sc_hd__dfxtp_1 _757_ (.CLK(_051_),
    .D(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_40.d ),
    .Q(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_40.s_currentState ));
 sky130_fd_sc_hd__dfxtp_2 _758_ (.CLK(_052_),
    .D(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_40.clock ),
    .Q(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_41.s_currentState ));
 sky130_fd_sc_hd__dfxtp_2 _759_ (.CLK(_053_),
    .D(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_41.clock ),
    .Q(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_42.s_currentState ));
 sky130_fd_sc_hd__dfxtp_1 _760_ (.CLK(net26),
    .D(_142_),
    .Q(\CIRCUIT_2223.tone_generator_2_2.GATES_8.input2 ));
 sky130_fd_sc_hd__dfxtp_1 _761_ (.CLK(net30),
    .D(_143_),
    .Q(\CIRCUIT_2223.tone_generator_2_2.GATES_9.input2 ));
 sky130_fd_sc_hd__dfxtp_1 _762_ (.CLK(net30),
    .D(_144_),
    .Q(\CIRCUIT_2223.tone_generator_2_2.GATES_10.input2 ));
 sky130_fd_sc_hd__dfxtp_1 _763_ (.CLK(net24),
    .D(_145_),
    .Q(\CIRCUIT_2223.triangle_wave_generator_1.GATES_11.input2 ));
 sky130_fd_sc_hd__dfxtp_1 _764_ (.CLK(net24),
    .D(_146_),
    .Q(\CIRCUIT_2223.triangle_wave_generator_1.GATES_12.input2 ));
 sky130_fd_sc_hd__dfxtp_1 _765_ (.CLK(net24),
    .D(_147_),
    .Q(\CIRCUIT_2223.triangle_wave_generator_1.GATES_13.input2 ));
 sky130_fd_sc_hd__dfxtp_1 _766_ (.CLK(net24),
    .D(_148_),
    .Q(\CIRCUIT_2223.triangle_wave_generator_1.GATES_14.input2 ));
 sky130_fd_sc_hd__dfxtp_1 _767_ (.CLK(net23),
    .D(_149_),
    .Q(\CIRCUIT_2223.triangle_wave_generator_1.GATES_15.input2 ));
 sky130_fd_sc_hd__dfxtp_1 _768_ (.CLK(net23),
    .D(_150_),
    .Q(\CIRCUIT_2223.triangle_wave_generator_1.GATES_16.input2 ));
 sky130_fd_sc_hd__dfxtp_1 _769_ (.CLK(net23),
    .D(_151_),
    .Q(\CIRCUIT_2223.triangle_wave_generator_1.GATES_17.input2 ));
 sky130_fd_sc_hd__dfxtp_1 _770_ (.CLK(net24),
    .D(_152_),
    .Q(\CIRCUIT_2223.triangle_wave_generator_1.GATES_7.input2 ));
 sky130_fd_sc_hd__dfrtp_2 _771_ (.CLK(_055_),
    .D(\CIRCUIT_2223.tone_generator_2_1.MEMORY_28.d ),
    .RESET_B(_054_),
    .Q(\CIRCUIT_2223.tone_generator_2_1.MEMORY_28.s_currentState ));
 sky130_fd_sc_hd__dfrtp_2 _772_ (.CLK(_057_),
    .D(\CIRCUIT_2223.tone_generator_2_1.MEMORY_29.d ),
    .RESET_B(_056_),
    .Q(\CIRCUIT_2223.tone_generator_2_1.MEMORY_29.s_currentState ));
 sky130_fd_sc_hd__dfrtp_2 _773_ (.CLK(_059_),
    .D(\CIRCUIT_2223.tone_generator_2_1.MEMORY_30.d ),
    .RESET_B(_058_),
    .Q(\CIRCUIT_2223.tone_generator_2_1.MEMORY_30.s_currentState ));
 sky130_fd_sc_hd__dfrtp_4 _774_ (.CLK(_061_),
    .D(\CIRCUIT_2223.tone_generator_2_1.MEMORY_31.d ),
    .RESET_B(_060_),
    .Q(\CIRCUIT_2223.tone_generator_2_1.MEMORY_31.s_currentState ));
 sky130_fd_sc_hd__dfrtp_2 _775_ (.CLK(\CIRCUIT_2223.MEMORY_18.s_currentState ),
    .D(\CIRCUIT_2223.tone_generator_2_1.MEMORY_32.d ),
    .RESET_B(_062_),
    .Q(\CIRCUIT_2223.tone_generator_2_1.MEMORY_32.s_currentState ));
 sky130_fd_sc_hd__dfrtp_2 _776_ (.CLK(_064_),
    .D(\CIRCUIT_2223.tone_generator_2_1.MEMORY_33.d ),
    .RESET_B(_063_),
    .Q(\CIRCUIT_2223.tone_generator_2_1.MEMORY_33.s_currentState ));
 sky130_fd_sc_hd__dfrtp_2 _777_ (.CLK(_066_),
    .D(\CIRCUIT_2223.tone_generator_2_1.MEMORY_34.d ),
    .RESET_B(_065_),
    .Q(\CIRCUIT_2223.tone_generator_2_1.MEMORY_34.s_currentState ));
 sky130_fd_sc_hd__dfrtp_2 _778_ (.CLK(_068_),
    .D(\CIRCUIT_2223.tone_generator_2_1.MEMORY_35.d ),
    .RESET_B(_067_),
    .Q(\CIRCUIT_2223.tone_generator_2_1.MEMORY_35.s_currentState ));
 sky130_fd_sc_hd__dfrtp_2 _779_ (.CLK(_070_),
    .D(\CIRCUIT_2223.tone_generator_2_1.MEMORY_36.d ),
    .RESET_B(_069_),
    .Q(\CIRCUIT_2223.tone_generator_2_1.MEMORY_36.s_currentState ));
 sky130_fd_sc_hd__dfrtp_2 _780_ (.CLK(_072_),
    .D(\CIRCUIT_2223.tone_generator_2_1.MEMORY_37.d ),
    .RESET_B(_071_),
    .Q(\CIRCUIT_2223.tone_generator_2_1.MEMORY_37.s_currentState ));
 sky130_fd_sc_hd__dfrtp_2 _781_ (.CLK(_074_),
    .D(\CIRCUIT_2223.tone_generator_2_1.MEMORY_28.clock ),
    .RESET_B(_073_),
    .Q(\CIRCUIT_2223.tone_generator_2_1.MEMORY_38.s_currentState ));
 sky130_fd_sc_hd__dfxtp_1 _782_ (.CLK(\CIRCUIT_2223.tone_generator_2_1.GATES_27.result ),
    .D(\CIRCUIT_2223.tone_generator_2_1.MEMORY_39.d ),
    .Q(\CIRCUIT_2223.tone_generator_2_1.MEMORY_39.s_currentState ));
 sky130_fd_sc_hd__dfxtp_1 _783_ (.CLK(net30),
    .D(_153_),
    .Q(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_8.input2 ));
 sky130_fd_sc_hd__dfxtp_1 _784_ (.CLK(net29),
    .D(_154_),
    .Q(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_9.input2 ));
 sky130_fd_sc_hd__dfxtp_1 _785_ (.CLK(net30),
    .D(_155_),
    .Q(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_10.input2 ));
 sky130_fd_sc_hd__dfxtp_1 _786_ (.CLK(net29),
    .D(_156_),
    .Q(\CIRCUIT_2223.tone_generator_2_1.GATES_11.input2 ));
 sky130_fd_sc_hd__dfxtp_1 _787_ (.CLK(net29),
    .D(_157_),
    .Q(\CIRCUIT_2223.tone_generator_2_1.GATES_12.input2 ));
 sky130_fd_sc_hd__dfxtp_1 _788_ (.CLK(net29),
    .D(_158_),
    .Q(\CIRCUIT_2223.tone_generator_2_1.GATES_13.input2 ));
 sky130_fd_sc_hd__dfxtp_1 _789_ (.CLK(net31),
    .D(_159_),
    .Q(\CIRCUIT_2223.tone_generator_2_1.GATES_14.input2 ));
 sky130_fd_sc_hd__dfxtp_1 _790_ (.CLK(net29),
    .D(_160_),
    .Q(\CIRCUIT_2223.tone_generator_2_1.GATES_15.input2 ));
 sky130_fd_sc_hd__dfxtp_1 _791_ (.CLK(net31),
    .D(_161_),
    .Q(\CIRCUIT_2223.tone_generator_2_1.GATES_16.input2 ));
 sky130_fd_sc_hd__dfxtp_1 _792_ (.CLK(net29),
    .D(_162_),
    .Q(\CIRCUIT_2223.tone_generator_2_1.GATES_17.input2 ));
 sky130_fd_sc_hd__dfxtp_1 _793_ (.CLK(net31),
    .D(_163_),
    .Q(\CIRCUIT_2223.tone_generator_2_1.GATES_7.input2 ));
 sky130_fd_sc_hd__dfrtp_2 _794_ (.CLK(_076_),
    .D(\CIRCUIT_2223.tone_generator_2_2.MEMORY_28.d ),
    .RESET_B(_075_),
    .Q(\CIRCUIT_2223.tone_generator_2_2.MEMORY_28.s_currentState ));
 sky130_fd_sc_hd__dfrtp_2 _795_ (.CLK(_078_),
    .D(\CIRCUIT_2223.tone_generator_2_2.MEMORY_29.d ),
    .RESET_B(_077_),
    .Q(\CIRCUIT_2223.tone_generator_2_2.MEMORY_29.s_currentState ));
 sky130_fd_sc_hd__dfrtp_2 _796_ (.CLK(_080_),
    .D(\CIRCUIT_2223.tone_generator_2_2.MEMORY_30.d ),
    .RESET_B(_079_),
    .Q(\CIRCUIT_2223.tone_generator_2_2.MEMORY_30.s_currentState ));
 sky130_fd_sc_hd__dfrtp_4 _797_ (.CLK(_082_),
    .D(\CIRCUIT_2223.tone_generator_2_2.MEMORY_31.d ),
    .RESET_B(_081_),
    .Q(\CIRCUIT_2223.tone_generator_2_2.MEMORY_31.s_currentState ));
 sky130_fd_sc_hd__dfrtp_2 _798_ (.CLK(\CIRCUIT_2223.MEMORY_18.s_currentState ),
    .D(\CIRCUIT_2223.tone_generator_2_2.MEMORY_32.d ),
    .RESET_B(_083_),
    .Q(\CIRCUIT_2223.tone_generator_2_2.MEMORY_32.s_currentState ));
 sky130_fd_sc_hd__dfrtp_2 _799_ (.CLK(_085_),
    .D(\CIRCUIT_2223.tone_generator_2_2.MEMORY_33.d ),
    .RESET_B(_084_),
    .Q(\CIRCUIT_2223.tone_generator_2_2.MEMORY_33.s_currentState ));
 sky130_fd_sc_hd__dfrtp_2 _800_ (.CLK(_087_),
    .D(\CIRCUIT_2223.tone_generator_2_2.MEMORY_34.d ),
    .RESET_B(_086_),
    .Q(\CIRCUIT_2223.tone_generator_2_2.MEMORY_34.s_currentState ));
 sky130_fd_sc_hd__dfrtp_2 _801_ (.CLK(_089_),
    .D(\CIRCUIT_2223.tone_generator_2_2.MEMORY_35.d ),
    .RESET_B(_088_),
    .Q(\CIRCUIT_2223.tone_generator_2_2.MEMORY_35.s_currentState ));
 sky130_fd_sc_hd__dfrtp_2 _802_ (.CLK(_091_),
    .D(\CIRCUIT_2223.tone_generator_2_2.MEMORY_36.d ),
    .RESET_B(_090_),
    .Q(\CIRCUIT_2223.tone_generator_2_2.MEMORY_36.s_currentState ));
 sky130_fd_sc_hd__dfrtp_2 _803_ (.CLK(_093_),
    .D(\CIRCUIT_2223.tone_generator_2_2.MEMORY_37.d ),
    .RESET_B(_092_),
    .Q(\CIRCUIT_2223.tone_generator_2_2.MEMORY_37.s_currentState ));
 sky130_fd_sc_hd__dfrtp_2 _804_ (.CLK(_095_),
    .D(\CIRCUIT_2223.tone_generator_2_2.MEMORY_28.clock ),
    .RESET_B(_094_),
    .Q(\CIRCUIT_2223.tone_generator_2_2.MEMORY_38.s_currentState ));
 sky130_fd_sc_hd__dfxtp_2 _805_ (.CLK(\CIRCUIT_2223.tone_generator_2_2.GATES_27.result ),
    .D(\CIRCUIT_2223.tone_generator_2_2.MEMORY_39.d ),
    .Q(\CIRCUIT_2223.tone_generator_2_2.MEMORY_39.s_currentState ));
 sky130_fd_sc_hd__dfxtp_1 _806_ (.CLK(net30),
    .D(_164_),
    .Q(\CIRCUIT_2223.tone_generator_2_1.GATES_8.input2 ));
 sky130_fd_sc_hd__dfxtp_1 _807_ (.CLK(net30),
    .D(_165_),
    .Q(\CIRCUIT_2223.tone_generator_2_1.GATES_9.input2 ));
 sky130_fd_sc_hd__dfxtp_1 _808_ (.CLK(net30),
    .D(_166_),
    .Q(\CIRCUIT_2223.tone_generator_2_1.GATES_10.input2 ));
 sky130_fd_sc_hd__dfxtp_1 _809_ (.CLK(net26),
    .D(_167_),
    .Q(\CIRCUIT_2223.tone_generator_2_2.GATES_11.input2 ));
 sky130_fd_sc_hd__dfxtp_1 _810_ (.CLK(net26),
    .D(_168_),
    .Q(\CIRCUIT_2223.tone_generator_2_2.GATES_12.input2 ));
 sky130_fd_sc_hd__dfxtp_1 _811_ (.CLK(net25),
    .D(_169_),
    .Q(\CIRCUIT_2223.tone_generator_2_2.GATES_13.input2 ));
 sky130_fd_sc_hd__dfxtp_1 _812_ (.CLK(net26),
    .D(_170_),
    .Q(\CIRCUIT_2223.tone_generator_2_2.GATES_14.input2 ));
 sky130_fd_sc_hd__dfxtp_1 _813_ (.CLK(net25),
    .D(_171_),
    .Q(\CIRCUIT_2223.tone_generator_2_2.GATES_15.input2 ));
 sky130_fd_sc_hd__dfxtp_1 _814_ (.CLK(net25),
    .D(_172_),
    .Q(\CIRCUIT_2223.tone_generator_2_2.GATES_16.input2 ));
 sky130_fd_sc_hd__dfxtp_1 _815_ (.CLK(net25),
    .D(_173_),
    .Q(\CIRCUIT_2223.tone_generator_2_2.GATES_17.input2 ));
 sky130_fd_sc_hd__dfxtp_1 _816_ (.CLK(net25),
    .D(_174_),
    .Q(\CIRCUIT_2223.tone_generator_2_2.GATES_7.input2 ));
 sky130_fd_sc_hd__dfxtp_1 _817_ (.CLK(_096_),
    .D(net38),
    .Q(net15));
 sky130_fd_sc_hd__dfxtp_1 _818_ (.CLK(_097_),
    .D(net38),
    .Q(net14));
 sky130_fd_sc_hd__dfrtp_4 _819_ (.CLK(net29),
    .D(_175_),
    .RESET_B(_098_),
    .Q(\CIRCUIT_2223.GATES_2.input2 ));
 sky130_fd_sc_hd__dfrtp_1 _820_ (.CLK(net29),
    .D(_176_),
    .RESET_B(_099_),
    .Q(\CIRCUIT_2223.GATES_3.input2 ));
 sky130_fd_sc_hd__dfrtp_2 _821_ (.CLK(net27),
    .D(_177_),
    .RESET_B(_100_),
    .Q(\CIRCUIT_2223.GATES_5.input2 ));
 sky130_fd_sc_hd__dfrtp_2 _822_ (.CLK(net27),
    .D(_178_),
    .RESET_B(_101_),
    .Q(\CIRCUIT_2223.s_logisimNet48 ));
 sky130_fd_sc_hd__dfrtp_4 _823_ (.CLK(_103_),
    .D(\CIRCUIT_2223.MEMORY_18.clock ),
    .RESET_B(_102_),
    .Q(\CIRCUIT_2223.MEMORY_26.s_currentState ));
 sky130_fd_sc_hd__dfrtp_4 _824_ (.CLK(_105_),
    .D(\CIRCUIT_2223.MEMORY_25.d ),
    .RESET_B(_104_),
    .Q(\CIRCUIT_2223.MEMORY_25.s_currentState ));
 sky130_fd_sc_hd__dfrtp_4 _825_ (.CLK(net39),
    .D(\CIRCUIT_2223.MEMORY_24.d ),
    .RESET_B(net44),
    .Q(\CIRCUIT_2223.MEMORY_24.s_currentState ));
 sky130_fd_sc_hd__dfrtp_1 _826_ (.CLK(_108_),
    .D(\CIRCUIT_2223.GATES_11.input2 ),
    .RESET_B(_107_),
    .Q(\CIRCUIT_2223.MEMORY_23.s_currentState ));
 sky130_fd_sc_hd__dfrtp_4 _827_ (.CLK(_110_),
    .D(\CIRCUIT_2223.MEMORY_22.d ),
    .RESET_B(_109_),
    .Q(\CIRCUIT_2223.MEMORY_22.s_currentState ));
 sky130_fd_sc_hd__dfrtp_4 _828_ (.CLK(_112_),
    .D(\CIRCUIT_2223.MEMORY_21.d ),
    .RESET_B(_111_),
    .Q(\CIRCUIT_2223.MEMORY_21.s_currentState ));
 sky130_fd_sc_hd__dfrtp_4 _829_ (.CLK(_114_),
    .D(\CIRCUIT_2223.MEMORY_20.d ),
    .RESET_B(_113_),
    .Q(\CIRCUIT_2223.MEMORY_20.s_currentState ));
 sky130_fd_sc_hd__dfrtp_4 _830_ (.CLK(_116_),
    .D(\CIRCUIT_2223.MEMORY_19.d ),
    .RESET_B(_115_),
    .Q(\CIRCUIT_2223.MEMORY_19.s_currentState ));
 sky130_fd_sc_hd__dfrtp_2 _831_ (.CLK(_118_),
    .D(\CIRCUIT_2223.MEMORY_18.d ),
    .RESET_B(_117_),
    .Q(\CIRCUIT_2223.MEMORY_18.s_currentState ));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__183_ (.A(_183_),
    .X(clknet_0__183_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__203_ (.A(_203_),
    .X(clknet_0__203_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__222_ (.A(_222_),
    .X(clknet_0__222_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__245_ (.A(_245_),
    .X(clknet_0__245_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__264_ (.A(_264_),
    .X(clknet_0__264_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__183_ (.A(clknet_0__183_),
    .X(clknet_1_0__leaf__183_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__203_ (.A(clknet_0__203_),
    .X(clknet_1_0__leaf__203_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__222_ (.A(clknet_0__222_),
    .X(clknet_1_0__leaf__222_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__245_ (.A(clknet_0__245_),
    .X(clknet_1_0__leaf__245_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__264_ (.A(clknet_0__264_),
    .X(clknet_1_0__leaf__264_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_clk (.A(clknet_0_clk),
    .X(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__183_ (.A(clknet_0__183_),
    .X(clknet_1_1__leaf__183_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__203_ (.A(clknet_0__203_),
    .X(clknet_1_1__leaf__203_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__222_ (.A(clknet_0__222_),
    .X(clknet_1_1__leaf__222_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__245_ (.A(clknet_0__245_),
    .X(clknet_1_1__leaf__245_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__264_ (.A(clknet_0__264_),
    .X(clknet_1_1__leaf__264_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_clk (.A(clknet_0_clk),
    .X(clknet_1_1__leaf_clk));
 sky130_fd_sc_hd__buf_4 fanout16 (.A(net17),
    .X(net16));
 sky130_fd_sc_hd__buf_4 fanout17 (.A(\CIRCUIT_2223.MEMORY_24.s_currentState ),
    .X(net17));
 sky130_fd_sc_hd__buf_12 fanout18 (.A(net20),
    .X(net18));
 sky130_fd_sc_hd__buf_12 fanout19 (.A(net20),
    .X(net19));
 sky130_fd_sc_hd__buf_12 fanout20 (.A(_000_),
    .X(net20));
 sky130_fd_sc_hd__buf_12 fanout21 (.A(net22),
    .X(net21));
 sky130_fd_sc_hd__buf_12 fanout22 (.A(_000_),
    .X(net22));
 sky130_fd_sc_hd__buf_6 fanout23 (.A(net32),
    .X(net23));
 sky130_fd_sc_hd__buf_4 fanout24 (.A(net42),
    .X(net24));
 sky130_fd_sc_hd__buf_4 fanout25 (.A(net32),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_2 fanout26 (.A(net32),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_4 fanout27 (.A(net28),
    .X(net27));
 sky130_fd_sc_hd__buf_4 fanout28 (.A(net31),
    .X(net28));
 sky130_fd_sc_hd__clkbuf_4 fanout29 (.A(net30),
    .X(net29));
 sky130_fd_sc_hd__buf_4 fanout30 (.A(net31),
    .X(net30));
 sky130_fd_sc_hd__buf_4 fanout31 (.A(net32),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_4 fanout32 (.A(net41),
    .X(net32));
 sky130_fd_sc_hd__buf_6 fanout33 (.A(net34),
    .X(net33));
 sky130_fd_sc_hd__buf_6 fanout34 (.A(net7),
    .X(net34));
 sky130_fd_sc_hd__buf_4 fanout35 (.A(net5),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_8 fanout36 (.A(net4),
    .X(net36));
 sky130_fd_sc_hd__clkbuf_8 fanout37 (.A(net3),
    .X(net37));
 sky130_fd_sc_hd__buf_2 fanout38 (.A(net3),
    .X(net38));
 sky130_fd_sc_hd__buf_2 hold1 (.A(net45),
    .X(net41));
 sky130_fd_sc_hd__buf_2 hold2 (.A(net32),
    .X(net42));
 sky130_fd_sc_hd__buf_2 hold3 (.A(net24),
    .X(net43));
 sky130_fd_sc_hd__buf_2 hold4 (.A(_106_),
    .X(net44));
 sky130_fd_sc_hd__buf_2 hold5 (.A(\CIRCUIT_2223.CLK ),
    .X(net45));
 sky130_fd_sc_hd__buf_6 input1 (.A(io_in[0]),
    .X(net1));
 sky130_fd_sc_hd__buf_6 input2 (.A(io_in[1]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_2 input3 (.A(io_in[2]),
    .X(net3));
 sky130_fd_sc_hd__buf_2 input4 (.A(io_in[3]),
    .X(net4));
 sky130_fd_sc_hd__buf_2 input5 (.A(io_in[4]),
    .X(net5));
 sky130_fd_sc_hd__buf_6 input6 (.A(io_in[5]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_4 input7 (.A(rst),
    .X(net7));
 sky130_fd_sc_hd__buf_4 output10 (.A(net10),
    .X(io_out[2]));
 sky130_fd_sc_hd__buf_4 output11 (.A(net11),
    .X(io_out[3]));
 sky130_fd_sc_hd__buf_4 output12 (.A(net12),
    .X(io_out[4]));
 sky130_fd_sc_hd__buf_4 output13 (.A(net13),
    .X(io_out[5]));
 sky130_fd_sc_hd__buf_4 output14 (.A(net14),
    .X(io_out[6]));
 sky130_fd_sc_hd__buf_4 output15 (.A(net15),
    .X(io_out[7]));
 sky130_fd_sc_hd__buf_4 output8 (.A(net8),
    .X(io_out[0]));
 sky130_fd_sc_hd__buf_4 output9 (.A(net9),
    .X(io_out[1]));
endmodule

