* NGSPICE file created from user_project_wrapper.ext - technology: sky130B

* Black-box entry subcircuit for tune_player abstract view
.subckt tune_player OP clk rst vccd1 vssd1
.ends

* Black-box entry subcircuit for posit_unit abstract view
.subckt posit_unit clk io_in[0] io_in[1] io_in[2] io_out[0] io_out[1] io_out[2] io_out[3]
+ rst vccd1 vssd1
.ends

* Black-box entry subcircuit for tt2_tholin_multiplexed_counter abstract view
.subckt tt2_tholin_multiplexed_counter clk io_out[0] io_out[10] io_out[11] io_out[1]
+ io_out[2] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7] io_out[8] io_out[9]
+ rst vccd1 vssd1
.ends

* Black-box entry subcircuit for wrapped_MC14500 abstract view
.subckt wrapped_MC14500 clk io_in[0] io_in[1] io_in[2] io_in[3] io_in[4] io_oeb io_out[0]
+ io_out[1] io_out[2] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7] io_out[8]
+ rst vccd1 vssd1
.ends

* Black-box entry subcircuit for multiplexer abstract view
.subckt multiplexer design_clk_o dsi_all[0] dsi_all[10] dsi_all[11] dsi_all[12] dsi_all[13]
+ dsi_all[14] dsi_all[15] dsi_all[16] dsi_all[17] dsi_all[18] dsi_all[19] dsi_all[1]
+ dsi_all[20] dsi_all[21] dsi_all[22] dsi_all[23] dsi_all[24] dsi_all[25] dsi_all[26]
+ dsi_all[27] dsi_all[2] dsi_all[3] dsi_all[4] dsi_all[5] dsi_all[6] dsi_all[7] dsi_all[8]
+ dsi_all[9] dso_6502[0] dso_6502[10] dso_6502[11] dso_6502[12] dso_6502[13] dso_6502[14]
+ dso_6502[15] dso_6502[16] dso_6502[17] dso_6502[18] dso_6502[19] dso_6502[1] dso_6502[20]
+ dso_6502[21] dso_6502[22] dso_6502[23] dso_6502[24] dso_6502[25] dso_6502[26] dso_6502[2]
+ dso_6502[3] dso_6502[4] dso_6502[5] dso_6502[6] dso_6502[7] dso_6502[8] dso_6502[9]
+ dso_LCD[0] dso_LCD[1] dso_LCD[2] dso_LCD[3] dso_LCD[4] dso_LCD[5] dso_LCD[6] dso_LCD[7]
+ dso_as1802[0] dso_as1802[10] dso_as1802[11] dso_as1802[12] dso_as1802[13] dso_as1802[14]
+ dso_as1802[15] dso_as1802[16] dso_as1802[17] dso_as1802[18] dso_as1802[19] dso_as1802[1]
+ dso_as1802[20] dso_as1802[21] dso_as1802[22] dso_as1802[23] dso_as1802[24] dso_as1802[25]
+ dso_as1802[26] dso_as1802[2] dso_as1802[3] dso_as1802[4] dso_as1802[5] dso_as1802[6]
+ dso_as1802[7] dso_as1802[8] dso_as1802[9] dso_as2650[0] dso_as2650[10] dso_as2650[11]
+ dso_as2650[12] dso_as2650[13] dso_as2650[14] dso_as2650[15] dso_as2650[16] dso_as2650[17]
+ dso_as2650[18] dso_as2650[19] dso_as2650[1] dso_as2650[20] dso_as2650[21] dso_as2650[22]
+ dso_as2650[23] dso_as2650[24] dso_as2650[25] dso_as2650[26] dso_as2650[2] dso_as2650[3]
+ dso_as2650[4] dso_as2650[5] dso_as2650[6] dso_as2650[7] dso_as2650[8] dso_as2650[9]
+ dso_as512512512[0] dso_as512512512[10] dso_as512512512[11] dso_as512512512[12] dso_as512512512[13]
+ dso_as512512512[14] dso_as512512512[15] dso_as512512512[16] dso_as512512512[17]
+ dso_as512512512[18] dso_as512512512[19] dso_as512512512[1] dso_as512512512[20] dso_as512512512[21]
+ dso_as512512512[22] dso_as512512512[23] dso_as512512512[24] dso_as512512512[25]
+ dso_as512512512[26] dso_as512512512[27] dso_as512512512[2] dso_as512512512[3] dso_as512512512[4]
+ dso_as512512512[5] dso_as512512512[6] dso_as512512512[7] dso_as512512512[8] dso_as512512512[9]
+ dso_as5401[0] dso_as5401[10] dso_as5401[11] dso_as5401[12] dso_as5401[13] dso_as5401[14]
+ dso_as5401[15] dso_as5401[16] dso_as5401[17] dso_as5401[18] dso_as5401[19] dso_as5401[1]
+ dso_as5401[20] dso_as5401[21] dso_as5401[22] dso_as5401[23] dso_as5401[24] dso_as5401[25]
+ dso_as5401[26] dso_as5401[2] dso_as5401[3] dso_as5401[4] dso_as5401[5] dso_as5401[6]
+ dso_as5401[7] dso_as5401[8] dso_as5401[9] dso_counter[0] dso_counter[10] dso_counter[11]
+ dso_counter[1] dso_counter[2] dso_counter[3] dso_counter[4] dso_counter[5] dso_counter[6]
+ dso_counter[7] dso_counter[8] dso_counter[9] dso_diceroll[0] dso_diceroll[1] dso_diceroll[2]
+ dso_diceroll[3] dso_diceroll[4] dso_diceroll[5] dso_diceroll[6] dso_diceroll[7]
+ dso_mc14500[0] dso_mc14500[1] dso_mc14500[2] dso_mc14500[3] dso_mc14500[4] dso_mc14500[5]
+ dso_mc14500[6] dso_mc14500[7] dso_mc14500[8] dso_multiplier[0] dso_multiplier[1]
+ dso_multiplier[2] dso_multiplier[3] dso_multiplier[4] dso_multiplier[5] dso_multiplier[6]
+ dso_multiplier[7] dso_posit[0] dso_posit[1] dso_posit[2] dso_posit[3] dso_tbb1143[0]
+ dso_tbb1143[1] dso_tbb1143[2] dso_tbb1143[3] dso_tbb1143[4] dso_tbb1143[5] dso_tbb1143[6]
+ dso_tbb1143[7] dso_tune io_in[0] io_in[10] io_in[11] io_in[12] io_in[13] io_in[14]
+ io_in[15] io_in[16] io_in[17] io_in[18] io_in[19] io_in[1] io_in[20] io_in[21] io_in[22]
+ io_in[23] io_in[24] io_in[25] io_in[26] io_in[27] io_in[28] io_in[29] io_in[2] io_in[30]
+ io_in[31] io_in[32] io_in[33] io_in[34] io_in[35] io_in[36] io_in[37] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_in[8] io_in[9] io_oeb[0] io_oeb[10] io_oeb[11] io_oeb[12]
+ io_oeb[13] io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18] io_oeb[19] io_oeb[1]
+ io_oeb[20] io_oeb[21] io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25] io_oeb[26] io_oeb[27]
+ io_oeb[28] io_oeb[29] io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32] io_oeb[33] io_oeb[34]
+ io_oeb[35] io_oeb[36] io_oeb[37] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7]
+ io_oeb[8] io_oeb[9] io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14]
+ io_out[15] io_out[16] io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21]
+ io_out[22] io_out[23] io_out[24] io_out[25] io_out[26] io_out[27] io_out[28] io_out[29]
+ io_out[2] io_out[30] io_out[31] io_out[32] io_out[33] io_out[34] io_out[35] io_out[36]
+ io_out[37] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7] io_out[8] io_out[9]
+ oeb_6502 oeb_as1802 oeb_as2650 oeb_as512512512 oeb_as5401 oeb_mc14500 rst_6502 rst_LCD
+ rst_as1802 rst_as2650 rst_as512512512 rst_as5401 rst_counter rst_diceroll rst_mc14500
+ rst_posit rst_tbb1143 rst_tune vccd1 vssd1 wb_clk_i wb_rst_i wbs_ack_o wbs_adr_i[0]
+ wbs_adr_i[10] wbs_adr_i[11] wbs_adr_i[12] wbs_adr_i[13] wbs_adr_i[14] wbs_adr_i[15]
+ wbs_adr_i[16] wbs_adr_i[17] wbs_adr_i[18] wbs_adr_i[19] wbs_adr_i[1] wbs_adr_i[20]
+ wbs_adr_i[21] wbs_adr_i[22] wbs_adr_i[23] wbs_adr_i[24] wbs_adr_i[25] wbs_adr_i[26]
+ wbs_adr_i[27] wbs_adr_i[28] wbs_adr_i[29] wbs_adr_i[2] wbs_adr_i[30] wbs_adr_i[31]
+ wbs_adr_i[3] wbs_adr_i[4] wbs_adr_i[5] wbs_adr_i[6] wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9]
+ wbs_cyc_i wbs_dat_i[0] wbs_dat_i[10] wbs_dat_i[11] wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14]
+ wbs_dat_i[15] wbs_dat_i[16] wbs_dat_i[17] wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1]
+ wbs_dat_i[20] wbs_dat_i[21] wbs_dat_i[22] wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25]
+ wbs_dat_i[26] wbs_dat_i[27] wbs_dat_i[28] wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30]
+ wbs_dat_i[31] wbs_dat_i[3] wbs_dat_i[4] wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8]
+ wbs_dat_i[9] wbs_dat_o[0] wbs_dat_o[10] wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13]
+ wbs_dat_o[14] wbs_dat_o[15] wbs_dat_o[16] wbs_dat_o[17] wbs_dat_o[18] wbs_dat_o[19]
+ wbs_dat_o[1] wbs_dat_o[20] wbs_dat_o[21] wbs_dat_o[22] wbs_dat_o[23] wbs_dat_o[24]
+ wbs_dat_o[25] wbs_dat_o[26] wbs_dat_o[27] wbs_dat_o[28] wbs_dat_o[29] wbs_dat_o[2]
+ wbs_dat_o[30] wbs_dat_o[31] wbs_dat_o[3] wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6]
+ wbs_dat_o[7] wbs_dat_o[8] wbs_dat_o[9] wbs_stb_i wbs_we_i
.ends

* Black-box entry subcircuit for tt2_tholin_multiplier abstract view
.subckt tt2_tholin_multiplier io_in[0] io_in[1] io_in[2] io_in[3] io_in[4] io_in[5]
+ io_in[6] io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5] io_out[6]
+ io_out[7] vccd1 vssd1
.ends

* Black-box entry subcircuit for tt2_tholin_diceroll abstract view
.subckt tt2_tholin_diceroll clk io_in io_out[0] io_out[1] io_out[2] io_out[3] io_out[4]
+ io_out[5] io_out[6] io_out[7] rst vccd1 vssd1
.ends

* Black-box entry subcircuit for tholin_avalonsemi_tbb1143 abstract view
.subckt tholin_avalonsemi_tbb1143 clk io_in[0] io_in[1] io_in[2] io_in[3] io_in[4]
+ io_in[5] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7]
+ rst vccd1 vssd1
.ends

* Black-box entry subcircuit for tholin_avalonsemi_5401 abstract view
.subckt tholin_avalonsemi_5401 clk io_in[0] io_in[1] io_in[2] io_in[3] io_in[4] io_in[5]
+ io_in[6] io_in[7] io_in[8] io_in[9] io_oeb io_out[0] io_out[10] io_out[11] io_out[12]
+ io_out[13] io_out[14] io_out[15] io_out[16] io_out[17] io_out[18] io_out[19] io_out[1]
+ io_out[20] io_out[21] io_out[22] io_out[23] io_out[24] io_out[25] io_out[26] io_out[2]
+ io_out[3] io_out[4] io_out[5] io_out[6] io_out[7] io_out[8] io_out[9] rst vccd1
+ vssd1
.ends

* Black-box entry subcircuit for wrapped_vgatest abstract view
.subckt wrapped_vgatest clk io_in io_out[0] io_out[1] io_out[2] io_out[3] io_out[4]
+ io_out[5] io_out[6] io_out[7] io_out[8] io_out[9] rst vccd1 vssd1
.ends

* Black-box entry subcircuit for wrapped_as512512512 abstract view
.subckt wrapped_as512512512 clk io_in[0] io_in[10] io_in[11] io_in[12] io_in[13] io_in[14]
+ io_in[15] io_in[16] io_in[17] io_in[18] io_in[19] io_in[1] io_in[20] io_in[21] io_in[22]
+ io_in[23] io_in[24] io_in[25] io_in[26] io_in[2] io_in[3] io_in[4] io_in[5] io_in[6]
+ io_in[7] io_in[8] io_in[9] io_oeb io_out[0] io_out[10] io_out[11] io_out[12] io_out[13]
+ io_out[14] io_out[15] io_out[16] io_out[17] io_out[18] io_out[19] io_out[1] io_out[20]
+ io_out[21] io_out[22] io_out[23] io_out[24] io_out[25] io_out[26] io_out[27] io_out[2]
+ io_out[3] io_out[4] io_out[5] io_out[6] io_out[7] io_out[8] io_out[9] rst vccd1
+ vssd1
.ends

* Black-box entry subcircuit for wrapped_as1802 abstract view
.subckt wrapped_as1802 clk io_in[0] io_in[10] io_in[11] io_in[12] io_in[1] io_in[2]
+ io_in[3] io_in[4] io_in[5] io_in[6] io_in[7] io_in[8] io_in[9] io_oeb io_out[0]
+ io_out[10] io_out[11] io_out[12] io_out[13] io_out[14] io_out[15] io_out[16] io_out[17]
+ io_out[18] io_out[19] io_out[1] io_out[20] io_out[21] io_out[22] io_out[23] io_out[24]
+ io_out[25] io_out[26] io_out[2] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7]
+ io_out[8] io_out[9] rst vccd1 vssd1
.ends

* Black-box entry subcircuit for wrapped_6502 abstract view
.subckt wrapped_6502 clk io_in[0] io_in[1] io_in[2] io_in[3] io_in[4] io_in[5] io_in[6]
+ io_in[7] io_in[8] io_in[9] io_oeb io_out[0] io_out[10] io_out[11] io_out[12] io_out[13]
+ io_out[14] io_out[15] io_out[16] io_out[17] io_out[18] io_out[19] io_out[1] io_out[20]
+ io_out[21] io_out[22] io_out[23] io_out[24] io_out[25] io_out[26] io_out[2] io_out[3]
+ io_out[4] io_out[5] io_out[6] io_out[7] io_out[8] io_out[9] rst vccd1 vssd1
.ends

* Black-box entry subcircuit for tt2_tholin_namebadge abstract view
.subckt tt2_tholin_namebadge clk io_in[0] io_in[1] io_in[2] io_oeb[0] io_oeb[10] io_oeb[11]
+ io_oeb[12] io_oeb[13] io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18] io_oeb[19]
+ io_oeb[1] io_oeb[20] io_oeb[21] io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25] io_oeb[26]
+ io_oeb[2] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7] io_oeb[8] io_oeb[9]
+ io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7]
+ rst vccd1 vssd1
.ends

* Black-box entry subcircuit for wrapped_as2650 abstract view
.subckt wrapped_as2650 clk io_in[0] io_in[1] io_in[2] io_in[3] io_in[4] io_in[5] io_in[6]
+ io_in[7] io_in[8] io_oeb io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14]
+ io_out[15] io_out[16] io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21]
+ io_out[22] io_out[23] io_out[24] io_out[25] io_out[26] io_out[2] io_out[3] io_out[4]
+ io_out[5] io_out[6] io_out[7] io_out[8] io_out[9] rst vccd1 vssd1
.ends

.subckt user_project_wrapper analog_io[0] analog_io[10] analog_io[11] analog_io[12]
+ analog_io[13] analog_io[14] analog_io[15] analog_io[16] analog_io[17] analog_io[18]
+ analog_io[19] analog_io[1] analog_io[20] analog_io[21] analog_io[22] analog_io[23]
+ analog_io[24] analog_io[25] analog_io[26] analog_io[27] analog_io[28] analog_io[2]
+ analog_io[3] analog_io[4] analog_io[5] analog_io[6] analog_io[7] analog_io[8] analog_io[9]
+ io_in[0] io_in[10] io_in[11] io_in[12] io_in[13] io_in[14] io_in[15] io_in[16] io_in[17]
+ io_in[18] io_in[19] io_in[1] io_in[20] io_in[21] io_in[22] io_in[23] io_in[24] io_in[25]
+ io_in[26] io_in[27] io_in[28] io_in[29] io_in[2] io_in[30] io_in[31] io_in[32] io_in[33]
+ io_in[34] io_in[35] io_in[36] io_in[37] io_in[3] io_in[4] io_in[5] io_in[6] io_in[7]
+ io_in[8] io_in[9] io_oeb[0] io_oeb[10] io_oeb[11] io_oeb[12] io_oeb[13] io_oeb[14]
+ io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18] io_oeb[19] io_oeb[1] io_oeb[20] io_oeb[21]
+ io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25] io_oeb[26] io_oeb[27] io_oeb[28] io_oeb[29]
+ io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32] io_oeb[33] io_oeb[34] io_oeb[35] io_oeb[36]
+ io_oeb[37] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7] io_oeb[8] io_oeb[9]
+ io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14] io_out[15] io_out[16]
+ io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21] io_out[22] io_out[23]
+ io_out[24] io_out[25] io_out[26] io_out[27] io_out[28] io_out[29] io_out[2] io_out[30]
+ io_out[31] io_out[32] io_out[33] io_out[34] io_out[35] io_out[36] io_out[37] io_out[3]
+ io_out[4] io_out[5] io_out[6] io_out[7] io_out[8] io_out[9] la_data_in[0] la_data_in[100]
+ la_data_in[101] la_data_in[102] la_data_in[103] la_data_in[104] la_data_in[105]
+ la_data_in[106] la_data_in[107] la_data_in[108] la_data_in[109] la_data_in[10] la_data_in[110]
+ la_data_in[111] la_data_in[112] la_data_in[113] la_data_in[114] la_data_in[115]
+ la_data_in[116] la_data_in[117] la_data_in[118] la_data_in[119] la_data_in[11] la_data_in[120]
+ la_data_in[121] la_data_in[122] la_data_in[123] la_data_in[124] la_data_in[125]
+ la_data_in[126] la_data_in[127] la_data_in[12] la_data_in[13] la_data_in[14] la_data_in[15]
+ la_data_in[16] la_data_in[17] la_data_in[18] la_data_in[19] la_data_in[1] la_data_in[20]
+ la_data_in[21] la_data_in[22] la_data_in[23] la_data_in[24] la_data_in[25] la_data_in[26]
+ la_data_in[27] la_data_in[28] la_data_in[29] la_data_in[2] la_data_in[30] la_data_in[31]
+ la_data_in[32] la_data_in[33] la_data_in[34] la_data_in[35] la_data_in[36] la_data_in[37]
+ la_data_in[38] la_data_in[39] la_data_in[3] la_data_in[40] la_data_in[41] la_data_in[42]
+ la_data_in[43] la_data_in[44] la_data_in[45] la_data_in[46] la_data_in[47] la_data_in[48]
+ la_data_in[49] la_data_in[4] la_data_in[50] la_data_in[51] la_data_in[52] la_data_in[53]
+ la_data_in[54] la_data_in[55] la_data_in[56] la_data_in[57] la_data_in[58] la_data_in[59]
+ la_data_in[5] la_data_in[60] la_data_in[61] la_data_in[62] la_data_in[63] la_data_in[64]
+ la_data_in[65] la_data_in[66] la_data_in[67] la_data_in[68] la_data_in[69] la_data_in[6]
+ la_data_in[70] la_data_in[71] la_data_in[72] la_data_in[73] la_data_in[74] la_data_in[75]
+ la_data_in[76] la_data_in[77] la_data_in[78] la_data_in[79] la_data_in[7] la_data_in[80]
+ la_data_in[81] la_data_in[82] la_data_in[83] la_data_in[84] la_data_in[85] la_data_in[86]
+ la_data_in[87] la_data_in[88] la_data_in[89] la_data_in[8] la_data_in[90] la_data_in[91]
+ la_data_in[92] la_data_in[93] la_data_in[94] la_data_in[95] la_data_in[96] la_data_in[97]
+ la_data_in[98] la_data_in[99] la_data_in[9] la_data_out[0] la_data_out[100] la_data_out[101]
+ la_data_out[102] la_data_out[103] la_data_out[104] la_data_out[105] la_data_out[106]
+ la_data_out[107] la_data_out[108] la_data_out[109] la_data_out[10] la_data_out[110]
+ la_data_out[111] la_data_out[112] la_data_out[113] la_data_out[114] la_data_out[115]
+ la_data_out[116] la_data_out[117] la_data_out[118] la_data_out[119] la_data_out[11]
+ la_data_out[120] la_data_out[121] la_data_out[122] la_data_out[123] la_data_out[124]
+ la_data_out[125] la_data_out[126] la_data_out[127] la_data_out[12] la_data_out[13]
+ la_data_out[14] la_data_out[15] la_data_out[16] la_data_out[17] la_data_out[18]
+ la_data_out[19] la_data_out[1] la_data_out[20] la_data_out[21] la_data_out[22] la_data_out[23]
+ la_data_out[24] la_data_out[25] la_data_out[26] la_data_out[27] la_data_out[28]
+ la_data_out[29] la_data_out[2] la_data_out[30] la_data_out[31] la_data_out[32] la_data_out[33]
+ la_data_out[34] la_data_out[35] la_data_out[36] la_data_out[37] la_data_out[38]
+ la_data_out[39] la_data_out[3] la_data_out[40] la_data_out[41] la_data_out[42] la_data_out[43]
+ la_data_out[44] la_data_out[45] la_data_out[46] la_data_out[47] la_data_out[48]
+ la_data_out[49] la_data_out[4] la_data_out[50] la_data_out[51] la_data_out[52] la_data_out[53]
+ la_data_out[54] la_data_out[55] la_data_out[56] la_data_out[57] la_data_out[58]
+ la_data_out[59] la_data_out[5] la_data_out[60] la_data_out[61] la_data_out[62] la_data_out[63]
+ la_data_out[64] la_data_out[65] la_data_out[66] la_data_out[67] la_data_out[68]
+ la_data_out[69] la_data_out[6] la_data_out[70] la_data_out[71] la_data_out[72] la_data_out[73]
+ la_data_out[74] la_data_out[75] la_data_out[76] la_data_out[77] la_data_out[78]
+ la_data_out[79] la_data_out[7] la_data_out[80] la_data_out[81] la_data_out[82] la_data_out[83]
+ la_data_out[84] la_data_out[85] la_data_out[86] la_data_out[87] la_data_out[88]
+ la_data_out[89] la_data_out[8] la_data_out[90] la_data_out[91] la_data_out[92] la_data_out[93]
+ la_data_out[94] la_data_out[95] la_data_out[96] la_data_out[97] la_data_out[98]
+ la_data_out[99] la_data_out[9] la_oenb[0] la_oenb[100] la_oenb[101] la_oenb[102]
+ la_oenb[103] la_oenb[104] la_oenb[105] la_oenb[106] la_oenb[107] la_oenb[108] la_oenb[109]
+ la_oenb[10] la_oenb[110] la_oenb[111] la_oenb[112] la_oenb[113] la_oenb[114] la_oenb[115]
+ la_oenb[116] la_oenb[117] la_oenb[118] la_oenb[119] la_oenb[11] la_oenb[120] la_oenb[121]
+ la_oenb[122] la_oenb[123] la_oenb[124] la_oenb[125] la_oenb[126] la_oenb[127] la_oenb[12]
+ la_oenb[13] la_oenb[14] la_oenb[15] la_oenb[16] la_oenb[17] la_oenb[18] la_oenb[19]
+ la_oenb[1] la_oenb[20] la_oenb[21] la_oenb[22] la_oenb[23] la_oenb[24] la_oenb[25]
+ la_oenb[26] la_oenb[27] la_oenb[28] la_oenb[29] la_oenb[2] la_oenb[30] la_oenb[31]
+ la_oenb[32] la_oenb[33] la_oenb[34] la_oenb[35] la_oenb[36] la_oenb[37] la_oenb[38]
+ la_oenb[39] la_oenb[3] la_oenb[40] la_oenb[41] la_oenb[42] la_oenb[43] la_oenb[44]
+ la_oenb[45] la_oenb[46] la_oenb[47] la_oenb[48] la_oenb[49] la_oenb[4] la_oenb[50]
+ la_oenb[51] la_oenb[52] la_oenb[53] la_oenb[54] la_oenb[55] la_oenb[56] la_oenb[57]
+ la_oenb[58] la_oenb[59] la_oenb[5] la_oenb[60] la_oenb[61] la_oenb[62] la_oenb[63]
+ la_oenb[64] la_oenb[65] la_oenb[66] la_oenb[67] la_oenb[68] la_oenb[69] la_oenb[6]
+ la_oenb[70] la_oenb[71] la_oenb[72] la_oenb[73] la_oenb[74] la_oenb[75] la_oenb[76]
+ la_oenb[77] la_oenb[78] la_oenb[79] la_oenb[7] la_oenb[80] la_oenb[81] la_oenb[82]
+ la_oenb[83] la_oenb[84] la_oenb[85] la_oenb[86] la_oenb[87] la_oenb[88] la_oenb[89]
+ la_oenb[8] la_oenb[90] la_oenb[91] la_oenb[92] la_oenb[93] la_oenb[94] la_oenb[95]
+ la_oenb[96] la_oenb[97] la_oenb[98] la_oenb[99] la_oenb[9] user_clock2 user_irq[0]
+ user_irq[1] user_irq[2] vccd1 vccd2 vdda1 vdda2 vssa1 vssa2 vssd1 vssd2 wb_clk_i
+ wb_rst_i wbs_ack_o wbs_adr_i[0] wbs_adr_i[10] wbs_adr_i[11] wbs_adr_i[12] wbs_adr_i[13]
+ wbs_adr_i[14] wbs_adr_i[15] wbs_adr_i[16] wbs_adr_i[17] wbs_adr_i[18] wbs_adr_i[19]
+ wbs_adr_i[1] wbs_adr_i[20] wbs_adr_i[21] wbs_adr_i[22] wbs_adr_i[23] wbs_adr_i[24]
+ wbs_adr_i[25] wbs_adr_i[26] wbs_adr_i[27] wbs_adr_i[28] wbs_adr_i[29] wbs_adr_i[2]
+ wbs_adr_i[30] wbs_adr_i[31] wbs_adr_i[3] wbs_adr_i[4] wbs_adr_i[5] wbs_adr_i[6]
+ wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9] wbs_cyc_i wbs_dat_i[0] wbs_dat_i[10] wbs_dat_i[11]
+ wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14] wbs_dat_i[15] wbs_dat_i[16] wbs_dat_i[17]
+ wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1] wbs_dat_i[20] wbs_dat_i[21] wbs_dat_i[22]
+ wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25] wbs_dat_i[26] wbs_dat_i[27] wbs_dat_i[28]
+ wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30] wbs_dat_i[31] wbs_dat_i[3] wbs_dat_i[4]
+ wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8] wbs_dat_i[9] wbs_dat_o[0] wbs_dat_o[10]
+ wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13] wbs_dat_o[14] wbs_dat_o[15] wbs_dat_o[16]
+ wbs_dat_o[17] wbs_dat_o[18] wbs_dat_o[19] wbs_dat_o[1] wbs_dat_o[20] wbs_dat_o[21]
+ wbs_dat_o[22] wbs_dat_o[23] wbs_dat_o[24] wbs_dat_o[25] wbs_dat_o[26] wbs_dat_o[27]
+ wbs_dat_o[28] wbs_dat_o[29] wbs_dat_o[2] wbs_dat_o[30] wbs_dat_o[31] wbs_dat_o[3]
+ wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6] wbs_dat_o[7] wbs_dat_o[8] wbs_dat_o[9] wbs_sel_i[0]
+ wbs_sel_i[1] wbs_sel_i[2] wbs_sel_i[3] wbs_stb_i wbs_we_i
Xtune_player dso_tune design_clk rst_tune vccd1 vssd1 tune_player
Xposit_unit design_clk dsi_all\[0\] dsi_all\[1\] dsi_all\[2\] dso_posit\[0\] dso_posit\[1\]
+ dso_posit\[2\] dso_posit\[3\] rst_posit vccd1 vssd1 posit_unit
Xtt2_tholin_multiplexed_counter design_clk dso_counter\[0\] dso_counter\[10\] dso_counter\[11\]
+ dso_counter\[1\] dso_counter\[2\] dso_counter\[3\] dso_counter\[4\] dso_counter\[5\]
+ dso_counter\[6\] dso_counter\[7\] dso_counter\[8\] dso_counter\[9\] rst_counter
+ vccd1 vssd1 tt2_tholin_multiplexed_counter
Xwrapped_MC14500 design_clk dsi_all\[0\] dsi_all\[1\] dsi_all\[2\] dsi_all\[3\] dsi_all\[4\]
+ oeb_mc14500 dso_mc14500\[0\] dso_mc14500\[1\] dso_mc14500\[2\] dso_mc14500\[3\]
+ dso_mc14500\[4\] dso_mc14500\[5\] dso_mc14500\[6\] dso_mc14500\[7\] dso_mc14500\[8\]
+ rst_mc14500 vccd1 vssd1 wrapped_MC14500
Xproj_multiplexer design_clk dsi_all\[0\] dsi_all\[10\] dsi_all\[11\] dsi_all\[12\]
+ dsi_all\[13\] dsi_all\[14\] dsi_all\[15\] dsi_all\[16\] dsi_all\[17\] dsi_all\[18\]
+ dsi_all\[19\] dsi_all\[1\] dsi_all\[20\] dsi_all\[21\] dsi_all\[22\] dsi_all\[23\]
+ dsi_all\[24\] dsi_all\[25\] dsi_all\[26\] dsi_all\[27\] dsi_all\[2\] dsi_all\[3\]
+ dsi_all\[4\] dsi_all\[5\] dsi_all\[6\] dsi_all\[7\] dsi_all\[8\] dsi_all\[9\] dso_6502\[0\]
+ dso_6502\[10\] dso_6502\[11\] dso_6502\[12\] dso_6502\[13\] dso_6502\[14\] dso_6502\[15\]
+ dso_6502\[16\] dso_6502\[17\] dso_6502\[18\] dso_6502\[19\] dso_6502\[1\] dso_6502\[20\]
+ dso_6502\[21\] dso_6502\[22\] dso_6502\[23\] dso_6502\[24\] dso_6502\[25\] dso_6502\[26\]
+ dso_6502\[2\] dso_6502\[3\] dso_6502\[4\] dso_6502\[5\] dso_6502\[6\] dso_6502\[7\]
+ dso_6502\[8\] dso_6502\[9\] dso_LCD\[0\] dso_LCD\[1\] dso_LCD\[2\] dso_LCD\[3\]
+ dso_LCD\[4\] dso_LCD\[5\] dso_LCD\[6\] dso_LCD\[7\] dso_as1802\[0\] dso_as1802\[10\]
+ dso_as1802\[11\] dso_as1802\[12\] dso_as1802\[13\] dso_as1802\[14\] dso_as1802\[15\]
+ dso_as1802\[16\] dso_as1802\[17\] dso_as1802\[18\] dso_as1802\[19\] dso_as1802\[1\]
+ dso_as1802\[20\] dso_as1802\[21\] dso_as1802\[22\] dso_as1802\[23\] dso_as1802\[24\]
+ dso_as1802\[25\] dso_as1802\[26\] dso_as1802\[2\] dso_as1802\[3\] dso_as1802\[4\]
+ dso_as1802\[5\] dso_as1802\[6\] dso_as1802\[7\] dso_as1802\[8\] dso_as1802\[9\]
+ dso_as2650\[0\] dso_as2650\[10\] dso_as2650\[11\] dso_as2650\[12\] dso_as2650\[13\]
+ dso_as2650\[14\] dso_as2650\[15\] dso_as2650\[16\] dso_as2650\[17\] dso_as2650\[18\]
+ dso_as2650\[19\] dso_as2650\[1\] dso_as2650\[20\] dso_as2650\[21\] dso_as2650\[22\]
+ dso_as2650\[23\] dso_as2650\[24\] dso_as2650\[25\] dso_as2650\[26\] dso_as2650\[2\]
+ dso_as2650\[3\] dso_as2650\[4\] dso_as2650\[5\] dso_as2650\[6\] dso_as2650\[7\]
+ dso_as2650\[8\] dso_as2650\[9\] dso_as512512512\[0\] dso_as512512512\[10\] dso_as512512512\[11\]
+ dso_as512512512\[12\] dso_as512512512\[13\] dso_as512512512\[14\] dso_as512512512\[15\]
+ dso_as512512512\[16\] dso_as512512512\[17\] dso_as512512512\[18\] dso_as512512512\[19\]
+ dso_as512512512\[1\] dso_as512512512\[20\] dso_as512512512\[21\] dso_as512512512\[22\]
+ dso_as512512512\[23\] dso_as512512512\[24\] dso_as512512512\[25\] dso_as512512512\[26\]
+ dso_as512512512\[27\] dso_as512512512\[2\] dso_as512512512\[3\] dso_as512512512\[4\]
+ dso_as512512512\[5\] dso_as512512512\[6\] dso_as512512512\[7\] dso_as512512512\[8\]
+ dso_as512512512\[9\] dso_as5401\[0\] dso_as5401\[10\] dso_as5401\[11\] dso_as5401\[12\]
+ dso_as5401\[13\] dso_as5401\[14\] dso_as5401\[15\] dso_as5401\[16\] dso_as5401\[17\]
+ dso_as5401\[18\] dso_as5401\[19\] dso_as5401\[1\] dso_as5401\[20\] dso_as5401\[21\]
+ dso_as5401\[22\] dso_as5401\[23\] dso_as5401\[24\] dso_as5401\[25\] dso_as5401\[26\]
+ dso_as5401\[2\] dso_as5401\[3\] dso_as5401\[4\] dso_as5401\[5\] dso_as5401\[6\]
+ dso_as5401\[7\] dso_as5401\[8\] dso_as5401\[9\] dso_counter\[0\] dso_counter\[10\]
+ dso_counter\[11\] dso_counter\[1\] dso_counter\[2\] dso_counter\[3\] dso_counter\[4\]
+ dso_counter\[5\] dso_counter\[6\] dso_counter\[7\] dso_counter\[8\] dso_counter\[9\]
+ dso_diceroll\[0\] dso_diceroll\[1\] dso_diceroll\[2\] dso_diceroll\[3\] dso_diceroll\[4\]
+ dso_diceroll\[5\] dso_diceroll\[6\] dso_diceroll\[7\] dso_mc14500\[0\] dso_mc14500\[1\]
+ dso_mc14500\[2\] dso_mc14500\[3\] dso_mc14500\[4\] dso_mc14500\[5\] dso_mc14500\[6\]
+ dso_mc14500\[7\] dso_mc14500\[8\] dso_multiplier\[0\] dso_multiplier\[1\] dso_multiplier\[2\]
+ dso_multiplier\[3\] dso_multiplier\[4\] dso_multiplier\[5\] dso_multiplier\[6\]
+ dso_multiplier\[7\] dso_posit\[0\] dso_posit\[1\] dso_posit\[2\] dso_posit\[3\]
+ dso_tbb1143\[0\] dso_tbb1143\[1\] dso_tbb1143\[2\] dso_tbb1143\[3\] dso_tbb1143\[4\]
+ dso_tbb1143\[5\] dso_tbb1143\[6\] dso_tbb1143\[7\] dso_tune io_in[0] io_in[10] io_in[11]
+ io_in[12] io_in[13] io_in[14] io_in[15] io_in[16] io_in[17] io_in[18] io_in[19]
+ io_in[1] io_in[20] io_in[21] io_in[22] io_in[23] io_in[24] io_in[25] io_in[26] io_in[27]
+ io_in[28] io_in[29] io_in[2] io_in[30] io_in[31] io_in[32] io_in[33] io_in[34] io_in[35]
+ io_in[36] io_in[37] io_in[3] io_in[4] io_in[5] io_in[6] io_in[7] io_in[8] io_in[9]
+ io_oeb[0] io_oeb[10] io_oeb[11] io_oeb[12] io_oeb[13] io_oeb[14] io_oeb[15] io_oeb[16]
+ io_oeb[17] io_oeb[18] io_oeb[19] io_oeb[1] io_oeb[20] io_oeb[21] io_oeb[22] io_oeb[23]
+ io_oeb[24] io_oeb[25] io_oeb[26] io_oeb[27] io_oeb[28] io_oeb[29] io_oeb[2] io_oeb[30]
+ io_oeb[31] io_oeb[32] io_oeb[33] io_oeb[34] io_oeb[35] io_oeb[36] io_oeb[37] io_oeb[3]
+ io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7] io_oeb[8] io_oeb[9] io_out[0] io_out[10]
+ io_out[11] io_out[12] io_out[13] io_out[14] io_out[15] io_out[16] io_out[17] io_out[18]
+ io_out[19] io_out[1] io_out[20] io_out[21] io_out[22] io_out[23] io_out[24] io_out[25]
+ io_out[26] io_out[27] io_out[28] io_out[29] io_out[2] io_out[30] io_out[31] io_out[32]
+ io_out[33] io_out[34] io_out[35] io_out[36] io_out[37] io_out[3] io_out[4] io_out[5]
+ io_out[6] io_out[7] io_out[8] io_out[9] oeb_6502 oeb_as1802 oeb_as2650 oeb_as512512512
+ oeb_as5401 oeb_mc14500 rst_6502 rst_LCD rst_as1802 rst_as2650 rst_as512512512 rst_as5401
+ rst_counter rst_diceroll rst_mc14500 rst_posit rst_tbb1143 rst_tune vccd1 vssd1
+ wb_clk_i wb_rst_i wbs_ack_o wbs_adr_i[0] wbs_adr_i[10] wbs_adr_i[11] wbs_adr_i[12]
+ wbs_adr_i[13] wbs_adr_i[14] wbs_adr_i[15] wbs_adr_i[16] wbs_adr_i[17] wbs_adr_i[18]
+ wbs_adr_i[19] wbs_adr_i[1] wbs_adr_i[20] wbs_adr_i[21] wbs_adr_i[22] wbs_adr_i[23]
+ wbs_adr_i[24] wbs_adr_i[25] wbs_adr_i[26] wbs_adr_i[27] wbs_adr_i[28] wbs_adr_i[29]
+ wbs_adr_i[2] wbs_adr_i[30] wbs_adr_i[31] wbs_adr_i[3] wbs_adr_i[4] wbs_adr_i[5]
+ wbs_adr_i[6] wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9] wbs_cyc_i wbs_dat_i[0] wbs_dat_i[10]
+ wbs_dat_i[11] wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14] wbs_dat_i[15] wbs_dat_i[16]
+ wbs_dat_i[17] wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1] wbs_dat_i[20] wbs_dat_i[21]
+ wbs_dat_i[22] wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25] wbs_dat_i[26] wbs_dat_i[27]
+ wbs_dat_i[28] wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30] wbs_dat_i[31] wbs_dat_i[3]
+ wbs_dat_i[4] wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8] wbs_dat_i[9] wbs_dat_o[0]
+ wbs_dat_o[10] wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13] wbs_dat_o[14] wbs_dat_o[15]
+ wbs_dat_o[16] wbs_dat_o[17] wbs_dat_o[18] wbs_dat_o[19] wbs_dat_o[1] wbs_dat_o[20]
+ wbs_dat_o[21] wbs_dat_o[22] wbs_dat_o[23] wbs_dat_o[24] wbs_dat_o[25] wbs_dat_o[26]
+ wbs_dat_o[27] wbs_dat_o[28] wbs_dat_o[29] wbs_dat_o[2] wbs_dat_o[30] wbs_dat_o[31]
+ wbs_dat_o[3] wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6] wbs_dat_o[7] wbs_dat_o[8] wbs_dat_o[9]
+ wbs_stb_i wbs_we_i multiplexer
Xtt2_tholin_multiplier dsi_all\[0\] dsi_all\[1\] dsi_all\[2\] dsi_all\[3\] dsi_all\[4\]
+ dsi_all\[5\] dsi_all\[6\] dsi_all\[7\] dso_multiplier\[0\] dso_multiplier\[1\] dso_multiplier\[2\]
+ dso_multiplier\[3\] dso_multiplier\[4\] dso_multiplier\[5\] dso_multiplier\[6\]
+ dso_multiplier\[7\] vccd1 vssd1 tt2_tholin_multiplier
Xtt2_tholin_diceroll design_clk dsi_all\[0\] dso_diceroll\[0\] dso_diceroll\[1\] dso_diceroll\[2\]
+ dso_diceroll\[3\] dso_diceroll\[4\] dso_diceroll\[5\] dso_diceroll\[6\] dso_diceroll\[7\]
+ rst_diceroll vccd1 vssd1 tt2_tholin_diceroll
Xtholin_avalonsemi_tbb1143 design_clk dsi_all\[0\] dsi_all\[1\] dsi_all\[2\] dsi_all\[3\]
+ dsi_all\[4\] dsi_all\[5\] dso_tbb1143\[0\] dso_tbb1143\[1\] dso_tbb1143\[2\] dso_tbb1143\[3\]
+ dso_tbb1143\[4\] dso_tbb1143\[5\] dso_tbb1143\[6\] dso_tbb1143\[7\] rst_tbb1143
+ vccd1 vssd1 tholin_avalonsemi_tbb1143
Xtholin_avalonsemi_5401 design_clk dsi_all\[0\] dsi_all\[1\] dsi_all\[2\] dsi_all\[3\]
+ dsi_all\[4\] dsi_all\[5\] dsi_all\[6\] dsi_all\[7\] dsi_all\[8\] dsi_all\[9\] oeb_as5401
+ dso_as5401\[0\] dso_as5401\[10\] dso_as5401\[11\] dso_as5401\[12\] dso_as5401\[13\]
+ dso_as5401\[14\] dso_as5401\[15\] dso_as5401\[16\] dso_as5401\[17\] dso_as5401\[18\]
+ dso_as5401\[19\] dso_as5401\[1\] dso_as5401\[20\] dso_as5401\[21\] dso_as5401\[22\]
+ dso_as5401\[23\] dso_as5401\[24\] dso_as5401\[25\] dso_as5401\[26\] dso_as5401\[2\]
+ dso_as5401\[3\] dso_as5401\[4\] dso_as5401\[5\] dso_as5401\[6\] dso_as5401\[7\]
+ dso_as5401\[8\] dso_as5401\[9\] rst_as5401 vccd1 vssd1 tholin_avalonsemi_5401
Xwrapped_vgatest design_clk dsi_all\[0\] wrapped_vgatest/io_out[0] wrapped_vgatest/io_out[1]
+ wrapped_vgatest/io_out[2] wrapped_vgatest/io_out[3] wrapped_vgatest/io_out[4] wrapped_vgatest/io_out[5]
+ wrapped_vgatest/io_out[6] wrapped_vgatest/io_out[7] wrapped_vgatest/io_out[8] wrapped_vgatest/io_out[9]
+ wrapped_vgatest/rst vccd1 vssd1 wrapped_vgatest
Xwrapped_as512512512 design_clk dsi_all\[0\] dsi_all\[10\] dsi_all\[11\] dsi_all\[12\]
+ dsi_all\[13\] dsi_all\[14\] dsi_all\[15\] dsi_all\[16\] dsi_all\[17\] dsi_all\[18\]
+ dsi_all\[19\] dsi_all\[1\] dsi_all\[20\] dsi_all\[21\] dsi_all\[22\] dsi_all\[23\]
+ dsi_all\[24\] dsi_all\[25\] dsi_all\[26\] dsi_all\[2\] dsi_all\[3\] dsi_all\[4\]
+ dsi_all\[5\] dsi_all\[6\] dsi_all\[7\] dsi_all\[8\] dsi_all\[9\] oeb_as512512512
+ dso_as512512512\[0\] dso_as512512512\[10\] dso_as512512512\[11\] dso_as512512512\[12\]
+ dso_as512512512\[13\] dso_as512512512\[14\] dso_as512512512\[15\] dso_as512512512\[16\]
+ dso_as512512512\[17\] dso_as512512512\[18\] dso_as512512512\[19\] dso_as512512512\[1\]
+ dso_as512512512\[20\] dso_as512512512\[21\] dso_as512512512\[22\] dso_as512512512\[23\]
+ dso_as512512512\[24\] dso_as512512512\[25\] dso_as512512512\[26\] dso_as512512512\[27\]
+ dso_as512512512\[2\] dso_as512512512\[3\] dso_as512512512\[4\] dso_as512512512\[5\]
+ dso_as512512512\[6\] dso_as512512512\[7\] dso_as512512512\[8\] dso_as512512512\[9\]
+ rst_as512512512 vccd1 vssd1 wrapped_as512512512
Xwrapped_as1802 design_clk dsi_all\[0\] dsi_all\[10\] dsi_all\[11\] dsi_all\[12\]
+ dsi_all\[1\] dsi_all\[2\] dsi_all\[3\] dsi_all\[4\] dsi_all\[5\] dsi_all\[6\] dsi_all\[7\]
+ dsi_all\[8\] dsi_all\[9\] oeb_as1802 dso_as1802\[0\] dso_as1802\[10\] dso_as1802\[11\]
+ dso_as1802\[12\] dso_as1802\[13\] dso_as1802\[14\] dso_as1802\[15\] dso_as1802\[16\]
+ dso_as1802\[17\] dso_as1802\[18\] dso_as1802\[19\] dso_as1802\[1\] dso_as1802\[20\]
+ dso_as1802\[21\] dso_as1802\[22\] dso_as1802\[23\] dso_as1802\[24\] dso_as1802\[25\]
+ dso_as1802\[26\] dso_as1802\[2\] dso_as1802\[3\] dso_as1802\[4\] dso_as1802\[5\]
+ dso_as1802\[6\] dso_as1802\[7\] dso_as1802\[8\] dso_as1802\[9\] rst_as1802 vccd1
+ vssd1 wrapped_as1802
Xwrapped_6502 design_clk dsi_all\[0\] dsi_all\[1\] dsi_all\[2\] dsi_all\[3\] dsi_all\[4\]
+ dsi_all\[5\] dsi_all\[6\] dsi_all\[7\] dsi_all\[8\] dsi_all\[9\] oeb_6502 dso_6502\[0\]
+ dso_6502\[10\] dso_6502\[11\] dso_6502\[12\] dso_6502\[13\] dso_6502\[14\] dso_6502\[15\]
+ dso_6502\[16\] dso_6502\[17\] dso_6502\[18\] dso_6502\[19\] dso_6502\[1\] dso_6502\[20\]
+ dso_6502\[21\] dso_6502\[22\] dso_6502\[23\] dso_6502\[24\] dso_6502\[25\] dso_6502\[26\]
+ dso_6502\[2\] dso_6502\[3\] dso_6502\[4\] dso_6502\[5\] dso_6502\[6\] dso_6502\[7\]
+ dso_6502\[8\] dso_6502\[9\] rst_6502 vccd1 vssd1 wrapped_6502
Xtt2_tholin_namebadge design_clk dsi_all\[8\] dsi_all\[9\] dsi_all\[10\] tt2_tholin_namebadge/io_oeb[0]
+ tt2_tholin_namebadge/io_oeb[10] tt2_tholin_namebadge/io_oeb[11] tt2_tholin_namebadge/io_oeb[12]
+ tt2_tholin_namebadge/io_oeb[13] tt2_tholin_namebadge/io_oeb[14] tt2_tholin_namebadge/io_oeb[15]
+ tt2_tholin_namebadge/io_oeb[16] tt2_tholin_namebadge/io_oeb[17] tt2_tholin_namebadge/io_oeb[18]
+ tt2_tholin_namebadge/io_oeb[19] tt2_tholin_namebadge/io_oeb[1] tt2_tholin_namebadge/io_oeb[20]
+ tt2_tholin_namebadge/io_oeb[21] tt2_tholin_namebadge/io_oeb[22] tt2_tholin_namebadge/io_oeb[23]
+ tt2_tholin_namebadge/io_oeb[24] tt2_tholin_namebadge/io_oeb[25] tt2_tholin_namebadge/io_oeb[26]
+ tt2_tholin_namebadge/io_oeb[2] tt2_tholin_namebadge/io_oeb[3] tt2_tholin_namebadge/io_oeb[4]
+ tt2_tholin_namebadge/io_oeb[5] tt2_tholin_namebadge/io_oeb[6] tt2_tholin_namebadge/io_oeb[7]
+ tt2_tholin_namebadge/io_oeb[8] tt2_tholin_namebadge/io_oeb[9] dso_LCD\[0\] dso_LCD\[1\]
+ dso_LCD\[2\] dso_LCD\[3\] dso_LCD\[4\] dso_LCD\[5\] dso_LCD\[6\] dso_LCD\[7\] rst_LCD
+ vccd1 vssd1 tt2_tholin_namebadge
Xwrapped_as2650 design_clk dsi_all\[0\] dsi_all\[1\] dsi_all\[2\] dsi_all\[3\] dsi_all\[4\]
+ dsi_all\[5\] dsi_all\[6\] dsi_all\[7\] dsi_all\[27\] oeb_as2650 dso_as2650\[0\]
+ dso_as2650\[10\] dso_as2650\[11\] dso_as2650\[12\] dso_as2650\[13\] dso_as2650\[14\]
+ dso_as2650\[15\] dso_as2650\[16\] dso_as2650\[17\] dso_as2650\[18\] dso_as2650\[19\]
+ dso_as2650\[1\] dso_as2650\[20\] dso_as2650\[21\] dso_as2650\[22\] dso_as2650\[23\]
+ dso_as2650\[24\] dso_as2650\[25\] dso_as2650\[26\] dso_as2650\[2\] dso_as2650\[3\]
+ dso_as2650\[4\] dso_as2650\[5\] dso_as2650\[6\] dso_as2650\[7\] dso_as2650\[8\]
+ dso_as2650\[9\] rst_as2650 vccd1 vssd1 wrapped_as2650
.ends

