magic
tech sky130B
magscale 1 2
timestamp 1674825087
<< obsli1 >>
rect 1104 2159 16836 15793
<< obsm1 >>
rect 1104 2128 16995 15904
<< metal2 >>
rect 4434 17200 4490 18000
rect 13450 17200 13506 18000
<< obsm2 >>
rect 1398 17144 4378 17354
rect 4546 17144 13394 17354
rect 13562 17144 16989 17354
rect 1398 711 16989 17144
<< metal3 >>
rect 0 17144 800 17264
rect 0 15648 800 15768
rect 0 14152 800 14272
rect 0 12656 800 12776
rect 0 11160 800 11280
rect 0 9664 800 9784
rect 0 8168 800 8288
rect 0 6672 800 6792
rect 0 5176 800 5296
rect 0 3680 800 3800
rect 0 2184 800 2304
rect 0 688 800 808
<< obsm3 >>
rect 880 17064 16993 17237
rect 800 15848 16993 17064
rect 880 15568 16993 15848
rect 800 14352 16993 15568
rect 880 14072 16993 14352
rect 800 12856 16993 14072
rect 880 12576 16993 12856
rect 800 11360 16993 12576
rect 880 11080 16993 11360
rect 800 9864 16993 11080
rect 880 9584 16993 9864
rect 800 8368 16993 9584
rect 880 8088 16993 8368
rect 800 6872 16993 8088
rect 880 6592 16993 6872
rect 800 5376 16993 6592
rect 880 5096 16993 5376
rect 800 3880 16993 5096
rect 880 3600 16993 3880
rect 800 2384 16993 3600
rect 880 2104 16993 2384
rect 800 888 16993 2104
rect 880 715 16993 888
<< metal4 >>
rect 2910 2128 3230 15824
rect 4876 2128 5196 15824
rect 6843 2128 7163 15824
rect 8809 2128 9129 15824
rect 10776 2128 11096 15824
rect 12742 2128 13062 15824
rect 14709 2128 15029 15824
rect 16675 2128 16995 15824
<< obsm4 >>
rect 3371 3979 3437 9757
<< labels >>
rlabel metal2 s 4434 17200 4490 18000 6 clk
port 1 nsew signal input
rlabel metal3 s 0 688 800 808 6 io_out[0]
port 2 nsew signal output
rlabel metal3 s 0 15648 800 15768 6 io_out[10]
port 3 nsew signal output
rlabel metal3 s 0 17144 800 17264 6 io_out[11]
port 4 nsew signal output
rlabel metal3 s 0 2184 800 2304 6 io_out[1]
port 5 nsew signal output
rlabel metal3 s 0 3680 800 3800 6 io_out[2]
port 6 nsew signal output
rlabel metal3 s 0 5176 800 5296 6 io_out[3]
port 7 nsew signal output
rlabel metal3 s 0 6672 800 6792 6 io_out[4]
port 8 nsew signal output
rlabel metal3 s 0 8168 800 8288 6 io_out[5]
port 9 nsew signal output
rlabel metal3 s 0 9664 800 9784 6 io_out[6]
port 10 nsew signal output
rlabel metal3 s 0 11160 800 11280 6 io_out[7]
port 11 nsew signal output
rlabel metal3 s 0 12656 800 12776 6 io_out[8]
port 12 nsew signal output
rlabel metal3 s 0 14152 800 14272 6 io_out[9]
port 13 nsew signal output
rlabel metal2 s 13450 17200 13506 18000 6 rst
port 14 nsew signal input
rlabel metal4 s 2910 2128 3230 15824 6 vccd1
port 15 nsew power bidirectional
rlabel metal4 s 6843 2128 7163 15824 6 vccd1
port 15 nsew power bidirectional
rlabel metal4 s 10776 2128 11096 15824 6 vccd1
port 15 nsew power bidirectional
rlabel metal4 s 14709 2128 15029 15824 6 vccd1
port 15 nsew power bidirectional
rlabel metal4 s 4876 2128 5196 15824 6 vssd1
port 16 nsew ground bidirectional
rlabel metal4 s 8809 2128 9129 15824 6 vssd1
port 16 nsew ground bidirectional
rlabel metal4 s 12742 2128 13062 15824 6 vssd1
port 16 nsew ground bidirectional
rlabel metal4 s 16675 2128 16995 15824 6 vssd1
port 16 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 18000 18000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 822340
string GDS_FILE /media/lucah/e6042058-84c8-448b-be8a-b40bc065b34b/TMBoC/openlane/MultiplexedCounter/runs/23_01_27_14_09/results/signoff/tt2_tholin_multiplexed_counter.magic.gds
string GDS_START 273440
<< end >>

