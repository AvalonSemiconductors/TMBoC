VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO wrapped_6502
  CLASS BLOCK ;
  FOREIGN wrapped_6502 ;
  ORIGIN 0.000 0.000 ;
  SIZE 225.000 BY 225.000 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 221.000 194.220 225.000 195.420 ;
    END
  END clk
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 221.000 10.620 225.000 11.820 ;
    END
  END io_in[0]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 221.000 28.980 225.000 30.180 ;
    END
  END io_in[1]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 221.000 47.340 225.000 48.540 ;
    END
  END io_in[2]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 221.000 65.700 225.000 66.900 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 221.000 84.060 225.000 85.260 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 221.000 102.420 225.000 103.620 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 221.000 120.780 225.000 121.980 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 221.000 139.140 225.000 140.340 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 221.000 157.500 225.000 158.700 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 221.000 175.860 225.000 177.060 ;
    END
  END io_in[9]
  PIN io_oeb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 217.530 221.000 218.090 225.000 ;
    END
  END io_oeb
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.390 221.000 6.950 225.000 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 84.590 221.000 85.150 225.000 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 92.410 221.000 92.970 225.000 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 100.230 221.000 100.790 225.000 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.050 221.000 108.610 225.000 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 115.870 221.000 116.430 225.000 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 123.690 221.000 124.250 225.000 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 131.510 221.000 132.070 225.000 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.330 221.000 139.890 225.000 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 147.150 221.000 147.710 225.000 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 154.970 221.000 155.530 225.000 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.210 221.000 14.770 225.000 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 162.790 221.000 163.350 225.000 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.610 221.000 171.170 225.000 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 178.430 221.000 178.990 225.000 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.250 221.000 186.810 225.000 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 194.070 221.000 194.630 225.000 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 201.890 221.000 202.450 225.000 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.710 221.000 210.270 225.000 ;
    END
  END io_out[26]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.030 221.000 22.590 225.000 ;
    END
  END io_out[2]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.850 221.000 30.410 225.000 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.670 221.000 38.230 225.000 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.490 221.000 46.050 225.000 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.310 221.000 53.870 225.000 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.130 221.000 61.690 225.000 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.950 221.000 69.510 225.000 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.770 221.000 77.330 225.000 ;
    END
  END io_out[9]
  PIN rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 221.000 212.580 225.000 213.780 ;
    END
  END rst
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 212.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 212.400 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 212.400 ;
    END
  END vssd1
  OBS
      LAYER nwell ;
        RECT 5.330 208.025 219.610 210.855 ;
        RECT 5.330 202.585 219.610 205.415 ;
        RECT 5.330 197.145 219.610 199.975 ;
        RECT 5.330 191.705 219.610 194.535 ;
        RECT 5.330 186.265 219.610 189.095 ;
        RECT 5.330 180.825 219.610 183.655 ;
        RECT 5.330 175.385 219.610 178.215 ;
        RECT 5.330 169.945 219.610 172.775 ;
        RECT 5.330 164.505 219.610 167.335 ;
        RECT 5.330 159.065 219.610 161.895 ;
        RECT 5.330 153.625 219.610 156.455 ;
        RECT 5.330 148.185 219.610 151.015 ;
        RECT 5.330 142.745 219.610 145.575 ;
        RECT 5.330 137.305 219.610 140.135 ;
        RECT 5.330 131.865 219.610 134.695 ;
        RECT 5.330 126.425 219.610 129.255 ;
        RECT 5.330 120.985 219.610 123.815 ;
        RECT 5.330 115.545 219.610 118.375 ;
        RECT 5.330 110.105 219.610 112.935 ;
        RECT 5.330 104.665 219.610 107.495 ;
        RECT 5.330 99.225 219.610 102.055 ;
        RECT 5.330 93.785 219.610 96.615 ;
        RECT 5.330 88.345 219.610 91.175 ;
        RECT 5.330 82.905 219.610 85.735 ;
        RECT 5.330 77.465 219.610 80.295 ;
        RECT 5.330 72.025 219.610 74.855 ;
        RECT 5.330 66.585 219.610 69.415 ;
        RECT 5.330 61.145 219.610 63.975 ;
        RECT 5.330 55.705 219.610 58.535 ;
        RECT 5.330 50.265 219.610 53.095 ;
        RECT 5.330 44.825 219.610 47.655 ;
        RECT 5.330 39.385 219.610 42.215 ;
        RECT 5.330 33.945 219.610 36.775 ;
        RECT 5.330 28.505 219.610 31.335 ;
        RECT 5.330 23.065 219.610 25.895 ;
        RECT 5.330 17.625 219.610 20.455 ;
        RECT 5.330 12.185 219.610 15.015 ;
      LAYER li1 ;
        RECT 5.520 10.795 219.420 212.245 ;
      LAYER met1 ;
        RECT 5.520 10.640 220.270 220.620 ;
      LAYER met2 ;
        RECT 7.230 220.720 13.930 221.000 ;
        RECT 15.050 220.720 21.750 221.000 ;
        RECT 22.870 220.720 29.570 221.000 ;
        RECT 30.690 220.720 37.390 221.000 ;
        RECT 38.510 220.720 45.210 221.000 ;
        RECT 46.330 220.720 53.030 221.000 ;
        RECT 54.150 220.720 60.850 221.000 ;
        RECT 61.970 220.720 68.670 221.000 ;
        RECT 69.790 220.720 76.490 221.000 ;
        RECT 77.610 220.720 84.310 221.000 ;
        RECT 85.430 220.720 92.130 221.000 ;
        RECT 93.250 220.720 99.950 221.000 ;
        RECT 101.070 220.720 107.770 221.000 ;
        RECT 108.890 220.720 115.590 221.000 ;
        RECT 116.710 220.720 123.410 221.000 ;
        RECT 124.530 220.720 131.230 221.000 ;
        RECT 132.350 220.720 139.050 221.000 ;
        RECT 140.170 220.720 146.870 221.000 ;
        RECT 147.990 220.720 154.690 221.000 ;
        RECT 155.810 220.720 162.510 221.000 ;
        RECT 163.630 220.720 170.330 221.000 ;
        RECT 171.450 220.720 178.150 221.000 ;
        RECT 179.270 220.720 185.970 221.000 ;
        RECT 187.090 220.720 193.790 221.000 ;
        RECT 194.910 220.720 201.610 221.000 ;
        RECT 202.730 220.720 209.430 221.000 ;
        RECT 210.550 220.720 217.250 221.000 ;
        RECT 218.370 220.720 220.250 221.000 ;
        RECT 6.540 10.695 220.250 220.720 ;
      LAYER met3 ;
        RECT 21.050 212.180 220.600 213.345 ;
        RECT 21.050 195.820 221.000 212.180 ;
        RECT 21.050 193.820 220.600 195.820 ;
        RECT 21.050 177.460 221.000 193.820 ;
        RECT 21.050 175.460 220.600 177.460 ;
        RECT 21.050 159.100 221.000 175.460 ;
        RECT 21.050 157.100 220.600 159.100 ;
        RECT 21.050 140.740 221.000 157.100 ;
        RECT 21.050 138.740 220.600 140.740 ;
        RECT 21.050 122.380 221.000 138.740 ;
        RECT 21.050 120.380 220.600 122.380 ;
        RECT 21.050 104.020 221.000 120.380 ;
        RECT 21.050 102.020 220.600 104.020 ;
        RECT 21.050 85.660 221.000 102.020 ;
        RECT 21.050 83.660 220.600 85.660 ;
        RECT 21.050 67.300 221.000 83.660 ;
        RECT 21.050 65.300 220.600 67.300 ;
        RECT 21.050 48.940 221.000 65.300 ;
        RECT 21.050 46.940 220.600 48.940 ;
        RECT 21.050 30.580 221.000 46.940 ;
        RECT 21.050 28.580 220.600 30.580 ;
        RECT 21.050 12.220 221.000 28.580 ;
        RECT 21.050 10.715 220.600 12.220 ;
      LAYER met4 ;
        RECT 122.655 56.615 174.240 199.745 ;
        RECT 176.640 56.615 206.705 199.745 ;
  END
END wrapped_6502
END LIBRARY

