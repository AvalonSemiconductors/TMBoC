magic
tech sky130B
magscale 1 2
timestamp 1674824561
<< viali >>
rect 9781 21981 9815 22015
rect 13093 21981 13127 22015
rect 13553 21981 13587 22015
rect 15117 21981 15151 22015
rect 17693 21981 17727 22015
rect 18153 21981 18187 22015
rect 22661 21981 22695 22015
rect 23121 21981 23155 22015
rect 7113 21913 7147 21947
rect 7757 21913 7791 21947
rect 9321 21913 9355 21947
rect 10048 21913 10082 21947
rect 12826 21913 12860 21947
rect 14289 21913 14323 21947
rect 14473 21913 14507 21947
rect 7665 21845 7699 21879
rect 11161 21845 11195 21879
rect 11713 21845 11747 21879
rect 13737 21845 13771 21879
rect 14657 21845 14691 21879
rect 17509 21845 17543 21879
rect 22477 21845 22511 21879
rect 12848 21573 12882 21607
rect 13553 21573 13587 21607
rect 7777 21505 7811 21539
rect 10048 21505 10082 21539
rect 13737 21505 13771 21539
rect 14657 21505 14691 21539
rect 14841 21505 14875 21539
rect 8033 21437 8067 21471
rect 9781 21437 9815 21471
rect 13093 21437 13127 21471
rect 13829 21437 13863 21471
rect 14197 21437 14231 21471
rect 11713 21369 11747 21403
rect 6653 21301 6687 21335
rect 11161 21301 11195 21335
rect 14749 21301 14783 21335
rect 11713 21097 11747 21131
rect 13001 21029 13035 21063
rect 13461 20961 13495 20995
rect 6285 20893 6319 20927
rect 6745 20893 6779 20927
rect 13369 20893 13403 20927
rect 6040 20825 6074 20859
rect 7012 20825 7046 20859
rect 10425 20825 10459 20859
rect 4905 20757 4939 20791
rect 8125 20757 8159 20791
rect 13093 20553 13127 20587
rect 10916 20485 10950 20519
rect 5374 20417 5408 20451
rect 5641 20417 5675 20451
rect 7205 20417 7239 20451
rect 7461 20417 7495 20451
rect 11161 20417 11195 20451
rect 12909 20417 12943 20451
rect 13093 20417 13127 20451
rect 4261 20213 4295 20247
rect 8585 20213 8619 20247
rect 9781 20213 9815 20247
rect 11713 20213 11747 20247
rect 11161 19873 11195 19907
rect 3985 19805 4019 19839
rect 8217 19805 8251 19839
rect 13001 19805 13035 19839
rect 4252 19737 4286 19771
rect 7972 19737 8006 19771
rect 10894 19737 10928 19771
rect 12756 19737 12790 19771
rect 5365 19669 5399 19703
rect 6837 19669 6871 19703
rect 9781 19669 9815 19703
rect 11621 19669 11655 19703
rect 3709 19465 3743 19499
rect 7113 19465 7147 19499
rect 4844 19397 4878 19431
rect 7665 19397 7699 19431
rect 5089 19329 5123 19363
rect 8953 19125 8987 19159
rect 2513 18921 2547 18955
rect 18245 18921 18279 18955
rect 6837 18785 6871 18819
rect 11713 18785 11747 18819
rect 2329 18717 2363 18751
rect 6377 18717 6411 18751
rect 9321 18717 9355 18751
rect 11437 18717 11471 18751
rect 18429 18717 18463 18751
rect 6110 18649 6144 18683
rect 7104 18649 7138 18683
rect 4997 18581 5031 18615
rect 8217 18581 8251 18615
rect 9137 18581 9171 18615
rect 10333 18581 10367 18615
rect 12265 18581 12299 18615
rect 4638 18241 4672 18275
rect 7380 18241 7414 18275
rect 9781 18241 9815 18275
rect 10048 18241 10082 18275
rect 12265 18241 12299 18275
rect 4905 18173 4939 18207
rect 7113 18173 7147 18207
rect 11161 18105 11195 18139
rect 3525 18037 3559 18071
rect 8493 18037 8527 18071
rect 11805 18037 11839 18071
rect 5549 17833 5583 17867
rect 8309 17833 8343 17867
rect 2053 17629 2087 17663
rect 7481 17629 7515 17663
rect 11253 17629 11287 17663
rect 11713 17629 11747 17663
rect 2320 17561 2354 17595
rect 7021 17561 7055 17595
rect 11008 17561 11042 17595
rect 11980 17561 12014 17595
rect 3433 17493 3467 17527
rect 7665 17493 7699 17527
rect 9873 17493 9907 17527
rect 13093 17493 13127 17527
rect 3258 17153 3292 17187
rect 3525 17153 3559 17187
rect 3985 17153 4019 17187
rect 4252 17153 4286 17187
rect 7021 17153 7055 17187
rect 7288 17153 7322 17187
rect 9781 17153 9815 17187
rect 10048 17153 10082 17187
rect 11161 17017 11195 17051
rect 2145 16949 2179 16983
rect 5365 16949 5399 16983
rect 8401 16949 8435 16983
rect 11805 16949 11839 16983
rect 2513 16745 2547 16779
rect 4629 16609 4663 16643
rect 8309 16609 8343 16643
rect 10057 16609 10091 16643
rect 2697 16541 2731 16575
rect 3433 16541 3467 16575
rect 16313 16541 16347 16575
rect 4874 16473 4908 16507
rect 8042 16473 8076 16507
rect 10324 16473 10358 16507
rect 3249 16405 3283 16439
rect 6009 16405 6043 16439
rect 6929 16405 6963 16439
rect 9229 16405 9263 16439
rect 11437 16405 11471 16439
rect 16129 16405 16163 16439
rect 2053 16201 2087 16235
rect 3065 16201 3099 16235
rect 5917 16201 5951 16235
rect 8309 16201 8343 16235
rect 4353 16133 4387 16167
rect 9597 16133 9631 16167
rect 1869 16065 1903 16099
rect 4997 16065 5031 16099
rect 5089 16065 5123 16099
rect 5181 16065 5215 16099
rect 5365 16065 5399 16099
rect 5825 16065 5859 16099
rect 6009 16065 6043 16099
rect 7021 16065 7055 16099
rect 7113 16065 7147 16099
rect 7389 16065 7423 16099
rect 12173 16065 12207 16099
rect 1685 15997 1719 16031
rect 7297 15997 7331 16031
rect 4813 15861 4847 15895
rect 6837 15861 6871 15895
rect 10241 15861 10275 15895
rect 11069 15861 11103 15895
rect 12081 15861 12115 15895
rect 14197 15861 14231 15895
rect 1593 15657 1627 15691
rect 2513 15657 2547 15691
rect 8401 15657 8435 15691
rect 12817 15657 12851 15691
rect 16589 15657 16623 15691
rect 3157 15521 3191 15555
rect 7205 15521 7239 15555
rect 7849 15521 7883 15555
rect 11161 15521 11195 15555
rect 12081 15521 12115 15555
rect 12173 15521 12207 15555
rect 14657 15521 14691 15555
rect 16129 15521 16163 15555
rect 17233 15521 17267 15555
rect 1777 15453 1811 15487
rect 2053 15453 2087 15487
rect 5365 15453 5399 15487
rect 5825 15453 5859 15487
rect 6009 15453 6043 15487
rect 6745 15453 6779 15487
rect 7021 15453 7055 15487
rect 9137 15453 9171 15487
rect 9321 15453 9355 15487
rect 11989 15453 12023 15487
rect 13001 15453 13035 15487
rect 13093 15453 13127 15487
rect 13277 15453 13311 15487
rect 13369 15453 13403 15487
rect 14473 15453 14507 15487
rect 14565 15453 14599 15487
rect 14749 15453 14783 15487
rect 2973 15385 3007 15419
rect 5098 15385 5132 15419
rect 7941 15385 7975 15419
rect 9229 15385 9263 15419
rect 10916 15385 10950 15419
rect 18061 15385 18095 15419
rect 1961 15317 1995 15351
rect 2881 15317 2915 15351
rect 3985 15317 4019 15351
rect 5917 15317 5951 15351
rect 8033 15317 8067 15351
rect 9781 15317 9815 15351
rect 11621 15317 11655 15351
rect 14289 15317 14323 15351
rect 16957 15317 16991 15351
rect 17049 15317 17083 15351
rect 19441 15317 19475 15351
rect 2053 15113 2087 15147
rect 3893 15113 3927 15147
rect 4353 15113 4387 15147
rect 7941 15113 7975 15147
rect 10977 15113 11011 15147
rect 12725 15113 12759 15147
rect 14565 15113 14599 15147
rect 15301 15113 15335 15147
rect 19441 15113 19475 15147
rect 2513 15045 2547 15079
rect 5365 15045 5399 15079
rect 6653 15045 6687 15079
rect 8309 15045 8343 15079
rect 10793 15045 10827 15079
rect 13737 15045 13771 15079
rect 15485 15045 15519 15079
rect 17049 15045 17083 15079
rect 17601 15045 17635 15079
rect 2743 15011 2777 15045
rect 1777 14977 1811 15011
rect 3341 14977 3375 15011
rect 3525 14977 3559 15011
rect 3617 14977 3651 15011
rect 3709 14977 3743 15011
rect 4537 14977 4571 15011
rect 4629 14977 4663 15011
rect 4767 14977 4801 15011
rect 4905 14977 4939 15011
rect 5549 14977 5583 15011
rect 5641 14977 5675 15011
rect 8125 14977 8159 15011
rect 8217 14977 8251 15011
rect 8493 14977 8527 15011
rect 9505 14977 9539 15011
rect 11713 14977 11747 15011
rect 12633 14977 12667 15011
rect 12817 14977 12851 15011
rect 13640 14967 13674 15001
rect 13829 14977 13863 15011
rect 14013 14977 14047 15011
rect 14473 14977 14507 15011
rect 14657 14977 14691 15011
rect 16865 14977 16899 15011
rect 17141 14977 17175 15011
rect 18521 14977 18555 15011
rect 18705 14977 18739 15011
rect 18797 14977 18831 15011
rect 19349 14977 19383 15011
rect 2053 14909 2087 14943
rect 11069 14909 11103 14943
rect 15853 14841 15887 14875
rect 16865 14841 16899 14875
rect 1869 14773 1903 14807
rect 2697 14773 2731 14807
rect 2881 14773 2915 14807
rect 5365 14773 5399 14807
rect 5825 14773 5859 14807
rect 6929 14773 6963 14807
rect 9045 14773 9079 14807
rect 9229 14773 9263 14807
rect 10517 14773 10551 14807
rect 11805 14773 11839 14807
rect 12173 14773 12207 14807
rect 14013 14773 14047 14807
rect 15485 14773 15519 14807
rect 18337 14773 18371 14807
rect 2145 14569 2179 14603
rect 2605 14569 2639 14603
rect 2789 14569 2823 14603
rect 4077 14569 4111 14603
rect 7113 14569 7147 14603
rect 7297 14569 7331 14603
rect 10793 14569 10827 14603
rect 11253 14569 11287 14603
rect 11713 14569 11747 14603
rect 12357 14569 12391 14603
rect 14289 14569 14323 14603
rect 15485 14569 15519 14603
rect 16589 14569 16623 14603
rect 18153 14569 18187 14603
rect 9137 14501 9171 14535
rect 10701 14501 10735 14535
rect 12541 14501 12575 14535
rect 15761 14501 15795 14535
rect 20453 14501 20487 14535
rect 5733 14433 5767 14467
rect 11437 14433 11471 14467
rect 13645 14433 13679 14467
rect 14657 14433 14691 14467
rect 15853 14433 15887 14467
rect 18797 14433 18831 14467
rect 4077 14365 4111 14399
rect 4353 14365 4387 14399
rect 5089 14365 5123 14399
rect 5457 14365 5491 14399
rect 5917 14365 5951 14399
rect 6469 14365 6503 14399
rect 8033 14365 8067 14399
rect 8125 14365 8159 14399
rect 8309 14365 8343 14399
rect 8401 14365 8435 14399
rect 9413 14365 9447 14399
rect 9873 14365 9907 14399
rect 10793 14365 10827 14399
rect 11253 14365 11287 14399
rect 11529 14365 11563 14399
rect 13553 14365 13587 14399
rect 13737 14365 13771 14399
rect 14381 14365 14415 14399
rect 14473 14365 14507 14399
rect 14749 14365 14783 14399
rect 15669 14365 15703 14399
rect 15945 14365 15979 14399
rect 16129 14365 16163 14399
rect 16865 14365 16899 14399
rect 16957 14365 16991 14399
rect 17049 14365 17083 14399
rect 17233 14365 17267 14399
rect 19625 14365 19659 14399
rect 20637 14365 20671 14399
rect 2973 14297 3007 14331
rect 6929 14297 6963 14331
rect 7129 14297 7163 14331
rect 9137 14297 9171 14331
rect 10517 14297 10551 14331
rect 12173 14297 12207 14331
rect 12357 14297 12391 14331
rect 2773 14229 2807 14263
rect 4261 14229 4295 14263
rect 7849 14229 7883 14263
rect 9321 14229 9355 14263
rect 9965 14229 9999 14263
rect 18521 14229 18555 14263
rect 18613 14229 18647 14263
rect 19533 14229 19567 14263
rect 2519 14025 2553 14059
rect 4905 14025 4939 14059
rect 7205 14025 7239 14059
rect 8309 14025 8343 14059
rect 9045 14025 9079 14059
rect 10977 14025 11011 14059
rect 12265 14025 12299 14059
rect 15209 14025 15243 14059
rect 16865 14025 16899 14059
rect 17233 14025 17267 14059
rect 19165 14025 19199 14059
rect 20269 14025 20303 14059
rect 2421 13957 2455 13991
rect 5181 13957 5215 13991
rect 5273 13957 5307 13991
rect 6837 13957 6871 13991
rect 7849 13957 7883 13991
rect 14749 13957 14783 13991
rect 17877 13957 17911 13991
rect 19533 13957 19567 13991
rect 1869 13889 1903 13923
rect 2605 13889 2639 13923
rect 2697 13889 2731 13923
rect 3157 13889 3191 13923
rect 3341 13889 3375 13923
rect 4169 13889 4203 13923
rect 4353 13889 4387 13923
rect 5089 13889 5123 13923
rect 5457 13889 5491 13923
rect 6653 13889 6687 13923
rect 6929 13889 6963 13923
rect 7021 13889 7055 13923
rect 9229 13889 9263 13923
rect 9873 13889 9907 13923
rect 11713 13889 11747 13923
rect 11989 13889 12023 13923
rect 14197 13889 14231 13923
rect 14473 13889 14507 13923
rect 14565 13889 14599 13923
rect 15485 13889 15519 13923
rect 17049 13889 17083 13923
rect 17325 13889 17359 13923
rect 18061 13889 18095 13923
rect 18153 13889 18187 13923
rect 18429 13889 18463 13923
rect 19349 13889 19383 13923
rect 19441 13889 19475 13923
rect 19717 13889 19751 13923
rect 20177 13889 20211 13923
rect 20361 13889 20395 13923
rect 10885 13821 10919 13855
rect 11069 13821 11103 13855
rect 12173 13821 12207 13855
rect 14289 13821 14323 13855
rect 15393 13821 15427 13855
rect 15577 13821 15611 13855
rect 15669 13821 15703 13855
rect 18337 13821 18371 13855
rect 4353 13753 4387 13787
rect 8125 13753 8159 13787
rect 3157 13685 3191 13719
rect 6009 13685 6043 13719
rect 10517 13685 10551 13719
rect 12909 13685 12943 13719
rect 16313 13685 16347 13719
rect 1961 13481 1995 13515
rect 4813 13481 4847 13515
rect 8033 13481 8067 13515
rect 10517 13481 10551 13515
rect 11437 13481 11471 13515
rect 11805 13481 11839 13515
rect 12449 13481 12483 13515
rect 15853 13481 15887 13515
rect 19441 13481 19475 13515
rect 20913 13481 20947 13515
rect 4353 13413 4387 13447
rect 13093 13413 13127 13447
rect 14841 13413 14875 13447
rect 17601 13413 17635 13447
rect 2697 13345 2731 13379
rect 6377 13345 6411 13379
rect 6469 13345 6503 13379
rect 11345 13345 11379 13379
rect 1869 13277 1903 13311
rect 2053 13277 2087 13311
rect 2513 13277 2547 13311
rect 2881 13277 2915 13311
rect 4997 13277 5031 13311
rect 5089 13277 5123 13311
rect 5457 13277 5491 13311
rect 6561 13277 6595 13311
rect 6653 13277 6687 13311
rect 7481 13277 7515 13311
rect 7941 13277 7975 13311
rect 8125 13277 8159 13311
rect 9321 13277 9355 13311
rect 10057 13277 10091 13311
rect 11621 13277 11655 13311
rect 12449 13277 12483 13311
rect 13001 13277 13035 13311
rect 16037 13277 16071 13311
rect 16313 13277 16347 13311
rect 16773 13277 16807 13311
rect 16957 13277 16991 13311
rect 17739 13277 17773 13311
rect 18152 13277 18186 13311
rect 18245 13277 18279 13311
rect 18705 13277 18739 13311
rect 18889 13277 18923 13311
rect 19579 13277 19613 13311
rect 19717 13277 19751 13311
rect 19992 13277 20026 13311
rect 20085 13277 20119 13311
rect 21649 13277 21683 13311
rect 3433 13209 3467 13243
rect 17877 13209 17911 13243
rect 17969 13209 18003 13243
rect 19809 13209 19843 13243
rect 20545 13209 20579 13243
rect 20729 13209 20763 13243
rect 2605 13141 2639 13175
rect 2789 13141 2823 13175
rect 5273 13141 5307 13175
rect 5365 13141 5399 13175
rect 6837 13141 6871 13175
rect 7389 13141 7423 13175
rect 9229 13141 9263 13175
rect 16221 13141 16255 13175
rect 16957 13141 16991 13175
rect 18797 13141 18831 13175
rect 21465 13141 21499 13175
rect 2329 12937 2363 12971
rect 3525 12937 3559 12971
rect 4537 12937 4571 12971
rect 5549 12937 5583 12971
rect 7849 12937 7883 12971
rect 15945 12937 15979 12971
rect 18245 12937 18279 12971
rect 19165 12937 19199 12971
rect 3893 12869 3927 12903
rect 8769 12869 8803 12903
rect 14381 12869 14415 12903
rect 16313 12869 16347 12903
rect 17141 12869 17175 12903
rect 17351 12869 17385 12903
rect 1593 12801 1627 12835
rect 2605 12801 2639 12835
rect 2697 12801 2731 12835
rect 2789 12801 2823 12835
rect 3709 12801 3743 12835
rect 3801 12801 3835 12835
rect 4077 12801 4111 12835
rect 5089 12801 5123 12835
rect 6837 12801 6871 12835
rect 6929 12801 6963 12835
rect 9597 12801 9631 12835
rect 10241 12801 10275 12835
rect 12541 12801 12575 12835
rect 12909 12801 12943 12835
rect 15117 12801 15151 12835
rect 15301 12801 15335 12835
rect 15853 12801 15887 12835
rect 16129 12801 16163 12835
rect 17049 12801 17083 12835
rect 17233 12801 17267 12835
rect 18429 12801 18463 12835
rect 18613 12801 18647 12835
rect 18705 12801 18739 12835
rect 19349 12801 19383 12835
rect 19533 12801 19567 12835
rect 20545 12801 20579 12835
rect 20637 12801 20671 12835
rect 20821 12801 20855 12835
rect 20913 12801 20947 12835
rect 2513 12733 2547 12767
rect 6653 12733 6687 12767
rect 6745 12733 6779 12767
rect 9229 12733 9263 12767
rect 9505 12733 9539 12767
rect 15025 12733 15059 12767
rect 15209 12733 15243 12767
rect 16865 12733 16899 12767
rect 17509 12733 17543 12767
rect 21373 12733 21407 12767
rect 10701 12665 10735 12699
rect 1777 12597 1811 12631
rect 5365 12597 5399 12631
rect 7113 12597 7147 12631
rect 10333 12597 10367 12631
rect 14841 12597 14875 12631
rect 20361 12597 20395 12631
rect 22109 12597 22143 12631
rect 2881 12393 2915 12427
rect 5733 12393 5767 12427
rect 6193 12393 6227 12427
rect 9137 12393 9171 12427
rect 11345 12393 11379 12427
rect 16313 12393 16347 12427
rect 18245 12393 18279 12427
rect 20177 12393 20211 12427
rect 4537 12325 4571 12359
rect 7297 12325 7331 12359
rect 13553 12325 13587 12359
rect 17693 12325 17727 12359
rect 4261 12257 4295 12291
rect 5365 12257 5399 12291
rect 7941 12257 7975 12291
rect 8493 12257 8527 12291
rect 11897 12257 11931 12291
rect 14473 12257 14507 12291
rect 14933 12257 14967 12291
rect 2237 12189 2271 12223
rect 4169 12189 4203 12223
rect 5273 12189 5307 12223
rect 5457 12189 5491 12223
rect 5549 12189 5583 12223
rect 6394 12199 6428 12233
rect 6837 12189 6871 12223
rect 7481 12189 7515 12223
rect 9321 12189 9355 12223
rect 9781 12189 9815 12223
rect 11805 12189 11839 12223
rect 11989 12189 12023 12223
rect 12633 12189 12667 12223
rect 12725 12189 12759 12223
rect 12909 12189 12943 12223
rect 13001 12189 13035 12223
rect 14565 12189 14599 12223
rect 15669 12189 15703 12223
rect 15853 12189 15887 12223
rect 16497 12189 16531 12223
rect 16773 12189 16807 12223
rect 17417 12189 17451 12223
rect 17509 12189 17543 12223
rect 17785 12167 17819 12201
rect 18429 12189 18463 12223
rect 18613 12189 18647 12223
rect 18889 12189 18923 12223
rect 19901 12189 19935 12223
rect 19993 12189 20027 12223
rect 21741 12189 21775 12223
rect 2789 12121 2823 12155
rect 6469 12121 6503 12155
rect 6561 12121 6595 12155
rect 6699 12121 6733 12155
rect 7573 12121 7607 12155
rect 7665 12121 7699 12155
rect 7803 12121 7837 12155
rect 9413 12121 9447 12155
rect 9505 12121 9539 12155
rect 9643 12121 9677 12155
rect 14841 12121 14875 12155
rect 15761 12121 15795 12155
rect 18521 12121 18555 12155
rect 18751 12121 18785 12155
rect 21189 12121 21223 12155
rect 2053 12053 2087 12087
rect 10333 12053 10367 12087
rect 12449 12053 12483 12087
rect 14289 12053 14323 12087
rect 16681 12053 16715 12087
rect 17417 12053 17451 12087
rect 21097 12053 21131 12087
rect 21833 12053 21867 12087
rect 22477 12053 22511 12087
rect 2973 11849 3007 11883
rect 4169 11849 4203 11883
rect 4721 11849 4755 11883
rect 5549 11849 5583 11883
rect 6009 11849 6043 11883
rect 7941 11849 7975 11883
rect 11713 11849 11747 11883
rect 13645 11849 13679 11883
rect 15485 11849 15519 11883
rect 16129 11849 16163 11883
rect 16865 11849 16899 11883
rect 17969 11849 18003 11883
rect 18429 11849 18463 11883
rect 2145 11781 2179 11815
rect 8217 11781 8251 11815
rect 11161 11781 11195 11815
rect 12081 11781 12115 11815
rect 19533 11781 19567 11815
rect 2053 11713 2087 11747
rect 2237 11713 2271 11747
rect 2697 11713 2731 11747
rect 3433 11713 3467 11747
rect 3525 11713 3559 11747
rect 3617 11713 3651 11747
rect 4629 11713 4663 11747
rect 4813 11713 4847 11747
rect 5641 11713 5675 11747
rect 6561 11713 6595 11747
rect 6745 11713 6779 11747
rect 6837 11713 6871 11747
rect 6929 11713 6963 11747
rect 8125 11713 8159 11747
rect 8309 11713 8343 11747
rect 8493 11713 8527 11747
rect 9505 11713 9539 11747
rect 9597 11713 9631 11747
rect 10149 11713 10183 11747
rect 11897 11713 11931 11747
rect 11989 11713 12023 11747
rect 12265 11713 12299 11747
rect 12725 11713 12759 11747
rect 12909 11713 12943 11747
rect 14013 11713 14047 11747
rect 14657 11713 14691 11747
rect 15393 11713 15427 11747
rect 15761 11713 15795 11747
rect 15853 11713 15887 11747
rect 17049 11713 17083 11747
rect 17233 11713 17267 11747
rect 18797 11713 18831 11747
rect 20269 11713 20303 11747
rect 20545 11713 20579 11747
rect 20729 11713 20763 11747
rect 21189 11713 21223 11747
rect 22017 11713 22051 11747
rect 22109 11713 22143 11747
rect 22293 11713 22327 11747
rect 2973 11645 3007 11679
rect 5457 11645 5491 11679
rect 7205 11645 7239 11679
rect 10425 11645 10459 11679
rect 13185 11645 13219 11679
rect 13921 11645 13955 11679
rect 14841 11645 14875 11679
rect 15669 11645 15703 11679
rect 17141 11645 17175 11679
rect 17325 11645 17359 11679
rect 18613 11645 18647 11679
rect 18705 11645 18739 11679
rect 18889 11645 18923 11679
rect 20085 11645 20119 11679
rect 2789 11577 2823 11611
rect 10241 11577 10275 11611
rect 14473 11577 14507 11611
rect 20361 11577 20395 11611
rect 20453 11577 20487 11611
rect 9321 11509 9355 11543
rect 10333 11509 10367 11543
rect 13093 11509 13127 11543
rect 14013 11509 14047 11543
rect 21373 11509 21407 11543
rect 22477 11509 22511 11543
rect 23029 11509 23063 11543
rect 2237 11305 2271 11339
rect 5181 11305 5215 11339
rect 5365 11305 5399 11339
rect 6285 11305 6319 11339
rect 6929 11305 6963 11339
rect 8401 11305 8435 11339
rect 8585 11305 8619 11339
rect 10333 11305 10367 11339
rect 14289 11305 14323 11339
rect 16497 11305 16531 11339
rect 17233 11305 17267 11339
rect 19809 11305 19843 11339
rect 20361 11305 20395 11339
rect 21465 11305 21499 11339
rect 21741 11305 21775 11339
rect 1685 11237 1719 11271
rect 15485 11237 15519 11271
rect 18429 11237 18463 11271
rect 18521 11237 18555 11271
rect 2605 11169 2639 11203
rect 8309 11169 8343 11203
rect 14565 11169 14599 11203
rect 18613 11169 18647 11203
rect 2145 11101 2179 11135
rect 3433 11101 3467 11135
rect 3985 11101 4019 11135
rect 4169 11101 4203 11135
rect 5917 11101 5951 11135
rect 6009 11101 6043 11135
rect 6101 11101 6135 11135
rect 7113 11101 7147 11135
rect 7205 11101 7239 11135
rect 7573 11101 7607 11135
rect 8217 11101 8251 11135
rect 9321 11101 9355 11135
rect 9413 11101 9447 11135
rect 9597 11101 9631 11135
rect 9689 11101 9723 11135
rect 10149 11101 10183 11135
rect 10333 11101 10367 11135
rect 11529 11101 11563 11135
rect 11989 11101 12023 11135
rect 13185 11101 13219 11135
rect 13461 11101 13495 11135
rect 14473 11101 14507 11135
rect 14657 11101 14691 11135
rect 14749 11101 14783 11135
rect 14933 11101 14967 11135
rect 15393 11101 15427 11135
rect 15577 11101 15611 11135
rect 16037 11101 16071 11135
rect 16313 11101 16347 11135
rect 16957 11101 16991 11135
rect 17049 11101 17083 11135
rect 18705 11101 18739 11135
rect 18889 11101 18923 11135
rect 19441 11101 19475 11135
rect 19625 11101 19659 11135
rect 19901 11101 19935 11135
rect 20637 11101 20671 11135
rect 20726 11098 20760 11132
rect 20821 11095 20855 11129
rect 21005 11101 21039 11135
rect 21741 11101 21775 11135
rect 21833 11101 21867 11135
rect 22293 11101 22327 11135
rect 3249 11033 3283 11067
rect 4997 11033 5031 11067
rect 5197 11033 5231 11067
rect 7297 11033 7331 11067
rect 7435 11033 7469 11067
rect 13277 11033 13311 11067
rect 16129 11033 16163 11067
rect 17233 11033 17267 11067
rect 22385 11033 22419 11067
rect 3065 10965 3099 10999
rect 4077 10965 4111 10999
rect 9137 10965 9171 10999
rect 13185 10965 13219 10999
rect 18153 10965 18187 10999
rect 4261 10761 4295 10795
rect 6561 10761 6595 10795
rect 8493 10761 8527 10795
rect 9597 10761 9631 10795
rect 12265 10761 12299 10795
rect 13093 10761 13127 10795
rect 16221 10761 16255 10795
rect 17693 10761 17727 10795
rect 18889 10761 18923 10795
rect 20361 10761 20395 10795
rect 20545 10761 20579 10795
rect 22017 10761 22051 10795
rect 6929 10693 6963 10727
rect 10885 10693 10919 10727
rect 12725 10693 12759 10727
rect 15301 10693 15335 10727
rect 15669 10693 15703 10727
rect 20729 10693 20763 10727
rect 1685 10625 1719 10659
rect 2605 10625 2639 10659
rect 2698 10625 2732 10659
rect 2881 10625 2915 10659
rect 2973 10625 3007 10659
rect 3070 10625 3104 10659
rect 3801 10625 3835 10659
rect 4077 10625 4111 10659
rect 4721 10625 4755 10659
rect 5457 10625 5491 10659
rect 5641 10625 5675 10659
rect 6745 10625 6779 10659
rect 7855 10625 7889 10659
rect 8033 10625 8067 10659
rect 8769 10625 8803 10659
rect 8861 10625 8895 10659
rect 8953 10625 8987 10659
rect 9137 10625 9171 10659
rect 9965 10625 9999 10659
rect 11161 10625 11195 10659
rect 11897 10625 11931 10659
rect 12081 10625 12115 10659
rect 13001 10625 13035 10659
rect 13185 10625 13219 10659
rect 14657 10625 14691 10659
rect 15485 10625 15519 10659
rect 16129 10625 16163 10659
rect 16313 10625 16347 10659
rect 17601 10625 17635 10659
rect 18337 10625 18371 10659
rect 18429 10625 18463 10659
rect 18613 10625 18647 10659
rect 18705 10625 18739 10659
rect 19625 10625 19659 10659
rect 19809 10625 19843 10659
rect 20637 10625 20671 10659
rect 2145 10557 2179 10591
rect 3893 10557 3927 10591
rect 9781 10557 9815 10591
rect 9873 10557 9907 10591
rect 10057 10557 10091 10591
rect 11805 10557 11839 10591
rect 11989 10557 12023 10591
rect 13461 10557 13495 10591
rect 19533 10557 19567 10591
rect 19717 10557 19751 10591
rect 3249 10489 3283 10523
rect 8033 10489 8067 10523
rect 11069 10489 11103 10523
rect 11161 10489 11195 10523
rect 16865 10489 16899 10523
rect 20913 10489 20947 10523
rect 1961 10421 1995 10455
rect 4077 10421 4111 10455
rect 4905 10421 4939 10455
rect 5641 10421 5675 10455
rect 13369 10421 13403 10455
rect 14013 10421 14047 10455
rect 14565 10421 14599 10455
rect 19349 10421 19383 10455
rect 21465 10421 21499 10455
rect 2237 10217 2271 10251
rect 2421 10217 2455 10251
rect 3985 10217 4019 10251
rect 5089 10217 5123 10251
rect 5917 10217 5951 10251
rect 6193 10217 6227 10251
rect 8401 10217 8435 10251
rect 9137 10217 9171 10251
rect 10885 10217 10919 10251
rect 11989 10217 12023 10251
rect 12449 10217 12483 10251
rect 13645 10217 13679 10251
rect 14657 10217 14691 10251
rect 17693 10217 17727 10251
rect 18797 10217 18831 10251
rect 19625 10217 19659 10251
rect 20720 10217 20754 10251
rect 20913 10217 20947 10251
rect 1777 10149 1811 10183
rect 3433 10149 3467 10183
rect 7021 10149 7055 10183
rect 10333 10149 10367 10183
rect 16037 10149 16071 10183
rect 2513 10081 2547 10115
rect 5181 10081 5215 10115
rect 5365 10081 5399 10115
rect 9597 10081 9631 10115
rect 11621 10081 11655 10115
rect 11713 10081 11747 10115
rect 12633 10081 12667 10115
rect 12725 10081 12759 10115
rect 12909 10081 12943 10115
rect 21373 10081 21407 10115
rect 2789 10013 2823 10047
rect 4169 10013 4203 10047
rect 4445 10013 4479 10047
rect 5089 10013 5123 10047
rect 5825 10013 5859 10047
rect 6009 10013 6043 10047
rect 6745 10013 6779 10047
rect 7757 10013 7791 10047
rect 7850 10013 7884 10047
rect 8033 10013 8067 10047
rect 8222 10013 8256 10047
rect 9321 10013 9355 10047
rect 9413 10013 9447 10047
rect 9505 10013 9539 10047
rect 10793 10013 10827 10047
rect 10977 10013 11011 10047
rect 11529 10013 11563 10047
rect 11805 10013 11839 10047
rect 12818 10013 12852 10047
rect 13461 10013 13495 10047
rect 14289 10013 14323 10047
rect 15393 10013 15427 10047
rect 15541 10013 15575 10047
rect 15761 10013 15795 10047
rect 15899 10013 15933 10047
rect 18337 10013 18371 10047
rect 18613 10013 18647 10047
rect 19441 10013 19475 10047
rect 19625 10013 19659 10047
rect 22477 10013 22511 10047
rect 4353 9945 4387 9979
rect 7021 9945 7055 9979
rect 8125 9945 8159 9979
rect 14473 9945 14507 9979
rect 15669 9945 15703 9979
rect 16497 9945 16531 9979
rect 17141 9945 17175 9979
rect 17417 9945 17451 9979
rect 17509 9945 17543 9979
rect 20545 9945 20579 9979
rect 6837 9877 6871 9911
rect 17325 9877 17359 9911
rect 18429 9877 18463 9911
rect 20745 9877 20779 9911
rect 21925 9877 21959 9911
rect 23121 9877 23155 9911
rect 1961 9673 1995 9707
rect 4537 9673 4571 9707
rect 6009 9673 6043 9707
rect 11161 9673 11195 9707
rect 17509 9673 17543 9707
rect 3341 9605 3375 9639
rect 12541 9605 12575 9639
rect 17785 9605 17819 9639
rect 19625 9605 19659 9639
rect 20453 9605 20487 9639
rect 2513 9537 2547 9571
rect 2605 9537 2639 9571
rect 4353 9537 4387 9571
rect 5365 9537 5399 9571
rect 5825 9537 5859 9571
rect 6745 9537 6779 9571
rect 7021 9537 7055 9571
rect 7113 9537 7147 9571
rect 7297 9537 7331 9571
rect 10149 9537 10183 9571
rect 10333 9537 10367 9571
rect 11805 9537 11839 9571
rect 12771 9537 12805 9571
rect 12890 9537 12924 9571
rect 13001 9537 13035 9571
rect 13185 9537 13219 9571
rect 13737 9537 13771 9571
rect 13921 9537 13955 9571
rect 14657 9537 14691 9571
rect 14749 9537 14783 9571
rect 14841 9537 14875 9571
rect 15025 9537 15059 9571
rect 15669 9537 15703 9571
rect 16129 9537 16163 9571
rect 17693 9537 17727 9571
rect 17877 9537 17911 9571
rect 18061 9537 18095 9571
rect 18153 9537 18187 9571
rect 19533 9537 19567 9571
rect 19717 9537 19751 9571
rect 20177 9537 20211 9571
rect 20325 9537 20359 9571
rect 20545 9537 20579 9571
rect 20683 9537 20717 9571
rect 22017 9537 22051 9571
rect 22109 9537 22143 9571
rect 23029 9537 23063 9571
rect 5641 9469 5675 9503
rect 6929 9469 6963 9503
rect 8861 9469 8895 9503
rect 10517 9469 10551 9503
rect 12081 9469 12115 9503
rect 15853 9469 15887 9503
rect 15945 9469 15979 9503
rect 16865 9469 16899 9503
rect 22293 9469 22327 9503
rect 2789 9401 2823 9435
rect 8309 9401 8343 9435
rect 15761 9401 15795 9435
rect 20821 9401 20855 9435
rect 22845 9401 22879 9435
rect 3617 9333 3651 9367
rect 5457 9333 5491 9367
rect 6561 9333 6595 9367
rect 7849 9333 7883 9367
rect 9689 9333 9723 9367
rect 11897 9333 11931 9367
rect 11989 9333 12023 9367
rect 13921 9333 13955 9367
rect 14381 9333 14415 9367
rect 15485 9333 15519 9367
rect 18613 9333 18647 9367
rect 21281 9333 21315 9367
rect 22201 9333 22235 9367
rect 4445 9129 4479 9163
rect 5457 9129 5491 9163
rect 6377 9129 6411 9163
rect 7113 9129 7147 9163
rect 8401 9129 8435 9163
rect 11253 9129 11287 9163
rect 11713 9129 11747 9163
rect 14289 9129 14323 9163
rect 18705 9129 18739 9163
rect 6561 9061 6595 9095
rect 8585 9061 8619 9095
rect 12541 9061 12575 9095
rect 13185 9061 13219 9095
rect 19993 9061 20027 9095
rect 2973 8993 3007 9027
rect 8217 8993 8251 9027
rect 14473 8993 14507 9027
rect 14749 8993 14783 9027
rect 15853 8993 15887 9027
rect 16405 8993 16439 9027
rect 16681 8993 16715 9027
rect 16865 8993 16899 9027
rect 17417 8993 17451 9027
rect 20637 8993 20671 9027
rect 20821 8993 20855 9027
rect 2697 8925 2731 8959
rect 2881 8925 2915 8959
rect 3065 8925 3099 8959
rect 3249 8925 3283 8959
rect 4445 8925 4479 8959
rect 4537 8925 4571 8959
rect 5273 8925 5307 8959
rect 5457 8925 5491 8959
rect 7941 8925 7975 8959
rect 8401 8925 8435 8959
rect 9137 8925 9171 8959
rect 9321 8925 9355 8959
rect 9413 8925 9447 8959
rect 9505 8925 9539 8959
rect 10241 8925 10275 8959
rect 11437 8925 11471 8959
rect 11529 8925 11563 8959
rect 11805 8925 11839 8959
rect 12265 8925 12299 8959
rect 12725 8925 12759 8959
rect 13369 8925 13403 8959
rect 13534 8925 13568 8959
rect 13645 8925 13679 8959
rect 13737 8925 13771 8959
rect 14566 8925 14600 8959
rect 14657 8925 14691 8959
rect 15669 8925 15703 8959
rect 15945 8925 15979 8959
rect 16589 8925 16623 8959
rect 16773 8925 16807 8959
rect 17693 8925 17727 8959
rect 17785 8925 17819 8959
rect 17877 8925 17911 8959
rect 18061 8925 18095 8959
rect 19717 8925 19751 8959
rect 19993 8925 20027 8959
rect 20729 8925 20763 8959
rect 20913 8925 20947 8959
rect 21557 8925 21591 8959
rect 22385 8925 22419 8959
rect 22477 8925 22511 8959
rect 22661 8925 22695 8959
rect 6423 8891 6457 8925
rect 6193 8857 6227 8891
rect 7205 8857 7239 8891
rect 10425 8857 10459 8891
rect 15485 8857 15519 8891
rect 18889 8857 18923 8891
rect 1685 8789 1719 8823
rect 2237 8789 2271 8823
rect 3433 8789 3467 8823
rect 4813 8789 4847 8823
rect 5641 8789 5675 8823
rect 9781 8789 9815 8823
rect 10609 8789 10643 8823
rect 12357 8789 12391 8823
rect 18521 8789 18555 8823
rect 18689 8789 18723 8823
rect 19809 8789 19843 8823
rect 20453 8789 20487 8823
rect 21649 8789 21683 8823
rect 22845 8789 22879 8823
rect 2053 8585 2087 8619
rect 4261 8585 4295 8619
rect 5181 8585 5215 8619
rect 7389 8585 7423 8619
rect 9505 8585 9539 8619
rect 12909 8585 12943 8619
rect 13369 8585 13403 8619
rect 14841 8585 14875 8619
rect 16145 8585 16179 8619
rect 16313 8585 16347 8619
rect 16957 8585 16991 8619
rect 18521 8585 18555 8619
rect 20545 8585 20579 8619
rect 22109 8585 22143 8619
rect 22477 8585 22511 8619
rect 23121 8585 23155 8619
rect 7757 8517 7791 8551
rect 9597 8517 9631 8551
rect 11805 8517 11839 8551
rect 12541 8517 12575 8551
rect 15945 8517 15979 8551
rect 1869 8449 1903 8483
rect 2697 8449 2731 8483
rect 3709 8449 3743 8483
rect 3801 8449 3835 8483
rect 3985 8449 4019 8483
rect 4077 8449 4111 8483
rect 5089 8449 5123 8483
rect 5365 8449 5399 8483
rect 6653 8449 6687 8483
rect 7573 8449 7607 8483
rect 7665 8449 7699 8483
rect 7875 8449 7909 8483
rect 8033 8449 8067 8483
rect 8485 8449 8519 8483
rect 9413 8449 9447 8483
rect 9781 8449 9815 8483
rect 10333 8449 10367 8483
rect 10517 8449 10551 8483
rect 12265 8449 12299 8483
rect 12358 8449 12392 8483
rect 12633 8449 12667 8483
rect 12771 8449 12805 8483
rect 13645 8449 13679 8483
rect 13737 8449 13771 8483
rect 14203 8449 14237 8483
rect 14381 8449 14415 8483
rect 15025 8449 15059 8483
rect 17141 8449 17175 8483
rect 17233 8449 17267 8483
rect 17417 8449 17451 8483
rect 17509 8449 17543 8483
rect 17969 8449 18003 8483
rect 18061 8449 18095 8483
rect 18245 8449 18279 8483
rect 18337 8449 18371 8483
rect 19717 8449 19751 8483
rect 19809 8449 19843 8483
rect 19901 8449 19935 8483
rect 20085 8449 20119 8483
rect 20729 8449 20763 8483
rect 20821 8449 20855 8483
rect 21005 8449 21039 8483
rect 21097 8449 21131 8483
rect 22017 8449 22051 8483
rect 22293 8449 22327 8483
rect 22937 8449 22971 8483
rect 1593 8381 1627 8415
rect 2513 8381 2547 8415
rect 2881 8381 2915 8415
rect 8585 8381 8619 8415
rect 9873 8381 9907 8415
rect 15117 8381 15151 8415
rect 15209 8381 15243 8415
rect 15301 8381 15335 8415
rect 5549 8313 5583 8347
rect 14289 8313 14323 8347
rect 1685 8245 1719 8279
rect 6745 8245 6779 8279
rect 9137 8245 9171 8279
rect 10333 8245 10367 8279
rect 10701 8245 10735 8279
rect 13553 8245 13587 8279
rect 16129 8245 16163 8279
rect 19441 8245 19475 8279
rect 1777 8041 1811 8075
rect 2697 8041 2731 8075
rect 3341 8041 3375 8075
rect 4261 8041 4295 8075
rect 5089 8041 5123 8075
rect 7297 8041 7331 8075
rect 7757 8041 7791 8075
rect 9689 8041 9723 8075
rect 10885 8041 10919 8075
rect 12909 8041 12943 8075
rect 14657 8041 14691 8075
rect 15761 8041 15795 8075
rect 16957 8041 16991 8075
rect 17785 8041 17819 8075
rect 19441 8041 19475 8075
rect 19809 8041 19843 8075
rect 20269 8041 20303 8075
rect 4721 7973 4755 8007
rect 5273 7973 5307 8007
rect 10241 7973 10275 8007
rect 16221 7973 16255 8007
rect 16865 7973 16899 8007
rect 3433 7905 3467 7939
rect 6561 7905 6595 7939
rect 12081 7905 12115 7939
rect 16773 7905 16807 7939
rect 20729 7905 20763 7939
rect 21281 7905 21315 7939
rect 2311 7837 2345 7871
rect 2421 7837 2455 7871
rect 2513 7837 2547 7871
rect 3157 7837 3191 7871
rect 3249 7837 3283 7871
rect 6285 7837 6319 7871
rect 6469 7837 6503 7871
rect 7205 7837 7239 7871
rect 7481 7837 7515 7871
rect 7573 7837 7607 7871
rect 7757 7837 7791 7871
rect 8217 7837 8251 7871
rect 8401 7837 8435 7871
rect 9137 7837 9171 7871
rect 9321 7837 9355 7871
rect 9413 7837 9447 7871
rect 9505 7837 9539 7871
rect 10701 7837 10735 7871
rect 11621 7837 11655 7871
rect 11897 7837 11931 7871
rect 13093 7837 13127 7871
rect 13185 7837 13219 7871
rect 13369 7837 13403 7871
rect 13461 7837 13495 7871
rect 14841 7837 14875 7871
rect 14933 7837 14967 7871
rect 15301 7837 15335 7871
rect 15945 7837 15979 7871
rect 16097 7837 16131 7871
rect 16313 7837 16347 7871
rect 17049 7837 17083 7871
rect 17969 7837 18003 7871
rect 18061 7837 18095 7871
rect 18245 7837 18279 7871
rect 18337 7837 18371 7871
rect 19441 7837 19475 7871
rect 19625 7837 19659 7871
rect 20453 7837 20487 7871
rect 20545 7837 20579 7871
rect 20821 7837 20855 7871
rect 21465 7837 21499 7871
rect 21741 7837 21775 7871
rect 5089 7769 5123 7803
rect 11713 7769 11747 7803
rect 15025 7769 15059 7803
rect 15163 7769 15197 7803
rect 22753 7769 22787 7803
rect 6101 7701 6135 7735
rect 8309 7701 8343 7735
rect 18889 7701 18923 7735
rect 21649 7701 21683 7735
rect 22293 7701 22327 7735
rect 2973 7497 3007 7531
rect 4997 7497 5031 7531
rect 8861 7497 8895 7531
rect 12265 7497 12299 7531
rect 12909 7497 12943 7531
rect 13001 7497 13035 7531
rect 15301 7497 15335 7531
rect 17417 7497 17451 7531
rect 20177 7497 20211 7531
rect 22017 7497 22051 7531
rect 23029 7497 23063 7531
rect 2513 7429 2547 7463
rect 3617 7429 3651 7463
rect 4629 7429 4663 7463
rect 10885 7429 10919 7463
rect 11989 7429 12023 7463
rect 12725 7429 12759 7463
rect 14841 7429 14875 7463
rect 19809 7429 19843 7463
rect 21005 7429 21039 7463
rect 2053 7361 2087 7395
rect 2789 7361 2823 7395
rect 3433 7361 3467 7395
rect 4813 7361 4847 7395
rect 5733 7361 5767 7395
rect 5825 7361 5859 7395
rect 7297 7361 7331 7395
rect 7849 7361 7883 7395
rect 9045 7361 9079 7395
rect 9321 7361 9355 7395
rect 9965 7361 9999 7395
rect 10149 7361 10183 7395
rect 10241 7361 10275 7395
rect 11161 7361 11195 7395
rect 11713 7361 11747 7395
rect 11897 7361 11931 7395
rect 12081 7361 12115 7395
rect 13093 7361 13127 7395
rect 14197 7361 14231 7395
rect 14381 7361 14415 7395
rect 14473 7361 14507 7395
rect 14565 7361 14599 7395
rect 15761 7361 15795 7395
rect 16865 7361 16899 7395
rect 16957 7361 16991 7395
rect 17141 7361 17175 7395
rect 17233 7361 17267 7395
rect 17877 7361 17911 7395
rect 18061 7361 18095 7395
rect 18981 7361 19015 7395
rect 19717 7361 19751 7395
rect 19993 7361 20027 7395
rect 20637 7361 20671 7395
rect 20821 7361 20855 7395
rect 22201 7361 22235 7395
rect 22293 7361 22327 7395
rect 22477 7361 22511 7395
rect 22569 7361 22603 7395
rect 2697 7293 2731 7327
rect 6009 7293 6043 7327
rect 7009 7293 7043 7327
rect 7757 7293 7791 7327
rect 9137 7293 9171 7327
rect 15485 7293 15519 7327
rect 15577 7293 15611 7327
rect 15669 7293 15703 7327
rect 18337 7293 18371 7327
rect 13277 7225 13311 7259
rect 18889 7225 18923 7259
rect 1869 7157 1903 7191
rect 2513 7157 2547 7191
rect 3709 7157 3743 7191
rect 5917 7157 5951 7191
rect 9137 7157 9171 7191
rect 9781 7157 9815 7191
rect 18245 7157 18279 7191
rect 2237 6953 2271 6987
rect 6653 6953 6687 6987
rect 10609 6953 10643 6987
rect 11161 6953 11195 6987
rect 13185 6953 13219 6987
rect 14933 6953 14967 6987
rect 15393 6953 15427 6987
rect 15577 6953 15611 6987
rect 2421 6885 2455 6919
rect 16497 6885 16531 6919
rect 18613 6885 18647 6919
rect 22017 6885 22051 6919
rect 5088 6817 5122 6851
rect 5365 6817 5399 6851
rect 6377 6817 6411 6851
rect 7849 6817 7883 6851
rect 7941 6817 7975 6851
rect 8033 6817 8067 6851
rect 9597 6817 9631 6851
rect 10885 6817 10919 6851
rect 14381 6817 14415 6851
rect 17969 6817 18003 6851
rect 20361 6817 20395 6851
rect 20821 6817 20855 6851
rect 2973 6749 3007 6783
rect 3985 6749 4019 6783
rect 4169 6749 4203 6783
rect 4537 6749 4571 6783
rect 5181 6749 5215 6783
rect 5272 6749 5306 6783
rect 6469 6749 6503 6783
rect 7757 6749 7791 6783
rect 9321 6749 9355 6783
rect 9413 6749 9447 6783
rect 9505 6749 9539 6783
rect 10977 6749 11011 6783
rect 11713 6749 11747 6783
rect 12541 6749 12575 6783
rect 13093 6749 13127 6783
rect 13277 6749 13311 6783
rect 16221 6749 16255 6783
rect 16405 6749 16439 6783
rect 16589 6749 16623 6783
rect 16681 6749 16715 6783
rect 17325 6749 17359 6783
rect 17509 6749 17543 6783
rect 17601 6749 17635 6783
rect 17693 6749 17727 6783
rect 18429 6749 18463 6783
rect 18521 6749 18555 6783
rect 19717 6749 19751 6783
rect 19901 6749 19935 6783
rect 19993 6749 20027 6783
rect 20085 6749 20119 6783
rect 21097 6749 21131 6783
rect 21189 6749 21223 6783
rect 21281 6749 21315 6783
rect 21465 6749 21499 6783
rect 22201 6749 22235 6783
rect 2053 6681 2087 6715
rect 4445 6681 4479 6715
rect 6009 6681 6043 6715
rect 10517 6681 10551 6715
rect 12449 6681 12483 6715
rect 15761 6681 15795 6715
rect 18889 6681 18923 6715
rect 2237 6613 2271 6647
rect 3157 6613 3191 6647
rect 5549 6613 5583 6647
rect 7113 6613 7147 6647
rect 8217 6613 8251 6647
rect 9137 6613 9171 6647
rect 11713 6613 11747 6647
rect 15561 6613 15595 6647
rect 16865 6613 16899 6647
rect 18797 6613 18831 6647
rect 4261 6409 4295 6443
rect 4353 6409 4387 6443
rect 5181 6409 5215 6443
rect 5273 6409 5307 6443
rect 7205 6409 7239 6443
rect 7941 6409 7975 6443
rect 9045 6409 9079 6443
rect 9505 6409 9539 6443
rect 11161 6409 11195 6443
rect 16221 6409 16255 6443
rect 17049 6409 17083 6443
rect 19809 6409 19843 6443
rect 21281 6409 21315 6443
rect 3801 6341 3835 6375
rect 4997 6341 5031 6375
rect 6837 6341 6871 6375
rect 6929 6341 6963 6375
rect 12725 6341 12759 6375
rect 13921 6341 13955 6375
rect 19349 6341 19383 6375
rect 1685 6273 1719 6307
rect 1777 6273 1811 6307
rect 1961 6273 1995 6307
rect 2605 6273 2639 6307
rect 2881 6273 2915 6307
rect 3249 6273 3283 6307
rect 5365 6273 5399 6307
rect 6561 6273 6595 6307
rect 6654 6273 6688 6307
rect 7067 6273 7101 6307
rect 8401 6273 8435 6307
rect 8585 6273 8619 6307
rect 8677 6273 8711 6307
rect 8769 6273 8803 6307
rect 9689 6273 9723 6307
rect 10701 6273 10735 6307
rect 10885 6273 10919 6307
rect 11989 6273 12023 6307
rect 13185 6273 13219 6307
rect 14473 6273 14507 6307
rect 14657 6273 14691 6307
rect 15393 6273 15427 6307
rect 16129 6273 16163 6307
rect 16313 6273 16347 6307
rect 16865 6273 16899 6307
rect 17049 6273 17083 6307
rect 18153 6273 18187 6307
rect 18245 6273 18279 6307
rect 18981 6273 19015 6307
rect 19257 6273 19291 6307
rect 20085 6273 20119 6307
rect 20177 6273 20211 6307
rect 20269 6273 20303 6307
rect 20465 6273 20499 6307
rect 21097 6273 21131 6307
rect 1869 6205 1903 6239
rect 3065 6205 3099 6239
rect 9965 6205 9999 6239
rect 10793 6205 10827 6239
rect 10977 6205 11011 6239
rect 12357 6205 12391 6239
rect 13553 6205 13587 6239
rect 18061 6205 18095 6239
rect 18337 6205 18371 6239
rect 20913 6205 20947 6239
rect 3801 6137 3835 6171
rect 5549 6137 5583 6171
rect 9873 6137 9907 6171
rect 12127 6137 12161 6171
rect 12265 6137 12299 6171
rect 14841 6137 14875 6171
rect 2145 6069 2179 6103
rect 4537 6069 4571 6103
rect 13323 6069 13357 6103
rect 13461 6069 13495 6103
rect 14657 6069 14691 6103
rect 15577 6069 15611 6103
rect 18521 6069 18555 6103
rect 22109 6069 22143 6103
rect 4077 5865 4111 5899
rect 7849 5865 7883 5899
rect 9137 5865 9171 5899
rect 10241 5865 10275 5899
rect 12265 5865 12299 5899
rect 14289 5865 14323 5899
rect 14657 5865 14691 5899
rect 16681 5865 16715 5899
rect 18245 5865 18279 5899
rect 20453 5865 20487 5899
rect 20545 5865 20579 5899
rect 2329 5797 2363 5831
rect 10425 5797 10459 5831
rect 11161 5797 11195 5831
rect 13461 5797 13495 5831
rect 16037 5797 16071 5831
rect 18521 5797 18555 5831
rect 21189 5797 21223 5831
rect 14381 5729 14415 5763
rect 15761 5729 15795 5763
rect 18705 5729 18739 5763
rect 1961 5661 1995 5695
rect 2145 5661 2179 5695
rect 2237 5661 2271 5695
rect 2421 5661 2455 5695
rect 3065 5661 3099 5695
rect 3249 5661 3283 5695
rect 3985 5661 4019 5695
rect 4905 5661 4939 5695
rect 5089 5661 5123 5695
rect 5457 5661 5491 5695
rect 6101 5661 6135 5695
rect 6285 5661 6319 5695
rect 7297 5661 7331 5695
rect 7389 5661 7423 5695
rect 7573 5661 7607 5695
rect 7665 5661 7699 5695
rect 9321 5661 9355 5695
rect 9505 5661 9539 5695
rect 9597 5661 9631 5695
rect 10057 5661 10091 5695
rect 10241 5661 10275 5695
rect 11069 5661 11103 5695
rect 11253 5661 11287 5695
rect 11345 5661 11379 5695
rect 11621 5661 11655 5695
rect 13553 5661 13587 5695
rect 13737 5661 13771 5695
rect 14289 5661 14323 5695
rect 15669 5661 15703 5695
rect 16497 5661 16531 5695
rect 16681 5661 16715 5695
rect 17325 5661 17359 5695
rect 18429 5661 18463 5695
rect 18613 5661 18647 5695
rect 18889 5661 18923 5695
rect 20361 5661 20395 5695
rect 20729 5661 20763 5695
rect 6561 5593 6595 5627
rect 12173 5593 12207 5627
rect 17601 5593 17635 5627
rect 19533 5593 19567 5627
rect 2605 5525 2639 5559
rect 3157 5525 3191 5559
rect 8493 5525 8527 5559
rect 19625 5525 19659 5559
rect 20637 5525 20671 5559
rect 3433 5321 3467 5355
rect 5181 5321 5215 5355
rect 7757 5321 7791 5355
rect 8861 5321 8895 5355
rect 11069 5321 11103 5355
rect 15025 5321 15059 5355
rect 16129 5321 16163 5355
rect 16957 5321 16991 5355
rect 18797 5321 18831 5355
rect 19441 5321 19475 5355
rect 20453 5321 20487 5355
rect 2513 5253 2547 5287
rect 5733 5253 5767 5287
rect 7481 5253 7515 5287
rect 9689 5253 9723 5287
rect 10701 5253 10735 5287
rect 10917 5253 10951 5287
rect 12265 5253 12299 5287
rect 15577 5253 15611 5287
rect 1961 5185 1995 5219
rect 2053 5185 2087 5219
rect 2237 5185 2271 5219
rect 2329 5185 2363 5219
rect 3249 5185 3283 5219
rect 4721 5185 4755 5219
rect 4905 5185 4939 5219
rect 4997 5185 5031 5219
rect 5825 5185 5859 5219
rect 7205 5185 7239 5219
rect 7389 5185 7423 5219
rect 7573 5185 7607 5219
rect 9873 5185 9907 5219
rect 11805 5185 11839 5219
rect 11897 5185 11931 5219
rect 12081 5185 12115 5219
rect 12817 5185 12851 5219
rect 13093 5185 13127 5219
rect 13829 5185 13863 5219
rect 13921 5185 13955 5219
rect 14657 5185 14691 5219
rect 14841 5185 14875 5219
rect 16865 5185 16899 5219
rect 17049 5185 17083 5219
rect 18337 5185 18371 5219
rect 18613 5185 18647 5219
rect 19625 5185 19659 5219
rect 19901 5185 19935 5219
rect 20361 5185 20395 5219
rect 20545 5185 20579 5219
rect 3617 5117 3651 5151
rect 4813 5117 4847 5151
rect 8585 5117 8619 5151
rect 8769 5117 8803 5151
rect 10057 5117 10091 5151
rect 13553 5117 13587 5151
rect 14105 5117 14139 5151
rect 4077 5049 4111 5083
rect 11989 5049 12023 5083
rect 12817 5049 12851 5083
rect 18429 5049 18463 5083
rect 3157 4981 3191 5015
rect 6653 4981 6687 5015
rect 9229 4981 9263 5015
rect 10885 4981 10919 5015
rect 13645 4981 13679 5015
rect 14657 4981 14691 5015
rect 17509 4981 17543 5015
rect 19809 4981 19843 5015
rect 1685 4777 1719 4811
rect 2513 4777 2547 4811
rect 4077 4777 4111 4811
rect 7389 4777 7423 4811
rect 8033 4777 8067 4811
rect 8401 4777 8435 4811
rect 11529 4777 11563 4811
rect 12265 4777 12299 4811
rect 13185 4777 13219 4811
rect 14381 4777 14415 4811
rect 15669 4777 15703 4811
rect 15853 4777 15887 4811
rect 18245 4777 18279 4811
rect 19533 4777 19567 4811
rect 2697 4709 2731 4743
rect 10333 4709 10367 4743
rect 12449 4709 12483 4743
rect 13553 4709 13587 4743
rect 16405 4709 16439 4743
rect 16957 4709 16991 4743
rect 17693 4709 17727 4743
rect 4261 4641 4295 4675
rect 4629 4641 4663 4675
rect 5825 4641 5859 4675
rect 7941 4641 7975 4675
rect 9597 4641 9631 4675
rect 12357 4641 12391 4675
rect 13277 4641 13311 4675
rect 14519 4641 14553 4675
rect 14933 4641 14967 4675
rect 18705 4641 18739 4675
rect 2145 4573 2179 4607
rect 2513 4573 2547 4607
rect 3249 4573 3283 4607
rect 3433 4573 3467 4607
rect 4353 4573 4387 4607
rect 5181 4573 5215 4607
rect 5549 4573 5583 4607
rect 5641 4573 5675 4607
rect 6745 4573 6779 4607
rect 6929 4573 6963 4607
rect 7021 4573 7055 4607
rect 7113 4573 7147 4607
rect 8217 4573 8251 4607
rect 9137 4573 9171 4607
rect 9229 4573 9263 4607
rect 9413 4573 9447 4607
rect 10057 4573 10091 4607
rect 10885 4573 10919 4607
rect 11048 4570 11082 4604
rect 11148 4570 11182 4604
rect 11253 4573 11287 4607
rect 11989 4573 12023 4607
rect 12173 4573 12207 4607
rect 13185 4573 13219 4607
rect 14657 4573 14691 4607
rect 3341 4505 3375 4539
rect 4721 4505 4755 4539
rect 10149 4505 10183 4539
rect 10333 4505 10367 4539
rect 15025 4505 15059 4539
rect 15485 4505 15519 4539
rect 5273 4437 5307 4471
rect 5365 4437 5399 4471
rect 12725 4437 12759 4471
rect 15685 4437 15719 4471
rect 1685 4233 1719 4267
rect 2145 4233 2179 4267
rect 4261 4233 4295 4267
rect 4353 4233 4387 4267
rect 7205 4233 7239 4267
rect 13017 4233 13051 4267
rect 15209 4233 15243 4267
rect 17141 4233 17175 4267
rect 18889 4233 18923 4267
rect 4997 4165 5031 4199
rect 6929 4165 6963 4199
rect 12817 4165 12851 4199
rect 15945 4165 15979 4199
rect 2697 4097 2731 4131
rect 2881 4097 2915 4131
rect 3341 4097 3375 4131
rect 3525 4097 3559 4131
rect 4445 4097 4479 4131
rect 4905 4097 4939 4131
rect 5089 4097 5123 4131
rect 5733 4097 5767 4131
rect 6719 4097 6753 4131
rect 6837 4097 6871 4131
rect 7021 4097 7055 4131
rect 7665 4097 7699 4131
rect 7849 4097 7883 4131
rect 8033 4097 8067 4131
rect 8125 4097 8159 4131
rect 9137 4097 9171 4131
rect 9413 4097 9447 4131
rect 9965 4097 9999 4131
rect 10149 4097 10183 4131
rect 11713 4097 11747 4131
rect 11897 4097 11931 4131
rect 11989 4097 12023 4131
rect 12081 4097 12115 4131
rect 13737 4097 13771 4131
rect 14381 4097 14415 4131
rect 15301 4097 15335 4131
rect 2789 4029 2823 4063
rect 3985 4029 4019 4063
rect 6009 4029 6043 4063
rect 6561 4029 6595 4063
rect 10517 4029 10551 4063
rect 12357 4029 12391 4063
rect 5549 3961 5583 3995
rect 10885 3961 10919 3995
rect 13185 3961 13219 3995
rect 3433 3893 3467 3927
rect 5917 3893 5951 3927
rect 13001 3893 13035 3927
rect 4445 3689 4479 3723
rect 4537 3689 4571 3723
rect 6653 3689 6687 3723
rect 8493 3689 8527 3723
rect 9781 3689 9815 3723
rect 11253 3689 11287 3723
rect 12449 3689 12483 3723
rect 13001 3689 13035 3723
rect 16037 3689 16071 3723
rect 16773 3689 16807 3723
rect 2145 3621 2179 3655
rect 4353 3621 4387 3655
rect 4905 3621 4939 3655
rect 7113 3621 7147 3655
rect 10793 3621 10827 3655
rect 6009 3553 6043 3587
rect 6101 3553 6135 3587
rect 9505 3553 9539 3587
rect 9597 3553 9631 3587
rect 12081 3553 12115 3587
rect 12265 3553 12299 3587
rect 1961 3485 1995 3519
rect 2145 3485 2179 3519
rect 2605 3485 2639 3519
rect 2789 3485 2823 3519
rect 3433 3485 3467 3519
rect 4169 3485 4203 3519
rect 4629 3485 4663 3519
rect 5549 3485 5583 3519
rect 6377 3485 6411 3519
rect 6469 3485 6503 3519
rect 7297 3485 7331 3519
rect 7481 3485 7515 3519
rect 7665 3485 7699 3519
rect 8125 3485 8159 3519
rect 9137 3485 9171 3519
rect 10241 3485 10275 3519
rect 10333 3485 10367 3519
rect 10517 3485 10551 3519
rect 10609 3485 10643 3519
rect 11253 3485 11287 3519
rect 11437 3485 11471 3519
rect 11989 3485 12023 3519
rect 12173 3485 12207 3519
rect 13553 3485 13587 3519
rect 15025 3485 15059 3519
rect 23305 3485 23339 3519
rect 7389 3417 7423 3451
rect 8309 3417 8343 3451
rect 9229 3417 9263 3451
rect 14289 3417 14323 3451
rect 15485 3417 15519 3451
rect 17969 3417 18003 3451
rect 2697 3349 2731 3383
rect 3249 3349 3283 3383
rect 9413 3349 9447 3383
rect 17325 3349 17359 3383
rect 1685 3145 1719 3179
rect 7113 3145 7147 3179
rect 7757 3145 7791 3179
rect 8217 3145 8251 3179
rect 11069 3145 11103 3179
rect 11913 3145 11947 3179
rect 12081 3145 12115 3179
rect 13921 3145 13955 3179
rect 14381 3145 14415 3179
rect 17417 3145 17451 3179
rect 8585 3077 8619 3111
rect 10425 3077 10459 3111
rect 11713 3077 11747 3111
rect 14933 3077 14967 3111
rect 2513 3009 2547 3043
rect 4813 3009 4847 3043
rect 5549 3009 5583 3043
rect 5733 3009 5767 3043
rect 8401 3009 8435 3043
rect 8677 3009 8711 3043
rect 9137 3009 9171 3043
rect 9321 3009 9355 3043
rect 10333 3009 10367 3043
rect 10517 3009 10551 3043
rect 10969 3015 11003 3049
rect 4169 2941 4203 2975
rect 7481 2941 7515 2975
rect 7573 2941 7607 2975
rect 9505 2941 9539 2975
rect 3525 2873 3559 2907
rect 6653 2873 6687 2907
rect 12541 2873 12575 2907
rect 13185 2873 13219 2907
rect 2329 2805 2363 2839
rect 5273 2805 5307 2839
rect 5549 2805 5583 2839
rect 11897 2805 11931 2839
rect 15761 2805 15795 2839
rect 16865 2805 16899 2839
rect 18337 2805 18371 2839
rect 20913 2805 20947 2839
rect 22845 2805 22879 2839
rect 7849 2601 7883 2635
rect 9137 2601 9171 2635
rect 11805 2601 11839 2635
rect 10517 2533 10551 2567
rect 9505 2465 9539 2499
rect 1869 2397 1903 2431
rect 2697 2397 2731 2431
rect 3433 2397 3467 2431
rect 4261 2397 4295 2431
rect 4997 2397 5031 2431
rect 5733 2397 5767 2431
rect 6837 2397 6871 2431
rect 7389 2397 7423 2431
rect 7481 2397 7515 2431
rect 7665 2397 7699 2431
rect 8585 2397 8619 2431
rect 9321 2397 9355 2431
rect 11161 2397 11195 2431
rect 11713 2397 11747 2431
rect 11897 2397 11931 2431
rect 12541 2397 12575 2431
rect 13185 2397 13219 2431
rect 14289 2397 14323 2431
rect 14933 2397 14967 2431
rect 15577 2397 15611 2431
rect 16865 2397 16899 2431
rect 17509 2397 17543 2431
rect 18153 2397 18187 2431
rect 19441 2397 19475 2431
rect 20085 2397 20119 2431
rect 20729 2397 20763 2431
rect 22017 2397 22051 2431
rect 22661 2397 22695 2431
rect 16221 2329 16255 2363
rect 18797 2329 18831 2363
rect 1685 2261 1719 2295
rect 2513 2261 2547 2295
rect 3249 2261 3283 2295
rect 4077 2261 4111 2295
rect 4813 2261 4847 2295
rect 5549 2261 5583 2295
rect 6653 2261 6687 2295
<< metal1 >>
rect 1104 22330 23828 22352
rect 1104 22278 3790 22330
rect 3842 22278 3854 22330
rect 3906 22278 3918 22330
rect 3970 22278 3982 22330
rect 4034 22278 4046 22330
rect 4098 22278 9471 22330
rect 9523 22278 9535 22330
rect 9587 22278 9599 22330
rect 9651 22278 9663 22330
rect 9715 22278 9727 22330
rect 9779 22278 15152 22330
rect 15204 22278 15216 22330
rect 15268 22278 15280 22330
rect 15332 22278 15344 22330
rect 15396 22278 15408 22330
rect 15460 22278 20833 22330
rect 20885 22278 20897 22330
rect 20949 22278 20961 22330
rect 21013 22278 21025 22330
rect 21077 22278 21089 22330
rect 21141 22278 23828 22330
rect 1104 22256 23828 22278
rect 9766 22012 9772 22024
rect 9727 21984 9772 22012
rect 9766 21972 9772 21984
rect 9824 21972 9830 22024
rect 12434 21972 12440 22024
rect 12492 22012 12498 22024
rect 13078 22012 13084 22024
rect 12492 21984 12940 22012
rect 13039 21984 13084 22012
rect 12492 21972 12498 21984
rect 7101 21947 7159 21953
rect 7101 21913 7113 21947
rect 7147 21944 7159 21947
rect 7466 21944 7472 21956
rect 7147 21916 7472 21944
rect 7147 21913 7159 21916
rect 7101 21907 7159 21913
rect 7466 21904 7472 21916
rect 7524 21944 7530 21956
rect 7745 21947 7803 21953
rect 7745 21944 7757 21947
rect 7524 21916 7757 21944
rect 7524 21904 7530 21916
rect 7745 21913 7757 21916
rect 7791 21913 7803 21947
rect 7745 21907 7803 21913
rect 9309 21947 9367 21953
rect 9309 21913 9321 21947
rect 9355 21944 9367 21947
rect 10036 21947 10094 21953
rect 10036 21944 10048 21947
rect 9355 21916 10048 21944
rect 9355 21913 9367 21916
rect 9309 21907 9367 21913
rect 10036 21913 10048 21916
rect 10082 21944 10094 21947
rect 10134 21944 10140 21956
rect 10082 21916 10140 21944
rect 10082 21913 10094 21916
rect 10036 21907 10094 21913
rect 10134 21904 10140 21916
rect 10192 21904 10198 21956
rect 11330 21904 11336 21956
rect 11388 21944 11394 21956
rect 12814 21947 12872 21953
rect 11388 21916 11744 21944
rect 11388 21904 11394 21916
rect 7558 21836 7564 21888
rect 7616 21876 7622 21888
rect 7653 21879 7711 21885
rect 7653 21876 7665 21879
rect 7616 21848 7665 21876
rect 7616 21836 7622 21848
rect 7653 21845 7665 21848
rect 7699 21845 7711 21879
rect 7653 21839 7711 21845
rect 11149 21879 11207 21885
rect 11149 21845 11161 21879
rect 11195 21876 11207 21879
rect 11422 21876 11428 21888
rect 11195 21848 11428 21876
rect 11195 21845 11207 21848
rect 11149 21839 11207 21845
rect 11422 21836 11428 21848
rect 11480 21836 11486 21888
rect 11716 21885 11744 21916
rect 12814 21913 12826 21947
rect 12860 21913 12872 21947
rect 12912 21944 12940 21984
rect 13078 21972 13084 21984
rect 13136 21972 13142 22024
rect 13541 22015 13599 22021
rect 13541 21981 13553 22015
rect 13587 22012 13599 22015
rect 15105 22015 15163 22021
rect 15105 22012 15117 22015
rect 13587 21984 15117 22012
rect 13587 21981 13599 21984
rect 13541 21975 13599 21981
rect 15105 21981 15117 21984
rect 15151 21981 15163 22015
rect 15105 21975 15163 21981
rect 13556 21944 13584 21975
rect 17402 21972 17408 22024
rect 17460 22012 17466 22024
rect 17681 22015 17739 22021
rect 17681 22012 17693 22015
rect 17460 21984 17693 22012
rect 17460 21972 17466 21984
rect 17681 21981 17693 21984
rect 17727 22012 17739 22015
rect 18141 22015 18199 22021
rect 18141 22012 18153 22015
rect 17727 21984 18153 22012
rect 17727 21981 17739 21984
rect 17681 21975 17739 21981
rect 18141 21981 18153 21984
rect 18187 21981 18199 22015
rect 18141 21975 18199 21981
rect 22370 21972 22376 22024
rect 22428 22012 22434 22024
rect 22649 22015 22707 22021
rect 22649 22012 22661 22015
rect 22428 21984 22661 22012
rect 22428 21972 22434 21984
rect 22649 21981 22661 21984
rect 22695 22012 22707 22015
rect 23109 22015 23167 22021
rect 23109 22012 23121 22015
rect 22695 21984 23121 22012
rect 22695 21981 22707 21984
rect 22649 21975 22707 21981
rect 23109 21981 23121 21984
rect 23155 21981 23167 22015
rect 23109 21975 23167 21981
rect 12912 21916 13584 21944
rect 14277 21947 14335 21953
rect 12814 21907 12872 21913
rect 14277 21913 14289 21947
rect 14323 21944 14335 21947
rect 14366 21944 14372 21956
rect 14323 21916 14372 21944
rect 14323 21913 14335 21916
rect 14277 21907 14335 21913
rect 11701 21879 11759 21885
rect 11701 21845 11713 21879
rect 11747 21845 11759 21879
rect 12820 21876 12848 21907
rect 14366 21904 14372 21916
rect 14424 21904 14430 21956
rect 14461 21947 14519 21953
rect 14461 21913 14473 21947
rect 14507 21913 14519 21947
rect 14461 21907 14519 21913
rect 13538 21876 13544 21888
rect 12820 21848 13544 21876
rect 11701 21839 11759 21845
rect 13538 21836 13544 21848
rect 13596 21836 13602 21888
rect 13722 21876 13728 21888
rect 13683 21848 13728 21876
rect 13722 21836 13728 21848
rect 13780 21876 13786 21888
rect 14476 21876 14504 21907
rect 14550 21904 14556 21956
rect 14608 21944 14614 21956
rect 14608 21916 22508 21944
rect 14608 21904 14614 21916
rect 14642 21876 14648 21888
rect 13780 21848 14504 21876
rect 14603 21848 14648 21876
rect 13780 21836 13786 21848
rect 14642 21836 14648 21848
rect 14700 21836 14706 21888
rect 17494 21876 17500 21888
rect 17455 21848 17500 21876
rect 17494 21836 17500 21848
rect 17552 21836 17558 21888
rect 22480 21885 22508 21916
rect 22465 21879 22523 21885
rect 22465 21845 22477 21879
rect 22511 21845 22523 21879
rect 22465 21839 22523 21845
rect 1104 21786 23987 21808
rect 1104 21734 6630 21786
rect 6682 21734 6694 21786
rect 6746 21734 6758 21786
rect 6810 21734 6822 21786
rect 6874 21734 6886 21786
rect 6938 21734 12311 21786
rect 12363 21734 12375 21786
rect 12427 21734 12439 21786
rect 12491 21734 12503 21786
rect 12555 21734 12567 21786
rect 12619 21734 17992 21786
rect 18044 21734 18056 21786
rect 18108 21734 18120 21786
rect 18172 21734 18184 21786
rect 18236 21734 18248 21786
rect 18300 21734 23673 21786
rect 23725 21734 23737 21786
rect 23789 21734 23801 21786
rect 23853 21734 23865 21786
rect 23917 21734 23929 21786
rect 23981 21734 23987 21786
rect 1104 21712 23987 21734
rect 12836 21607 12894 21613
rect 12836 21573 12848 21607
rect 12882 21604 12894 21607
rect 13541 21607 13599 21613
rect 13541 21604 13553 21607
rect 12882 21576 13553 21604
rect 12882 21573 12894 21576
rect 12836 21567 12894 21573
rect 13541 21573 13553 21576
rect 13587 21573 13599 21607
rect 13541 21567 13599 21573
rect 7765 21539 7823 21545
rect 7765 21505 7777 21539
rect 7811 21536 7823 21539
rect 9306 21536 9312 21548
rect 7811 21508 9312 21536
rect 7811 21505 7823 21508
rect 7765 21499 7823 21505
rect 9306 21496 9312 21508
rect 9364 21496 9370 21548
rect 10036 21539 10094 21545
rect 10036 21505 10048 21539
rect 10082 21536 10094 21539
rect 11238 21536 11244 21548
rect 10082 21508 11244 21536
rect 10082 21505 10094 21508
rect 10036 21499 10094 21505
rect 11238 21496 11244 21508
rect 11296 21496 11302 21548
rect 13725 21539 13783 21545
rect 13725 21505 13737 21539
rect 13771 21536 13783 21539
rect 14642 21536 14648 21548
rect 13771 21508 14648 21536
rect 13771 21505 13783 21508
rect 13725 21499 13783 21505
rect 14642 21496 14648 21508
rect 14700 21496 14706 21548
rect 14829 21539 14887 21545
rect 14829 21505 14841 21539
rect 14875 21505 14887 21539
rect 14829 21499 14887 21505
rect 8021 21471 8079 21477
rect 8021 21437 8033 21471
rect 8067 21468 8079 21471
rect 9766 21468 9772 21480
rect 8067 21440 9772 21468
rect 8067 21437 8079 21440
rect 8021 21431 8079 21437
rect 9766 21428 9772 21440
rect 9824 21428 9830 21480
rect 13078 21428 13084 21480
rect 13136 21468 13142 21480
rect 13817 21471 13875 21477
rect 13136 21440 13229 21468
rect 13136 21428 13142 21440
rect 13817 21437 13829 21471
rect 13863 21437 13875 21471
rect 14182 21468 14188 21480
rect 14143 21440 14188 21468
rect 13817 21431 13875 21437
rect 11054 21360 11060 21412
rect 11112 21400 11118 21412
rect 11701 21403 11759 21409
rect 11701 21400 11713 21403
rect 11112 21372 11713 21400
rect 11112 21360 11118 21372
rect 11701 21369 11713 21372
rect 11747 21369 11759 21403
rect 11701 21363 11759 21369
rect 6641 21335 6699 21341
rect 6641 21301 6653 21335
rect 6687 21332 6699 21335
rect 7098 21332 7104 21344
rect 6687 21304 7104 21332
rect 6687 21301 6699 21304
rect 6641 21295 6699 21301
rect 7098 21292 7104 21304
rect 7156 21292 7162 21344
rect 11149 21335 11207 21341
rect 11149 21301 11161 21335
rect 11195 21332 11207 21335
rect 11514 21332 11520 21344
rect 11195 21304 11520 21332
rect 11195 21301 11207 21304
rect 11149 21295 11207 21301
rect 11514 21292 11520 21304
rect 11572 21292 11578 21344
rect 11790 21292 11796 21344
rect 11848 21332 11854 21344
rect 13096 21332 13124 21428
rect 13354 21360 13360 21412
rect 13412 21400 13418 21412
rect 13832 21400 13860 21431
rect 14182 21428 14188 21440
rect 14240 21468 14246 21480
rect 14844 21468 14872 21499
rect 14240 21440 14872 21468
rect 14240 21428 14246 21440
rect 17494 21400 17500 21412
rect 13412 21372 17500 21400
rect 13412 21360 13418 21372
rect 17494 21360 17500 21372
rect 17552 21360 17558 21412
rect 11848 21304 13124 21332
rect 11848 21292 11854 21304
rect 13446 21292 13452 21344
rect 13504 21332 13510 21344
rect 14737 21335 14795 21341
rect 14737 21332 14749 21335
rect 13504 21304 14749 21332
rect 13504 21292 13510 21304
rect 14737 21301 14749 21304
rect 14783 21301 14795 21335
rect 14737 21295 14795 21301
rect 1104 21242 23828 21264
rect 1104 21190 3790 21242
rect 3842 21190 3854 21242
rect 3906 21190 3918 21242
rect 3970 21190 3982 21242
rect 4034 21190 4046 21242
rect 4098 21190 9471 21242
rect 9523 21190 9535 21242
rect 9587 21190 9599 21242
rect 9651 21190 9663 21242
rect 9715 21190 9727 21242
rect 9779 21190 15152 21242
rect 15204 21190 15216 21242
rect 15268 21190 15280 21242
rect 15332 21190 15344 21242
rect 15396 21190 15408 21242
rect 15460 21190 20833 21242
rect 20885 21190 20897 21242
rect 20949 21190 20961 21242
rect 21013 21190 21025 21242
rect 21077 21190 21089 21242
rect 21141 21190 23828 21242
rect 1104 21168 23828 21190
rect 2498 21088 2504 21140
rect 2556 21128 2562 21140
rect 7098 21128 7104 21140
rect 2556 21100 7104 21128
rect 2556 21088 2562 21100
rect 7098 21088 7104 21100
rect 7156 21088 7162 21140
rect 9858 21088 9864 21140
rect 9916 21128 9922 21140
rect 11146 21128 11152 21140
rect 9916 21100 11152 21128
rect 9916 21088 9922 21100
rect 11146 21088 11152 21100
rect 11204 21128 11210 21140
rect 11701 21131 11759 21137
rect 11701 21128 11713 21131
rect 11204 21100 11713 21128
rect 11204 21088 11210 21100
rect 11701 21097 11713 21100
rect 11747 21128 11759 21131
rect 11790 21128 11796 21140
rect 11747 21100 11796 21128
rect 11747 21097 11759 21100
rect 11701 21091 11759 21097
rect 11790 21088 11796 21100
rect 11848 21088 11854 21140
rect 9306 21020 9312 21072
rect 9364 21060 9370 21072
rect 12989 21063 13047 21069
rect 12989 21060 13001 21063
rect 9364 21032 13001 21060
rect 9364 21020 9370 21032
rect 12989 21029 13001 21032
rect 13035 21029 13047 21063
rect 12989 21023 13047 21029
rect 13446 20992 13452 21004
rect 13407 20964 13452 20992
rect 13446 20952 13452 20964
rect 13504 20952 13510 21004
rect 5534 20884 5540 20936
rect 5592 20924 5598 20936
rect 6273 20927 6331 20933
rect 6273 20924 6285 20927
rect 5592 20896 6285 20924
rect 5592 20884 5598 20896
rect 6273 20893 6285 20896
rect 6319 20924 6331 20927
rect 6733 20927 6791 20933
rect 6733 20924 6745 20927
rect 6319 20896 6745 20924
rect 6319 20893 6331 20896
rect 6273 20887 6331 20893
rect 6733 20893 6745 20896
rect 6779 20893 6791 20927
rect 13354 20924 13360 20936
rect 13315 20896 13360 20924
rect 6733 20887 6791 20893
rect 13354 20884 13360 20896
rect 13412 20884 13418 20936
rect 6028 20859 6086 20865
rect 6028 20825 6040 20859
rect 6074 20856 6086 20859
rect 6178 20856 6184 20868
rect 6074 20828 6184 20856
rect 6074 20825 6086 20828
rect 6028 20819 6086 20825
rect 6178 20816 6184 20828
rect 6236 20816 6242 20868
rect 7000 20859 7058 20865
rect 7000 20825 7012 20859
rect 7046 20856 7058 20859
rect 7650 20856 7656 20868
rect 7046 20828 7656 20856
rect 7046 20825 7058 20828
rect 7000 20819 7058 20825
rect 7650 20816 7656 20828
rect 7708 20816 7714 20868
rect 8938 20816 8944 20868
rect 8996 20856 9002 20868
rect 10413 20859 10471 20865
rect 10413 20856 10425 20859
rect 8996 20828 10425 20856
rect 8996 20816 9002 20828
rect 10413 20825 10425 20828
rect 10459 20825 10471 20859
rect 10413 20819 10471 20825
rect 4890 20788 4896 20800
rect 4851 20760 4896 20788
rect 4890 20748 4896 20760
rect 4948 20748 4954 20800
rect 8110 20788 8116 20800
rect 8071 20760 8116 20788
rect 8110 20748 8116 20760
rect 8168 20748 8174 20800
rect 1104 20698 23987 20720
rect 1104 20646 6630 20698
rect 6682 20646 6694 20698
rect 6746 20646 6758 20698
rect 6810 20646 6822 20698
rect 6874 20646 6886 20698
rect 6938 20646 12311 20698
rect 12363 20646 12375 20698
rect 12427 20646 12439 20698
rect 12491 20646 12503 20698
rect 12555 20646 12567 20698
rect 12619 20646 17992 20698
rect 18044 20646 18056 20698
rect 18108 20646 18120 20698
rect 18172 20646 18184 20698
rect 18236 20646 18248 20698
rect 18300 20646 23673 20698
rect 23725 20646 23737 20698
rect 23789 20646 23801 20698
rect 23853 20646 23865 20698
rect 23917 20646 23929 20698
rect 23981 20646 23987 20698
rect 1104 20624 23987 20646
rect 13081 20587 13139 20593
rect 13081 20553 13093 20587
rect 13127 20584 13139 20587
rect 14182 20584 14188 20596
rect 13127 20556 14188 20584
rect 13127 20553 13139 20556
rect 13081 20547 13139 20553
rect 14182 20544 14188 20556
rect 14240 20544 14246 20596
rect 10904 20519 10962 20525
rect 10904 20485 10916 20519
rect 10950 20516 10962 20519
rect 12710 20516 12716 20528
rect 10950 20488 12716 20516
rect 10950 20485 10962 20488
rect 10904 20479 10962 20485
rect 12710 20476 12716 20488
rect 12768 20476 12774 20528
rect 14366 20516 14372 20528
rect 12912 20488 14372 20516
rect 4890 20408 4896 20460
rect 4948 20448 4954 20460
rect 5362 20451 5420 20457
rect 5362 20448 5374 20451
rect 4948 20420 5374 20448
rect 4948 20408 4954 20420
rect 5362 20417 5374 20420
rect 5408 20417 5420 20451
rect 5362 20411 5420 20417
rect 5534 20408 5540 20460
rect 5592 20448 5598 20460
rect 5629 20451 5687 20457
rect 5629 20448 5641 20451
rect 5592 20420 5641 20448
rect 5592 20408 5598 20420
rect 5629 20417 5641 20420
rect 5675 20448 5687 20451
rect 7193 20451 7251 20457
rect 7193 20448 7205 20451
rect 5675 20420 7205 20448
rect 5675 20417 5687 20420
rect 5629 20411 5687 20417
rect 7193 20417 7205 20420
rect 7239 20417 7251 20451
rect 7193 20411 7251 20417
rect 7282 20408 7288 20460
rect 7340 20448 7346 20460
rect 7449 20451 7507 20457
rect 7449 20448 7461 20451
rect 7340 20420 7461 20448
rect 7340 20408 7346 20420
rect 7449 20417 7461 20420
rect 7495 20417 7507 20451
rect 11146 20448 11152 20460
rect 11107 20420 11152 20448
rect 7449 20411 7507 20417
rect 11146 20408 11152 20420
rect 11204 20408 11210 20460
rect 12912 20457 12940 20488
rect 14366 20476 14372 20488
rect 14424 20476 14430 20528
rect 12897 20451 12955 20457
rect 12897 20417 12909 20451
rect 12943 20417 12955 20451
rect 12897 20411 12955 20417
rect 13081 20451 13139 20457
rect 13081 20417 13093 20451
rect 13127 20448 13139 20451
rect 13722 20448 13728 20460
rect 13127 20420 13728 20448
rect 13127 20417 13139 20420
rect 13081 20411 13139 20417
rect 13722 20408 13728 20420
rect 13780 20408 13786 20460
rect 4249 20247 4307 20253
rect 4249 20213 4261 20247
rect 4295 20244 4307 20247
rect 4430 20244 4436 20256
rect 4295 20216 4436 20244
rect 4295 20213 4307 20216
rect 4249 20207 4307 20213
rect 4430 20204 4436 20216
rect 4488 20204 4494 20256
rect 8110 20204 8116 20256
rect 8168 20244 8174 20256
rect 8573 20247 8631 20253
rect 8573 20244 8585 20247
rect 8168 20216 8585 20244
rect 8168 20204 8174 20216
rect 8573 20213 8585 20216
rect 8619 20213 8631 20247
rect 8573 20207 8631 20213
rect 9769 20247 9827 20253
rect 9769 20213 9781 20247
rect 9815 20244 9827 20247
rect 10410 20244 10416 20256
rect 9815 20216 10416 20244
rect 9815 20213 9827 20216
rect 9769 20207 9827 20213
rect 10410 20204 10416 20216
rect 10468 20204 10474 20256
rect 11238 20204 11244 20256
rect 11296 20244 11302 20256
rect 11701 20247 11759 20253
rect 11701 20244 11713 20247
rect 11296 20216 11713 20244
rect 11296 20204 11302 20216
rect 11701 20213 11713 20216
rect 11747 20213 11759 20247
rect 11701 20207 11759 20213
rect 1104 20154 23828 20176
rect 1104 20102 3790 20154
rect 3842 20102 3854 20154
rect 3906 20102 3918 20154
rect 3970 20102 3982 20154
rect 4034 20102 4046 20154
rect 4098 20102 9471 20154
rect 9523 20102 9535 20154
rect 9587 20102 9599 20154
rect 9651 20102 9663 20154
rect 9715 20102 9727 20154
rect 9779 20102 15152 20154
rect 15204 20102 15216 20154
rect 15268 20102 15280 20154
rect 15332 20102 15344 20154
rect 15396 20102 15408 20154
rect 15460 20102 20833 20154
rect 20885 20102 20897 20154
rect 20949 20102 20961 20154
rect 21013 20102 21025 20154
rect 21077 20102 21089 20154
rect 21141 20102 23828 20154
rect 1104 20080 23828 20102
rect 11146 19904 11152 19916
rect 11107 19876 11152 19904
rect 11146 19864 11152 19876
rect 11204 19864 11210 19916
rect 3973 19839 4031 19845
rect 3973 19805 3985 19839
rect 4019 19836 4031 19839
rect 5534 19836 5540 19848
rect 4019 19808 5540 19836
rect 4019 19805 4031 19808
rect 3973 19799 4031 19805
rect 5534 19796 5540 19808
rect 5592 19796 5598 19848
rect 8205 19839 8263 19845
rect 8205 19805 8217 19839
rect 8251 19836 8263 19839
rect 8294 19836 8300 19848
rect 8251 19808 8300 19836
rect 8251 19805 8263 19808
rect 8205 19799 8263 19805
rect 8294 19796 8300 19808
rect 8352 19796 8358 19848
rect 11164 19836 11192 19864
rect 11698 19836 11704 19848
rect 11164 19808 11704 19836
rect 11698 19796 11704 19808
rect 11756 19836 11762 19848
rect 12989 19839 13047 19845
rect 12989 19836 13001 19839
rect 11756 19808 13001 19836
rect 11756 19796 11762 19808
rect 12989 19805 13001 19808
rect 13035 19805 13047 19839
rect 12989 19799 13047 19805
rect 4246 19777 4252 19780
rect 4240 19731 4252 19777
rect 4304 19768 4310 19780
rect 7960 19771 8018 19777
rect 4304 19740 4340 19768
rect 4246 19728 4252 19731
rect 4304 19728 4310 19740
rect 7960 19737 7972 19771
rect 8006 19768 8018 19771
rect 10882 19771 10940 19777
rect 8006 19740 8248 19768
rect 8006 19737 8018 19740
rect 7960 19731 8018 19737
rect 8220 19712 8248 19740
rect 10882 19737 10894 19771
rect 10928 19737 10940 19771
rect 10882 19731 10940 19737
rect 12744 19771 12802 19777
rect 12744 19737 12756 19771
rect 12790 19768 12802 19771
rect 18322 19768 18328 19780
rect 12790 19740 18328 19768
rect 12790 19737 12802 19740
rect 12744 19731 12802 19737
rect 2130 19660 2136 19712
rect 2188 19700 2194 19712
rect 5353 19703 5411 19709
rect 5353 19700 5365 19703
rect 2188 19672 5365 19700
rect 2188 19660 2194 19672
rect 5353 19669 5365 19672
rect 5399 19669 5411 19703
rect 5353 19663 5411 19669
rect 6362 19660 6368 19712
rect 6420 19700 6426 19712
rect 6825 19703 6883 19709
rect 6825 19700 6837 19703
rect 6420 19672 6837 19700
rect 6420 19660 6426 19672
rect 6825 19669 6837 19672
rect 6871 19669 6883 19703
rect 6825 19663 6883 19669
rect 8202 19660 8208 19712
rect 8260 19660 8266 19712
rect 9769 19703 9827 19709
rect 9769 19669 9781 19703
rect 9815 19700 9827 19703
rect 10778 19700 10784 19712
rect 9815 19672 10784 19700
rect 9815 19669 9827 19672
rect 9769 19663 9827 19669
rect 10778 19660 10784 19672
rect 10836 19660 10842 19712
rect 10888 19700 10916 19731
rect 18322 19728 18328 19740
rect 18380 19728 18386 19780
rect 10962 19700 10968 19712
rect 10888 19672 10968 19700
rect 10962 19660 10968 19672
rect 11020 19660 11026 19712
rect 11606 19700 11612 19712
rect 11567 19672 11612 19700
rect 11606 19660 11612 19672
rect 11664 19660 11670 19712
rect 1104 19610 23987 19632
rect 1104 19558 6630 19610
rect 6682 19558 6694 19610
rect 6746 19558 6758 19610
rect 6810 19558 6822 19610
rect 6874 19558 6886 19610
rect 6938 19558 12311 19610
rect 12363 19558 12375 19610
rect 12427 19558 12439 19610
rect 12491 19558 12503 19610
rect 12555 19558 12567 19610
rect 12619 19558 17992 19610
rect 18044 19558 18056 19610
rect 18108 19558 18120 19610
rect 18172 19558 18184 19610
rect 18236 19558 18248 19610
rect 18300 19558 23673 19610
rect 23725 19558 23737 19610
rect 23789 19558 23801 19610
rect 23853 19558 23865 19610
rect 23917 19558 23929 19610
rect 23981 19558 23987 19610
rect 1104 19536 23987 19558
rect 3694 19496 3700 19508
rect 3655 19468 3700 19496
rect 3694 19456 3700 19468
rect 3752 19456 3758 19508
rect 7098 19496 7104 19508
rect 7059 19468 7104 19496
rect 7098 19456 7104 19468
rect 7156 19456 7162 19508
rect 4832 19431 4890 19437
rect 4832 19397 4844 19431
rect 4878 19428 4890 19431
rect 5902 19428 5908 19440
rect 4878 19400 5908 19428
rect 4878 19397 4890 19400
rect 4832 19391 4890 19397
rect 5902 19388 5908 19400
rect 5960 19388 5966 19440
rect 7116 19428 7144 19456
rect 7653 19431 7711 19437
rect 7653 19428 7665 19431
rect 7116 19400 7665 19428
rect 7653 19397 7665 19400
rect 7699 19397 7711 19431
rect 7653 19391 7711 19397
rect 5077 19363 5135 19369
rect 5077 19329 5089 19363
rect 5123 19360 5135 19363
rect 5534 19360 5540 19372
rect 5123 19332 5540 19360
rect 5123 19329 5135 19332
rect 5077 19323 5135 19329
rect 5534 19320 5540 19332
rect 5592 19320 5598 19372
rect 8938 19156 8944 19168
rect 8899 19128 8944 19156
rect 8938 19116 8944 19128
rect 8996 19116 9002 19168
rect 1104 19066 23828 19088
rect 1104 19014 3790 19066
rect 3842 19014 3854 19066
rect 3906 19014 3918 19066
rect 3970 19014 3982 19066
rect 4034 19014 4046 19066
rect 4098 19014 9471 19066
rect 9523 19014 9535 19066
rect 9587 19014 9599 19066
rect 9651 19014 9663 19066
rect 9715 19014 9727 19066
rect 9779 19014 15152 19066
rect 15204 19014 15216 19066
rect 15268 19014 15280 19066
rect 15332 19014 15344 19066
rect 15396 19014 15408 19066
rect 15460 19014 20833 19066
rect 20885 19014 20897 19066
rect 20949 19014 20961 19066
rect 21013 19014 21025 19066
rect 21077 19014 21089 19066
rect 21141 19014 23828 19066
rect 1104 18992 23828 19014
rect 2501 18955 2559 18961
rect 2501 18921 2513 18955
rect 2547 18952 2559 18955
rect 4246 18952 4252 18964
rect 2547 18924 4252 18952
rect 2547 18921 2559 18924
rect 2501 18915 2559 18921
rect 4246 18912 4252 18924
rect 4304 18912 4310 18964
rect 18233 18955 18291 18961
rect 18233 18921 18245 18955
rect 18279 18952 18291 18955
rect 18322 18952 18328 18964
rect 18279 18924 18328 18952
rect 18279 18921 18291 18924
rect 18233 18915 18291 18921
rect 18322 18912 18328 18924
rect 18380 18912 18386 18964
rect 6825 18819 6883 18825
rect 6825 18816 6837 18819
rect 6288 18788 6837 18816
rect 2314 18748 2320 18760
rect 2275 18720 2320 18748
rect 2314 18708 2320 18720
rect 2372 18708 2378 18760
rect 5534 18708 5540 18760
rect 5592 18748 5598 18760
rect 6288 18748 6316 18788
rect 6825 18785 6837 18788
rect 6871 18785 6883 18819
rect 11698 18816 11704 18828
rect 11659 18788 11704 18816
rect 6825 18779 6883 18785
rect 11698 18776 11704 18788
rect 11756 18776 11762 18828
rect 5592 18720 6316 18748
rect 6365 18751 6423 18757
rect 5592 18708 5598 18720
rect 6365 18717 6377 18751
rect 6411 18748 6423 18751
rect 8294 18748 8300 18760
rect 6411 18720 8300 18748
rect 6411 18717 6423 18720
rect 6365 18711 6423 18717
rect 8294 18708 8300 18720
rect 8352 18708 8358 18760
rect 8386 18708 8392 18760
rect 8444 18748 8450 18760
rect 9309 18751 9367 18757
rect 9309 18748 9321 18751
rect 8444 18720 9321 18748
rect 8444 18708 8450 18720
rect 9309 18717 9321 18720
rect 9355 18717 9367 18751
rect 9309 18711 9367 18717
rect 11425 18751 11483 18757
rect 11425 18717 11437 18751
rect 11471 18748 11483 18751
rect 18414 18748 18420 18760
rect 11471 18720 12296 18748
rect 18375 18720 18420 18748
rect 11471 18717 11483 18720
rect 11425 18711 11483 18717
rect 6086 18680 6092 18692
rect 6144 18689 6150 18692
rect 6056 18652 6092 18680
rect 6086 18640 6092 18652
rect 6144 18643 6156 18689
rect 7092 18683 7150 18689
rect 7092 18649 7104 18683
rect 7138 18680 7150 18683
rect 7138 18652 9168 18680
rect 7138 18649 7150 18652
rect 7092 18643 7150 18649
rect 6144 18640 6150 18643
rect 4985 18615 5043 18621
rect 4985 18581 4997 18615
rect 5031 18612 5043 18615
rect 5074 18612 5080 18624
rect 5031 18584 5080 18612
rect 5031 18581 5043 18584
rect 4985 18575 5043 18581
rect 5074 18572 5080 18584
rect 5132 18572 5138 18624
rect 8018 18572 8024 18624
rect 8076 18612 8082 18624
rect 9140 18621 9168 18652
rect 8205 18615 8263 18621
rect 8205 18612 8217 18615
rect 8076 18584 8217 18612
rect 8076 18572 8082 18584
rect 8205 18581 8217 18584
rect 8251 18581 8263 18615
rect 8205 18575 8263 18581
rect 9125 18615 9183 18621
rect 9125 18581 9137 18615
rect 9171 18581 9183 18615
rect 9125 18575 9183 18581
rect 10321 18615 10379 18621
rect 10321 18581 10333 18615
rect 10367 18612 10379 18615
rect 11698 18612 11704 18624
rect 10367 18584 11704 18612
rect 10367 18581 10379 18584
rect 10321 18575 10379 18581
rect 11698 18572 11704 18584
rect 11756 18572 11762 18624
rect 12268 18621 12296 18720
rect 18414 18708 18420 18720
rect 18472 18708 18478 18760
rect 12253 18615 12311 18621
rect 12253 18581 12265 18615
rect 12299 18612 12311 18615
rect 13446 18612 13452 18624
rect 12299 18584 13452 18612
rect 12299 18581 12311 18584
rect 12253 18575 12311 18581
rect 13446 18572 13452 18584
rect 13504 18572 13510 18624
rect 1104 18522 23987 18544
rect 1104 18470 6630 18522
rect 6682 18470 6694 18522
rect 6746 18470 6758 18522
rect 6810 18470 6822 18522
rect 6874 18470 6886 18522
rect 6938 18470 12311 18522
rect 12363 18470 12375 18522
rect 12427 18470 12439 18522
rect 12491 18470 12503 18522
rect 12555 18470 12567 18522
rect 12619 18470 17992 18522
rect 18044 18470 18056 18522
rect 18108 18470 18120 18522
rect 18172 18470 18184 18522
rect 18236 18470 18248 18522
rect 18300 18470 23673 18522
rect 23725 18470 23737 18522
rect 23789 18470 23801 18522
rect 23853 18470 23865 18522
rect 23917 18470 23929 18522
rect 23981 18470 23987 18522
rect 1104 18448 23987 18470
rect 4338 18232 4344 18284
rect 4396 18272 4402 18284
rect 7374 18281 7380 18284
rect 4626 18275 4684 18281
rect 4626 18272 4638 18275
rect 4396 18244 4638 18272
rect 4396 18232 4402 18244
rect 4626 18241 4638 18244
rect 4672 18241 4684 18275
rect 4626 18235 4684 18241
rect 7368 18235 7380 18281
rect 7432 18272 7438 18284
rect 7432 18244 7468 18272
rect 7374 18232 7380 18235
rect 7432 18232 7438 18244
rect 8294 18232 8300 18284
rect 8352 18272 8358 18284
rect 9306 18272 9312 18284
rect 8352 18244 9312 18272
rect 8352 18232 8358 18244
rect 9306 18232 9312 18244
rect 9364 18272 9370 18284
rect 9769 18275 9827 18281
rect 9769 18272 9781 18275
rect 9364 18244 9781 18272
rect 9364 18232 9370 18244
rect 9769 18241 9781 18244
rect 9815 18241 9827 18275
rect 9769 18235 9827 18241
rect 10036 18275 10094 18281
rect 10036 18241 10048 18275
rect 10082 18272 10094 18275
rect 12066 18272 12072 18284
rect 10082 18244 12072 18272
rect 10082 18241 10094 18244
rect 10036 18235 10094 18241
rect 12066 18232 12072 18244
rect 12124 18272 12130 18284
rect 12253 18275 12311 18281
rect 12253 18272 12265 18275
rect 12124 18244 12265 18272
rect 12124 18232 12130 18244
rect 12253 18241 12265 18244
rect 12299 18241 12311 18275
rect 12253 18235 12311 18241
rect 4893 18207 4951 18213
rect 4893 18173 4905 18207
rect 4939 18204 4951 18207
rect 7098 18204 7104 18216
rect 4939 18176 7104 18204
rect 4939 18173 4951 18176
rect 4893 18167 4951 18173
rect 3510 18068 3516 18080
rect 3471 18040 3516 18068
rect 3510 18028 3516 18040
rect 3568 18028 3574 18080
rect 4614 18028 4620 18080
rect 4672 18068 4678 18080
rect 4908 18068 4936 18167
rect 7098 18164 7104 18176
rect 7156 18164 7162 18216
rect 11149 18139 11207 18145
rect 11149 18105 11161 18139
rect 11195 18136 11207 18139
rect 11882 18136 11888 18148
rect 11195 18108 11888 18136
rect 11195 18105 11207 18108
rect 11149 18099 11207 18105
rect 11882 18096 11888 18108
rect 11940 18096 11946 18148
rect 4672 18040 4936 18068
rect 8481 18071 8539 18077
rect 4672 18028 4678 18040
rect 8481 18037 8493 18071
rect 8527 18068 8539 18071
rect 9122 18068 9128 18080
rect 8527 18040 9128 18068
rect 8527 18037 8539 18040
rect 8481 18031 8539 18037
rect 9122 18028 9128 18040
rect 9180 18028 9186 18080
rect 11790 18068 11796 18080
rect 11751 18040 11796 18068
rect 11790 18028 11796 18040
rect 11848 18028 11854 18080
rect 1104 17978 23828 18000
rect 1104 17926 3790 17978
rect 3842 17926 3854 17978
rect 3906 17926 3918 17978
rect 3970 17926 3982 17978
rect 4034 17926 4046 17978
rect 4098 17926 9471 17978
rect 9523 17926 9535 17978
rect 9587 17926 9599 17978
rect 9651 17926 9663 17978
rect 9715 17926 9727 17978
rect 9779 17926 15152 17978
rect 15204 17926 15216 17978
rect 15268 17926 15280 17978
rect 15332 17926 15344 17978
rect 15396 17926 15408 17978
rect 15460 17926 20833 17978
rect 20885 17926 20897 17978
rect 20949 17926 20961 17978
rect 21013 17926 21025 17978
rect 21077 17926 21089 17978
rect 21141 17926 23828 17978
rect 1104 17904 23828 17926
rect 5534 17864 5540 17876
rect 5495 17836 5540 17864
rect 5534 17824 5540 17836
rect 5592 17824 5598 17876
rect 8110 17824 8116 17876
rect 8168 17864 8174 17876
rect 8297 17867 8355 17873
rect 8297 17864 8309 17867
rect 8168 17836 8309 17864
rect 8168 17824 8174 17836
rect 8297 17833 8309 17836
rect 8343 17833 8355 17867
rect 8297 17827 8355 17833
rect 2041 17663 2099 17669
rect 2041 17629 2053 17663
rect 2087 17660 2099 17663
rect 4614 17660 4620 17672
rect 2087 17632 4620 17660
rect 2087 17629 2099 17632
rect 2041 17623 2099 17629
rect 4614 17620 4620 17632
rect 4672 17620 4678 17672
rect 7466 17660 7472 17672
rect 7427 17632 7472 17660
rect 7466 17620 7472 17632
rect 7524 17620 7530 17672
rect 9306 17620 9312 17672
rect 9364 17660 9370 17672
rect 11146 17660 11152 17672
rect 9364 17632 11152 17660
rect 9364 17620 9370 17632
rect 11146 17620 11152 17632
rect 11204 17660 11210 17672
rect 11241 17663 11299 17669
rect 11241 17660 11253 17663
rect 11204 17632 11253 17660
rect 11204 17620 11210 17632
rect 11241 17629 11253 17632
rect 11287 17660 11299 17663
rect 11701 17663 11759 17669
rect 11701 17660 11713 17663
rect 11287 17632 11713 17660
rect 11287 17629 11299 17632
rect 11241 17623 11299 17629
rect 11701 17629 11713 17632
rect 11747 17629 11759 17663
rect 11701 17623 11759 17629
rect 2308 17595 2366 17601
rect 2308 17561 2320 17595
rect 2354 17592 2366 17595
rect 2498 17592 2504 17604
rect 2354 17564 2504 17592
rect 2354 17561 2366 17564
rect 2308 17555 2366 17561
rect 2498 17552 2504 17564
rect 2556 17552 2562 17604
rect 7006 17592 7012 17604
rect 6967 17564 7012 17592
rect 7006 17552 7012 17564
rect 7064 17552 7070 17604
rect 10996 17595 11054 17601
rect 10996 17561 11008 17595
rect 11042 17592 11054 17595
rect 11790 17592 11796 17604
rect 11042 17564 11796 17592
rect 11042 17561 11054 17564
rect 10996 17555 11054 17561
rect 11790 17552 11796 17564
rect 11848 17552 11854 17604
rect 11968 17595 12026 17601
rect 11968 17561 11980 17595
rect 12014 17592 12026 17595
rect 12986 17592 12992 17604
rect 12014 17564 12992 17592
rect 12014 17561 12026 17564
rect 11968 17555 12026 17561
rect 12986 17552 12992 17564
rect 13044 17552 13050 17604
rect 3418 17524 3424 17536
rect 3379 17496 3424 17524
rect 3418 17484 3424 17496
rect 3476 17484 3482 17536
rect 5994 17484 6000 17536
rect 6052 17524 6058 17536
rect 7653 17527 7711 17533
rect 7653 17524 7665 17527
rect 6052 17496 7665 17524
rect 6052 17484 6058 17496
rect 7653 17493 7665 17496
rect 7699 17493 7711 17527
rect 7653 17487 7711 17493
rect 9861 17527 9919 17533
rect 9861 17493 9873 17527
rect 9907 17524 9919 17527
rect 10870 17524 10876 17536
rect 9907 17496 10876 17524
rect 9907 17493 9919 17496
rect 9861 17487 9919 17493
rect 10870 17484 10876 17496
rect 10928 17484 10934 17536
rect 13081 17527 13139 17533
rect 13081 17493 13093 17527
rect 13127 17524 13139 17527
rect 16022 17524 16028 17536
rect 13127 17496 16028 17524
rect 13127 17493 13139 17496
rect 13081 17487 13139 17493
rect 16022 17484 16028 17496
rect 16080 17484 16086 17536
rect 1104 17434 23987 17456
rect 1104 17382 6630 17434
rect 6682 17382 6694 17434
rect 6746 17382 6758 17434
rect 6810 17382 6822 17434
rect 6874 17382 6886 17434
rect 6938 17382 12311 17434
rect 12363 17382 12375 17434
rect 12427 17382 12439 17434
rect 12491 17382 12503 17434
rect 12555 17382 12567 17434
rect 12619 17382 17992 17434
rect 18044 17382 18056 17434
rect 18108 17382 18120 17434
rect 18172 17382 18184 17434
rect 18236 17382 18248 17434
rect 18300 17382 23673 17434
rect 23725 17382 23737 17434
rect 23789 17382 23801 17434
rect 23853 17382 23865 17434
rect 23917 17382 23929 17434
rect 23981 17382 23987 17434
rect 1104 17360 23987 17382
rect 11790 17280 11796 17332
rect 11848 17320 11854 17332
rect 13998 17320 14004 17332
rect 11848 17292 14004 17320
rect 11848 17280 11854 17292
rect 13998 17280 14004 17292
rect 14056 17280 14062 17332
rect 4614 17252 4620 17264
rect 3988 17224 4620 17252
rect 3234 17184 3240 17196
rect 3292 17193 3298 17196
rect 3988 17193 4016 17224
rect 4614 17212 4620 17224
rect 4672 17212 4678 17264
rect 4246 17193 4252 17196
rect 3204 17156 3240 17184
rect 3234 17144 3240 17156
rect 3292 17147 3304 17193
rect 3513 17187 3571 17193
rect 3513 17153 3525 17187
rect 3559 17184 3571 17187
rect 3973 17187 4031 17193
rect 3973 17184 3985 17187
rect 3559 17156 3985 17184
rect 3559 17153 3571 17156
rect 3513 17147 3571 17153
rect 3973 17153 3985 17156
rect 4019 17153 4031 17187
rect 3973 17147 4031 17153
rect 4240 17147 4252 17193
rect 4304 17184 4310 17196
rect 7009 17187 7067 17193
rect 4304 17156 4340 17184
rect 3292 17144 3298 17147
rect 4246 17144 4252 17147
rect 4304 17144 4310 17156
rect 7009 17153 7021 17187
rect 7055 17184 7067 17187
rect 7098 17184 7104 17196
rect 7055 17156 7104 17184
rect 7055 17153 7067 17156
rect 7009 17147 7067 17153
rect 7098 17144 7104 17156
rect 7156 17144 7162 17196
rect 7276 17187 7334 17193
rect 7276 17153 7288 17187
rect 7322 17184 7334 17187
rect 7742 17184 7748 17196
rect 7322 17156 7748 17184
rect 7322 17153 7334 17156
rect 7276 17147 7334 17153
rect 7742 17144 7748 17156
rect 7800 17144 7806 17196
rect 9306 17144 9312 17196
rect 9364 17184 9370 17196
rect 9769 17187 9827 17193
rect 9769 17184 9781 17187
rect 9364 17156 9781 17184
rect 9364 17144 9370 17156
rect 9769 17153 9781 17156
rect 9815 17153 9827 17187
rect 9769 17147 9827 17153
rect 10036 17187 10094 17193
rect 10036 17153 10048 17187
rect 10082 17184 10094 17187
rect 11790 17184 11796 17196
rect 10082 17156 11796 17184
rect 10082 17153 10094 17156
rect 10036 17147 10094 17153
rect 11790 17144 11796 17156
rect 11848 17144 11854 17196
rect 11149 17051 11207 17057
rect 11149 17017 11161 17051
rect 11195 17048 11207 17051
rect 13078 17048 13084 17060
rect 11195 17020 13084 17048
rect 11195 17017 11207 17020
rect 11149 17011 11207 17017
rect 13078 17008 13084 17020
rect 13136 17008 13142 17060
rect 2133 16983 2191 16989
rect 2133 16949 2145 16983
rect 2179 16980 2191 16983
rect 2222 16980 2228 16992
rect 2179 16952 2228 16980
rect 2179 16949 2191 16952
rect 2133 16943 2191 16949
rect 2222 16940 2228 16952
rect 2280 16940 2286 16992
rect 5350 16980 5356 16992
rect 5311 16952 5356 16980
rect 5350 16940 5356 16952
rect 5408 16940 5414 16992
rect 8389 16983 8447 16989
rect 8389 16949 8401 16983
rect 8435 16980 8447 16983
rect 8478 16980 8484 16992
rect 8435 16952 8484 16980
rect 8435 16949 8447 16952
rect 8389 16943 8447 16949
rect 8478 16940 8484 16952
rect 8536 16940 8542 16992
rect 11790 16980 11796 16992
rect 11751 16952 11796 16980
rect 11790 16940 11796 16952
rect 11848 16940 11854 16992
rect 1104 16890 23828 16912
rect 1104 16838 3790 16890
rect 3842 16838 3854 16890
rect 3906 16838 3918 16890
rect 3970 16838 3982 16890
rect 4034 16838 4046 16890
rect 4098 16838 9471 16890
rect 9523 16838 9535 16890
rect 9587 16838 9599 16890
rect 9651 16838 9663 16890
rect 9715 16838 9727 16890
rect 9779 16838 15152 16890
rect 15204 16838 15216 16890
rect 15268 16838 15280 16890
rect 15332 16838 15344 16890
rect 15396 16838 15408 16890
rect 15460 16838 20833 16890
rect 20885 16838 20897 16890
rect 20949 16838 20961 16890
rect 21013 16838 21025 16890
rect 21077 16838 21089 16890
rect 21141 16838 23828 16890
rect 1104 16816 23828 16838
rect 2498 16776 2504 16788
rect 2459 16748 2504 16776
rect 2498 16736 2504 16748
rect 2556 16736 2562 16788
rect 5534 16776 5540 16788
rect 2746 16748 5540 16776
rect 2222 16668 2228 16720
rect 2280 16708 2286 16720
rect 2746 16708 2774 16748
rect 5534 16736 5540 16748
rect 5592 16736 5598 16788
rect 2280 16680 2774 16708
rect 2280 16668 2286 16680
rect 4614 16640 4620 16652
rect 4575 16612 4620 16640
rect 4614 16600 4620 16612
rect 4672 16600 4678 16652
rect 8294 16600 8300 16652
rect 8352 16640 8358 16652
rect 9306 16640 9312 16652
rect 8352 16612 9312 16640
rect 8352 16600 8358 16612
rect 9306 16600 9312 16612
rect 9364 16640 9370 16652
rect 10045 16643 10103 16649
rect 10045 16640 10057 16643
rect 9364 16612 10057 16640
rect 9364 16600 9370 16612
rect 10045 16609 10057 16612
rect 10091 16609 10103 16643
rect 10045 16603 10103 16609
rect 2498 16532 2504 16584
rect 2556 16572 2562 16584
rect 2685 16575 2743 16581
rect 2685 16572 2697 16575
rect 2556 16544 2697 16572
rect 2556 16532 2562 16544
rect 2685 16541 2697 16544
rect 2731 16541 2743 16575
rect 2685 16535 2743 16541
rect 3050 16532 3056 16584
rect 3108 16572 3114 16584
rect 3421 16575 3479 16581
rect 3421 16572 3433 16575
rect 3108 16544 3433 16572
rect 3108 16532 3114 16544
rect 3421 16541 3433 16544
rect 3467 16572 3479 16575
rect 3510 16572 3516 16584
rect 3467 16544 3516 16572
rect 3467 16541 3479 16544
rect 3421 16535 3479 16541
rect 3510 16532 3516 16544
rect 3568 16532 3574 16584
rect 16301 16575 16359 16581
rect 16301 16541 16313 16575
rect 16347 16572 16359 16575
rect 16574 16572 16580 16584
rect 16347 16544 16580 16572
rect 16347 16541 16359 16544
rect 16301 16535 16359 16541
rect 16574 16532 16580 16544
rect 16632 16532 16638 16584
rect 3694 16464 3700 16516
rect 3752 16504 3758 16516
rect 4862 16507 4920 16513
rect 4862 16504 4874 16507
rect 3752 16476 4874 16504
rect 3752 16464 3758 16476
rect 4862 16473 4874 16476
rect 4908 16473 4920 16507
rect 7466 16504 7472 16516
rect 4862 16467 4920 16473
rect 6012 16476 7472 16504
rect 3237 16439 3295 16445
rect 3237 16405 3249 16439
rect 3283 16436 3295 16439
rect 4706 16436 4712 16448
rect 3283 16408 4712 16436
rect 3283 16405 3295 16408
rect 3237 16399 3295 16405
rect 4706 16396 4712 16408
rect 4764 16396 4770 16448
rect 6012 16445 6040 16476
rect 7466 16464 7472 16476
rect 7524 16464 7530 16516
rect 7926 16464 7932 16516
rect 7984 16504 7990 16516
rect 8030 16507 8088 16513
rect 8030 16504 8042 16507
rect 7984 16476 8042 16504
rect 7984 16464 7990 16476
rect 8030 16473 8042 16476
rect 8076 16473 8088 16507
rect 8030 16467 8088 16473
rect 10312 16507 10370 16513
rect 10312 16473 10324 16507
rect 10358 16504 10370 16507
rect 10358 16476 12434 16504
rect 10358 16473 10370 16476
rect 10312 16467 10370 16473
rect 5997 16439 6055 16445
rect 5997 16405 6009 16439
rect 6043 16405 6055 16439
rect 5997 16399 6055 16405
rect 6917 16439 6975 16445
rect 6917 16405 6929 16439
rect 6963 16436 6975 16439
rect 7834 16436 7840 16448
rect 6963 16408 7840 16436
rect 6963 16405 6975 16408
rect 6917 16399 6975 16405
rect 7834 16396 7840 16408
rect 7892 16396 7898 16448
rect 9217 16439 9275 16445
rect 9217 16405 9229 16439
rect 9263 16436 9275 16439
rect 9306 16436 9312 16448
rect 9263 16408 9312 16436
rect 9263 16405 9275 16408
rect 9217 16399 9275 16405
rect 9306 16396 9312 16408
rect 9364 16396 9370 16448
rect 11425 16439 11483 16445
rect 11425 16405 11437 16439
rect 11471 16436 11483 16439
rect 11974 16436 11980 16448
rect 11471 16408 11980 16436
rect 11471 16405 11483 16408
rect 11425 16399 11483 16405
rect 11974 16396 11980 16408
rect 12032 16396 12038 16448
rect 12406 16436 12434 16476
rect 16117 16439 16175 16445
rect 16117 16436 16129 16439
rect 12406 16408 16129 16436
rect 16117 16405 16129 16408
rect 16163 16405 16175 16439
rect 16117 16399 16175 16405
rect 1104 16346 23987 16368
rect 1104 16294 6630 16346
rect 6682 16294 6694 16346
rect 6746 16294 6758 16346
rect 6810 16294 6822 16346
rect 6874 16294 6886 16346
rect 6938 16294 12311 16346
rect 12363 16294 12375 16346
rect 12427 16294 12439 16346
rect 12491 16294 12503 16346
rect 12555 16294 12567 16346
rect 12619 16294 17992 16346
rect 18044 16294 18056 16346
rect 18108 16294 18120 16346
rect 18172 16294 18184 16346
rect 18236 16294 18248 16346
rect 18300 16294 23673 16346
rect 23725 16294 23737 16346
rect 23789 16294 23801 16346
rect 23853 16294 23865 16346
rect 23917 16294 23929 16346
rect 23981 16294 23987 16346
rect 1104 16272 23987 16294
rect 2041 16235 2099 16241
rect 2041 16201 2053 16235
rect 2087 16232 2099 16235
rect 2314 16232 2320 16244
rect 2087 16204 2320 16232
rect 2087 16201 2099 16204
rect 2041 16195 2099 16201
rect 2314 16192 2320 16204
rect 2372 16192 2378 16244
rect 3053 16235 3111 16241
rect 3053 16201 3065 16235
rect 3099 16232 3111 16235
rect 4614 16232 4620 16244
rect 3099 16204 4620 16232
rect 3099 16201 3111 16204
rect 3053 16195 3111 16201
rect 4614 16192 4620 16204
rect 4672 16192 4678 16244
rect 5902 16232 5908 16244
rect 5863 16204 5908 16232
rect 5902 16192 5908 16204
rect 5960 16192 5966 16244
rect 7006 16192 7012 16244
rect 7064 16192 7070 16244
rect 8294 16232 8300 16244
rect 8255 16204 8300 16232
rect 8294 16192 8300 16204
rect 8352 16192 8358 16244
rect 4341 16167 4399 16173
rect 4341 16133 4353 16167
rect 4387 16164 4399 16167
rect 7024 16164 7052 16192
rect 8938 16164 8944 16176
rect 4387 16136 8944 16164
rect 4387 16133 4399 16136
rect 4341 16127 4399 16133
rect 8938 16124 8944 16136
rect 8996 16164 9002 16176
rect 9585 16167 9643 16173
rect 9585 16164 9597 16167
rect 8996 16136 9597 16164
rect 8996 16124 9002 16136
rect 9585 16133 9597 16136
rect 9631 16133 9643 16167
rect 9585 16127 9643 16133
rect 1578 16056 1584 16108
rect 1636 16096 1642 16108
rect 1857 16099 1915 16105
rect 1857 16096 1869 16099
rect 1636 16068 1869 16096
rect 1636 16056 1642 16068
rect 1857 16065 1869 16068
rect 1903 16065 1915 16099
rect 1857 16059 1915 16065
rect 3694 16056 3700 16108
rect 3752 16096 3758 16108
rect 4985 16099 5043 16105
rect 4985 16096 4997 16099
rect 3752 16068 4997 16096
rect 3752 16056 3758 16068
rect 4985 16065 4997 16068
rect 5031 16065 5043 16099
rect 4985 16059 5043 16065
rect 5077 16099 5135 16105
rect 5077 16065 5089 16099
rect 5123 16065 5135 16099
rect 5077 16059 5135 16065
rect 1673 16031 1731 16037
rect 1673 15997 1685 16031
rect 1719 16028 1731 16031
rect 4154 16028 4160 16040
rect 1719 16000 4160 16028
rect 1719 15997 1731 16000
rect 1673 15991 1731 15997
rect 4154 15988 4160 16000
rect 4212 15988 4218 16040
rect 2958 15920 2964 15972
rect 3016 15960 3022 15972
rect 5092 15960 5120 16059
rect 5166 16056 5172 16108
rect 5224 16096 5230 16108
rect 5353 16099 5411 16105
rect 5224 16068 5269 16096
rect 5224 16056 5230 16068
rect 5353 16065 5365 16099
rect 5399 16096 5411 16099
rect 5718 16096 5724 16108
rect 5399 16068 5724 16096
rect 5399 16065 5411 16068
rect 5353 16059 5411 16065
rect 5718 16056 5724 16068
rect 5776 16056 5782 16108
rect 5813 16099 5871 16105
rect 5813 16065 5825 16099
rect 5859 16065 5871 16099
rect 5994 16096 6000 16108
rect 5955 16068 6000 16096
rect 5813 16059 5871 16065
rect 5828 15972 5856 16059
rect 5994 16056 6000 16068
rect 6052 16056 6058 16108
rect 7009 16099 7067 16105
rect 7009 16065 7021 16099
rect 7055 16065 7067 16099
rect 7009 16059 7067 16065
rect 7024 16028 7052 16059
rect 7098 16056 7104 16108
rect 7156 16096 7162 16108
rect 7374 16096 7380 16108
rect 7156 16068 7201 16096
rect 7287 16068 7380 16096
rect 7156 16056 7162 16068
rect 7374 16056 7380 16068
rect 7432 16096 7438 16108
rect 8110 16096 8116 16108
rect 7432 16068 8116 16096
rect 7432 16056 7438 16068
rect 8110 16056 8116 16068
rect 8168 16056 8174 16108
rect 12161 16099 12219 16105
rect 12161 16065 12173 16099
rect 12207 16096 12219 16099
rect 12802 16096 12808 16108
rect 12207 16068 12808 16096
rect 12207 16065 12219 16068
rect 12161 16059 12219 16065
rect 12802 16056 12808 16068
rect 12860 16056 12866 16108
rect 7190 16028 7196 16040
rect 7024 16000 7196 16028
rect 7190 15988 7196 16000
rect 7248 15988 7254 16040
rect 7285 16031 7343 16037
rect 7285 15997 7297 16031
rect 7331 16028 7343 16031
rect 11054 16028 11060 16040
rect 7331 16000 11060 16028
rect 7331 15997 7343 16000
rect 7285 15991 7343 15997
rect 11054 15988 11060 16000
rect 11112 15988 11118 16040
rect 5810 15960 5816 15972
rect 3016 15932 5120 15960
rect 5723 15932 5816 15960
rect 3016 15920 3022 15932
rect 5810 15920 5816 15932
rect 5868 15960 5874 15972
rect 7558 15960 7564 15972
rect 5868 15932 7564 15960
rect 5868 15920 5874 15932
rect 7558 15920 7564 15932
rect 7616 15920 7622 15972
rect 4798 15892 4804 15904
rect 4759 15864 4804 15892
rect 4798 15852 4804 15864
rect 4856 15852 4862 15904
rect 6546 15852 6552 15904
rect 6604 15892 6610 15904
rect 6825 15895 6883 15901
rect 6825 15892 6837 15895
rect 6604 15864 6837 15892
rect 6604 15852 6610 15864
rect 6825 15861 6837 15864
rect 6871 15861 6883 15895
rect 6825 15855 6883 15861
rect 9306 15852 9312 15904
rect 9364 15892 9370 15904
rect 10229 15895 10287 15901
rect 10229 15892 10241 15895
rect 9364 15864 10241 15892
rect 9364 15852 9370 15864
rect 10229 15861 10241 15864
rect 10275 15892 10287 15895
rect 11054 15892 11060 15904
rect 10275 15864 11060 15892
rect 10275 15861 10287 15864
rect 10229 15855 10287 15861
rect 11054 15852 11060 15864
rect 11112 15852 11118 15904
rect 11790 15852 11796 15904
rect 11848 15892 11854 15904
rect 12069 15895 12127 15901
rect 12069 15892 12081 15895
rect 11848 15864 12081 15892
rect 11848 15852 11854 15864
rect 12069 15861 12081 15864
rect 12115 15892 12127 15895
rect 14182 15892 14188 15904
rect 12115 15864 14188 15892
rect 12115 15861 12127 15864
rect 12069 15855 12127 15861
rect 14182 15852 14188 15864
rect 14240 15852 14246 15904
rect 1104 15802 23828 15824
rect 1104 15750 3790 15802
rect 3842 15750 3854 15802
rect 3906 15750 3918 15802
rect 3970 15750 3982 15802
rect 4034 15750 4046 15802
rect 4098 15750 9471 15802
rect 9523 15750 9535 15802
rect 9587 15750 9599 15802
rect 9651 15750 9663 15802
rect 9715 15750 9727 15802
rect 9779 15750 15152 15802
rect 15204 15750 15216 15802
rect 15268 15750 15280 15802
rect 15332 15750 15344 15802
rect 15396 15750 15408 15802
rect 15460 15750 20833 15802
rect 20885 15750 20897 15802
rect 20949 15750 20961 15802
rect 21013 15750 21025 15802
rect 21077 15750 21089 15802
rect 21141 15750 23828 15802
rect 1104 15728 23828 15750
rect 1578 15688 1584 15700
rect 1539 15660 1584 15688
rect 1578 15648 1584 15660
rect 1636 15648 1642 15700
rect 2498 15688 2504 15700
rect 2459 15660 2504 15688
rect 2498 15648 2504 15660
rect 2556 15648 2562 15700
rect 4706 15648 4712 15700
rect 4764 15688 4770 15700
rect 7098 15688 7104 15700
rect 4764 15660 7104 15688
rect 4764 15648 4770 15660
rect 7098 15648 7104 15660
rect 7156 15648 7162 15700
rect 8386 15688 8392 15700
rect 8347 15660 8392 15688
rect 8386 15648 8392 15660
rect 8444 15648 8450 15700
rect 12802 15688 12808 15700
rect 12763 15660 12808 15688
rect 12802 15648 12808 15660
rect 12860 15648 12866 15700
rect 16574 15688 16580 15700
rect 16535 15660 16580 15688
rect 16574 15648 16580 15660
rect 16632 15648 16638 15700
rect 5442 15580 5448 15632
rect 5500 15620 5506 15632
rect 7374 15620 7380 15632
rect 5500 15592 7380 15620
rect 5500 15580 5506 15592
rect 7374 15580 7380 15592
rect 7432 15580 7438 15632
rect 11256 15592 12204 15620
rect 1946 15552 1952 15564
rect 1780 15524 1952 15552
rect 1780 15493 1808 15524
rect 1946 15512 1952 15524
rect 2004 15512 2010 15564
rect 3145 15555 3203 15561
rect 3145 15521 3157 15555
rect 3191 15552 3203 15555
rect 3418 15552 3424 15564
rect 3191 15524 3424 15552
rect 3191 15521 3203 15524
rect 3145 15515 3203 15521
rect 3418 15512 3424 15524
rect 3476 15512 3482 15564
rect 7190 15552 7196 15564
rect 7151 15524 7196 15552
rect 7190 15512 7196 15524
rect 7248 15512 7254 15564
rect 7837 15555 7895 15561
rect 7837 15521 7849 15555
rect 7883 15552 7895 15555
rect 8018 15552 8024 15564
rect 7883 15524 8024 15552
rect 7883 15521 7895 15524
rect 7837 15515 7895 15521
rect 8018 15512 8024 15524
rect 8076 15552 8082 15564
rect 9214 15552 9220 15564
rect 8076 15524 9220 15552
rect 8076 15512 8082 15524
rect 9214 15512 9220 15524
rect 9272 15512 9278 15564
rect 11146 15552 11152 15564
rect 11107 15524 11152 15552
rect 11146 15512 11152 15524
rect 11204 15512 11210 15564
rect 1765 15487 1823 15493
rect 1765 15453 1777 15487
rect 1811 15453 1823 15487
rect 1765 15447 1823 15453
rect 1854 15444 1860 15496
rect 1912 15484 1918 15496
rect 2041 15487 2099 15493
rect 2041 15484 2053 15487
rect 1912 15456 2053 15484
rect 1912 15444 1918 15456
rect 2041 15453 2053 15456
rect 2087 15453 2099 15487
rect 2041 15447 2099 15453
rect 3050 15444 3056 15496
rect 3108 15484 3114 15496
rect 4522 15484 4528 15496
rect 3108 15456 4528 15484
rect 3108 15444 3114 15456
rect 4522 15444 4528 15456
rect 4580 15444 4586 15496
rect 4614 15444 4620 15496
rect 4672 15484 4678 15496
rect 5353 15487 5411 15493
rect 5353 15484 5365 15487
rect 4672 15456 5365 15484
rect 4672 15444 4678 15456
rect 5353 15453 5365 15456
rect 5399 15453 5411 15487
rect 5353 15447 5411 15453
rect 5813 15487 5871 15493
rect 5813 15453 5825 15487
rect 5859 15453 5871 15487
rect 5813 15447 5871 15453
rect 5997 15487 6055 15493
rect 5997 15453 6009 15487
rect 6043 15484 6055 15487
rect 6270 15484 6276 15496
rect 6043 15456 6276 15484
rect 6043 15453 6055 15456
rect 5997 15447 6055 15453
rect 2961 15419 3019 15425
rect 2961 15385 2973 15419
rect 3007 15416 3019 15419
rect 4154 15416 4160 15428
rect 3007 15388 4160 15416
rect 3007 15385 3019 15388
rect 2961 15379 3019 15385
rect 4154 15376 4160 15388
rect 4212 15376 4218 15428
rect 4798 15376 4804 15428
rect 4856 15416 4862 15428
rect 5086 15419 5144 15425
rect 5086 15416 5098 15419
rect 4856 15388 5098 15416
rect 4856 15376 4862 15388
rect 5086 15385 5098 15388
rect 5132 15385 5144 15419
rect 5086 15379 5144 15385
rect 5258 15376 5264 15428
rect 5316 15416 5322 15428
rect 5828 15416 5856 15447
rect 6270 15444 6276 15456
rect 6328 15444 6334 15496
rect 6733 15487 6791 15493
rect 6733 15453 6745 15487
rect 6779 15453 6791 15487
rect 6733 15447 6791 15453
rect 7009 15487 7067 15493
rect 7009 15453 7021 15487
rect 7055 15484 7067 15487
rect 7558 15484 7564 15496
rect 7055 15456 7564 15484
rect 7055 15453 7067 15456
rect 7009 15447 7067 15453
rect 5316 15388 5856 15416
rect 6748 15416 6776 15447
rect 7558 15444 7564 15456
rect 7616 15444 7622 15496
rect 9122 15484 9128 15496
rect 9083 15456 9128 15484
rect 9122 15444 9128 15456
rect 9180 15444 9186 15496
rect 9309 15487 9367 15493
rect 9309 15453 9321 15487
rect 9355 15484 9367 15487
rect 9398 15484 9404 15496
rect 9355 15456 9404 15484
rect 9355 15453 9367 15456
rect 9309 15447 9367 15453
rect 9398 15444 9404 15456
rect 9456 15444 9462 15496
rect 11054 15444 11060 15496
rect 11112 15484 11118 15496
rect 11256 15484 11284 15592
rect 11422 15512 11428 15564
rect 11480 15552 11486 15564
rect 12176 15561 12204 15592
rect 12069 15555 12127 15561
rect 12069 15552 12081 15555
rect 11480 15524 12081 15552
rect 11480 15512 11486 15524
rect 12069 15521 12081 15524
rect 12115 15521 12127 15555
rect 12069 15515 12127 15521
rect 12161 15555 12219 15561
rect 12161 15521 12173 15555
rect 12207 15521 12219 15555
rect 12161 15515 12219 15521
rect 12250 15512 12256 15564
rect 12308 15552 12314 15564
rect 12308 15524 13400 15552
rect 12308 15512 12314 15524
rect 11974 15484 11980 15496
rect 11112 15456 11284 15484
rect 11935 15456 11980 15484
rect 11112 15444 11118 15456
rect 11974 15444 11980 15456
rect 12032 15444 12038 15496
rect 12802 15444 12808 15496
rect 12860 15484 12866 15496
rect 12989 15487 13047 15493
rect 12989 15484 13001 15487
rect 12860 15456 13001 15484
rect 12860 15444 12866 15456
rect 12989 15453 13001 15456
rect 13035 15453 13047 15487
rect 12989 15447 13047 15453
rect 13078 15444 13084 15496
rect 13136 15484 13142 15496
rect 13262 15484 13268 15496
rect 13136 15456 13181 15484
rect 13223 15456 13268 15484
rect 13136 15444 13142 15456
rect 13262 15444 13268 15456
rect 13320 15444 13326 15496
rect 13372 15493 13400 15524
rect 13630 15512 13636 15564
rect 13688 15552 13694 15564
rect 14182 15552 14188 15564
rect 13688 15524 14188 15552
rect 13688 15512 13694 15524
rect 14182 15512 14188 15524
rect 14240 15552 14246 15564
rect 14645 15555 14703 15561
rect 14645 15552 14657 15555
rect 14240 15524 14657 15552
rect 14240 15512 14246 15524
rect 14645 15521 14657 15524
rect 14691 15552 14703 15555
rect 16117 15555 16175 15561
rect 16117 15552 16129 15555
rect 14691 15524 16129 15552
rect 14691 15521 14703 15524
rect 14645 15515 14703 15521
rect 16117 15521 16129 15524
rect 16163 15552 16175 15555
rect 17221 15555 17279 15561
rect 17221 15552 17233 15555
rect 16163 15524 17233 15552
rect 16163 15521 16175 15524
rect 16117 15515 16175 15521
rect 17221 15521 17233 15524
rect 17267 15552 17279 15555
rect 17267 15524 18092 15552
rect 17267 15521 17279 15524
rect 17221 15515 17279 15521
rect 13357 15487 13415 15493
rect 13357 15453 13369 15487
rect 13403 15453 13415 15487
rect 13357 15447 13415 15453
rect 13906 15444 13912 15496
rect 13964 15484 13970 15496
rect 14461 15487 14519 15493
rect 14461 15484 14473 15487
rect 13964 15456 14473 15484
rect 13964 15444 13970 15456
rect 14461 15453 14473 15456
rect 14507 15453 14519 15487
rect 14461 15447 14519 15453
rect 14550 15444 14556 15496
rect 14608 15484 14614 15496
rect 14737 15487 14795 15493
rect 14608 15456 14653 15484
rect 14608 15444 14614 15456
rect 14737 15453 14749 15487
rect 14783 15484 14795 15487
rect 15286 15484 15292 15496
rect 14783 15456 15292 15484
rect 14783 15453 14795 15456
rect 14737 15447 14795 15453
rect 15286 15444 15292 15456
rect 15344 15444 15350 15496
rect 7466 15416 7472 15428
rect 6748 15388 7472 15416
rect 5316 15376 5322 15388
rect 7466 15376 7472 15388
rect 7524 15376 7530 15428
rect 7929 15419 7987 15425
rect 7929 15385 7941 15419
rect 7975 15416 7987 15419
rect 8294 15416 8300 15428
rect 7975 15388 8300 15416
rect 7975 15385 7987 15388
rect 7929 15379 7987 15385
rect 8294 15376 8300 15388
rect 8352 15376 8358 15428
rect 9217 15419 9275 15425
rect 9217 15385 9229 15419
rect 9263 15416 9275 15419
rect 9858 15416 9864 15428
rect 9263 15388 9864 15416
rect 9263 15385 9275 15388
rect 9217 15379 9275 15385
rect 9858 15376 9864 15388
rect 9916 15376 9922 15428
rect 18064 15425 18092 15524
rect 10904 15419 10962 15425
rect 10904 15385 10916 15419
rect 10950 15416 10962 15419
rect 18049 15419 18107 15425
rect 10950 15388 14320 15416
rect 10950 15385 10962 15388
rect 10904 15379 10962 15385
rect 1949 15351 2007 15357
rect 1949 15317 1961 15351
rect 1995 15348 2007 15351
rect 2498 15348 2504 15360
rect 1995 15320 2504 15348
rect 1995 15317 2007 15320
rect 1949 15311 2007 15317
rect 2498 15308 2504 15320
rect 2556 15308 2562 15360
rect 2866 15348 2872 15360
rect 2827 15320 2872 15348
rect 2866 15308 2872 15320
rect 2924 15308 2930 15360
rect 3970 15348 3976 15360
rect 3931 15320 3976 15348
rect 3970 15308 3976 15320
rect 4028 15308 4034 15360
rect 4982 15308 4988 15360
rect 5040 15348 5046 15360
rect 5442 15348 5448 15360
rect 5040 15320 5448 15348
rect 5040 15308 5046 15320
rect 5442 15308 5448 15320
rect 5500 15308 5506 15360
rect 5902 15348 5908 15360
rect 5863 15320 5908 15348
rect 5902 15308 5908 15320
rect 5960 15308 5966 15360
rect 8018 15308 8024 15360
rect 8076 15348 8082 15360
rect 9769 15351 9827 15357
rect 8076 15320 8121 15348
rect 8076 15308 8082 15320
rect 9769 15317 9781 15351
rect 9815 15348 9827 15351
rect 10686 15348 10692 15360
rect 9815 15320 10692 15348
rect 9815 15317 9827 15320
rect 9769 15311 9827 15317
rect 10686 15308 10692 15320
rect 10744 15308 10750 15360
rect 11146 15308 11152 15360
rect 11204 15348 11210 15360
rect 14292 15357 14320 15388
rect 18049 15385 18061 15419
rect 18095 15416 18107 15419
rect 19058 15416 19064 15428
rect 18095 15388 19064 15416
rect 18095 15385 18107 15388
rect 18049 15379 18107 15385
rect 19058 15376 19064 15388
rect 19116 15376 19122 15428
rect 11609 15351 11667 15357
rect 11609 15348 11621 15351
rect 11204 15320 11621 15348
rect 11204 15308 11210 15320
rect 11609 15317 11621 15320
rect 11655 15317 11667 15351
rect 11609 15311 11667 15317
rect 14277 15351 14335 15357
rect 14277 15317 14289 15351
rect 14323 15317 14335 15351
rect 16942 15348 16948 15360
rect 16903 15320 16948 15348
rect 14277 15311 14335 15317
rect 16942 15308 16948 15320
rect 17000 15308 17006 15360
rect 17034 15308 17040 15360
rect 17092 15348 17098 15360
rect 17092 15320 17137 15348
rect 17092 15308 17098 15320
rect 18690 15308 18696 15360
rect 18748 15348 18754 15360
rect 19429 15351 19487 15357
rect 19429 15348 19441 15351
rect 18748 15320 19441 15348
rect 18748 15308 18754 15320
rect 19429 15317 19441 15320
rect 19475 15317 19487 15351
rect 19429 15311 19487 15317
rect 1104 15258 23987 15280
rect 1104 15206 6630 15258
rect 6682 15206 6694 15258
rect 6746 15206 6758 15258
rect 6810 15206 6822 15258
rect 6874 15206 6886 15258
rect 6938 15206 12311 15258
rect 12363 15206 12375 15258
rect 12427 15206 12439 15258
rect 12491 15206 12503 15258
rect 12555 15206 12567 15258
rect 12619 15206 17992 15258
rect 18044 15206 18056 15258
rect 18108 15206 18120 15258
rect 18172 15206 18184 15258
rect 18236 15206 18248 15258
rect 18300 15206 23673 15258
rect 23725 15206 23737 15258
rect 23789 15206 23801 15258
rect 23853 15206 23865 15258
rect 23917 15206 23929 15258
rect 23981 15206 23987 15258
rect 1104 15184 23987 15206
rect 2041 15147 2099 15153
rect 2041 15113 2053 15147
rect 2087 15144 2099 15147
rect 3881 15147 3939 15153
rect 2087 15116 3832 15144
rect 2087 15113 2099 15116
rect 2041 15107 2099 15113
rect 2498 15076 2504 15088
rect 2459 15048 2504 15076
rect 2498 15036 2504 15048
rect 2556 15036 2562 15088
rect 3804 15076 3832 15116
rect 3881 15113 3893 15147
rect 3927 15144 3939 15147
rect 4246 15144 4252 15156
rect 3927 15116 4252 15144
rect 3927 15113 3939 15116
rect 3881 15107 3939 15113
rect 4246 15104 4252 15116
rect 4304 15104 4310 15156
rect 4338 15104 4344 15156
rect 4396 15144 4402 15156
rect 4396 15116 4441 15144
rect 4396 15104 4402 15116
rect 4522 15104 4528 15156
rect 4580 15144 4586 15156
rect 4580 15116 5396 15144
rect 4580 15104 4586 15116
rect 5166 15076 5172 15088
rect 2731 15045 2789 15051
rect 3804 15048 5172 15076
rect 1765 15011 1823 15017
rect 1765 14977 1777 15011
rect 1811 15008 1823 15011
rect 1854 15008 1860 15020
rect 1811 14980 1860 15008
rect 1811 14977 1823 14980
rect 1765 14971 1823 14977
rect 1854 14968 1860 14980
rect 1912 15008 1918 15020
rect 2590 15008 2596 15020
rect 1912 14980 2596 15008
rect 1912 14968 1918 14980
rect 2590 14968 2596 14980
rect 2648 15008 2654 15020
rect 2731 15011 2743 15045
rect 2777 15011 2789 15045
rect 5166 15036 5172 15048
rect 5224 15036 5230 15088
rect 5368 15085 5396 15116
rect 5534 15104 5540 15156
rect 5592 15104 5598 15156
rect 7742 15104 7748 15156
rect 7800 15144 7806 15156
rect 7929 15147 7987 15153
rect 7929 15144 7941 15147
rect 7800 15116 7941 15144
rect 7800 15104 7806 15116
rect 7929 15113 7941 15116
rect 7975 15113 7987 15147
rect 7929 15107 7987 15113
rect 10965 15147 11023 15153
rect 10965 15113 10977 15147
rect 11011 15144 11023 15147
rect 11606 15144 11612 15156
rect 11011 15116 11612 15144
rect 11011 15113 11023 15116
rect 10965 15107 11023 15113
rect 11606 15104 11612 15116
rect 11664 15104 11670 15156
rect 12713 15147 12771 15153
rect 12713 15113 12725 15147
rect 12759 15144 12771 15147
rect 13262 15144 13268 15156
rect 12759 15116 13268 15144
rect 12759 15113 12771 15116
rect 12713 15107 12771 15113
rect 13262 15104 13268 15116
rect 13320 15104 13326 15156
rect 14550 15144 14556 15156
rect 14511 15116 14556 15144
rect 14550 15104 14556 15116
rect 14608 15104 14614 15156
rect 15286 15144 15292 15156
rect 15247 15116 15292 15144
rect 15286 15104 15292 15116
rect 15344 15104 15350 15156
rect 19242 15144 19248 15156
rect 17604 15116 19248 15144
rect 5353 15079 5411 15085
rect 5353 15045 5365 15079
rect 5399 15045 5411 15079
rect 5353 15039 5411 15045
rect 2731 15008 2789 15011
rect 2648 15005 2789 15008
rect 2648 14980 2774 15005
rect 2648 14968 2654 14980
rect 3142 14968 3148 15020
rect 3200 15008 3206 15020
rect 3329 15011 3387 15017
rect 3329 15008 3341 15011
rect 3200 14980 3341 15008
rect 3200 14968 3206 14980
rect 3329 14977 3341 14980
rect 3375 14977 3387 15011
rect 3510 15008 3516 15020
rect 3471 14980 3516 15008
rect 3329 14971 3387 14977
rect 3510 14968 3516 14980
rect 3568 14968 3574 15020
rect 3605 15011 3663 15017
rect 3605 14977 3617 15011
rect 3651 14977 3663 15011
rect 3605 14971 3663 14977
rect 2038 14940 2044 14952
rect 1999 14912 2044 14940
rect 2038 14900 2044 14912
rect 2096 14900 2102 14952
rect 2682 14900 2688 14952
rect 2740 14940 2746 14952
rect 3620 14940 3648 14971
rect 3694 14968 3700 15020
rect 3752 15008 3758 15020
rect 4522 15008 4528 15020
rect 3752 14980 4528 15008
rect 3752 14968 3758 14980
rect 4522 14968 4528 14980
rect 4580 14968 4586 15020
rect 4614 14968 4620 15020
rect 4672 15008 4678 15020
rect 4798 15017 4804 15020
rect 4755 15011 4804 15017
rect 4672 14980 4717 15008
rect 4672 14968 4678 14980
rect 4755 14977 4767 15011
rect 4801 14977 4804 15011
rect 4755 14971 4804 14977
rect 4798 14968 4804 14971
rect 4856 14968 4862 15020
rect 4893 15011 4951 15017
rect 4893 14977 4905 15011
rect 4939 15008 4951 15011
rect 5442 15008 5448 15020
rect 4939 14980 5448 15008
rect 4939 14977 4951 14980
rect 4893 14971 4951 14977
rect 5442 14968 5448 14980
rect 5500 14968 5506 15020
rect 5552 15017 5580 15104
rect 6638 15076 6644 15088
rect 6599 15048 6644 15076
rect 6638 15036 6644 15048
rect 6696 15036 6702 15088
rect 8294 15076 8300 15088
rect 8255 15048 8300 15076
rect 8294 15036 8300 15048
rect 8352 15036 8358 15088
rect 10778 15076 10784 15088
rect 10739 15048 10784 15076
rect 10778 15036 10784 15048
rect 10836 15036 10842 15088
rect 13078 15076 13084 15088
rect 12636 15048 13084 15076
rect 5537 15011 5595 15017
rect 5537 14977 5549 15011
rect 5583 14977 5595 15011
rect 5537 14971 5595 14977
rect 5629 15011 5687 15017
rect 5629 14977 5641 15011
rect 5675 14977 5687 15011
rect 5629 14971 5687 14977
rect 2740 14912 3648 14940
rect 2740 14900 2746 14912
rect 3970 14900 3976 14952
rect 4028 14940 4034 14952
rect 5644 14940 5672 14971
rect 8018 14968 8024 15020
rect 8076 15008 8082 15020
rect 8113 15011 8171 15017
rect 8113 15008 8125 15011
rect 8076 14980 8125 15008
rect 8076 14968 8082 14980
rect 8113 14977 8125 14980
rect 8159 14977 8171 15011
rect 8113 14971 8171 14977
rect 8205 15011 8263 15017
rect 8205 14977 8217 15011
rect 8251 15008 8263 15011
rect 8386 15008 8392 15020
rect 8251 14980 8392 15008
rect 8251 14977 8263 14980
rect 8205 14971 8263 14977
rect 8386 14968 8392 14980
rect 8444 14968 8450 15020
rect 8478 14968 8484 15020
rect 8536 15008 8542 15020
rect 9306 15008 9312 15020
rect 8536 14980 9312 15008
rect 8536 14968 8542 14980
rect 9306 14968 9312 14980
rect 9364 15008 9370 15020
rect 9493 15011 9551 15017
rect 9493 15008 9505 15011
rect 9364 14980 9505 15008
rect 9364 14968 9370 14980
rect 9493 14977 9505 14980
rect 9539 14977 9551 15011
rect 9493 14971 9551 14977
rect 11514 14968 11520 15020
rect 11572 15008 11578 15020
rect 12636 15017 12664 15048
rect 13078 15036 13084 15048
rect 13136 15036 13142 15088
rect 13725 15079 13783 15085
rect 13725 15045 13737 15079
rect 13771 15076 13783 15079
rect 14090 15076 14096 15088
rect 13771 15048 14096 15076
rect 13771 15045 13783 15048
rect 13725 15039 13783 15045
rect 14090 15036 14096 15048
rect 14148 15076 14154 15088
rect 15470 15076 15476 15088
rect 14148 15048 14688 15076
rect 15431 15048 15476 15076
rect 14148 15036 14154 15048
rect 11701 15011 11759 15017
rect 11701 15008 11713 15011
rect 11572 14980 11713 15008
rect 11572 14968 11578 14980
rect 11701 14977 11713 14980
rect 11747 14977 11759 15011
rect 11701 14971 11759 14977
rect 12621 15011 12679 15017
rect 12621 14977 12633 15011
rect 12667 14977 12679 15011
rect 12802 15008 12808 15020
rect 12763 14980 12808 15008
rect 12621 14971 12679 14977
rect 12802 14968 12808 14980
rect 12860 14968 12866 15020
rect 13628 15001 13686 15007
rect 13628 14967 13640 15001
rect 13674 14967 13686 15001
rect 13814 14968 13820 15020
rect 13872 15008 13878 15020
rect 14001 15011 14059 15017
rect 13872 14980 13917 15008
rect 13872 14968 13878 14980
rect 14001 14977 14013 15011
rect 14047 14977 14059 15011
rect 14001 14971 14059 14977
rect 13628 14961 13686 14967
rect 11054 14940 11060 14952
rect 4028 14912 5672 14940
rect 11015 14912 11060 14940
rect 4028 14900 4034 14912
rect 11054 14900 11060 14912
rect 11112 14900 11118 14952
rect 2498 14832 2504 14884
rect 2556 14872 2562 14884
rect 3142 14872 3148 14884
rect 2556 14844 3148 14872
rect 2556 14832 2562 14844
rect 3142 14832 3148 14844
rect 3200 14832 3206 14884
rect 3326 14832 3332 14884
rect 3384 14872 3390 14884
rect 3988 14872 4016 14900
rect 8846 14872 8852 14884
rect 3384 14844 4016 14872
rect 7024 14844 8852 14872
rect 3384 14832 3390 14844
rect 7024 14816 7052 14844
rect 8846 14832 8852 14844
rect 8904 14872 8910 14884
rect 9398 14872 9404 14884
rect 8904 14844 9404 14872
rect 8904 14832 8910 14844
rect 9398 14832 9404 14844
rect 9456 14832 9462 14884
rect 11238 14832 11244 14884
rect 11296 14872 11302 14884
rect 11422 14872 11428 14884
rect 11296 14844 11428 14872
rect 11296 14832 11302 14844
rect 11422 14832 11428 14844
rect 11480 14832 11486 14884
rect 13648 14872 13676 14961
rect 14016 14940 14044 14971
rect 14274 14968 14280 15020
rect 14332 15008 14338 15020
rect 14660 15017 14688 15048
rect 15470 15036 15476 15048
rect 15528 15036 15534 15088
rect 16758 15036 16764 15088
rect 16816 15076 16822 15088
rect 17604 15085 17632 15116
rect 19242 15104 19248 15116
rect 19300 15144 19306 15156
rect 19429 15147 19487 15153
rect 19429 15144 19441 15147
rect 19300 15116 19441 15144
rect 19300 15104 19306 15116
rect 19429 15113 19441 15116
rect 19475 15113 19487 15147
rect 19429 15107 19487 15113
rect 17037 15079 17095 15085
rect 17037 15076 17049 15079
rect 16816 15048 17049 15076
rect 16816 15036 16822 15048
rect 17037 15045 17049 15048
rect 17083 15076 17095 15079
rect 17589 15079 17647 15085
rect 17589 15076 17601 15079
rect 17083 15048 17601 15076
rect 17083 15045 17095 15048
rect 17037 15039 17095 15045
rect 17589 15045 17601 15048
rect 17635 15045 17647 15079
rect 17589 15039 17647 15045
rect 18524 15048 19380 15076
rect 14461 15011 14519 15017
rect 14461 15008 14473 15011
rect 14332 14980 14473 15008
rect 14332 14968 14338 14980
rect 14461 14977 14473 14980
rect 14507 14977 14519 15011
rect 14461 14971 14519 14977
rect 14645 15011 14703 15017
rect 14645 14977 14657 15011
rect 14691 15008 14703 15011
rect 16206 15008 16212 15020
rect 14691 14980 16212 15008
rect 14691 14977 14703 14980
rect 14645 14971 14703 14977
rect 16206 14968 16212 14980
rect 16264 14968 16270 15020
rect 16574 14968 16580 15020
rect 16632 15008 16638 15020
rect 16853 15011 16911 15017
rect 16853 15008 16865 15011
rect 16632 14980 16865 15008
rect 16632 14968 16638 14980
rect 16853 14977 16865 14980
rect 16899 14977 16911 15011
rect 16853 14971 16911 14977
rect 17126 14968 17132 15020
rect 17184 15008 17190 15020
rect 18524 15017 18552 15048
rect 18509 15011 18567 15017
rect 17184 14980 17229 15008
rect 17184 14968 17190 14980
rect 18509 14977 18521 15011
rect 18555 14977 18567 15011
rect 18690 15008 18696 15020
rect 18651 14980 18696 15008
rect 18509 14971 18567 14977
rect 18690 14968 18696 14980
rect 18748 14968 18754 15020
rect 19352 15017 19380 15048
rect 18785 15011 18843 15017
rect 18785 14977 18797 15011
rect 18831 14977 18843 15011
rect 18785 14971 18843 14977
rect 19337 15011 19395 15017
rect 19337 14977 19349 15011
rect 19383 15008 19395 15011
rect 19610 15008 19616 15020
rect 19383 14980 19616 15008
rect 19383 14977 19395 14980
rect 19337 14971 19395 14977
rect 18598 14940 18604 14952
rect 14016 14912 18604 14940
rect 18598 14900 18604 14912
rect 18656 14900 18662 14952
rect 14182 14872 14188 14884
rect 13648 14844 14188 14872
rect 14182 14832 14188 14844
rect 14240 14832 14246 14884
rect 14550 14832 14556 14884
rect 14608 14872 14614 14884
rect 15838 14872 15844 14884
rect 14608 14844 15608 14872
rect 15799 14844 15844 14872
rect 14608 14832 14614 14844
rect 1854 14804 1860 14816
rect 1815 14776 1860 14804
rect 1854 14764 1860 14776
rect 1912 14764 1918 14816
rect 1946 14764 1952 14816
rect 2004 14804 2010 14816
rect 2685 14807 2743 14813
rect 2685 14804 2697 14807
rect 2004 14776 2697 14804
rect 2004 14764 2010 14776
rect 2685 14773 2697 14776
rect 2731 14773 2743 14807
rect 2866 14804 2872 14816
rect 2827 14776 2872 14804
rect 2685 14767 2743 14773
rect 2866 14764 2872 14776
rect 2924 14764 2930 14816
rect 3694 14764 3700 14816
rect 3752 14804 3758 14816
rect 5350 14804 5356 14816
rect 3752 14776 5356 14804
rect 3752 14764 3758 14776
rect 5350 14764 5356 14776
rect 5408 14764 5414 14816
rect 5813 14807 5871 14813
rect 5813 14773 5825 14807
rect 5859 14804 5871 14807
rect 6454 14804 6460 14816
rect 5859 14776 6460 14804
rect 5859 14773 5871 14776
rect 5813 14767 5871 14773
rect 6454 14764 6460 14776
rect 6512 14764 6518 14816
rect 6917 14807 6975 14813
rect 6917 14773 6929 14807
rect 6963 14804 6975 14807
rect 7006 14804 7012 14816
rect 6963 14776 7012 14804
rect 6963 14773 6975 14776
rect 6917 14767 6975 14773
rect 7006 14764 7012 14776
rect 7064 14764 7070 14816
rect 8938 14764 8944 14816
rect 8996 14804 9002 14816
rect 9033 14807 9091 14813
rect 9033 14804 9045 14807
rect 8996 14776 9045 14804
rect 8996 14764 9002 14776
rect 9033 14773 9045 14776
rect 9079 14773 9091 14807
rect 9214 14804 9220 14816
rect 9175 14776 9220 14804
rect 9033 14767 9091 14773
rect 9214 14764 9220 14776
rect 9272 14764 9278 14816
rect 10502 14804 10508 14816
rect 10463 14776 10508 14804
rect 10502 14764 10508 14776
rect 10560 14764 10566 14816
rect 10778 14764 10784 14816
rect 10836 14804 10842 14816
rect 11793 14807 11851 14813
rect 11793 14804 11805 14807
rect 10836 14776 11805 14804
rect 10836 14764 10842 14776
rect 11793 14773 11805 14776
rect 11839 14773 11851 14807
rect 11793 14767 11851 14773
rect 12161 14807 12219 14813
rect 12161 14773 12173 14807
rect 12207 14804 12219 14807
rect 12342 14804 12348 14816
rect 12207 14776 12348 14804
rect 12207 14773 12219 14776
rect 12161 14767 12219 14773
rect 12342 14764 12348 14776
rect 12400 14764 12406 14816
rect 13538 14764 13544 14816
rect 13596 14804 13602 14816
rect 14001 14807 14059 14813
rect 14001 14804 14013 14807
rect 13596 14776 14013 14804
rect 13596 14764 13602 14776
rect 14001 14773 14013 14776
rect 14047 14773 14059 14807
rect 14001 14767 14059 14773
rect 14366 14764 14372 14816
rect 14424 14804 14430 14816
rect 15473 14807 15531 14813
rect 15473 14804 15485 14807
rect 14424 14776 15485 14804
rect 14424 14764 14430 14776
rect 15473 14773 15485 14776
rect 15519 14773 15531 14807
rect 15580 14804 15608 14844
rect 15838 14832 15844 14844
rect 15896 14832 15902 14884
rect 16853 14875 16911 14881
rect 16853 14841 16865 14875
rect 16899 14872 16911 14875
rect 17034 14872 17040 14884
rect 16899 14844 17040 14872
rect 16899 14841 16911 14844
rect 16853 14835 16911 14841
rect 17034 14832 17040 14844
rect 17092 14832 17098 14884
rect 18800 14872 18828 14971
rect 19610 14968 19616 14980
rect 19668 14968 19674 15020
rect 17144 14844 18828 14872
rect 17144 14804 17172 14844
rect 18322 14804 18328 14816
rect 15580 14776 17172 14804
rect 18283 14776 18328 14804
rect 15473 14767 15531 14773
rect 18322 14764 18328 14776
rect 18380 14764 18386 14816
rect 1104 14714 23828 14736
rect 1104 14662 3790 14714
rect 3842 14662 3854 14714
rect 3906 14662 3918 14714
rect 3970 14662 3982 14714
rect 4034 14662 4046 14714
rect 4098 14662 9471 14714
rect 9523 14662 9535 14714
rect 9587 14662 9599 14714
rect 9651 14662 9663 14714
rect 9715 14662 9727 14714
rect 9779 14662 15152 14714
rect 15204 14662 15216 14714
rect 15268 14662 15280 14714
rect 15332 14662 15344 14714
rect 15396 14662 15408 14714
rect 15460 14662 20833 14714
rect 20885 14662 20897 14714
rect 20949 14662 20961 14714
rect 21013 14662 21025 14714
rect 21077 14662 21089 14714
rect 21141 14662 23828 14714
rect 1104 14640 23828 14662
rect 1762 14560 1768 14612
rect 1820 14600 1826 14612
rect 2130 14600 2136 14612
rect 1820 14572 2136 14600
rect 1820 14560 1826 14572
rect 2130 14560 2136 14572
rect 2188 14560 2194 14612
rect 2590 14600 2596 14612
rect 2551 14572 2596 14600
rect 2590 14560 2596 14572
rect 2648 14560 2654 14612
rect 2682 14560 2688 14612
rect 2740 14600 2746 14612
rect 2777 14603 2835 14609
rect 2777 14600 2789 14603
rect 2740 14572 2789 14600
rect 2740 14560 2746 14572
rect 2777 14569 2789 14572
rect 2823 14569 2835 14603
rect 2777 14563 2835 14569
rect 3142 14560 3148 14612
rect 3200 14600 3206 14612
rect 4065 14603 4123 14609
rect 3200 14572 4016 14600
rect 3200 14560 3206 14572
rect 2608 14532 2636 14560
rect 3988 14544 4016 14572
rect 4065 14569 4077 14603
rect 4111 14600 4123 14603
rect 4154 14600 4160 14612
rect 4111 14572 4160 14600
rect 4111 14569 4123 14572
rect 4065 14563 4123 14569
rect 4154 14560 4160 14572
rect 4212 14560 4218 14612
rect 5626 14600 5632 14612
rect 4264 14572 5632 14600
rect 2608 14504 3924 14532
rect 1578 14424 1584 14476
rect 1636 14464 1642 14476
rect 3694 14464 3700 14476
rect 1636 14436 3700 14464
rect 1636 14424 1642 14436
rect 3694 14424 3700 14436
rect 3752 14424 3758 14476
rect 3896 14464 3924 14504
rect 3970 14492 3976 14544
rect 4028 14532 4034 14544
rect 4264 14532 4292 14572
rect 5626 14560 5632 14572
rect 5684 14600 5690 14612
rect 6362 14600 6368 14612
rect 5684 14572 6368 14600
rect 5684 14560 5690 14572
rect 6362 14560 6368 14572
rect 6420 14600 6426 14612
rect 6822 14600 6828 14612
rect 6420 14572 6828 14600
rect 6420 14560 6426 14572
rect 6822 14560 6828 14572
rect 6880 14560 6886 14612
rect 7101 14603 7159 14609
rect 7101 14569 7113 14603
rect 7147 14569 7159 14603
rect 7101 14563 7159 14569
rect 7285 14603 7343 14609
rect 7285 14569 7297 14603
rect 7331 14600 7343 14603
rect 8018 14600 8024 14612
rect 7331 14572 8024 14600
rect 7331 14569 7343 14572
rect 7285 14563 7343 14569
rect 4028 14504 4292 14532
rect 4028 14492 4034 14504
rect 4338 14492 4344 14544
rect 4396 14532 4402 14544
rect 4982 14532 4988 14544
rect 4396 14504 4988 14532
rect 4396 14492 4402 14504
rect 4982 14492 4988 14504
rect 5040 14492 5046 14544
rect 5258 14492 5264 14544
rect 5316 14532 5322 14544
rect 7116 14532 7144 14563
rect 8018 14560 8024 14572
rect 8076 14560 8082 14612
rect 10778 14600 10784 14612
rect 10739 14572 10784 14600
rect 10778 14560 10784 14572
rect 10836 14560 10842 14612
rect 11241 14603 11299 14609
rect 11241 14569 11253 14603
rect 11287 14600 11299 14603
rect 11606 14600 11612 14612
rect 11287 14572 11612 14600
rect 11287 14569 11299 14572
rect 11241 14563 11299 14569
rect 5316 14504 7144 14532
rect 9125 14535 9183 14541
rect 5316 14492 5322 14504
rect 5718 14464 5724 14476
rect 3896 14436 5580 14464
rect 5679 14436 5724 14464
rect 2866 14356 2872 14408
rect 2924 14396 2930 14408
rect 4065 14399 4123 14405
rect 4065 14396 4077 14399
rect 2924 14368 4077 14396
rect 2924 14356 2930 14368
rect 4065 14365 4077 14368
rect 4111 14365 4123 14399
rect 4065 14359 4123 14365
rect 4341 14399 4399 14405
rect 4341 14365 4353 14399
rect 4387 14365 4399 14399
rect 4341 14359 4399 14365
rect 5077 14399 5135 14405
rect 5077 14365 5089 14399
rect 5123 14365 5135 14399
rect 5442 14396 5448 14408
rect 5403 14368 5448 14396
rect 5077 14359 5135 14365
rect 2406 14288 2412 14340
rect 2464 14328 2470 14340
rect 2958 14328 2964 14340
rect 2464 14300 2964 14328
rect 2464 14288 2470 14300
rect 2958 14288 2964 14300
rect 3016 14328 3022 14340
rect 3694 14328 3700 14340
rect 3016 14300 3700 14328
rect 3016 14288 3022 14300
rect 3694 14288 3700 14300
rect 3752 14288 3758 14340
rect 2761 14263 2819 14269
rect 2761 14229 2773 14263
rect 2807 14260 2819 14263
rect 2866 14260 2872 14272
rect 2807 14232 2872 14260
rect 2807 14229 2819 14232
rect 2761 14223 2819 14229
rect 2866 14220 2872 14232
rect 2924 14220 2930 14272
rect 4246 14260 4252 14272
rect 4207 14232 4252 14260
rect 4246 14220 4252 14232
rect 4304 14220 4310 14272
rect 4356 14260 4384 14359
rect 5092 14328 5120 14359
rect 5442 14356 5448 14368
rect 5500 14356 5506 14408
rect 5350 14328 5356 14340
rect 5092 14300 5356 14328
rect 5350 14288 5356 14300
rect 5408 14288 5414 14340
rect 5552 14328 5580 14436
rect 5718 14424 5724 14436
rect 5776 14424 5782 14476
rect 5905 14399 5963 14405
rect 5905 14365 5917 14399
rect 5951 14396 5963 14399
rect 6012 14396 6040 14504
rect 9125 14501 9137 14535
rect 9171 14501 9183 14535
rect 9125 14495 9183 14501
rect 6822 14424 6828 14476
rect 6880 14464 6886 14476
rect 9140 14464 9168 14495
rect 10410 14492 10416 14544
rect 10468 14532 10474 14544
rect 10689 14535 10747 14541
rect 10689 14532 10701 14535
rect 10468 14504 10701 14532
rect 10468 14492 10474 14504
rect 10689 14501 10701 14504
rect 10735 14532 10747 14535
rect 11256 14532 11284 14563
rect 11606 14560 11612 14572
rect 11664 14560 11670 14612
rect 11701 14603 11759 14609
rect 11701 14569 11713 14603
rect 11747 14600 11759 14603
rect 12345 14603 12403 14609
rect 12345 14600 12357 14603
rect 11747 14572 12357 14600
rect 11747 14569 11759 14572
rect 11701 14563 11759 14569
rect 12345 14569 12357 14572
rect 12391 14600 12403 14603
rect 12802 14600 12808 14612
rect 12391 14572 12808 14600
rect 12391 14569 12403 14572
rect 12345 14563 12403 14569
rect 12802 14560 12808 14572
rect 12860 14560 12866 14612
rect 13814 14560 13820 14612
rect 13872 14600 13878 14612
rect 14277 14603 14335 14609
rect 14277 14600 14289 14603
rect 13872 14572 14289 14600
rect 13872 14560 13878 14572
rect 14277 14569 14289 14572
rect 14323 14569 14335 14603
rect 14277 14563 14335 14569
rect 15473 14603 15531 14609
rect 15473 14569 15485 14603
rect 15519 14600 15531 14603
rect 15838 14600 15844 14612
rect 15519 14572 15844 14600
rect 15519 14569 15531 14572
rect 15473 14563 15531 14569
rect 15838 14560 15844 14572
rect 15896 14560 15902 14612
rect 15930 14560 15936 14612
rect 15988 14600 15994 14612
rect 16574 14600 16580 14612
rect 15988 14572 16436 14600
rect 16535 14572 16580 14600
rect 15988 14560 15994 14572
rect 11514 14532 11520 14544
rect 10735 14504 11284 14532
rect 11440 14504 11520 14532
rect 10735 14501 10747 14504
rect 10689 14495 10747 14501
rect 11440 14473 11468 14504
rect 11514 14492 11520 14504
rect 11572 14492 11578 14544
rect 12529 14535 12587 14541
rect 12529 14501 12541 14535
rect 12575 14532 12587 14535
rect 15749 14535 15807 14541
rect 12575 14504 15148 14532
rect 12575 14501 12587 14504
rect 12529 14495 12587 14501
rect 6880 14436 8156 14464
rect 6880 14424 6886 14436
rect 6454 14396 6460 14408
rect 5951 14368 6040 14396
rect 6415 14368 6460 14396
rect 5951 14365 5963 14368
rect 5905 14359 5963 14365
rect 6454 14356 6460 14368
rect 6512 14356 6518 14408
rect 6564 14368 7052 14396
rect 6564 14328 6592 14368
rect 5552 14300 5948 14328
rect 5810 14260 5816 14272
rect 4356 14232 5816 14260
rect 5810 14220 5816 14232
rect 5868 14220 5874 14272
rect 5920 14260 5948 14300
rect 6104 14300 6592 14328
rect 6104 14260 6132 14300
rect 6822 14288 6828 14340
rect 6880 14328 6886 14340
rect 6917 14331 6975 14337
rect 6917 14328 6929 14331
rect 6880 14300 6929 14328
rect 6880 14288 6886 14300
rect 6917 14297 6929 14300
rect 6963 14297 6975 14331
rect 7024 14328 7052 14368
rect 7374 14356 7380 14408
rect 7432 14396 7438 14408
rect 8128 14405 8156 14436
rect 8312 14436 9168 14464
rect 11425 14467 11483 14473
rect 8312 14405 8340 14436
rect 11425 14433 11437 14467
rect 11471 14433 11483 14467
rect 11425 14427 11483 14433
rect 13633 14467 13691 14473
rect 13633 14433 13645 14467
rect 13679 14464 13691 14467
rect 14645 14467 14703 14473
rect 14645 14464 14657 14467
rect 13679 14436 14657 14464
rect 13679 14433 13691 14436
rect 13633 14427 13691 14433
rect 14645 14433 14657 14436
rect 14691 14433 14703 14467
rect 14645 14427 14703 14433
rect 8021 14399 8079 14405
rect 8021 14396 8033 14399
rect 7432 14368 8033 14396
rect 7432 14356 7438 14368
rect 8021 14365 8033 14368
rect 8067 14365 8079 14399
rect 8021 14359 8079 14365
rect 8113 14399 8171 14405
rect 8113 14365 8125 14399
rect 8159 14365 8171 14399
rect 8113 14359 8171 14365
rect 8297 14399 8355 14405
rect 8297 14365 8309 14399
rect 8343 14365 8355 14399
rect 8297 14359 8355 14365
rect 8389 14399 8447 14405
rect 8389 14365 8401 14399
rect 8435 14365 8447 14399
rect 8389 14359 8447 14365
rect 7117 14331 7175 14337
rect 7117 14328 7129 14331
rect 7024 14300 7129 14328
rect 6917 14291 6975 14297
rect 7117 14297 7129 14300
rect 7163 14297 7175 14331
rect 7117 14291 7175 14297
rect 7742 14288 7748 14340
rect 7800 14328 7806 14340
rect 8404 14328 8432 14359
rect 9306 14356 9312 14408
rect 9364 14396 9370 14408
rect 9401 14399 9459 14405
rect 9401 14396 9413 14399
rect 9364 14368 9413 14396
rect 9364 14356 9370 14368
rect 9401 14365 9413 14368
rect 9447 14365 9459 14399
rect 9858 14396 9864 14408
rect 9819 14368 9864 14396
rect 9401 14359 9459 14365
rect 9858 14356 9864 14368
rect 9916 14356 9922 14408
rect 10781 14399 10839 14405
rect 10781 14365 10793 14399
rect 10827 14396 10839 14399
rect 11238 14396 11244 14408
rect 10827 14368 11244 14396
rect 10827 14365 10839 14368
rect 10781 14359 10839 14365
rect 11238 14356 11244 14368
rect 11296 14356 11302 14408
rect 11517 14399 11575 14405
rect 11517 14365 11529 14399
rect 11563 14396 11575 14399
rect 11698 14396 11704 14408
rect 11563 14368 11704 14396
rect 11563 14365 11575 14368
rect 11517 14359 11575 14365
rect 9122 14328 9128 14340
rect 7800 14300 8432 14328
rect 9083 14300 9128 14328
rect 7800 14288 7806 14300
rect 9122 14288 9128 14300
rect 9180 14288 9186 14340
rect 10505 14331 10563 14337
rect 10505 14297 10517 14331
rect 10551 14328 10563 14331
rect 11054 14328 11060 14340
rect 10551 14300 11060 14328
rect 10551 14297 10563 14300
rect 10505 14291 10563 14297
rect 11054 14288 11060 14300
rect 11112 14328 11118 14340
rect 11532 14328 11560 14359
rect 11698 14356 11704 14368
rect 11756 14356 11762 14408
rect 12710 14356 12716 14408
rect 12768 14396 12774 14408
rect 13078 14396 13084 14408
rect 12768 14368 13084 14396
rect 12768 14356 12774 14368
rect 13078 14356 13084 14368
rect 13136 14396 13142 14408
rect 13541 14399 13599 14405
rect 13541 14396 13553 14399
rect 13136 14368 13553 14396
rect 13136 14356 13142 14368
rect 13541 14365 13553 14368
rect 13587 14365 13599 14399
rect 13541 14359 13599 14365
rect 13725 14399 13783 14405
rect 13725 14365 13737 14399
rect 13771 14365 13783 14399
rect 14366 14396 14372 14408
rect 14327 14368 14372 14396
rect 13725 14359 13783 14365
rect 11112 14300 11560 14328
rect 11112 14288 11118 14300
rect 11790 14288 11796 14340
rect 11848 14328 11854 14340
rect 12161 14331 12219 14337
rect 12161 14328 12173 14331
rect 11848 14300 12173 14328
rect 11848 14288 11854 14300
rect 12161 14297 12173 14300
rect 12207 14297 12219 14331
rect 12342 14328 12348 14340
rect 12303 14300 12348 14328
rect 12161 14291 12219 14297
rect 12342 14288 12348 14300
rect 12400 14288 12406 14340
rect 13740 14328 13768 14359
rect 14366 14356 14372 14368
rect 14424 14356 14430 14408
rect 14458 14356 14464 14408
rect 14516 14396 14522 14408
rect 14734 14396 14740 14408
rect 14516 14368 14561 14396
rect 14695 14368 14740 14396
rect 14516 14356 14522 14368
rect 14734 14356 14740 14368
rect 14792 14356 14798 14408
rect 15120 14396 15148 14504
rect 15749 14501 15761 14535
rect 15795 14532 15807 14535
rect 16114 14532 16120 14544
rect 15795 14504 16120 14532
rect 15795 14501 15807 14504
rect 15749 14495 15807 14501
rect 15562 14424 15568 14476
rect 15620 14464 15626 14476
rect 15841 14467 15899 14473
rect 15841 14464 15853 14467
rect 15620 14436 15853 14464
rect 15620 14424 15626 14436
rect 15841 14433 15853 14436
rect 15887 14433 15899 14467
rect 15948 14464 15976 14504
rect 16114 14492 16120 14504
rect 16172 14492 16178 14544
rect 16408 14532 16436 14572
rect 16574 14560 16580 14572
rect 16632 14560 16638 14612
rect 16666 14560 16672 14612
rect 16724 14600 16730 14612
rect 18141 14603 18199 14609
rect 16724 14572 17356 14600
rect 16724 14560 16730 14572
rect 17328 14532 17356 14572
rect 18141 14569 18153 14603
rect 18187 14600 18199 14603
rect 18414 14600 18420 14612
rect 18187 14572 18420 14600
rect 18187 14569 18199 14572
rect 18141 14563 18199 14569
rect 18414 14560 18420 14572
rect 18472 14560 18478 14612
rect 19978 14532 19984 14544
rect 16408 14504 17264 14532
rect 17328 14504 19984 14532
rect 15948 14436 16896 14464
rect 15841 14427 15899 14433
rect 15120 14368 15608 14396
rect 15378 14328 15384 14340
rect 13740 14300 15384 14328
rect 15378 14288 15384 14300
rect 15436 14288 15442 14340
rect 15580 14328 15608 14368
rect 15654 14356 15660 14408
rect 15712 14396 15718 14408
rect 15930 14396 15936 14408
rect 15712 14368 15757 14396
rect 15891 14368 15936 14396
rect 15712 14356 15718 14368
rect 15930 14356 15936 14368
rect 15988 14356 15994 14408
rect 16117 14399 16175 14405
rect 16117 14365 16129 14399
rect 16163 14396 16175 14399
rect 16206 14396 16212 14408
rect 16163 14368 16212 14396
rect 16163 14365 16175 14368
rect 16117 14359 16175 14365
rect 16206 14356 16212 14368
rect 16264 14396 16270 14408
rect 16666 14396 16672 14408
rect 16264 14368 16672 14396
rect 16264 14356 16270 14368
rect 16666 14356 16672 14368
rect 16724 14356 16730 14408
rect 16868 14405 16896 14436
rect 16853 14399 16911 14405
rect 16853 14365 16865 14399
rect 16899 14365 16911 14399
rect 16853 14359 16911 14365
rect 16945 14399 17003 14405
rect 16945 14365 16957 14399
rect 16991 14365 17003 14399
rect 16945 14359 17003 14365
rect 15838 14328 15844 14340
rect 15580 14300 15844 14328
rect 15838 14288 15844 14300
rect 15896 14288 15902 14340
rect 15948 14328 15976 14356
rect 16960 14328 16988 14359
rect 17034 14356 17040 14408
rect 17092 14396 17098 14408
rect 17236 14405 17264 14504
rect 19978 14492 19984 14504
rect 20036 14532 20042 14544
rect 20441 14535 20499 14541
rect 20441 14532 20453 14535
rect 20036 14504 20453 14532
rect 20036 14492 20042 14504
rect 20441 14501 20453 14504
rect 20487 14501 20499 14535
rect 20441 14495 20499 14501
rect 18785 14467 18843 14473
rect 18785 14433 18797 14467
rect 18831 14464 18843 14467
rect 19058 14464 19064 14476
rect 18831 14436 19064 14464
rect 18831 14433 18843 14436
rect 18785 14427 18843 14433
rect 19058 14424 19064 14436
rect 19116 14424 19122 14476
rect 17221 14399 17279 14405
rect 17092 14368 17137 14396
rect 17092 14356 17098 14368
rect 17221 14365 17233 14399
rect 17267 14396 17279 14399
rect 18414 14396 18420 14408
rect 17267 14368 18420 14396
rect 17267 14365 17279 14368
rect 17221 14359 17279 14365
rect 18414 14356 18420 14368
rect 18472 14396 18478 14408
rect 19613 14399 19671 14405
rect 19613 14396 19625 14399
rect 18472 14368 19625 14396
rect 18472 14356 18478 14368
rect 19613 14365 19625 14368
rect 19659 14396 19671 14399
rect 19702 14396 19708 14408
rect 19659 14368 19708 14396
rect 19659 14365 19671 14368
rect 19613 14359 19671 14365
rect 19702 14356 19708 14368
rect 19760 14396 19766 14408
rect 20438 14396 20444 14408
rect 19760 14368 20444 14396
rect 19760 14356 19766 14368
rect 20438 14356 20444 14368
rect 20496 14396 20502 14408
rect 20625 14399 20683 14405
rect 20625 14396 20637 14399
rect 20496 14368 20637 14396
rect 20496 14356 20502 14368
rect 20625 14365 20637 14368
rect 20671 14365 20683 14399
rect 20625 14359 20683 14365
rect 21634 14328 21640 14340
rect 15948 14300 16988 14328
rect 18340 14300 21640 14328
rect 5920 14232 6132 14260
rect 7837 14263 7895 14269
rect 7837 14229 7849 14263
rect 7883 14260 7895 14263
rect 8110 14260 8116 14272
rect 7883 14232 8116 14260
rect 7883 14229 7895 14232
rect 7837 14223 7895 14229
rect 8110 14220 8116 14232
rect 8168 14220 8174 14272
rect 9214 14220 9220 14272
rect 9272 14260 9278 14272
rect 9309 14263 9367 14269
rect 9309 14260 9321 14263
rect 9272 14232 9321 14260
rect 9272 14220 9278 14232
rect 9309 14229 9321 14232
rect 9355 14229 9367 14263
rect 9950 14260 9956 14272
rect 9911 14232 9956 14260
rect 9309 14223 9367 14229
rect 9950 14220 9956 14232
rect 10008 14220 10014 14272
rect 13814 14220 13820 14272
rect 13872 14260 13878 14272
rect 15286 14260 15292 14272
rect 13872 14232 15292 14260
rect 13872 14220 13878 14232
rect 15286 14220 15292 14232
rect 15344 14220 15350 14272
rect 15654 14220 15660 14272
rect 15712 14260 15718 14272
rect 16206 14260 16212 14272
rect 15712 14232 16212 14260
rect 15712 14220 15718 14232
rect 16206 14220 16212 14232
rect 16264 14220 16270 14272
rect 16666 14220 16672 14272
rect 16724 14260 16730 14272
rect 18340 14260 18368 14300
rect 21634 14288 21640 14300
rect 21692 14288 21698 14340
rect 18506 14260 18512 14272
rect 16724 14232 18368 14260
rect 18467 14232 18512 14260
rect 16724 14220 16730 14232
rect 18506 14220 18512 14232
rect 18564 14220 18570 14272
rect 18601 14263 18659 14269
rect 18601 14229 18613 14263
rect 18647 14260 18659 14263
rect 19150 14260 19156 14272
rect 18647 14232 19156 14260
rect 18647 14229 18659 14232
rect 18601 14223 18659 14229
rect 19150 14220 19156 14232
rect 19208 14220 19214 14272
rect 19521 14263 19579 14269
rect 19521 14229 19533 14263
rect 19567 14260 19579 14263
rect 19610 14260 19616 14272
rect 19567 14232 19616 14260
rect 19567 14229 19579 14232
rect 19521 14223 19579 14229
rect 19610 14220 19616 14232
rect 19668 14220 19674 14272
rect 1104 14170 23987 14192
rect 1104 14118 6630 14170
rect 6682 14118 6694 14170
rect 6746 14118 6758 14170
rect 6810 14118 6822 14170
rect 6874 14118 6886 14170
rect 6938 14118 12311 14170
rect 12363 14118 12375 14170
rect 12427 14118 12439 14170
rect 12491 14118 12503 14170
rect 12555 14118 12567 14170
rect 12619 14118 17992 14170
rect 18044 14118 18056 14170
rect 18108 14118 18120 14170
rect 18172 14118 18184 14170
rect 18236 14118 18248 14170
rect 18300 14118 23673 14170
rect 23725 14118 23737 14170
rect 23789 14118 23801 14170
rect 23853 14118 23865 14170
rect 23917 14118 23929 14170
rect 23981 14118 23987 14170
rect 1104 14096 23987 14118
rect 1854 14016 1860 14068
rect 1912 14056 1918 14068
rect 2507 14059 2565 14065
rect 2507 14056 2519 14059
rect 1912 14028 2519 14056
rect 1912 14016 1918 14028
rect 2507 14025 2519 14028
rect 2553 14025 2565 14059
rect 2507 14019 2565 14025
rect 2682 14016 2688 14068
rect 2740 14016 2746 14068
rect 4890 14056 4896 14068
rect 4851 14028 4896 14056
rect 4890 14016 4896 14028
rect 4948 14016 4954 14068
rect 7193 14059 7251 14065
rect 5000 14028 7052 14056
rect 2406 13988 2412 14000
rect 2367 13960 2412 13988
rect 2406 13948 2412 13960
rect 2464 13948 2470 14000
rect 2700 13988 2728 14016
rect 2608 13960 3372 13988
rect 1762 13880 1768 13932
rect 1820 13920 1826 13932
rect 1857 13923 1915 13929
rect 1857 13920 1869 13923
rect 1820 13892 1869 13920
rect 1820 13880 1826 13892
rect 1857 13889 1869 13892
rect 1903 13889 1915 13923
rect 1857 13883 1915 13889
rect 2130 13880 2136 13932
rect 2188 13920 2194 13932
rect 2608 13929 2636 13960
rect 2593 13923 2651 13929
rect 2593 13920 2605 13923
rect 2188 13892 2605 13920
rect 2188 13880 2194 13892
rect 2593 13889 2605 13892
rect 2639 13889 2651 13923
rect 2593 13883 2651 13889
rect 2685 13923 2743 13929
rect 2685 13889 2697 13923
rect 2731 13920 2743 13923
rect 2866 13920 2872 13932
rect 2731 13892 2872 13920
rect 2731 13889 2743 13892
rect 2685 13883 2743 13889
rect 2866 13880 2872 13892
rect 2924 13920 2930 13932
rect 3344 13929 3372 13960
rect 3602 13948 3608 14000
rect 3660 13988 3666 14000
rect 4522 13988 4528 14000
rect 3660 13960 4528 13988
rect 3660 13948 3666 13960
rect 4522 13948 4528 13960
rect 4580 13988 4586 14000
rect 5000 13988 5028 14028
rect 5166 13988 5172 14000
rect 4580 13960 5028 13988
rect 5127 13960 5172 13988
rect 4580 13948 4586 13960
rect 3145 13923 3203 13929
rect 3145 13920 3157 13923
rect 2924 13892 3157 13920
rect 2924 13880 2930 13892
rect 3145 13889 3157 13892
rect 3191 13889 3203 13923
rect 3145 13883 3203 13889
rect 3329 13923 3387 13929
rect 3329 13889 3341 13923
rect 3375 13889 3387 13923
rect 4154 13920 4160 13932
rect 4115 13892 4160 13920
rect 3329 13883 3387 13889
rect 4154 13880 4160 13892
rect 4212 13880 4218 13932
rect 4341 13923 4399 13929
rect 4341 13889 4353 13923
rect 4387 13920 4399 13923
rect 4430 13920 4436 13932
rect 4387 13892 4436 13920
rect 4387 13889 4399 13892
rect 4341 13883 4399 13889
rect 4430 13880 4436 13892
rect 4488 13880 4494 13932
rect 5000 13920 5028 13960
rect 5166 13948 5172 13960
rect 5224 13948 5230 14000
rect 5261 13991 5319 13997
rect 5261 13957 5273 13991
rect 5307 13988 5319 13991
rect 5718 13988 5724 14000
rect 5307 13960 5724 13988
rect 5307 13957 5319 13960
rect 5261 13951 5319 13957
rect 5077 13923 5135 13929
rect 5077 13920 5089 13923
rect 5000 13892 5089 13920
rect 5077 13889 5089 13892
rect 5123 13889 5135 13923
rect 5077 13883 5135 13889
rect 5276 13852 5304 13951
rect 5718 13948 5724 13960
rect 5776 13948 5782 14000
rect 6822 13988 6828 14000
rect 6783 13960 6828 13988
rect 6822 13948 6828 13960
rect 6880 13948 6886 14000
rect 5445 13923 5503 13929
rect 5445 13889 5457 13923
rect 5491 13920 5503 13923
rect 5902 13920 5908 13932
rect 5491 13892 5908 13920
rect 5491 13889 5503 13892
rect 5445 13883 5503 13889
rect 5902 13880 5908 13892
rect 5960 13880 5966 13932
rect 6362 13880 6368 13932
rect 6420 13920 6426 13932
rect 6641 13923 6699 13929
rect 6641 13920 6653 13923
rect 6420 13892 6653 13920
rect 6420 13880 6426 13892
rect 6641 13889 6653 13892
rect 6687 13889 6699 13923
rect 6914 13920 6920 13932
rect 6875 13892 6920 13920
rect 6641 13883 6699 13889
rect 6914 13880 6920 13892
rect 6972 13880 6978 13932
rect 7024 13929 7052 14028
rect 7193 14025 7205 14059
rect 7239 14056 7251 14059
rect 7282 14056 7288 14068
rect 7239 14028 7288 14056
rect 7239 14025 7251 14028
rect 7193 14019 7251 14025
rect 7282 14016 7288 14028
rect 7340 14016 7346 14068
rect 8294 14056 8300 14068
rect 8255 14028 8300 14056
rect 8294 14016 8300 14028
rect 8352 14016 8358 14068
rect 9030 14056 9036 14068
rect 8991 14028 9036 14056
rect 9030 14016 9036 14028
rect 9088 14016 9094 14068
rect 10965 14059 11023 14065
rect 10965 14025 10977 14059
rect 11011 14056 11023 14059
rect 11330 14056 11336 14068
rect 11011 14028 11336 14056
rect 11011 14025 11023 14028
rect 10965 14019 11023 14025
rect 11330 14016 11336 14028
rect 11388 14016 11394 14068
rect 12253 14059 12311 14065
rect 12253 14025 12265 14059
rect 12299 14056 12311 14059
rect 13814 14056 13820 14068
rect 12299 14028 13820 14056
rect 12299 14025 12311 14028
rect 12253 14019 12311 14025
rect 13814 14016 13820 14028
rect 13872 14016 13878 14068
rect 14458 14016 14464 14068
rect 14516 14056 14522 14068
rect 15197 14059 15255 14065
rect 15197 14056 15209 14059
rect 14516 14028 15209 14056
rect 14516 14016 14522 14028
rect 15197 14025 15209 14028
rect 15243 14025 15255 14059
rect 15197 14019 15255 14025
rect 15286 14016 15292 14068
rect 15344 14056 15350 14068
rect 16666 14056 16672 14068
rect 15344 14028 16672 14056
rect 15344 14016 15350 14028
rect 16666 14016 16672 14028
rect 16724 14016 16730 14068
rect 16853 14059 16911 14065
rect 16853 14025 16865 14059
rect 16899 14056 16911 14059
rect 17034 14056 17040 14068
rect 16899 14028 17040 14056
rect 16899 14025 16911 14028
rect 16853 14019 16911 14025
rect 17034 14016 17040 14028
rect 17092 14016 17098 14068
rect 17221 14059 17279 14065
rect 17221 14025 17233 14059
rect 17267 14056 17279 14059
rect 18782 14056 18788 14068
rect 17267 14028 18788 14056
rect 17267 14025 17279 14028
rect 17221 14019 17279 14025
rect 18782 14016 18788 14028
rect 18840 14016 18846 14068
rect 19150 14056 19156 14068
rect 19111 14028 19156 14056
rect 19150 14016 19156 14028
rect 19208 14016 19214 14068
rect 20257 14059 20315 14065
rect 20257 14056 20269 14059
rect 19260 14028 20269 14056
rect 7098 13948 7104 14000
rect 7156 13988 7162 14000
rect 7374 13988 7380 14000
rect 7156 13960 7380 13988
rect 7156 13948 7162 13960
rect 7374 13948 7380 13960
rect 7432 13948 7438 14000
rect 7837 13991 7895 13997
rect 7837 13957 7849 13991
rect 7883 13988 7895 13991
rect 8018 13988 8024 14000
rect 7883 13960 8024 13988
rect 7883 13957 7895 13960
rect 7837 13951 7895 13957
rect 8018 13948 8024 13960
rect 8076 13948 8082 14000
rect 12158 13948 12164 14000
rect 12216 13948 12222 14000
rect 14734 13988 14740 14000
rect 12406 13960 14504 13988
rect 14647 13960 14740 13988
rect 7009 13923 7067 13929
rect 7009 13889 7021 13923
rect 7055 13920 7067 13923
rect 7282 13920 7288 13932
rect 7055 13892 7288 13920
rect 7055 13889 7067 13892
rect 7009 13883 7067 13889
rect 7282 13880 7288 13892
rect 7340 13920 7346 13932
rect 7742 13920 7748 13932
rect 7340 13892 7748 13920
rect 7340 13880 7346 13892
rect 7742 13880 7748 13892
rect 7800 13880 7806 13932
rect 9214 13920 9220 13932
rect 9175 13892 9220 13920
rect 9214 13880 9220 13892
rect 9272 13880 9278 13932
rect 9306 13880 9312 13932
rect 9364 13920 9370 13932
rect 9861 13923 9919 13929
rect 9861 13920 9873 13923
rect 9364 13892 9873 13920
rect 9364 13880 9370 13892
rect 9861 13889 9873 13892
rect 9907 13889 9919 13923
rect 9861 13883 9919 13889
rect 10778 13880 10784 13932
rect 10836 13920 10842 13932
rect 11701 13923 11759 13929
rect 11701 13920 11713 13923
rect 10836 13892 11713 13920
rect 10836 13880 10842 13892
rect 11701 13889 11713 13892
rect 11747 13889 11759 13923
rect 11701 13883 11759 13889
rect 11977 13923 12035 13929
rect 11977 13889 11989 13923
rect 12023 13920 12035 13923
rect 12176 13920 12204 13948
rect 12406 13920 12434 13960
rect 12023 13892 12434 13920
rect 12023 13889 12035 13892
rect 11977 13883 12035 13889
rect 9030 13852 9036 13864
rect 2746 13824 5304 13852
rect 5460 13824 9036 13852
rect 2746 13796 2774 13824
rect 5460 13796 5488 13824
rect 9030 13812 9036 13824
rect 9088 13812 9094 13864
rect 10686 13812 10692 13864
rect 10744 13852 10750 13864
rect 10873 13855 10931 13861
rect 10873 13852 10885 13855
rect 10744 13824 10885 13852
rect 10744 13812 10750 13824
rect 10873 13821 10885 13824
rect 10919 13821 10931 13855
rect 10873 13815 10931 13821
rect 11057 13855 11115 13861
rect 11057 13821 11069 13855
rect 11103 13821 11115 13855
rect 11057 13815 11115 13821
rect 2682 13744 2688 13796
rect 2740 13756 2774 13796
rect 4341 13787 4399 13793
rect 2740 13744 2746 13756
rect 4341 13753 4353 13787
rect 4387 13784 4399 13787
rect 5350 13784 5356 13796
rect 4387 13756 5356 13784
rect 4387 13753 4399 13756
rect 4341 13747 4399 13753
rect 5350 13744 5356 13756
rect 5408 13744 5414 13796
rect 5442 13744 5448 13796
rect 5500 13744 5506 13796
rect 7006 13784 7012 13796
rect 5644 13756 7012 13784
rect 3142 13716 3148 13728
rect 3103 13688 3148 13716
rect 3142 13676 3148 13688
rect 3200 13676 3206 13728
rect 4798 13676 4804 13728
rect 4856 13716 4862 13728
rect 5644 13716 5672 13756
rect 7006 13744 7012 13756
rect 7064 13744 7070 13796
rect 8110 13784 8116 13796
rect 8071 13756 8116 13784
rect 8110 13744 8116 13756
rect 8168 13744 8174 13796
rect 10778 13744 10784 13796
rect 10836 13784 10842 13796
rect 11072 13784 11100 13815
rect 11514 13812 11520 13864
rect 11572 13852 11578 13864
rect 11992 13852 12020 13883
rect 13354 13880 13360 13932
rect 13412 13920 13418 13932
rect 14476 13929 14504 13960
rect 14734 13948 14740 13960
rect 14792 13988 14798 14000
rect 16758 13988 16764 14000
rect 14792 13960 16764 13988
rect 14792 13948 14798 13960
rect 16758 13948 16764 13960
rect 16816 13948 16822 14000
rect 16942 13948 16948 14000
rect 17000 13988 17006 14000
rect 17865 13991 17923 13997
rect 17865 13988 17877 13991
rect 17000 13960 17877 13988
rect 17000 13948 17006 13960
rect 17865 13957 17877 13960
rect 17911 13957 17923 13991
rect 18322 13988 18328 14000
rect 17865 13951 17923 13957
rect 18156 13960 18328 13988
rect 14185 13923 14243 13929
rect 14185 13920 14197 13923
rect 13412 13892 14197 13920
rect 13412 13880 13418 13892
rect 14185 13889 14197 13892
rect 14231 13889 14243 13923
rect 14185 13883 14243 13889
rect 14461 13923 14519 13929
rect 14461 13889 14473 13923
rect 14507 13889 14519 13923
rect 14461 13883 14519 13889
rect 14550 13880 14556 13932
rect 14608 13920 14614 13932
rect 15473 13923 15531 13929
rect 14608 13892 14653 13920
rect 14608 13880 14614 13892
rect 15473 13889 15485 13923
rect 15519 13920 15531 13923
rect 15746 13920 15752 13932
rect 15519 13892 15752 13920
rect 15519 13889 15531 13892
rect 15473 13883 15531 13889
rect 15746 13880 15752 13892
rect 15804 13880 15810 13932
rect 18156 13929 18184 13960
rect 18322 13948 18328 13960
rect 18380 13948 18386 14000
rect 18598 13948 18604 14000
rect 18656 13988 18662 14000
rect 19260 13988 19288 14028
rect 20257 14025 20269 14028
rect 20303 14025 20315 14059
rect 20257 14019 20315 14025
rect 19518 13988 19524 14000
rect 18656 13960 19288 13988
rect 19479 13960 19524 13988
rect 18656 13948 18662 13960
rect 19518 13948 19524 13960
rect 19576 13948 19582 14000
rect 17037 13923 17095 13929
rect 17037 13889 17049 13923
rect 17083 13889 17095 13923
rect 17037 13883 17095 13889
rect 17313 13923 17371 13929
rect 17313 13889 17325 13923
rect 17359 13920 17371 13923
rect 18049 13923 18107 13929
rect 17359 13892 17908 13920
rect 17359 13889 17371 13892
rect 17313 13883 17371 13889
rect 12158 13852 12164 13864
rect 11572 13824 12020 13852
rect 12119 13824 12164 13852
rect 11572 13812 11578 13824
rect 12158 13812 12164 13824
rect 12216 13812 12222 13864
rect 13998 13812 14004 13864
rect 14056 13852 14062 13864
rect 14277 13855 14335 13861
rect 14277 13852 14289 13855
rect 14056 13824 14289 13852
rect 14056 13812 14062 13824
rect 14277 13821 14289 13824
rect 14323 13821 14335 13855
rect 15378 13852 15384 13864
rect 15339 13824 15384 13852
rect 14277 13815 14335 13821
rect 15378 13812 15384 13824
rect 15436 13812 15442 13864
rect 15565 13855 15623 13861
rect 15565 13821 15577 13855
rect 15611 13821 15623 13855
rect 15565 13815 15623 13821
rect 15657 13855 15715 13861
rect 15657 13821 15669 13855
rect 15703 13852 15715 13855
rect 16298 13852 16304 13864
rect 15703 13824 16304 13852
rect 15703 13821 15715 13824
rect 15657 13815 15715 13821
rect 10836 13756 11100 13784
rect 10836 13744 10842 13756
rect 12986 13744 12992 13796
rect 13044 13784 13050 13796
rect 15580 13784 15608 13815
rect 16298 13812 16304 13824
rect 16356 13812 16362 13864
rect 17052 13852 17080 13883
rect 17880 13864 17908 13892
rect 18049 13889 18061 13923
rect 18095 13889 18107 13923
rect 18049 13883 18107 13889
rect 18141 13923 18199 13929
rect 18141 13889 18153 13923
rect 18187 13889 18199 13923
rect 18414 13920 18420 13932
rect 18375 13892 18420 13920
rect 18141 13883 18199 13889
rect 17770 13852 17776 13864
rect 17052 13824 17776 13852
rect 17770 13812 17776 13824
rect 17828 13812 17834 13864
rect 17862 13812 17868 13864
rect 17920 13812 17926 13864
rect 13044 13756 15608 13784
rect 18064 13784 18092 13883
rect 18414 13880 18420 13892
rect 18472 13880 18478 13932
rect 19334 13920 19340 13932
rect 19295 13892 19340 13920
rect 19334 13880 19340 13892
rect 19392 13880 19398 13932
rect 19426 13880 19432 13932
rect 19484 13920 19490 13932
rect 19702 13920 19708 13932
rect 19484 13892 19529 13920
rect 19663 13892 19708 13920
rect 19484 13880 19490 13892
rect 19702 13880 19708 13892
rect 19760 13880 19766 13932
rect 19978 13880 19984 13932
rect 20036 13920 20042 13932
rect 20165 13923 20223 13929
rect 20165 13920 20177 13923
rect 20036 13892 20177 13920
rect 20036 13880 20042 13892
rect 20165 13889 20177 13892
rect 20211 13889 20223 13923
rect 20346 13920 20352 13932
rect 20307 13892 20352 13920
rect 20165 13883 20223 13889
rect 20346 13880 20352 13892
rect 20404 13880 20410 13932
rect 18322 13852 18328 13864
rect 18283 13824 18328 13852
rect 18322 13812 18328 13824
rect 18380 13812 18386 13864
rect 18414 13784 18420 13796
rect 18064 13756 18420 13784
rect 13044 13744 13050 13756
rect 4856 13688 5672 13716
rect 5997 13719 6055 13725
rect 4856 13676 4862 13688
rect 5997 13685 6009 13719
rect 6043 13716 6055 13719
rect 6270 13716 6276 13728
rect 6043 13688 6276 13716
rect 6043 13685 6055 13688
rect 5997 13679 6055 13685
rect 6270 13676 6276 13688
rect 6328 13716 6334 13728
rect 6730 13716 6736 13728
rect 6328 13688 6736 13716
rect 6328 13676 6334 13688
rect 6730 13676 6736 13688
rect 6788 13676 6794 13728
rect 10410 13676 10416 13728
rect 10468 13716 10474 13728
rect 10505 13719 10563 13725
rect 10505 13716 10517 13719
rect 10468 13688 10517 13716
rect 10468 13676 10474 13688
rect 10505 13685 10517 13688
rect 10551 13685 10563 13719
rect 10505 13679 10563 13685
rect 12434 13676 12440 13728
rect 12492 13716 12498 13728
rect 12897 13719 12955 13725
rect 12897 13716 12909 13719
rect 12492 13688 12909 13716
rect 12492 13676 12498 13688
rect 12897 13685 12909 13688
rect 12943 13716 12955 13719
rect 13630 13716 13636 13728
rect 12943 13688 13636 13716
rect 12943 13685 12955 13688
rect 12897 13679 12955 13685
rect 13630 13676 13636 13688
rect 13688 13676 13694 13728
rect 15580 13716 15608 13756
rect 18414 13744 18420 13756
rect 18472 13744 18478 13796
rect 15654 13716 15660 13728
rect 15580 13688 15660 13716
rect 15654 13676 15660 13688
rect 15712 13676 15718 13728
rect 16206 13676 16212 13728
rect 16264 13716 16270 13728
rect 16301 13719 16359 13725
rect 16301 13716 16313 13719
rect 16264 13688 16313 13716
rect 16264 13676 16270 13688
rect 16301 13685 16313 13688
rect 16347 13716 16359 13719
rect 17218 13716 17224 13728
rect 16347 13688 17224 13716
rect 16347 13685 16359 13688
rect 16301 13679 16359 13685
rect 17218 13676 17224 13688
rect 17276 13716 17282 13728
rect 18690 13716 18696 13728
rect 17276 13688 18696 13716
rect 17276 13676 17282 13688
rect 18690 13676 18696 13688
rect 18748 13676 18754 13728
rect 1104 13626 23828 13648
rect 1104 13574 3790 13626
rect 3842 13574 3854 13626
rect 3906 13574 3918 13626
rect 3970 13574 3982 13626
rect 4034 13574 4046 13626
rect 4098 13574 9471 13626
rect 9523 13574 9535 13626
rect 9587 13574 9599 13626
rect 9651 13574 9663 13626
rect 9715 13574 9727 13626
rect 9779 13574 15152 13626
rect 15204 13574 15216 13626
rect 15268 13574 15280 13626
rect 15332 13574 15344 13626
rect 15396 13574 15408 13626
rect 15460 13574 20833 13626
rect 20885 13574 20897 13626
rect 20949 13574 20961 13626
rect 21013 13574 21025 13626
rect 21077 13574 21089 13626
rect 21141 13574 23828 13626
rect 1104 13552 23828 13574
rect 1949 13515 2007 13521
rect 1949 13481 1961 13515
rect 1995 13512 2007 13515
rect 3510 13512 3516 13524
rect 1995 13484 3516 13512
rect 1995 13481 2007 13484
rect 1949 13475 2007 13481
rect 3510 13472 3516 13484
rect 3568 13472 3574 13524
rect 4430 13512 4436 13524
rect 4172 13484 4436 13512
rect 4172 13444 4200 13484
rect 4430 13472 4436 13484
rect 4488 13512 4494 13524
rect 4614 13512 4620 13524
rect 4488 13484 4620 13512
rect 4488 13472 4494 13484
rect 4614 13472 4620 13484
rect 4672 13472 4678 13524
rect 4706 13472 4712 13524
rect 4764 13512 4770 13524
rect 4801 13515 4859 13521
rect 4801 13512 4813 13515
rect 4764 13484 4813 13512
rect 4764 13472 4770 13484
rect 4801 13481 4813 13484
rect 4847 13481 4859 13515
rect 6270 13512 6276 13524
rect 4801 13475 4859 13481
rect 4908 13484 6276 13512
rect 2700 13416 4200 13444
rect 2700 13385 2728 13416
rect 4246 13404 4252 13456
rect 4304 13444 4310 13456
rect 4341 13447 4399 13453
rect 4341 13444 4353 13447
rect 4304 13416 4353 13444
rect 4304 13404 4310 13416
rect 4341 13413 4353 13416
rect 4387 13444 4399 13447
rect 4908 13444 4936 13484
rect 6270 13472 6276 13484
rect 6328 13472 6334 13524
rect 6822 13472 6828 13524
rect 6880 13512 6886 13524
rect 8021 13515 8079 13521
rect 8021 13512 8033 13515
rect 6880 13484 8033 13512
rect 6880 13472 6886 13484
rect 8021 13481 8033 13484
rect 8067 13481 8079 13515
rect 8021 13475 8079 13481
rect 8846 13472 8852 13524
rect 8904 13512 8910 13524
rect 10505 13515 10563 13521
rect 10505 13512 10517 13515
rect 8904 13484 10517 13512
rect 8904 13472 8910 13484
rect 10505 13481 10517 13484
rect 10551 13512 10563 13515
rect 10778 13512 10784 13524
rect 10551 13484 10784 13512
rect 10551 13481 10563 13484
rect 10505 13475 10563 13481
rect 10778 13472 10784 13484
rect 10836 13472 10842 13524
rect 11238 13472 11244 13524
rect 11296 13512 11302 13524
rect 11425 13515 11483 13521
rect 11425 13512 11437 13515
rect 11296 13484 11437 13512
rect 11296 13472 11302 13484
rect 11425 13481 11437 13484
rect 11471 13512 11483 13515
rect 11698 13512 11704 13524
rect 11471 13484 11704 13512
rect 11471 13481 11483 13484
rect 11425 13475 11483 13481
rect 11698 13472 11704 13484
rect 11756 13472 11762 13524
rect 11793 13515 11851 13521
rect 11793 13481 11805 13515
rect 11839 13512 11851 13515
rect 12158 13512 12164 13524
rect 11839 13484 12164 13512
rect 11839 13481 11851 13484
rect 11793 13475 11851 13481
rect 12158 13472 12164 13484
rect 12216 13472 12222 13524
rect 12437 13515 12495 13521
rect 12437 13481 12449 13515
rect 12483 13512 12495 13515
rect 14366 13512 14372 13524
rect 12483 13484 14372 13512
rect 12483 13481 12495 13484
rect 12437 13475 12495 13481
rect 4387 13416 4936 13444
rect 4387 13413 4399 13416
rect 4341 13407 4399 13413
rect 5718 13404 5724 13456
rect 5776 13444 5782 13456
rect 5776 13416 8156 13444
rect 5776 13404 5782 13416
rect 2685 13379 2743 13385
rect 2685 13345 2697 13379
rect 2731 13345 2743 13379
rect 4890 13376 4896 13388
rect 2685 13339 2743 13345
rect 2776 13348 4896 13376
rect 1854 13308 1860 13320
rect 1815 13280 1860 13308
rect 1854 13268 1860 13280
rect 1912 13268 1918 13320
rect 2038 13268 2044 13320
rect 2096 13308 2102 13320
rect 2498 13308 2504 13320
rect 2096 13280 2189 13308
rect 2411 13280 2504 13308
rect 2096 13268 2102 13280
rect 2498 13268 2504 13280
rect 2556 13308 2562 13320
rect 2776 13308 2804 13348
rect 4890 13336 4896 13348
rect 4948 13336 4954 13388
rect 6362 13376 6368 13388
rect 6323 13348 6368 13376
rect 6362 13336 6368 13348
rect 6420 13336 6426 13388
rect 6454 13336 6460 13388
rect 6512 13376 6518 13388
rect 6512 13348 6557 13376
rect 6512 13336 6518 13348
rect 8128 13320 8156 13416
rect 9214 13336 9220 13388
rect 9272 13376 9278 13388
rect 9582 13376 9588 13388
rect 9272 13348 9588 13376
rect 9272 13336 9278 13348
rect 9582 13336 9588 13348
rect 9640 13376 9646 13388
rect 9640 13348 10088 13376
rect 9640 13336 9646 13348
rect 2556 13280 2804 13308
rect 2869 13311 2927 13317
rect 2556 13268 2562 13280
rect 2869 13277 2881 13311
rect 2915 13308 2927 13311
rect 3786 13308 3792 13320
rect 2915 13280 3792 13308
rect 2915 13277 2927 13280
rect 2869 13271 2927 13277
rect 3786 13268 3792 13280
rect 3844 13268 3850 13320
rect 4985 13311 5043 13317
rect 4985 13277 4997 13311
rect 5031 13277 5043 13311
rect 4985 13271 5043 13277
rect 2056 13240 2084 13268
rect 2682 13240 2688 13252
rect 2056 13212 2688 13240
rect 2682 13200 2688 13212
rect 2740 13200 2746 13252
rect 3421 13243 3479 13249
rect 3421 13209 3433 13243
rect 3467 13240 3479 13243
rect 4338 13240 4344 13252
rect 3467 13212 4344 13240
rect 3467 13209 3479 13212
rect 3421 13203 3479 13209
rect 4338 13200 4344 13212
rect 4396 13200 4402 13252
rect 5000 13240 5028 13271
rect 5074 13268 5080 13320
rect 5132 13308 5138 13320
rect 5132 13280 5177 13308
rect 5132 13268 5138 13280
rect 5350 13268 5356 13320
rect 5408 13308 5414 13320
rect 5445 13311 5503 13317
rect 5445 13308 5457 13311
rect 5408 13280 5457 13308
rect 5408 13268 5414 13280
rect 5445 13277 5457 13280
rect 5491 13277 5503 13311
rect 5445 13271 5503 13277
rect 6270 13268 6276 13320
rect 6328 13308 6334 13320
rect 6549 13311 6607 13317
rect 6328 13286 6409 13308
rect 6549 13302 6561 13311
rect 6472 13286 6561 13302
rect 6328 13280 6561 13286
rect 6328 13268 6334 13280
rect 6381 13277 6561 13280
rect 6595 13277 6607 13311
rect 6381 13274 6607 13277
rect 6381 13258 6500 13274
rect 6549 13271 6607 13274
rect 6638 13268 6644 13320
rect 6696 13308 6702 13320
rect 7466 13308 7472 13320
rect 6696 13280 6741 13308
rect 7427 13280 7472 13308
rect 6696 13268 6702 13280
rect 7466 13268 7472 13280
rect 7524 13268 7530 13320
rect 7558 13268 7564 13320
rect 7616 13308 7622 13320
rect 7929 13311 7987 13317
rect 7929 13308 7941 13311
rect 7616 13280 7941 13308
rect 7616 13268 7622 13280
rect 7929 13277 7941 13280
rect 7975 13277 7987 13311
rect 8110 13308 8116 13320
rect 8071 13280 8116 13308
rect 7929 13271 7987 13277
rect 8110 13268 8116 13280
rect 8168 13268 8174 13320
rect 9306 13308 9312 13320
rect 9267 13280 9312 13308
rect 9306 13268 9312 13280
rect 9364 13268 9370 13320
rect 10060 13317 10088 13348
rect 11054 13336 11060 13388
rect 11112 13376 11118 13388
rect 11330 13376 11336 13388
rect 11112 13348 11336 13376
rect 11112 13336 11118 13348
rect 11330 13336 11336 13348
rect 11388 13336 11394 13388
rect 12158 13336 12164 13388
rect 12216 13376 12222 13388
rect 12452 13376 12480 13475
rect 14366 13472 14372 13484
rect 14424 13472 14430 13524
rect 15470 13472 15476 13524
rect 15528 13512 15534 13524
rect 15841 13515 15899 13521
rect 15841 13512 15853 13515
rect 15528 13484 15853 13512
rect 15528 13472 15534 13484
rect 15841 13481 15853 13484
rect 15887 13481 15899 13515
rect 15841 13475 15899 13481
rect 16758 13472 16764 13524
rect 16816 13512 16822 13524
rect 18966 13512 18972 13524
rect 16816 13484 18972 13512
rect 16816 13472 16822 13484
rect 18966 13472 18972 13484
rect 19024 13472 19030 13524
rect 19426 13512 19432 13524
rect 19387 13484 19432 13512
rect 19426 13472 19432 13484
rect 19484 13472 19490 13524
rect 19794 13472 19800 13524
rect 19852 13512 19858 13524
rect 20901 13515 20959 13521
rect 20901 13512 20913 13515
rect 19852 13484 20913 13512
rect 19852 13472 19858 13484
rect 20901 13481 20913 13484
rect 20947 13481 20959 13515
rect 20901 13475 20959 13481
rect 12986 13404 12992 13456
rect 13044 13444 13050 13456
rect 13081 13447 13139 13453
rect 13081 13444 13093 13447
rect 13044 13416 13093 13444
rect 13044 13404 13050 13416
rect 13081 13413 13093 13416
rect 13127 13413 13139 13447
rect 13081 13407 13139 13413
rect 13998 13404 14004 13456
rect 14056 13444 14062 13456
rect 14829 13447 14887 13453
rect 14829 13444 14841 13447
rect 14056 13416 14841 13444
rect 14056 13404 14062 13416
rect 14829 13413 14841 13416
rect 14875 13444 14887 13447
rect 14918 13444 14924 13456
rect 14875 13416 14924 13444
rect 14875 13413 14887 13416
rect 14829 13407 14887 13413
rect 14918 13404 14924 13416
rect 14976 13404 14982 13456
rect 15746 13404 15752 13456
rect 15804 13444 15810 13456
rect 17310 13444 17316 13456
rect 15804 13416 17316 13444
rect 15804 13404 15810 13416
rect 17310 13404 17316 13416
rect 17368 13404 17374 13456
rect 17589 13447 17647 13453
rect 17589 13413 17601 13447
rect 17635 13413 17647 13447
rect 19886 13444 19892 13456
rect 17589 13407 17647 13413
rect 18156 13416 19892 13444
rect 17604 13376 17632 13407
rect 12216 13348 12480 13376
rect 16316 13348 17632 13376
rect 12216 13336 12222 13348
rect 10045 13311 10103 13317
rect 10045 13277 10057 13311
rect 10091 13277 10103 13311
rect 11606 13308 11612 13320
rect 11567 13280 11612 13308
rect 10045 13271 10103 13277
rect 11606 13268 11612 13280
rect 11664 13268 11670 13320
rect 12434 13308 12440 13320
rect 12395 13280 12440 13308
rect 12434 13268 12440 13280
rect 12492 13268 12498 13320
rect 12989 13311 13047 13317
rect 12989 13277 13001 13311
rect 13035 13308 13047 13311
rect 13354 13308 13360 13320
rect 13035 13280 13360 13308
rect 13035 13277 13047 13280
rect 12989 13271 13047 13277
rect 13354 13268 13360 13280
rect 13412 13268 13418 13320
rect 15838 13268 15844 13320
rect 15896 13308 15902 13320
rect 16316 13317 16344 13348
rect 16025 13311 16083 13317
rect 16025 13308 16037 13311
rect 15896 13280 16037 13308
rect 15896 13268 15902 13280
rect 16025 13277 16037 13280
rect 16071 13277 16083 13311
rect 16025 13271 16083 13277
rect 16301 13311 16359 13317
rect 16301 13277 16313 13311
rect 16347 13277 16359 13311
rect 16758 13308 16764 13320
rect 16719 13280 16764 13308
rect 16301 13271 16359 13277
rect 16758 13268 16764 13280
rect 16816 13268 16822 13320
rect 16945 13311 17003 13317
rect 16945 13277 16957 13311
rect 16991 13308 17003 13311
rect 17494 13308 17500 13320
rect 16991 13280 17500 13308
rect 16991 13277 17003 13280
rect 16945 13271 17003 13277
rect 17494 13268 17500 13280
rect 17552 13308 17558 13320
rect 18156 13317 18184 13416
rect 19886 13404 19892 13416
rect 19944 13404 19950 13456
rect 18248 13348 20116 13376
rect 18248 13320 18276 13348
rect 17727 13311 17785 13317
rect 17727 13308 17739 13311
rect 17552 13280 17739 13308
rect 17552 13268 17558 13280
rect 17727 13277 17739 13280
rect 17773 13277 17785 13311
rect 17727 13271 17785 13277
rect 18140 13311 18198 13317
rect 18140 13277 18152 13311
rect 18186 13277 18198 13311
rect 18140 13271 18198 13277
rect 18230 13268 18236 13320
rect 18288 13308 18294 13320
rect 18288 13280 18333 13308
rect 18288 13268 18294 13280
rect 18598 13268 18604 13320
rect 18656 13308 18662 13320
rect 18693 13311 18751 13317
rect 18693 13308 18705 13311
rect 18656 13280 18705 13308
rect 18656 13268 18662 13280
rect 18693 13277 18705 13280
rect 18739 13277 18751 13311
rect 18874 13308 18880 13320
rect 18835 13280 18880 13308
rect 18693 13271 18751 13277
rect 18874 13268 18880 13280
rect 18932 13268 18938 13320
rect 18966 13268 18972 13320
rect 19024 13308 19030 13320
rect 19567 13311 19625 13317
rect 19567 13308 19579 13311
rect 19024 13280 19579 13308
rect 19024 13268 19030 13280
rect 19567 13277 19579 13280
rect 19613 13277 19625 13311
rect 19567 13271 19625 13277
rect 19702 13268 19708 13320
rect 19760 13308 19766 13320
rect 20088 13317 20116 13348
rect 19980 13311 20038 13317
rect 19760 13280 19805 13308
rect 19760 13268 19766 13280
rect 19980 13277 19992 13311
rect 20026 13277 20038 13311
rect 19980 13271 20038 13277
rect 20073 13311 20131 13317
rect 20073 13277 20085 13311
rect 20119 13308 20131 13311
rect 20254 13308 20260 13320
rect 20119 13280 20260 13308
rect 20119 13277 20131 13280
rect 20073 13271 20131 13277
rect 5166 13240 5172 13252
rect 5000 13212 5172 13240
rect 5166 13200 5172 13212
rect 5224 13200 5230 13252
rect 6730 13200 6736 13252
rect 6788 13240 6794 13252
rect 6788 13212 7236 13240
rect 6788 13200 6794 13212
rect 2590 13172 2596 13184
rect 2551 13144 2596 13172
rect 2590 13132 2596 13144
rect 2648 13132 2654 13184
rect 2774 13132 2780 13184
rect 2832 13172 2838 13184
rect 5258 13172 5264 13184
rect 2832 13144 2877 13172
rect 5219 13144 5264 13172
rect 2832 13132 2838 13144
rect 5258 13132 5264 13144
rect 5316 13132 5322 13184
rect 5353 13175 5411 13181
rect 5353 13141 5365 13175
rect 5399 13172 5411 13175
rect 5442 13172 5448 13184
rect 5399 13144 5448 13172
rect 5399 13141 5411 13144
rect 5353 13135 5411 13141
rect 5442 13132 5448 13144
rect 5500 13132 5506 13184
rect 6825 13175 6883 13181
rect 6825 13141 6837 13175
rect 6871 13172 6883 13175
rect 7098 13172 7104 13184
rect 6871 13144 7104 13172
rect 6871 13141 6883 13144
rect 6825 13135 6883 13141
rect 7098 13132 7104 13144
rect 7156 13132 7162 13184
rect 7208 13172 7236 13212
rect 7742 13200 7748 13252
rect 7800 13240 7806 13252
rect 7800 13212 9260 13240
rect 7800 13200 7806 13212
rect 7377 13175 7435 13181
rect 7377 13172 7389 13175
rect 7208 13144 7389 13172
rect 7377 13141 7389 13144
rect 7423 13172 7435 13175
rect 9122 13172 9128 13184
rect 7423 13144 9128 13172
rect 7423 13141 7435 13144
rect 7377 13135 7435 13141
rect 9122 13132 9128 13144
rect 9180 13132 9186 13184
rect 9232 13181 9260 13212
rect 17310 13200 17316 13252
rect 17368 13240 17374 13252
rect 17865 13243 17923 13249
rect 17865 13240 17877 13243
rect 17368 13212 17877 13240
rect 17368 13200 17374 13212
rect 17865 13209 17877 13212
rect 17911 13209 17923 13243
rect 17865 13203 17923 13209
rect 17957 13243 18015 13249
rect 17957 13209 17969 13243
rect 18003 13240 18015 13243
rect 19797 13243 19855 13249
rect 18003 13212 18644 13240
rect 18003 13209 18015 13212
rect 17957 13203 18015 13209
rect 18616 13184 18644 13212
rect 19797 13209 19809 13243
rect 19843 13209 19855 13243
rect 19995 13240 20023 13271
rect 20254 13268 20260 13280
rect 20312 13268 20318 13320
rect 21266 13308 21272 13320
rect 20456 13280 21272 13308
rect 20456 13240 20484 13280
rect 21266 13268 21272 13280
rect 21324 13268 21330 13320
rect 21634 13308 21640 13320
rect 21595 13280 21640 13308
rect 21634 13268 21640 13280
rect 21692 13268 21698 13320
rect 19995 13212 20484 13240
rect 19797 13203 19855 13209
rect 9217 13175 9275 13181
rect 9217 13141 9229 13175
rect 9263 13141 9275 13175
rect 16206 13172 16212 13184
rect 16167 13144 16212 13172
rect 9217 13135 9275 13141
rect 16206 13132 16212 13144
rect 16264 13132 16270 13184
rect 16945 13175 17003 13181
rect 16945 13141 16957 13175
rect 16991 13172 17003 13175
rect 17034 13172 17040 13184
rect 16991 13144 17040 13172
rect 16991 13141 17003 13144
rect 16945 13135 17003 13141
rect 17034 13132 17040 13144
rect 17092 13132 17098 13184
rect 18598 13132 18604 13184
rect 18656 13132 18662 13184
rect 18785 13175 18843 13181
rect 18785 13141 18797 13175
rect 18831 13172 18843 13175
rect 18966 13172 18972 13184
rect 18831 13144 18972 13172
rect 18831 13141 18843 13144
rect 18785 13135 18843 13141
rect 18966 13132 18972 13144
rect 19024 13172 19030 13184
rect 19812 13172 19840 13203
rect 20530 13200 20536 13252
rect 20588 13240 20594 13252
rect 20717 13243 20775 13249
rect 20588 13212 20633 13240
rect 20588 13200 20594 13212
rect 20717 13209 20729 13243
rect 20763 13240 20775 13243
rect 20763 13212 21496 13240
rect 20763 13209 20775 13212
rect 20717 13203 20775 13209
rect 19024 13144 19840 13172
rect 19024 13132 19030 13144
rect 20254 13132 20260 13184
rect 20312 13172 20318 13184
rect 20732 13172 20760 13203
rect 21468 13181 21496 13212
rect 20312 13144 20760 13172
rect 21453 13175 21511 13181
rect 20312 13132 20318 13144
rect 21453 13141 21465 13175
rect 21499 13141 21511 13175
rect 21453 13135 21511 13141
rect 1104 13082 23987 13104
rect 1104 13030 6630 13082
rect 6682 13030 6694 13082
rect 6746 13030 6758 13082
rect 6810 13030 6822 13082
rect 6874 13030 6886 13082
rect 6938 13030 12311 13082
rect 12363 13030 12375 13082
rect 12427 13030 12439 13082
rect 12491 13030 12503 13082
rect 12555 13030 12567 13082
rect 12619 13030 17992 13082
rect 18044 13030 18056 13082
rect 18108 13030 18120 13082
rect 18172 13030 18184 13082
rect 18236 13030 18248 13082
rect 18300 13030 23673 13082
rect 23725 13030 23737 13082
rect 23789 13030 23801 13082
rect 23853 13030 23865 13082
rect 23917 13030 23929 13082
rect 23981 13030 23987 13082
rect 1104 13008 23987 13030
rect 1854 12928 1860 12980
rect 1912 12968 1918 12980
rect 2317 12971 2375 12977
rect 2317 12968 2329 12971
rect 1912 12940 2329 12968
rect 1912 12928 1918 12940
rect 2317 12937 2329 12940
rect 2363 12937 2375 12971
rect 2317 12931 2375 12937
rect 2590 12928 2596 12980
rect 2648 12968 2654 12980
rect 2648 12940 2728 12968
rect 2648 12928 2654 12940
rect 2498 12860 2504 12912
rect 2556 12900 2562 12912
rect 2556 12872 2636 12900
rect 2556 12860 2562 12872
rect 1578 12832 1584 12844
rect 1539 12804 1584 12832
rect 1578 12792 1584 12804
rect 1636 12792 1642 12844
rect 2608 12841 2636 12872
rect 2700 12841 2728 12940
rect 3234 12928 3240 12980
rect 3292 12968 3298 12980
rect 3513 12971 3571 12977
rect 3513 12968 3525 12971
rect 3292 12940 3525 12968
rect 3292 12928 3298 12940
rect 3513 12937 3525 12940
rect 3559 12937 3571 12971
rect 4522 12968 4528 12980
rect 4483 12940 4528 12968
rect 3513 12931 3571 12937
rect 4522 12928 4528 12940
rect 4580 12928 4586 12980
rect 5537 12971 5595 12977
rect 5537 12937 5549 12971
rect 5583 12968 5595 12971
rect 7834 12968 7840 12980
rect 5583 12940 6960 12968
rect 7795 12940 7840 12968
rect 5583 12937 5595 12940
rect 5537 12931 5595 12937
rect 2958 12860 2964 12912
rect 3016 12900 3022 12912
rect 3881 12903 3939 12909
rect 3881 12900 3893 12903
rect 3016 12872 3893 12900
rect 3016 12860 3022 12872
rect 3881 12869 3893 12872
rect 3927 12869 3939 12903
rect 3881 12863 3939 12869
rect 6454 12860 6460 12912
rect 6512 12900 6518 12912
rect 6730 12900 6736 12912
rect 6512 12872 6736 12900
rect 6512 12860 6518 12872
rect 6730 12860 6736 12872
rect 6788 12860 6794 12912
rect 2593 12835 2651 12841
rect 2593 12801 2605 12835
rect 2639 12801 2651 12835
rect 2593 12795 2651 12801
rect 2685 12835 2743 12841
rect 2685 12801 2697 12835
rect 2731 12801 2743 12835
rect 2685 12795 2743 12801
rect 2777 12835 2835 12841
rect 2777 12801 2789 12835
rect 2823 12832 2835 12835
rect 3142 12832 3148 12844
rect 2823 12804 3148 12832
rect 2823 12801 2835 12804
rect 2777 12795 2835 12801
rect 2501 12767 2559 12773
rect 2501 12733 2513 12767
rect 2547 12733 2559 12767
rect 2700 12764 2728 12795
rect 3142 12792 3148 12804
rect 3200 12792 3206 12844
rect 3602 12792 3608 12844
rect 3660 12832 3666 12844
rect 3697 12835 3755 12841
rect 3697 12832 3709 12835
rect 3660 12804 3709 12832
rect 3660 12792 3666 12804
rect 3697 12801 3709 12804
rect 3743 12801 3755 12835
rect 3697 12795 3755 12801
rect 3786 12792 3792 12844
rect 3844 12832 3850 12844
rect 4062 12832 4068 12844
rect 3844 12804 3889 12832
rect 4023 12804 4068 12832
rect 3844 12792 3850 12804
rect 4062 12792 4068 12804
rect 4120 12792 4126 12844
rect 4706 12792 4712 12844
rect 4764 12832 4770 12844
rect 5077 12835 5135 12841
rect 5077 12832 5089 12835
rect 4764 12804 5089 12832
rect 4764 12792 4770 12804
rect 5077 12801 5089 12804
rect 5123 12801 5135 12835
rect 5077 12795 5135 12801
rect 6270 12792 6276 12844
rect 6328 12832 6334 12844
rect 6932 12841 6960 12940
rect 7834 12928 7840 12940
rect 7892 12968 7898 12980
rect 8018 12968 8024 12980
rect 7892 12940 8024 12968
rect 7892 12928 7898 12940
rect 8018 12928 8024 12940
rect 8076 12928 8082 12980
rect 15654 12928 15660 12980
rect 15712 12968 15718 12980
rect 15933 12971 15991 12977
rect 15933 12968 15945 12971
rect 15712 12940 15945 12968
rect 15712 12928 15718 12940
rect 15933 12937 15945 12940
rect 15979 12937 15991 12971
rect 15933 12931 15991 12937
rect 16482 12928 16488 12980
rect 16540 12968 16546 12980
rect 18233 12971 18291 12977
rect 16540 12940 17264 12968
rect 16540 12928 16546 12940
rect 7098 12860 7104 12912
rect 7156 12900 7162 12912
rect 8570 12900 8576 12912
rect 7156 12872 8576 12900
rect 7156 12860 7162 12872
rect 8570 12860 8576 12872
rect 8628 12860 8634 12912
rect 8757 12903 8815 12909
rect 8757 12869 8769 12903
rect 8803 12900 8815 12903
rect 9122 12900 9128 12912
rect 8803 12872 9128 12900
rect 8803 12869 8815 12872
rect 8757 12863 8815 12869
rect 9122 12860 9128 12872
rect 9180 12900 9186 12912
rect 10042 12900 10048 12912
rect 9180 12872 10048 12900
rect 9180 12860 9186 12872
rect 10042 12860 10048 12872
rect 10100 12860 10106 12912
rect 11330 12860 11336 12912
rect 11388 12900 11394 12912
rect 14369 12903 14427 12909
rect 11388 12872 12940 12900
rect 11388 12860 11394 12872
rect 6825 12835 6883 12841
rect 6825 12832 6837 12835
rect 6328 12804 6837 12832
rect 6328 12792 6334 12804
rect 6825 12801 6837 12804
rect 6871 12801 6883 12835
rect 6825 12795 6883 12801
rect 6917 12835 6975 12841
rect 6917 12801 6929 12835
rect 6963 12832 6975 12835
rect 7558 12832 7564 12844
rect 6963 12804 7564 12832
rect 6963 12801 6975 12804
rect 6917 12795 6975 12801
rect 7558 12792 7564 12804
rect 7616 12792 7622 12844
rect 9582 12832 9588 12844
rect 9543 12804 9588 12832
rect 9582 12792 9588 12804
rect 9640 12832 9646 12844
rect 10229 12835 10287 12841
rect 10229 12832 10241 12835
rect 9640 12804 10241 12832
rect 9640 12792 9646 12804
rect 10229 12801 10241 12804
rect 10275 12801 10287 12835
rect 10229 12795 10287 12801
rect 11698 12792 11704 12844
rect 11756 12832 11762 12844
rect 12912 12841 12940 12872
rect 14369 12869 14381 12903
rect 14415 12900 14427 12903
rect 14550 12900 14556 12912
rect 14415 12872 14556 12900
rect 14415 12869 14427 12872
rect 14369 12863 14427 12869
rect 14550 12860 14556 12872
rect 14608 12860 14614 12912
rect 15746 12900 15752 12912
rect 15120 12872 15752 12900
rect 15120 12841 15148 12872
rect 15746 12860 15752 12872
rect 15804 12860 15810 12912
rect 16301 12903 16359 12909
rect 16301 12869 16313 12903
rect 16347 12900 16359 12903
rect 17129 12903 17187 12909
rect 17129 12900 17141 12903
rect 16347 12872 17141 12900
rect 16347 12869 16359 12872
rect 16301 12863 16359 12869
rect 17129 12869 17141 12872
rect 17175 12869 17187 12903
rect 17236 12900 17264 12940
rect 18233 12937 18245 12971
rect 18279 12968 18291 12971
rect 18414 12968 18420 12980
rect 18279 12940 18420 12968
rect 18279 12937 18291 12940
rect 18233 12931 18291 12937
rect 18414 12928 18420 12940
rect 18472 12928 18478 12980
rect 19153 12971 19211 12977
rect 19153 12937 19165 12971
rect 19199 12968 19211 12971
rect 19334 12968 19340 12980
rect 19199 12940 19340 12968
rect 19199 12937 19211 12940
rect 19153 12931 19211 12937
rect 19334 12928 19340 12940
rect 19392 12928 19398 12980
rect 17339 12903 17397 12909
rect 17339 12900 17351 12903
rect 17236 12872 17351 12900
rect 17129 12863 17187 12869
rect 17339 12869 17351 12872
rect 17385 12869 17397 12903
rect 17339 12863 17397 12869
rect 18432 12872 20944 12900
rect 12529 12835 12587 12841
rect 12529 12832 12541 12835
rect 11756 12804 12541 12832
rect 11756 12792 11762 12804
rect 12529 12801 12541 12804
rect 12575 12801 12587 12835
rect 12529 12795 12587 12801
rect 12897 12835 12955 12841
rect 12897 12801 12909 12835
rect 12943 12801 12955 12835
rect 12897 12795 12955 12801
rect 15105 12835 15163 12841
rect 15105 12801 15117 12835
rect 15151 12801 15163 12835
rect 15286 12832 15292 12844
rect 15247 12804 15292 12832
rect 15105 12795 15163 12801
rect 15286 12792 15292 12804
rect 15344 12832 15350 12844
rect 15562 12832 15568 12844
rect 15344 12804 15568 12832
rect 15344 12792 15350 12804
rect 15562 12792 15568 12804
rect 15620 12792 15626 12844
rect 15841 12835 15899 12841
rect 15841 12801 15853 12835
rect 15887 12801 15899 12835
rect 15841 12795 15899 12801
rect 16117 12835 16175 12841
rect 16117 12801 16129 12835
rect 16163 12832 16175 12835
rect 17034 12832 17040 12844
rect 16163 12804 16528 12832
rect 16995 12804 17040 12832
rect 16163 12801 16175 12804
rect 16117 12795 16175 12801
rect 2700 12736 3464 12764
rect 2501 12727 2559 12733
rect 2516 12696 2544 12727
rect 3142 12696 3148 12708
rect 2516 12668 3148 12696
rect 3142 12656 3148 12668
rect 3200 12656 3206 12708
rect 3436 12696 3464 12736
rect 3510 12724 3516 12776
rect 3568 12764 3574 12776
rect 3804 12764 3832 12792
rect 3568 12736 3832 12764
rect 3568 12724 3574 12736
rect 5718 12724 5724 12776
rect 5776 12764 5782 12776
rect 6362 12764 6368 12776
rect 5776 12736 6368 12764
rect 5776 12724 5782 12736
rect 6362 12724 6368 12736
rect 6420 12764 6426 12776
rect 6641 12767 6699 12773
rect 6641 12764 6653 12767
rect 6420 12736 6653 12764
rect 6420 12724 6426 12736
rect 6641 12733 6653 12736
rect 6687 12733 6699 12767
rect 6641 12727 6699 12733
rect 6730 12724 6736 12776
rect 6788 12764 6794 12776
rect 7098 12764 7104 12776
rect 6788 12736 7104 12764
rect 6788 12724 6794 12736
rect 7098 12724 7104 12736
rect 7156 12764 7162 12776
rect 7742 12764 7748 12776
rect 7156 12736 7748 12764
rect 7156 12724 7162 12736
rect 7742 12724 7748 12736
rect 7800 12724 7806 12776
rect 8386 12724 8392 12776
rect 8444 12764 8450 12776
rect 8662 12764 8668 12776
rect 8444 12736 8668 12764
rect 8444 12724 8450 12736
rect 8662 12724 8668 12736
rect 8720 12764 8726 12776
rect 9217 12767 9275 12773
rect 9217 12764 9229 12767
rect 8720 12736 9229 12764
rect 8720 12724 8726 12736
rect 9217 12733 9229 12736
rect 9263 12733 9275 12767
rect 9217 12727 9275 12733
rect 9306 12724 9312 12776
rect 9364 12764 9370 12776
rect 9493 12767 9551 12773
rect 9493 12764 9505 12767
rect 9364 12736 9505 12764
rect 9364 12724 9370 12736
rect 9493 12733 9505 12736
rect 9539 12733 9551 12767
rect 9493 12727 9551 12733
rect 13814 12724 13820 12776
rect 13872 12764 13878 12776
rect 15013 12767 15071 12773
rect 15013 12764 15025 12767
rect 13872 12736 15025 12764
rect 13872 12724 13878 12736
rect 15013 12733 15025 12736
rect 15059 12733 15071 12767
rect 15013 12727 15071 12733
rect 15197 12767 15255 12773
rect 15197 12733 15209 12767
rect 15243 12764 15255 12767
rect 15654 12764 15660 12776
rect 15243 12736 15660 12764
rect 15243 12733 15255 12736
rect 15197 12727 15255 12733
rect 4154 12696 4160 12708
rect 3436 12668 4160 12696
rect 4154 12656 4160 12668
rect 4212 12656 4218 12708
rect 4522 12656 4528 12708
rect 4580 12696 4586 12708
rect 7834 12696 7840 12708
rect 4580 12668 7840 12696
rect 4580 12656 4586 12668
rect 7834 12656 7840 12668
rect 7892 12656 7898 12708
rect 8754 12656 8760 12708
rect 8812 12696 8818 12708
rect 10689 12699 10747 12705
rect 10689 12696 10701 12699
rect 8812 12668 10701 12696
rect 8812 12656 8818 12668
rect 10689 12665 10701 12668
rect 10735 12665 10747 12699
rect 10689 12659 10747 12665
rect 13354 12656 13360 12708
rect 13412 12696 13418 12708
rect 15028 12696 15056 12727
rect 15654 12724 15660 12736
rect 15712 12724 15718 12776
rect 15856 12696 15884 12795
rect 13412 12668 14964 12696
rect 15028 12668 15884 12696
rect 13412 12656 13418 12668
rect 1765 12631 1823 12637
rect 1765 12597 1777 12631
rect 1811 12628 1823 12631
rect 2130 12628 2136 12640
rect 1811 12600 2136 12628
rect 1811 12597 1823 12600
rect 1765 12591 1823 12597
rect 2130 12588 2136 12600
rect 2188 12588 2194 12640
rect 2498 12588 2504 12640
rect 2556 12628 2562 12640
rect 4338 12628 4344 12640
rect 2556 12600 4344 12628
rect 2556 12588 2562 12600
rect 4338 12588 4344 12600
rect 4396 12588 4402 12640
rect 5350 12628 5356 12640
rect 5311 12600 5356 12628
rect 5350 12588 5356 12600
rect 5408 12588 5414 12640
rect 7101 12631 7159 12637
rect 7101 12597 7113 12631
rect 7147 12628 7159 12631
rect 7466 12628 7472 12640
rect 7147 12600 7472 12628
rect 7147 12597 7159 12600
rect 7101 12591 7159 12597
rect 7466 12588 7472 12600
rect 7524 12588 7530 12640
rect 9306 12588 9312 12640
rect 9364 12628 9370 12640
rect 10321 12631 10379 12637
rect 10321 12628 10333 12631
rect 9364 12600 10333 12628
rect 9364 12588 9370 12600
rect 10321 12597 10333 12600
rect 10367 12597 10379 12631
rect 14826 12628 14832 12640
rect 14787 12600 14832 12628
rect 10321 12591 10379 12597
rect 14826 12588 14832 12600
rect 14884 12588 14890 12640
rect 14936 12628 14964 12668
rect 15746 12628 15752 12640
rect 14936 12600 15752 12628
rect 15746 12588 15752 12600
rect 15804 12588 15810 12640
rect 16390 12588 16396 12640
rect 16448 12628 16454 12640
rect 16500 12628 16528 12804
rect 17034 12792 17040 12804
rect 17092 12792 17098 12844
rect 17218 12832 17224 12844
rect 17179 12804 17224 12832
rect 17218 12792 17224 12804
rect 17276 12832 17282 12844
rect 18230 12832 18236 12844
rect 17276 12804 18236 12832
rect 17276 12792 17282 12804
rect 18230 12792 18236 12804
rect 18288 12792 18294 12844
rect 18432 12841 18460 12872
rect 18417 12835 18475 12841
rect 18417 12801 18429 12835
rect 18463 12801 18475 12835
rect 18598 12832 18604 12844
rect 18559 12804 18604 12832
rect 18417 12795 18475 12801
rect 16853 12767 16911 12773
rect 16853 12733 16865 12767
rect 16899 12764 16911 12767
rect 17126 12764 17132 12776
rect 16899 12736 17132 12764
rect 16899 12733 16911 12736
rect 16853 12727 16911 12733
rect 17126 12724 17132 12736
rect 17184 12724 17190 12776
rect 17497 12767 17555 12773
rect 17497 12764 17509 12767
rect 17236 12736 17509 12764
rect 17236 12708 17264 12736
rect 17497 12733 17509 12736
rect 17543 12733 17555 12767
rect 17497 12727 17555 12733
rect 17678 12724 17684 12776
rect 17736 12764 17742 12776
rect 18432 12764 18460 12795
rect 18598 12792 18604 12804
rect 18656 12792 18662 12844
rect 18693 12835 18751 12841
rect 18693 12801 18705 12835
rect 18739 12832 18751 12835
rect 18966 12832 18972 12844
rect 18739 12804 18972 12832
rect 18739 12801 18751 12804
rect 18693 12795 18751 12801
rect 18966 12792 18972 12804
rect 19024 12792 19030 12844
rect 19334 12832 19340 12844
rect 19295 12804 19340 12832
rect 19334 12792 19340 12804
rect 19392 12792 19398 12844
rect 19521 12835 19579 12841
rect 19521 12801 19533 12835
rect 19567 12832 19579 12835
rect 19610 12832 19616 12844
rect 19567 12804 19616 12832
rect 19567 12801 19579 12804
rect 19521 12795 19579 12801
rect 19610 12792 19616 12804
rect 19668 12792 19674 12844
rect 20162 12792 20168 12844
rect 20220 12832 20226 12844
rect 20533 12835 20591 12841
rect 20533 12832 20545 12835
rect 20220 12804 20545 12832
rect 20220 12792 20226 12804
rect 20533 12801 20545 12804
rect 20579 12801 20591 12835
rect 20533 12795 20591 12801
rect 20625 12835 20683 12841
rect 20625 12801 20637 12835
rect 20671 12801 20683 12835
rect 20806 12832 20812 12844
rect 20767 12804 20812 12832
rect 20625 12795 20683 12801
rect 17736 12736 18460 12764
rect 20640 12764 20668 12795
rect 20806 12792 20812 12804
rect 20864 12792 20870 12844
rect 20916 12841 20944 12872
rect 20901 12835 20959 12841
rect 20901 12801 20913 12835
rect 20947 12801 20959 12835
rect 20901 12795 20959 12801
rect 21361 12767 21419 12773
rect 21361 12764 21373 12767
rect 20640 12736 21373 12764
rect 17736 12724 17742 12736
rect 21361 12733 21373 12736
rect 21407 12764 21419 12767
rect 21407 12736 22094 12764
rect 21407 12733 21419 12736
rect 21361 12727 21419 12733
rect 17218 12656 17224 12708
rect 17276 12656 17282 12708
rect 18966 12656 18972 12708
rect 19024 12696 19030 12708
rect 20530 12696 20536 12708
rect 19024 12668 20536 12696
rect 19024 12656 19030 12668
rect 20530 12656 20536 12668
rect 20588 12656 20594 12708
rect 22066 12640 22094 12736
rect 18874 12628 18880 12640
rect 16448 12600 18880 12628
rect 16448 12588 16454 12600
rect 18874 12588 18880 12600
rect 18932 12588 18938 12640
rect 19426 12588 19432 12640
rect 19484 12628 19490 12640
rect 20349 12631 20407 12637
rect 20349 12628 20361 12631
rect 19484 12600 20361 12628
rect 19484 12588 19490 12600
rect 20349 12597 20361 12600
rect 20395 12597 20407 12631
rect 20349 12591 20407 12597
rect 20806 12588 20812 12640
rect 20864 12628 20870 12640
rect 21726 12628 21732 12640
rect 20864 12600 21732 12628
rect 20864 12588 20870 12600
rect 21726 12588 21732 12600
rect 21784 12588 21790 12640
rect 22066 12628 22100 12640
rect 22055 12600 22100 12628
rect 22094 12588 22100 12600
rect 22152 12588 22158 12640
rect 1104 12538 23828 12560
rect 1104 12486 3790 12538
rect 3842 12486 3854 12538
rect 3906 12486 3918 12538
rect 3970 12486 3982 12538
rect 4034 12486 4046 12538
rect 4098 12486 9471 12538
rect 9523 12486 9535 12538
rect 9587 12486 9599 12538
rect 9651 12486 9663 12538
rect 9715 12486 9727 12538
rect 9779 12486 15152 12538
rect 15204 12486 15216 12538
rect 15268 12486 15280 12538
rect 15332 12486 15344 12538
rect 15396 12486 15408 12538
rect 15460 12486 20833 12538
rect 20885 12486 20897 12538
rect 20949 12486 20961 12538
rect 21013 12486 21025 12538
rect 21077 12486 21089 12538
rect 21141 12486 23828 12538
rect 1104 12464 23828 12486
rect 1946 12384 1952 12436
rect 2004 12424 2010 12436
rect 2869 12427 2927 12433
rect 2869 12424 2881 12427
rect 2004 12396 2881 12424
rect 2004 12384 2010 12396
rect 2869 12393 2881 12396
rect 2915 12393 2927 12427
rect 5718 12424 5724 12436
rect 5679 12396 5724 12424
rect 2869 12387 2927 12393
rect 5718 12384 5724 12396
rect 5776 12384 5782 12436
rect 6178 12424 6184 12436
rect 6139 12396 6184 12424
rect 6178 12384 6184 12396
rect 6236 12384 6242 12436
rect 7834 12384 7840 12436
rect 7892 12384 7898 12436
rect 8202 12384 8208 12436
rect 8260 12424 8266 12436
rect 9125 12427 9183 12433
rect 9125 12424 9137 12427
rect 8260 12396 9137 12424
rect 8260 12384 8266 12396
rect 9125 12393 9137 12396
rect 9171 12393 9183 12427
rect 9125 12387 9183 12393
rect 11238 12384 11244 12436
rect 11296 12424 11302 12436
rect 11333 12427 11391 12433
rect 11333 12424 11345 12427
rect 11296 12396 11345 12424
rect 11296 12384 11302 12396
rect 11333 12393 11345 12396
rect 11379 12424 11391 12427
rect 12066 12424 12072 12436
rect 11379 12396 12072 12424
rect 11379 12393 11391 12396
rect 11333 12387 11391 12393
rect 4525 12359 4583 12365
rect 4525 12325 4537 12359
rect 4571 12356 4583 12359
rect 5166 12356 5172 12368
rect 4571 12328 5172 12356
rect 4571 12325 4583 12328
rect 4525 12319 4583 12325
rect 5166 12316 5172 12328
rect 5224 12316 5230 12368
rect 6086 12316 6092 12368
rect 6144 12356 6150 12368
rect 7285 12359 7343 12365
rect 7285 12356 7297 12359
rect 6144 12328 7297 12356
rect 6144 12316 6150 12328
rect 7285 12325 7297 12328
rect 7331 12325 7343 12359
rect 7285 12319 7343 12325
rect 4249 12291 4307 12297
rect 4249 12257 4261 12291
rect 4295 12288 4307 12291
rect 4706 12288 4712 12300
rect 4295 12260 4712 12288
rect 4295 12257 4307 12260
rect 4249 12251 4307 12257
rect 4706 12248 4712 12260
rect 4764 12248 4770 12300
rect 5350 12288 5356 12300
rect 5263 12260 5356 12288
rect 5350 12248 5356 12260
rect 5408 12288 5414 12300
rect 7190 12288 7196 12300
rect 5408 12260 5672 12288
rect 5408 12248 5414 12260
rect 2222 12220 2228 12232
rect 2183 12192 2228 12220
rect 2222 12180 2228 12192
rect 2280 12180 2286 12232
rect 4157 12223 4215 12229
rect 4157 12189 4169 12223
rect 4203 12220 4215 12223
rect 4338 12220 4344 12232
rect 4203 12192 4344 12220
rect 4203 12189 4215 12192
rect 4157 12183 4215 12189
rect 4338 12180 4344 12192
rect 4396 12180 4402 12232
rect 5166 12180 5172 12232
rect 5224 12220 5230 12232
rect 5261 12223 5319 12229
rect 5261 12220 5273 12223
rect 5224 12192 5273 12220
rect 5224 12180 5230 12192
rect 5261 12189 5273 12192
rect 5307 12189 5319 12223
rect 5442 12220 5448 12232
rect 5403 12192 5448 12220
rect 5261 12183 5319 12189
rect 5442 12180 5448 12192
rect 5500 12180 5506 12232
rect 5537 12223 5595 12229
rect 5537 12189 5549 12223
rect 5583 12189 5595 12223
rect 5537 12183 5595 12189
rect 1762 12112 1768 12164
rect 1820 12152 1826 12164
rect 2777 12155 2835 12161
rect 2777 12152 2789 12155
rect 1820 12124 2789 12152
rect 1820 12112 1826 12124
rect 2777 12121 2789 12124
rect 2823 12121 2835 12155
rect 2777 12115 2835 12121
rect 2038 12084 2044 12096
rect 1999 12056 2044 12084
rect 2038 12044 2044 12056
rect 2096 12044 2102 12096
rect 2590 12044 2596 12096
rect 2648 12084 2654 12096
rect 3050 12084 3056 12096
rect 2648 12056 3056 12084
rect 2648 12044 2654 12056
rect 3050 12044 3056 12056
rect 3108 12044 3114 12096
rect 5442 12044 5448 12096
rect 5500 12084 5506 12096
rect 5552 12084 5580 12183
rect 5500 12056 5580 12084
rect 5644 12084 5672 12260
rect 6472 12260 7196 12288
rect 6382 12233 6440 12239
rect 6382 12199 6394 12233
rect 6428 12230 6440 12233
rect 6472 12230 6500 12260
rect 7190 12248 7196 12260
rect 7248 12248 7254 12300
rect 7852 12288 7880 12384
rect 7929 12291 7987 12297
rect 7929 12288 7941 12291
rect 7300 12260 7788 12288
rect 7852 12260 7941 12288
rect 6428 12202 6500 12230
rect 6428 12199 6440 12202
rect 6382 12193 6440 12199
rect 6822 12180 6828 12232
rect 6880 12220 6886 12232
rect 6880 12192 6925 12220
rect 6880 12180 6886 12192
rect 5994 12112 6000 12164
rect 6052 12152 6058 12164
rect 6457 12155 6515 12161
rect 6457 12152 6469 12155
rect 6052 12124 6469 12152
rect 6052 12112 6058 12124
rect 6457 12121 6469 12124
rect 6503 12121 6515 12155
rect 6457 12115 6515 12121
rect 6546 12112 6552 12164
rect 6604 12152 6610 12164
rect 6687 12155 6745 12161
rect 6604 12124 6649 12152
rect 6604 12112 6610 12124
rect 6687 12121 6699 12155
rect 6733 12152 6745 12155
rect 7300 12152 7328 12260
rect 7760 12254 7788 12260
rect 7929 12257 7941 12260
rect 7975 12257 7987 12291
rect 8478 12288 8484 12300
rect 8439 12260 8484 12288
rect 7466 12220 7472 12232
rect 7427 12192 7472 12220
rect 7466 12180 7472 12192
rect 7524 12180 7530 12232
rect 7760 12226 7814 12254
rect 7929 12251 7987 12257
rect 8478 12248 8484 12260
rect 8536 12248 8542 12300
rect 8570 12248 8576 12300
rect 8628 12288 8634 12300
rect 8628 12260 9352 12288
rect 8628 12248 8634 12260
rect 9324 12229 9352 12260
rect 7558 12152 7564 12164
rect 6733 12124 7328 12152
rect 7519 12124 7564 12152
rect 6733 12121 6745 12124
rect 6687 12115 6745 12121
rect 7558 12112 7564 12124
rect 7616 12112 7622 12164
rect 7786 12161 7814 12226
rect 9309 12223 9367 12229
rect 9309 12189 9321 12223
rect 9355 12189 9367 12223
rect 9766 12220 9772 12232
rect 9727 12192 9772 12220
rect 9309 12183 9367 12189
rect 9766 12180 9772 12192
rect 9824 12180 9830 12232
rect 11808 12229 11836 12396
rect 12066 12384 12072 12396
rect 12124 12384 12130 12436
rect 12710 12384 12716 12436
rect 12768 12424 12774 12436
rect 12768 12396 15884 12424
rect 12768 12384 12774 12396
rect 13541 12359 13599 12365
rect 13541 12325 13553 12359
rect 13587 12356 13599 12359
rect 13630 12356 13636 12368
rect 13587 12328 13636 12356
rect 13587 12325 13599 12328
rect 13541 12319 13599 12325
rect 13630 12316 13636 12328
rect 13688 12316 13694 12368
rect 15856 12356 15884 12396
rect 15930 12384 15936 12436
rect 15988 12424 15994 12436
rect 16301 12427 16359 12433
rect 16301 12424 16313 12427
rect 15988 12396 16313 12424
rect 15988 12384 15994 12396
rect 16301 12393 16313 12396
rect 16347 12393 16359 12427
rect 16301 12387 16359 12393
rect 16574 12384 16580 12436
rect 16632 12424 16638 12436
rect 17402 12424 17408 12436
rect 16632 12396 17408 12424
rect 16632 12384 16638 12396
rect 17402 12384 17408 12396
rect 17460 12384 17466 12436
rect 18233 12427 18291 12433
rect 18233 12393 18245 12427
rect 18279 12424 18291 12427
rect 18322 12424 18328 12436
rect 18279 12396 18328 12424
rect 18279 12393 18291 12396
rect 18233 12387 18291 12393
rect 18322 12384 18328 12396
rect 18380 12384 18386 12436
rect 18966 12424 18972 12436
rect 18432 12396 18972 12424
rect 16666 12356 16672 12368
rect 15856 12328 16672 12356
rect 11885 12291 11943 12297
rect 11885 12257 11897 12291
rect 11931 12288 11943 12291
rect 13814 12288 13820 12300
rect 11931 12260 13820 12288
rect 11931 12257 11943 12260
rect 11885 12251 11943 12257
rect 11793 12223 11851 12229
rect 11793 12189 11805 12223
rect 11839 12189 11851 12223
rect 11793 12183 11851 12189
rect 11977 12223 12035 12229
rect 11977 12189 11989 12223
rect 12023 12220 12035 12223
rect 12066 12220 12072 12232
rect 12023 12192 12072 12220
rect 12023 12189 12035 12192
rect 11977 12183 12035 12189
rect 12066 12180 12072 12192
rect 12124 12180 12130 12232
rect 12636 12229 12664 12260
rect 13814 12248 13820 12260
rect 13872 12248 13878 12300
rect 14461 12291 14519 12297
rect 13924 12260 14412 12288
rect 12621 12223 12679 12229
rect 12621 12189 12633 12223
rect 12667 12189 12679 12223
rect 12621 12183 12679 12189
rect 12710 12180 12716 12232
rect 12768 12220 12774 12232
rect 12894 12220 12900 12232
rect 12768 12192 12813 12220
rect 12855 12192 12900 12220
rect 12768 12180 12774 12192
rect 12894 12180 12900 12192
rect 12952 12180 12958 12232
rect 12989 12223 13047 12229
rect 12989 12189 13001 12223
rect 13035 12220 13047 12223
rect 13078 12220 13084 12232
rect 13035 12192 13084 12220
rect 13035 12189 13047 12192
rect 12989 12183 13047 12189
rect 13078 12180 13084 12192
rect 13136 12220 13142 12232
rect 13924 12220 13952 12260
rect 13136 12192 13952 12220
rect 13136 12180 13142 12192
rect 14274 12180 14280 12232
rect 14332 12180 14338 12232
rect 7653 12155 7711 12161
rect 7653 12121 7665 12155
rect 7699 12121 7711 12155
rect 7786 12155 7849 12161
rect 7786 12124 7803 12155
rect 7653 12115 7711 12121
rect 7791 12121 7803 12124
rect 7837 12152 7849 12155
rect 8202 12152 8208 12164
rect 7837 12124 8208 12152
rect 7837 12121 7849 12124
rect 7791 12115 7849 12121
rect 7006 12084 7012 12096
rect 5644 12056 7012 12084
rect 5500 12044 5506 12056
rect 7006 12044 7012 12056
rect 7064 12044 7070 12096
rect 7190 12044 7196 12096
rect 7248 12084 7254 12096
rect 7668 12084 7696 12115
rect 8202 12112 8208 12124
rect 8260 12112 8266 12164
rect 8570 12112 8576 12164
rect 8628 12152 8634 12164
rect 9674 12161 9680 12164
rect 9401 12155 9459 12161
rect 9401 12152 9413 12155
rect 8628 12124 9413 12152
rect 8628 12112 8634 12124
rect 9401 12121 9413 12124
rect 9447 12121 9459 12155
rect 9401 12115 9459 12121
rect 9493 12155 9551 12161
rect 9493 12121 9505 12155
rect 9539 12121 9551 12155
rect 9631 12155 9680 12161
rect 9631 12152 9643 12155
rect 9587 12124 9643 12152
rect 9493 12115 9551 12121
rect 9631 12121 9643 12124
rect 9677 12121 9680 12155
rect 9631 12115 9680 12121
rect 9508 12084 9536 12115
rect 9674 12112 9680 12115
rect 9732 12112 9738 12164
rect 9858 12084 9864 12096
rect 7248 12056 9864 12084
rect 7248 12044 7254 12056
rect 9858 12044 9864 12056
rect 9916 12044 9922 12096
rect 10042 12044 10048 12096
rect 10100 12084 10106 12096
rect 10321 12087 10379 12093
rect 10321 12084 10333 12087
rect 10100 12056 10333 12084
rect 10100 12044 10106 12056
rect 10321 12053 10333 12056
rect 10367 12084 10379 12087
rect 10594 12084 10600 12096
rect 10367 12056 10600 12084
rect 10367 12053 10379 12056
rect 10321 12047 10379 12053
rect 10594 12044 10600 12056
rect 10652 12044 10658 12096
rect 11790 12044 11796 12096
rect 11848 12084 11854 12096
rect 12066 12084 12072 12096
rect 11848 12056 12072 12084
rect 11848 12044 11854 12056
rect 12066 12044 12072 12056
rect 12124 12044 12130 12096
rect 12437 12087 12495 12093
rect 12437 12053 12449 12087
rect 12483 12084 12495 12087
rect 12802 12084 12808 12096
rect 12483 12056 12808 12084
rect 12483 12053 12495 12056
rect 12437 12047 12495 12053
rect 12802 12044 12808 12056
rect 12860 12044 12866 12096
rect 14292 12093 14320 12180
rect 14384 12152 14412 12260
rect 14461 12257 14473 12291
rect 14507 12288 14519 12291
rect 14507 12260 14780 12288
rect 14507 12257 14519 12260
rect 14461 12251 14519 12257
rect 14550 12180 14556 12232
rect 14608 12220 14614 12232
rect 14752 12220 14780 12260
rect 14826 12248 14832 12300
rect 14884 12288 14890 12300
rect 14921 12291 14979 12297
rect 14921 12288 14933 12291
rect 14884 12260 14933 12288
rect 14884 12248 14890 12260
rect 14921 12257 14933 12260
rect 14967 12257 14979 12291
rect 14921 12251 14979 12257
rect 15562 12220 15568 12232
rect 14608 12192 14653 12220
rect 14752 12192 15568 12220
rect 14608 12180 14614 12192
rect 15562 12180 15568 12192
rect 15620 12180 15626 12232
rect 15654 12180 15660 12232
rect 15712 12220 15718 12232
rect 15856 12229 15884 12328
rect 16666 12316 16672 12328
rect 16724 12316 16730 12368
rect 17310 12316 17316 12368
rect 17368 12356 17374 12368
rect 17681 12359 17739 12365
rect 17681 12356 17693 12359
rect 17368 12328 17693 12356
rect 17368 12316 17374 12328
rect 17681 12325 17693 12328
rect 17727 12325 17739 12359
rect 17681 12319 17739 12325
rect 17862 12288 17868 12300
rect 16408 12260 17868 12288
rect 15841 12223 15899 12229
rect 15712 12192 15757 12220
rect 15712 12180 15718 12192
rect 15841 12189 15853 12223
rect 15887 12189 15899 12223
rect 15841 12183 15899 12189
rect 14829 12155 14887 12161
rect 14829 12152 14841 12155
rect 14384 12124 14841 12152
rect 14829 12121 14841 12124
rect 14875 12121 14887 12155
rect 14829 12115 14887 12121
rect 15749 12155 15807 12161
rect 15749 12121 15761 12155
rect 15795 12152 15807 12155
rect 16408 12152 16436 12260
rect 16776 12229 16804 12260
rect 17862 12248 17868 12260
rect 17920 12288 17926 12300
rect 18432 12288 18460 12396
rect 18966 12384 18972 12396
rect 19024 12384 19030 12436
rect 20162 12424 20168 12436
rect 20123 12396 20168 12424
rect 20162 12384 20168 12396
rect 20220 12384 20226 12436
rect 18874 12356 18880 12368
rect 17920 12260 18460 12288
rect 18616 12328 18880 12356
rect 17920 12248 17926 12260
rect 16485 12223 16543 12229
rect 16485 12189 16497 12223
rect 16531 12189 16543 12223
rect 16485 12183 16543 12189
rect 16761 12223 16819 12229
rect 16761 12189 16773 12223
rect 16807 12189 16819 12223
rect 16761 12183 16819 12189
rect 15795 12124 16436 12152
rect 16500 12152 16528 12183
rect 17218 12180 17224 12232
rect 17276 12220 17282 12232
rect 17405 12223 17463 12229
rect 17405 12220 17417 12223
rect 17276 12192 17417 12220
rect 17276 12180 17282 12192
rect 17405 12189 17417 12192
rect 17451 12189 17463 12223
rect 17405 12183 17463 12189
rect 17497 12223 17555 12229
rect 17497 12189 17509 12223
rect 17543 12220 17555 12223
rect 17586 12220 17592 12232
rect 17543 12192 17592 12220
rect 17543 12189 17555 12192
rect 17497 12183 17555 12189
rect 17586 12180 17592 12192
rect 17644 12180 17650 12232
rect 18414 12220 18420 12232
rect 17773 12201 17831 12207
rect 17773 12167 17785 12201
rect 17819 12167 17831 12201
rect 18375 12192 18420 12220
rect 18414 12180 18420 12192
rect 18472 12180 18478 12232
rect 18616 12229 18644 12328
rect 18874 12316 18880 12328
rect 18932 12316 18938 12368
rect 18601 12223 18659 12229
rect 18601 12189 18613 12223
rect 18647 12189 18659 12223
rect 18601 12183 18659 12189
rect 18877 12223 18935 12229
rect 18877 12189 18889 12223
rect 18923 12220 18935 12223
rect 19426 12220 19432 12232
rect 18923 12192 19432 12220
rect 18923 12189 18935 12192
rect 18877 12183 18935 12189
rect 19426 12180 19432 12192
rect 19484 12180 19490 12232
rect 19886 12220 19892 12232
rect 19847 12192 19892 12220
rect 19886 12180 19892 12192
rect 19944 12180 19950 12232
rect 19981 12223 20039 12229
rect 19981 12189 19993 12223
rect 20027 12220 20039 12223
rect 20070 12220 20076 12232
rect 20027 12192 20076 12220
rect 20027 12189 20039 12192
rect 19981 12183 20039 12189
rect 20070 12180 20076 12192
rect 20128 12180 20134 12232
rect 21082 12180 21088 12232
rect 21140 12220 21146 12232
rect 21634 12220 21640 12232
rect 21140 12192 21640 12220
rect 21140 12180 21146 12192
rect 21634 12180 21640 12192
rect 21692 12220 21698 12232
rect 21729 12223 21787 12229
rect 21729 12220 21741 12223
rect 21692 12192 21741 12220
rect 21692 12180 21698 12192
rect 21729 12189 21741 12192
rect 21775 12189 21787 12223
rect 21729 12183 21787 12189
rect 16942 12152 16948 12164
rect 16500 12124 16948 12152
rect 15795 12121 15807 12124
rect 15749 12115 15807 12121
rect 16942 12112 16948 12124
rect 17000 12112 17006 12164
rect 17773 12161 17831 12167
rect 14277 12087 14335 12093
rect 14277 12053 14289 12087
rect 14323 12053 14335 12087
rect 14277 12047 14335 12053
rect 15378 12044 15384 12096
rect 15436 12084 15442 12096
rect 16390 12084 16396 12096
rect 15436 12056 16396 12084
rect 15436 12044 15442 12056
rect 16390 12044 16396 12056
rect 16448 12044 16454 12096
rect 16669 12087 16727 12093
rect 16669 12053 16681 12087
rect 16715 12084 16727 12087
rect 16850 12084 16856 12096
rect 16715 12056 16856 12084
rect 16715 12053 16727 12056
rect 16669 12047 16727 12053
rect 16850 12044 16856 12056
rect 16908 12044 16914 12096
rect 17402 12084 17408 12096
rect 17363 12056 17408 12084
rect 17402 12044 17408 12056
rect 17460 12044 17466 12096
rect 17494 12044 17500 12096
rect 17552 12084 17558 12096
rect 17788 12084 17816 12161
rect 17862 12112 17868 12164
rect 17920 12152 17926 12164
rect 18509 12155 18567 12161
rect 18509 12152 18521 12155
rect 17920 12124 18521 12152
rect 17920 12112 17926 12124
rect 18509 12121 18521 12124
rect 18555 12121 18567 12155
rect 18509 12115 18567 12121
rect 18739 12155 18797 12161
rect 18739 12121 18751 12155
rect 18785 12152 18797 12155
rect 20714 12152 20720 12164
rect 18785 12124 20720 12152
rect 18785 12121 18797 12124
rect 18739 12115 18797 12121
rect 20714 12112 20720 12124
rect 20772 12112 20778 12164
rect 21174 12152 21180 12164
rect 21135 12124 21180 12152
rect 21174 12112 21180 12124
rect 21232 12112 21238 12164
rect 22094 12152 22100 12164
rect 21284 12124 22100 12152
rect 21085 12087 21143 12093
rect 21085 12084 21097 12087
rect 17552 12056 21097 12084
rect 17552 12044 17558 12056
rect 21085 12053 21097 12056
rect 21131 12084 21143 12087
rect 21284 12084 21312 12124
rect 22094 12112 22100 12124
rect 22152 12152 22158 12164
rect 23106 12152 23112 12164
rect 22152 12124 23112 12152
rect 22152 12112 22158 12124
rect 23106 12112 23112 12124
rect 23164 12112 23170 12164
rect 21131 12056 21312 12084
rect 21131 12053 21143 12056
rect 21085 12047 21143 12053
rect 21358 12044 21364 12096
rect 21416 12084 21422 12096
rect 21821 12087 21879 12093
rect 21821 12084 21833 12087
rect 21416 12056 21833 12084
rect 21416 12044 21422 12056
rect 21821 12053 21833 12056
rect 21867 12053 21879 12087
rect 21821 12047 21879 12053
rect 22465 12087 22523 12093
rect 22465 12053 22477 12087
rect 22511 12084 22523 12087
rect 22554 12084 22560 12096
rect 22511 12056 22560 12084
rect 22511 12053 22523 12056
rect 22465 12047 22523 12053
rect 22554 12044 22560 12056
rect 22612 12044 22618 12096
rect 1104 11994 23987 12016
rect 1104 11942 6630 11994
rect 6682 11942 6694 11994
rect 6746 11942 6758 11994
rect 6810 11942 6822 11994
rect 6874 11942 6886 11994
rect 6938 11942 12311 11994
rect 12363 11942 12375 11994
rect 12427 11942 12439 11994
rect 12491 11942 12503 11994
rect 12555 11942 12567 11994
rect 12619 11942 17992 11994
rect 18044 11942 18056 11994
rect 18108 11942 18120 11994
rect 18172 11942 18184 11994
rect 18236 11942 18248 11994
rect 18300 11942 23673 11994
rect 23725 11942 23737 11994
rect 23789 11942 23801 11994
rect 23853 11942 23865 11994
rect 23917 11942 23929 11994
rect 23981 11942 23987 11994
rect 1104 11920 23987 11942
rect 2958 11880 2964 11892
rect 2919 11852 2964 11880
rect 2958 11840 2964 11852
rect 3016 11840 3022 11892
rect 4157 11883 4215 11889
rect 4157 11849 4169 11883
rect 4203 11880 4215 11883
rect 4246 11880 4252 11892
rect 4203 11852 4252 11880
rect 4203 11849 4215 11852
rect 4157 11843 4215 11849
rect 4246 11840 4252 11852
rect 4304 11840 4310 11892
rect 4706 11880 4712 11892
rect 4667 11852 4712 11880
rect 4706 11840 4712 11852
rect 4764 11840 4770 11892
rect 5350 11840 5356 11892
rect 5408 11880 5414 11892
rect 5537 11883 5595 11889
rect 5537 11880 5549 11883
rect 5408 11852 5549 11880
rect 5408 11840 5414 11852
rect 5537 11849 5549 11852
rect 5583 11849 5595 11883
rect 5994 11880 6000 11892
rect 5955 11852 6000 11880
rect 5537 11843 5595 11849
rect 5994 11840 6000 11852
rect 6052 11840 6058 11892
rect 7190 11880 7196 11892
rect 6748 11852 7196 11880
rect 2133 11815 2191 11821
rect 2133 11781 2145 11815
rect 2179 11812 2191 11815
rect 3234 11812 3240 11824
rect 2179 11784 3240 11812
rect 2179 11781 2191 11784
rect 2133 11775 2191 11781
rect 3234 11772 3240 11784
rect 3292 11812 3298 11824
rect 4724 11812 4752 11840
rect 3292 11784 3464 11812
rect 3292 11772 3298 11784
rect 2038 11744 2044 11756
rect 1951 11716 2044 11744
rect 2038 11704 2044 11716
rect 2096 11744 2102 11756
rect 2225 11747 2283 11753
rect 2096 11716 2176 11744
rect 2096 11704 2102 11716
rect 2148 11540 2176 11716
rect 2225 11713 2237 11747
rect 2271 11744 2283 11747
rect 2590 11744 2596 11756
rect 2271 11716 2596 11744
rect 2271 11713 2283 11716
rect 2225 11707 2283 11713
rect 2590 11704 2596 11716
rect 2648 11704 2654 11756
rect 3436 11753 3464 11784
rect 3620 11784 4752 11812
rect 3620 11753 3648 11784
rect 2685 11747 2743 11753
rect 2685 11713 2697 11747
rect 2731 11713 2743 11747
rect 3421 11747 3479 11753
rect 2685 11707 2743 11713
rect 2884 11716 3188 11744
rect 2700 11676 2728 11707
rect 2884 11688 2912 11716
rect 2866 11676 2872 11688
rect 2700 11648 2872 11676
rect 2866 11636 2872 11648
rect 2924 11636 2930 11688
rect 2958 11636 2964 11688
rect 3016 11676 3022 11688
rect 3160 11676 3188 11716
rect 3421 11713 3433 11747
rect 3467 11713 3479 11747
rect 3421 11707 3479 11713
rect 3513 11747 3571 11753
rect 3513 11713 3525 11747
rect 3559 11713 3571 11747
rect 3513 11707 3571 11713
rect 3605 11747 3663 11753
rect 3605 11713 3617 11747
rect 3651 11713 3663 11747
rect 3605 11707 3663 11713
rect 3528 11676 3556 11707
rect 4154 11704 4160 11756
rect 4212 11744 4218 11756
rect 4617 11747 4675 11753
rect 4617 11744 4629 11747
rect 4212 11716 4629 11744
rect 4212 11704 4218 11716
rect 4617 11713 4629 11716
rect 4663 11713 4675 11747
rect 4798 11744 4804 11756
rect 4759 11716 4804 11744
rect 4617 11707 4675 11713
rect 3016 11648 3061 11676
rect 3160 11648 3556 11676
rect 4632 11676 4660 11707
rect 4798 11704 4804 11716
rect 4856 11704 4862 11756
rect 5368 11744 5396 11840
rect 5626 11744 5632 11756
rect 4908 11716 5396 11744
rect 5587 11716 5632 11744
rect 4908 11676 4936 11716
rect 5626 11704 5632 11716
rect 5684 11744 5690 11756
rect 6748 11753 6776 11852
rect 7190 11840 7196 11852
rect 7248 11840 7254 11892
rect 7926 11840 7932 11892
rect 7984 11880 7990 11892
rect 7984 11852 8029 11880
rect 7984 11840 7990 11852
rect 8110 11840 8116 11892
rect 8168 11880 8174 11892
rect 8168 11852 8248 11880
rect 8168 11840 8174 11852
rect 8220 11821 8248 11852
rect 8294 11840 8300 11892
rect 8352 11880 8358 11892
rect 8352 11852 10180 11880
rect 8352 11840 8358 11852
rect 8205 11815 8263 11821
rect 8205 11781 8217 11815
rect 8251 11781 8263 11815
rect 8205 11775 8263 11781
rect 9030 11772 9036 11824
rect 9088 11812 9094 11824
rect 9088 11784 9628 11812
rect 9088 11772 9094 11784
rect 6549 11747 6607 11753
rect 6549 11744 6561 11747
rect 5684 11716 6561 11744
rect 5684 11704 5690 11716
rect 6549 11713 6561 11716
rect 6595 11713 6607 11747
rect 6549 11707 6607 11713
rect 6733 11747 6791 11753
rect 6733 11713 6745 11747
rect 6779 11713 6791 11747
rect 6733 11707 6791 11713
rect 6825 11747 6883 11753
rect 6825 11713 6837 11747
rect 6871 11713 6883 11747
rect 6825 11707 6883 11713
rect 6917 11747 6975 11753
rect 6917 11713 6929 11747
rect 6963 11744 6975 11747
rect 7098 11744 7104 11756
rect 6963 11716 7104 11744
rect 6963 11713 6975 11716
rect 6917 11707 6975 11713
rect 5442 11676 5448 11688
rect 4632 11648 4936 11676
rect 5403 11648 5448 11676
rect 3016 11636 3022 11648
rect 5442 11636 5448 11648
rect 5500 11636 5506 11688
rect 6178 11636 6184 11688
rect 6236 11676 6242 11688
rect 6840 11676 6868 11707
rect 7098 11704 7104 11716
rect 7156 11744 7162 11756
rect 7742 11744 7748 11756
rect 7156 11716 7748 11744
rect 7156 11704 7162 11716
rect 7742 11704 7748 11716
rect 7800 11704 7806 11756
rect 8110 11744 8116 11756
rect 8071 11716 8116 11744
rect 8110 11704 8116 11716
rect 8168 11704 8174 11756
rect 8294 11744 8300 11756
rect 8255 11716 8300 11744
rect 8294 11704 8300 11716
rect 8352 11704 8358 11756
rect 8481 11747 8539 11753
rect 8481 11713 8493 11747
rect 8527 11713 8539 11747
rect 8481 11707 8539 11713
rect 6236 11648 6868 11676
rect 7193 11679 7251 11685
rect 6236 11636 6242 11648
rect 7193 11645 7205 11679
rect 7239 11676 7251 11679
rect 8496 11676 8524 11707
rect 9306 11704 9312 11756
rect 9364 11744 9370 11756
rect 9600 11753 9628 11784
rect 10152 11753 10180 11852
rect 10962 11840 10968 11892
rect 11020 11880 11026 11892
rect 11701 11883 11759 11889
rect 11701 11880 11713 11883
rect 11020 11852 11713 11880
rect 11020 11840 11026 11852
rect 11701 11849 11713 11852
rect 11747 11849 11759 11883
rect 11701 11843 11759 11849
rect 13633 11883 13691 11889
rect 13633 11849 13645 11883
rect 13679 11880 13691 11883
rect 13906 11880 13912 11892
rect 13679 11852 13912 11880
rect 13679 11849 13691 11852
rect 13633 11843 13691 11849
rect 13906 11840 13912 11852
rect 13964 11840 13970 11892
rect 15470 11880 15476 11892
rect 15431 11852 15476 11880
rect 15470 11840 15476 11852
rect 15528 11840 15534 11892
rect 16117 11883 16175 11889
rect 16117 11849 16129 11883
rect 16163 11880 16175 11883
rect 16206 11880 16212 11892
rect 16163 11852 16212 11880
rect 16163 11849 16175 11852
rect 16117 11843 16175 11849
rect 16206 11840 16212 11852
rect 16264 11840 16270 11892
rect 16298 11840 16304 11892
rect 16356 11880 16362 11892
rect 16853 11883 16911 11889
rect 16853 11880 16865 11883
rect 16356 11852 16865 11880
rect 16356 11840 16362 11852
rect 16853 11849 16865 11852
rect 16899 11849 16911 11883
rect 17310 11880 17316 11892
rect 16853 11843 16911 11849
rect 17052 11852 17316 11880
rect 11149 11815 11207 11821
rect 11149 11781 11161 11815
rect 11195 11812 11207 11815
rect 11422 11812 11428 11824
rect 11195 11784 11428 11812
rect 11195 11781 11207 11784
rect 11149 11775 11207 11781
rect 9493 11747 9551 11753
rect 9493 11744 9505 11747
rect 9364 11716 9505 11744
rect 9364 11704 9370 11716
rect 9493 11713 9505 11716
rect 9539 11713 9551 11747
rect 9493 11707 9551 11713
rect 9585 11747 9643 11753
rect 9585 11713 9597 11747
rect 9631 11713 9643 11747
rect 9585 11707 9643 11713
rect 10137 11747 10195 11753
rect 10137 11713 10149 11747
rect 10183 11713 10195 11747
rect 10137 11707 10195 11713
rect 10962 11704 10968 11756
rect 11020 11744 11026 11756
rect 11164 11744 11192 11775
rect 11422 11772 11428 11784
rect 11480 11772 11486 11824
rect 12069 11815 12127 11821
rect 12069 11781 12081 11815
rect 12115 11812 12127 11815
rect 13262 11812 13268 11824
rect 12115 11784 13268 11812
rect 12115 11781 12127 11784
rect 12069 11775 12127 11781
rect 13262 11772 13268 11784
rect 13320 11772 13326 11824
rect 14090 11772 14096 11824
rect 14148 11812 14154 11824
rect 16942 11812 16948 11824
rect 14148 11784 16948 11812
rect 14148 11772 14154 11784
rect 11882 11744 11888 11756
rect 11020 11716 11192 11744
rect 11843 11716 11888 11744
rect 11020 11704 11026 11716
rect 11882 11704 11888 11716
rect 11940 11704 11946 11756
rect 11977 11747 12035 11753
rect 11977 11713 11989 11747
rect 12023 11744 12035 11747
rect 12158 11744 12164 11756
rect 12023 11716 12164 11744
rect 12023 11713 12035 11716
rect 11977 11707 12035 11713
rect 12158 11704 12164 11716
rect 12216 11704 12222 11756
rect 12253 11747 12311 11753
rect 12253 11713 12265 11747
rect 12299 11744 12311 11747
rect 12713 11747 12771 11753
rect 12713 11744 12725 11747
rect 12299 11716 12725 11744
rect 12299 11713 12311 11716
rect 12253 11707 12311 11713
rect 12713 11713 12725 11716
rect 12759 11713 12771 11747
rect 12713 11707 12771 11713
rect 12894 11704 12900 11756
rect 12952 11744 12958 11756
rect 13630 11744 13636 11756
rect 12952 11716 13636 11744
rect 12952 11704 12958 11716
rect 13630 11704 13636 11716
rect 13688 11704 13694 11756
rect 14001 11747 14059 11753
rect 14001 11713 14013 11747
rect 14047 11744 14059 11747
rect 14366 11744 14372 11756
rect 14047 11716 14372 11744
rect 14047 11713 14059 11716
rect 14001 11707 14059 11713
rect 14366 11704 14372 11716
rect 14424 11704 14430 11756
rect 14550 11704 14556 11756
rect 14608 11744 14614 11756
rect 14645 11747 14703 11753
rect 14645 11744 14657 11747
rect 14608 11716 14657 11744
rect 14608 11704 14614 11716
rect 14645 11713 14657 11716
rect 14691 11744 14703 11747
rect 15378 11744 15384 11756
rect 14691 11716 14964 11744
rect 15339 11716 15384 11744
rect 14691 11713 14703 11716
rect 14645 11707 14703 11713
rect 10413 11679 10471 11685
rect 7239 11648 8524 11676
rect 9692 11648 10364 11676
rect 7239 11645 7251 11648
rect 7193 11639 7251 11645
rect 9692 11620 9720 11648
rect 2774 11568 2780 11620
rect 2832 11608 2838 11620
rect 2832 11580 2877 11608
rect 2832 11568 2838 11580
rect 5166 11568 5172 11620
rect 5224 11608 5230 11620
rect 7282 11608 7288 11620
rect 5224 11580 7288 11608
rect 5224 11568 5230 11580
rect 7282 11568 7288 11580
rect 7340 11568 7346 11620
rect 8110 11568 8116 11620
rect 8168 11608 8174 11620
rect 9674 11608 9680 11620
rect 8168 11580 9680 11608
rect 8168 11568 8174 11580
rect 9674 11568 9680 11580
rect 9732 11568 9738 11620
rect 10226 11608 10232 11620
rect 10187 11580 10232 11608
rect 10226 11568 10232 11580
rect 10284 11568 10290 11620
rect 10336 11608 10364 11648
rect 10413 11645 10425 11679
rect 10459 11676 10471 11679
rect 10594 11676 10600 11688
rect 10459 11648 10600 11676
rect 10459 11645 10471 11648
rect 10413 11639 10471 11645
rect 10594 11636 10600 11648
rect 10652 11636 10658 11688
rect 13173 11679 13231 11685
rect 13173 11645 13185 11679
rect 13219 11645 13231 11679
rect 13173 11639 13231 11645
rect 13909 11679 13967 11685
rect 13909 11645 13921 11679
rect 13955 11676 13967 11679
rect 14274 11676 14280 11688
rect 13955 11648 14280 11676
rect 13955 11645 13967 11648
rect 13909 11639 13967 11645
rect 10778 11608 10784 11620
rect 10336 11580 10784 11608
rect 10778 11568 10784 11580
rect 10836 11568 10842 11620
rect 13188 11608 13216 11639
rect 14274 11636 14280 11648
rect 14332 11636 14338 11688
rect 14826 11676 14832 11688
rect 14787 11648 14832 11676
rect 14826 11636 14832 11648
rect 14884 11636 14890 11688
rect 14936 11676 14964 11716
rect 15378 11704 15384 11716
rect 15436 11704 15442 11756
rect 15562 11704 15568 11756
rect 15620 11744 15626 11756
rect 15856 11753 15884 11784
rect 16942 11772 16948 11784
rect 17000 11772 17006 11824
rect 17052 11753 17080 11852
rect 17310 11840 17316 11852
rect 17368 11840 17374 11892
rect 17954 11880 17960 11892
rect 17867 11852 17960 11880
rect 17954 11840 17960 11852
rect 18012 11880 18018 11892
rect 18322 11880 18328 11892
rect 18012 11852 18328 11880
rect 18012 11840 18018 11852
rect 18322 11840 18328 11852
rect 18380 11840 18386 11892
rect 18417 11883 18475 11889
rect 18417 11849 18429 11883
rect 18463 11880 18475 11883
rect 18506 11880 18512 11892
rect 18463 11852 18512 11880
rect 18463 11849 18475 11852
rect 18417 11843 18475 11849
rect 18506 11840 18512 11852
rect 18564 11840 18570 11892
rect 17494 11812 17500 11824
rect 17236 11784 17500 11812
rect 17236 11753 17264 11784
rect 17494 11772 17500 11784
rect 17552 11772 17558 11824
rect 18340 11812 18368 11840
rect 19058 11812 19064 11824
rect 18340 11784 19064 11812
rect 19058 11772 19064 11784
rect 19116 11772 19122 11824
rect 19521 11815 19579 11821
rect 19521 11781 19533 11815
rect 19567 11812 19579 11815
rect 20070 11812 20076 11824
rect 19567 11784 20076 11812
rect 19567 11781 19579 11784
rect 19521 11775 19579 11781
rect 20070 11772 20076 11784
rect 20128 11772 20134 11824
rect 20162 11772 20168 11824
rect 20220 11812 20226 11824
rect 21818 11812 21824 11824
rect 20220 11784 21824 11812
rect 20220 11772 20226 11784
rect 21818 11772 21824 11784
rect 21876 11812 21882 11824
rect 21876 11784 22048 11812
rect 21876 11772 21882 11784
rect 15749 11747 15807 11753
rect 15749 11744 15761 11747
rect 15620 11716 15761 11744
rect 15620 11704 15626 11716
rect 15749 11713 15761 11716
rect 15795 11713 15807 11747
rect 15749 11707 15807 11713
rect 15841 11747 15899 11753
rect 15841 11713 15853 11747
rect 15887 11713 15899 11747
rect 15841 11707 15899 11713
rect 17037 11747 17095 11753
rect 17037 11713 17049 11747
rect 17083 11713 17095 11747
rect 17037 11707 17095 11713
rect 17221 11747 17279 11753
rect 17221 11713 17233 11747
rect 17267 11713 17279 11747
rect 17221 11707 17279 11713
rect 17402 11704 17408 11756
rect 17460 11744 17466 11756
rect 18785 11747 18843 11753
rect 18785 11744 18797 11747
rect 17460 11716 18797 11744
rect 17460 11704 17466 11716
rect 18785 11713 18797 11716
rect 18831 11713 18843 11747
rect 20254 11744 20260 11756
rect 20167 11716 20260 11744
rect 18785 11707 18843 11713
rect 20180 11688 20208 11716
rect 20254 11704 20260 11716
rect 20312 11704 20318 11756
rect 20438 11704 20444 11756
rect 20496 11744 20502 11756
rect 20533 11747 20591 11753
rect 20533 11744 20545 11747
rect 20496 11716 20545 11744
rect 20496 11704 20502 11716
rect 20533 11713 20545 11716
rect 20579 11713 20591 11747
rect 20533 11707 20591 11713
rect 20717 11747 20775 11753
rect 20717 11713 20729 11747
rect 20763 11713 20775 11747
rect 21174 11744 21180 11756
rect 21087 11716 21180 11744
rect 20717 11707 20775 11713
rect 15657 11679 15715 11685
rect 15657 11676 15669 11679
rect 14936 11648 15669 11676
rect 15657 11645 15669 11648
rect 15703 11676 15715 11679
rect 16942 11676 16948 11688
rect 15703 11648 16948 11676
rect 15703 11645 15715 11648
rect 15657 11639 15715 11645
rect 16942 11636 16948 11648
rect 17000 11636 17006 11688
rect 17126 11676 17132 11688
rect 17087 11648 17132 11676
rect 17126 11636 17132 11648
rect 17184 11636 17190 11688
rect 17313 11679 17371 11685
rect 17313 11645 17325 11679
rect 17359 11645 17371 11679
rect 18598 11676 18604 11688
rect 18559 11648 18604 11676
rect 17313 11639 17371 11645
rect 13446 11608 13452 11620
rect 13188 11580 13452 11608
rect 13446 11568 13452 11580
rect 13504 11608 13510 11620
rect 14461 11611 14519 11617
rect 13504 11580 14044 11608
rect 13504 11568 13510 11580
rect 14016 11552 14044 11580
rect 14461 11577 14473 11611
rect 14507 11608 14519 11611
rect 15010 11608 15016 11620
rect 14507 11580 15016 11608
rect 14507 11577 14519 11580
rect 14461 11571 14519 11577
rect 15010 11568 15016 11580
rect 15068 11568 15074 11620
rect 16022 11568 16028 11620
rect 16080 11608 16086 11620
rect 17328 11608 17356 11639
rect 18598 11636 18604 11648
rect 18656 11636 18662 11688
rect 18693 11679 18751 11685
rect 18693 11645 18705 11679
rect 18739 11645 18751 11679
rect 18693 11639 18751 11645
rect 18877 11679 18935 11685
rect 18877 11645 18889 11679
rect 18923 11676 18935 11679
rect 20073 11679 20131 11685
rect 20073 11676 20085 11679
rect 18923 11648 20085 11676
rect 18923 11645 18935 11648
rect 18877 11639 18935 11645
rect 20073 11645 20085 11648
rect 20119 11645 20131 11679
rect 20073 11639 20131 11645
rect 17678 11608 17684 11620
rect 16080 11580 17684 11608
rect 16080 11568 16086 11580
rect 17678 11568 17684 11580
rect 17736 11608 17742 11620
rect 18322 11608 18328 11620
rect 17736 11580 18328 11608
rect 17736 11568 17742 11580
rect 18322 11568 18328 11580
rect 18380 11568 18386 11620
rect 18708 11608 18736 11639
rect 20162 11636 20168 11688
rect 20220 11636 20226 11688
rect 20732 11676 20760 11707
rect 21174 11704 21180 11716
rect 21232 11744 21238 11756
rect 21634 11744 21640 11756
rect 21232 11716 21640 11744
rect 21232 11704 21238 11716
rect 21634 11704 21640 11716
rect 21692 11704 21698 11756
rect 22020 11753 22048 11784
rect 22005 11747 22063 11753
rect 22005 11713 22017 11747
rect 22051 11713 22063 11747
rect 22005 11707 22063 11713
rect 22097 11747 22155 11753
rect 22097 11713 22109 11747
rect 22143 11713 22155 11747
rect 22097 11707 22155 11713
rect 21910 11676 21916 11688
rect 20732 11648 21916 11676
rect 21910 11636 21916 11648
rect 21968 11636 21974 11688
rect 19242 11608 19248 11620
rect 18708 11580 19248 11608
rect 19242 11568 19248 11580
rect 19300 11568 19306 11620
rect 19610 11568 19616 11620
rect 19668 11608 19674 11620
rect 20349 11611 20407 11617
rect 20349 11608 20361 11611
rect 19668 11580 20361 11608
rect 19668 11568 19674 11580
rect 20349 11577 20361 11580
rect 20395 11577 20407 11611
rect 20349 11571 20407 11577
rect 20438 11568 20444 11620
rect 20496 11608 20502 11620
rect 20496 11580 20541 11608
rect 20496 11568 20502 11580
rect 3602 11540 3608 11552
rect 2148 11512 3608 11540
rect 3602 11500 3608 11512
rect 3660 11500 3666 11552
rect 7558 11500 7564 11552
rect 7616 11540 7622 11552
rect 7834 11540 7840 11552
rect 7616 11512 7840 11540
rect 7616 11500 7622 11512
rect 7834 11500 7840 11512
rect 7892 11500 7898 11552
rect 8386 11500 8392 11552
rect 8444 11540 8450 11552
rect 9309 11543 9367 11549
rect 9309 11540 9321 11543
rect 8444 11512 9321 11540
rect 8444 11500 8450 11512
rect 9309 11509 9321 11512
rect 9355 11509 9367 11543
rect 10318 11540 10324 11552
rect 10279 11512 10324 11540
rect 9309 11503 9367 11509
rect 10318 11500 10324 11512
rect 10376 11500 10382 11552
rect 13078 11540 13084 11552
rect 13039 11512 13084 11540
rect 13078 11500 13084 11512
rect 13136 11500 13142 11552
rect 13998 11540 14004 11552
rect 13959 11512 14004 11540
rect 13998 11500 14004 11512
rect 14056 11500 14062 11552
rect 16666 11500 16672 11552
rect 16724 11540 16730 11552
rect 17402 11540 17408 11552
rect 16724 11512 17408 11540
rect 16724 11500 16730 11512
rect 17402 11500 17408 11512
rect 17460 11500 17466 11552
rect 21361 11543 21419 11549
rect 21361 11509 21373 11543
rect 21407 11540 21419 11543
rect 22002 11540 22008 11552
rect 21407 11512 22008 11540
rect 21407 11509 21419 11512
rect 21361 11503 21419 11509
rect 22002 11500 22008 11512
rect 22060 11540 22066 11552
rect 22112 11540 22140 11707
rect 22186 11704 22192 11756
rect 22244 11744 22250 11756
rect 22281 11747 22339 11753
rect 22281 11744 22293 11747
rect 22244 11716 22293 11744
rect 22244 11704 22250 11716
rect 22281 11713 22293 11716
rect 22327 11744 22339 11747
rect 22554 11744 22560 11756
rect 22327 11716 22560 11744
rect 22327 11713 22339 11716
rect 22281 11707 22339 11713
rect 22554 11704 22560 11716
rect 22612 11704 22618 11756
rect 22060 11512 22140 11540
rect 22060 11500 22066 11512
rect 22186 11500 22192 11552
rect 22244 11540 22250 11552
rect 22465 11543 22523 11549
rect 22465 11540 22477 11543
rect 22244 11512 22477 11540
rect 22244 11500 22250 11512
rect 22465 11509 22477 11512
rect 22511 11509 22523 11543
rect 22465 11503 22523 11509
rect 23017 11543 23075 11549
rect 23017 11509 23029 11543
rect 23063 11540 23075 11543
rect 23106 11540 23112 11552
rect 23063 11512 23112 11540
rect 23063 11509 23075 11512
rect 23017 11503 23075 11509
rect 23106 11500 23112 11512
rect 23164 11500 23170 11552
rect 1104 11450 23828 11472
rect 1104 11398 3790 11450
rect 3842 11398 3854 11450
rect 3906 11398 3918 11450
rect 3970 11398 3982 11450
rect 4034 11398 4046 11450
rect 4098 11398 9471 11450
rect 9523 11398 9535 11450
rect 9587 11398 9599 11450
rect 9651 11398 9663 11450
rect 9715 11398 9727 11450
rect 9779 11398 15152 11450
rect 15204 11398 15216 11450
rect 15268 11398 15280 11450
rect 15332 11398 15344 11450
rect 15396 11398 15408 11450
rect 15460 11398 20833 11450
rect 20885 11398 20897 11450
rect 20949 11398 20961 11450
rect 21013 11398 21025 11450
rect 21077 11398 21089 11450
rect 21141 11398 23828 11450
rect 1104 11376 23828 11398
rect 1578 11296 1584 11348
rect 1636 11336 1642 11348
rect 2225 11339 2283 11345
rect 2225 11336 2237 11339
rect 1636 11308 2237 11336
rect 1636 11296 1642 11308
rect 2225 11305 2237 11308
rect 2271 11305 2283 11339
rect 2225 11299 2283 11305
rect 5169 11339 5227 11345
rect 5169 11305 5181 11339
rect 5215 11336 5227 11339
rect 5353 11339 5411 11345
rect 5215 11308 5304 11336
rect 5215 11305 5227 11308
rect 5169 11299 5227 11305
rect 1673 11271 1731 11277
rect 1673 11237 1685 11271
rect 1719 11268 1731 11271
rect 1762 11268 1768 11280
rect 1719 11240 1768 11268
rect 1719 11237 1731 11240
rect 1673 11231 1731 11237
rect 1762 11228 1768 11240
rect 1820 11268 1826 11280
rect 2406 11268 2412 11280
rect 1820 11240 2412 11268
rect 1820 11228 1826 11240
rect 2406 11228 2412 11240
rect 2464 11228 2470 11280
rect 3142 11228 3148 11280
rect 3200 11268 3206 11280
rect 3418 11268 3424 11280
rect 3200 11240 3424 11268
rect 3200 11228 3206 11240
rect 3418 11228 3424 11240
rect 3476 11228 3482 11280
rect 2593 11203 2651 11209
rect 2593 11169 2605 11203
rect 2639 11200 2651 11203
rect 2866 11200 2872 11212
rect 2639 11172 2872 11200
rect 2639 11169 2651 11172
rect 2593 11163 2651 11169
rect 2866 11160 2872 11172
rect 2924 11160 2930 11212
rect 3050 11160 3056 11212
rect 3108 11200 3114 11212
rect 3234 11200 3240 11212
rect 3108 11172 3240 11200
rect 3108 11160 3114 11172
rect 3234 11160 3240 11172
rect 3292 11160 3298 11212
rect 2133 11135 2191 11141
rect 2133 11101 2145 11135
rect 2179 11132 2191 11135
rect 2498 11132 2504 11144
rect 2179 11104 2504 11132
rect 2179 11101 2191 11104
rect 2133 11095 2191 11101
rect 2498 11092 2504 11104
rect 2556 11092 2562 11144
rect 2774 11092 2780 11144
rect 2832 11132 2838 11144
rect 3418 11132 3424 11144
rect 2832 11104 3424 11132
rect 2832 11092 2838 11104
rect 3418 11092 3424 11104
rect 3476 11092 3482 11144
rect 3973 11135 4031 11141
rect 3973 11101 3985 11135
rect 4019 11132 4031 11135
rect 4062 11132 4068 11144
rect 4019 11104 4068 11132
rect 4019 11101 4031 11104
rect 3973 11095 4031 11101
rect 4062 11092 4068 11104
rect 4120 11092 4126 11144
rect 4157 11135 4215 11141
rect 4157 11101 4169 11135
rect 4203 11132 4215 11135
rect 4338 11132 4344 11144
rect 4203 11104 4344 11132
rect 4203 11101 4215 11104
rect 4157 11095 4215 11101
rect 4338 11092 4344 11104
rect 4396 11092 4402 11144
rect 1486 11024 1492 11076
rect 1544 11064 1550 11076
rect 2222 11064 2228 11076
rect 1544 11036 2228 11064
rect 1544 11024 1550 11036
rect 2222 11024 2228 11036
rect 2280 11064 2286 11076
rect 3237 11067 3295 11073
rect 3237 11064 3249 11067
rect 2280 11036 3249 11064
rect 2280 11024 2286 11036
rect 3237 11033 3249 11036
rect 3283 11033 3295 11067
rect 4982 11064 4988 11076
rect 4943 11036 4988 11064
rect 3237 11027 3295 11033
rect 4982 11024 4988 11036
rect 5040 11024 5046 11076
rect 5074 11024 5080 11076
rect 5132 11064 5138 11076
rect 5185 11067 5243 11073
rect 5185 11064 5197 11067
rect 5132 11036 5197 11064
rect 5132 11024 5138 11036
rect 5185 11033 5197 11036
rect 5231 11033 5243 11067
rect 5276 11064 5304 11308
rect 5353 11305 5365 11339
rect 5399 11336 5411 11339
rect 5442 11336 5448 11348
rect 5399 11308 5448 11336
rect 5399 11305 5411 11308
rect 5353 11299 5411 11305
rect 5442 11296 5448 11308
rect 5500 11296 5506 11348
rect 6270 11336 6276 11348
rect 6231 11308 6276 11336
rect 6270 11296 6276 11308
rect 6328 11296 6334 11348
rect 6917 11339 6975 11345
rect 6917 11305 6929 11339
rect 6963 11336 6975 11339
rect 7650 11336 7656 11348
rect 6963 11308 7656 11336
rect 6963 11305 6975 11308
rect 6917 11299 6975 11305
rect 7650 11296 7656 11308
rect 7708 11296 7714 11348
rect 8386 11336 8392 11348
rect 8347 11308 8392 11336
rect 8386 11296 8392 11308
rect 8444 11296 8450 11348
rect 8570 11336 8576 11348
rect 8531 11308 8576 11336
rect 8570 11296 8576 11308
rect 8628 11296 8634 11348
rect 9858 11296 9864 11348
rect 9916 11336 9922 11348
rect 10321 11339 10379 11345
rect 10321 11336 10333 11339
rect 9916 11308 10333 11336
rect 9916 11296 9922 11308
rect 10321 11305 10333 11308
rect 10367 11305 10379 11339
rect 10321 11299 10379 11305
rect 13078 11296 13084 11348
rect 13136 11336 13142 11348
rect 14277 11339 14335 11345
rect 14277 11336 14289 11339
rect 13136 11308 14289 11336
rect 13136 11296 13142 11308
rect 14277 11305 14289 11308
rect 14323 11305 14335 11339
rect 14277 11299 14335 11305
rect 14366 11296 14372 11348
rect 14424 11336 14430 11348
rect 14826 11336 14832 11348
rect 14424 11308 14832 11336
rect 14424 11296 14430 11308
rect 14826 11296 14832 11308
rect 14884 11296 14890 11348
rect 16482 11336 16488 11348
rect 16443 11308 16488 11336
rect 16482 11296 16488 11308
rect 16540 11296 16546 11348
rect 17218 11336 17224 11348
rect 17179 11308 17224 11336
rect 17218 11296 17224 11308
rect 17276 11296 17282 11348
rect 17586 11296 17592 11348
rect 17644 11336 17650 11348
rect 19797 11339 19855 11345
rect 19797 11336 19809 11339
rect 17644 11308 19809 11336
rect 17644 11296 17650 11308
rect 19797 11305 19809 11308
rect 19843 11305 19855 11339
rect 20346 11336 20352 11348
rect 20307 11308 20352 11336
rect 19797 11299 19855 11305
rect 20346 11296 20352 11308
rect 20404 11296 20410 11348
rect 20714 11296 20720 11348
rect 20772 11336 20778 11348
rect 21453 11339 21511 11345
rect 21453 11336 21465 11339
rect 20772 11308 21465 11336
rect 20772 11296 20778 11308
rect 21453 11305 21465 11308
rect 21499 11305 21511 11339
rect 21726 11336 21732 11348
rect 21687 11308 21732 11336
rect 21453 11299 21511 11305
rect 21726 11296 21732 11308
rect 21784 11296 21790 11348
rect 5460 11132 5488 11296
rect 9030 11228 9036 11280
rect 9088 11268 9094 11280
rect 9214 11268 9220 11280
rect 9088 11240 9220 11268
rect 9088 11228 9094 11240
rect 9214 11228 9220 11240
rect 9272 11268 9278 11280
rect 9398 11268 9404 11280
rect 9272 11240 9404 11268
rect 9272 11228 9278 11240
rect 9398 11228 9404 11240
rect 9456 11228 9462 11280
rect 11330 11228 11336 11280
rect 11388 11268 11394 11280
rect 11606 11268 11612 11280
rect 11388 11240 11612 11268
rect 11388 11228 11394 11240
rect 11606 11228 11612 11240
rect 11664 11228 11670 11280
rect 15473 11271 15531 11277
rect 15473 11268 15485 11271
rect 13464 11240 15485 11268
rect 5626 11160 5632 11212
rect 5684 11200 5690 11212
rect 5684 11172 6132 11200
rect 5684 11160 5690 11172
rect 6104 11141 6132 11172
rect 6270 11160 6276 11212
rect 6328 11200 6334 11212
rect 8297 11203 8355 11209
rect 8297 11200 8309 11203
rect 6328 11172 8309 11200
rect 6328 11160 6334 11172
rect 8297 11169 8309 11172
rect 8343 11169 8355 11203
rect 10226 11200 10232 11212
rect 8297 11163 8355 11169
rect 8588 11172 10232 11200
rect 5905 11135 5963 11141
rect 5905 11132 5917 11135
rect 5460 11104 5917 11132
rect 5905 11101 5917 11104
rect 5951 11101 5963 11135
rect 5905 11095 5963 11101
rect 5997 11135 6055 11141
rect 5997 11101 6009 11135
rect 6043 11101 6055 11135
rect 5997 11095 6055 11101
rect 6089 11135 6147 11141
rect 6089 11101 6101 11135
rect 6135 11101 6147 11135
rect 7098 11132 7104 11144
rect 7059 11104 7104 11132
rect 6089 11095 6147 11101
rect 5718 11064 5724 11076
rect 5276 11036 5724 11064
rect 5185 11027 5243 11033
rect 5718 11024 5724 11036
rect 5776 11024 5782 11076
rect 6012 11064 6040 11095
rect 7098 11092 7104 11104
rect 7156 11092 7162 11144
rect 7190 11092 7196 11144
rect 7248 11132 7254 11144
rect 7558 11132 7564 11144
rect 7248 11104 7293 11132
rect 7519 11104 7564 11132
rect 7248 11092 7254 11104
rect 7558 11092 7564 11104
rect 7616 11092 7622 11144
rect 8205 11135 8263 11141
rect 8205 11101 8217 11135
rect 8251 11101 8263 11135
rect 8312 11132 8340 11163
rect 8588 11132 8616 11172
rect 8312 11104 8616 11132
rect 8205 11095 8263 11101
rect 6178 11064 6184 11076
rect 6012 11036 6184 11064
rect 6178 11024 6184 11036
rect 6236 11024 6242 11076
rect 7006 11024 7012 11076
rect 7064 11064 7070 11076
rect 7282 11064 7288 11076
rect 7064 11036 7288 11064
rect 7064 11024 7070 11036
rect 7282 11024 7288 11036
rect 7340 11024 7346 11076
rect 7423 11067 7481 11073
rect 7423 11033 7435 11067
rect 7469 11064 7481 11067
rect 8110 11064 8116 11076
rect 7469 11036 8116 11064
rect 7469 11033 7481 11036
rect 7423 11027 7481 11033
rect 8110 11024 8116 11036
rect 8168 11024 8174 11076
rect 8220 11064 8248 11095
rect 9122 11092 9128 11144
rect 9180 11132 9186 11144
rect 9309 11135 9367 11141
rect 9309 11132 9321 11135
rect 9180 11104 9321 11132
rect 9180 11092 9186 11104
rect 9309 11101 9321 11104
rect 9355 11101 9367 11135
rect 9309 11095 9367 11101
rect 9398 11092 9404 11144
rect 9456 11132 9462 11144
rect 9692 11141 9720 11172
rect 10226 11160 10232 11172
rect 10284 11160 10290 11212
rect 9585 11135 9643 11141
rect 9456 11104 9501 11132
rect 9456 11092 9462 11104
rect 9585 11101 9597 11135
rect 9631 11101 9643 11135
rect 9585 11095 9643 11101
rect 9677 11135 9735 11141
rect 9677 11101 9689 11135
rect 9723 11101 9735 11135
rect 9677 11095 9735 11101
rect 10137 11135 10195 11141
rect 10137 11101 10149 11135
rect 10183 11101 10195 11135
rect 10318 11132 10324 11144
rect 10279 11104 10324 11132
rect 10137 11095 10195 11101
rect 8478 11064 8484 11076
rect 8220 11036 8484 11064
rect 8478 11024 8484 11036
rect 8536 11024 8542 11076
rect 9030 11024 9036 11076
rect 9088 11064 9094 11076
rect 9600 11064 9628 11095
rect 9088 11036 9628 11064
rect 10152 11064 10180 11095
rect 10318 11092 10324 11104
rect 10376 11092 10382 11144
rect 11517 11135 11575 11141
rect 11517 11101 11529 11135
rect 11563 11101 11575 11135
rect 11517 11095 11575 11101
rect 10594 11064 10600 11076
rect 10152 11036 10600 11064
rect 9088 11024 9094 11036
rect 10594 11024 10600 11036
rect 10652 11024 10658 11076
rect 11532 11064 11560 11095
rect 11606 11092 11612 11144
rect 11664 11132 11670 11144
rect 11977 11135 12035 11141
rect 11977 11132 11989 11135
rect 11664 11104 11989 11132
rect 11664 11092 11670 11104
rect 11977 11101 11989 11104
rect 12023 11101 12035 11135
rect 13170 11132 13176 11144
rect 13131 11104 13176 11132
rect 11977 11095 12035 11101
rect 13170 11092 13176 11104
rect 13228 11132 13234 11144
rect 13464 11141 13492 11240
rect 15473 11237 15485 11240
rect 15519 11268 15531 11271
rect 17862 11268 17868 11280
rect 15519 11240 17868 11268
rect 15519 11237 15531 11240
rect 15473 11231 15531 11237
rect 17862 11228 17868 11240
rect 17920 11228 17926 11280
rect 18322 11228 18328 11280
rect 18380 11268 18386 11280
rect 18417 11271 18475 11277
rect 18417 11268 18429 11271
rect 18380 11240 18429 11268
rect 18380 11228 18386 11240
rect 18417 11237 18429 11240
rect 18463 11237 18475 11271
rect 18417 11231 18475 11237
rect 18509 11271 18567 11277
rect 18509 11237 18521 11271
rect 18555 11268 18567 11271
rect 19610 11268 19616 11280
rect 18555 11240 19616 11268
rect 18555 11237 18567 11240
rect 18509 11231 18567 11237
rect 13814 11160 13820 11212
rect 13872 11200 13878 11212
rect 14550 11200 14556 11212
rect 13872 11172 14556 11200
rect 13872 11160 13878 11172
rect 14550 11160 14556 11172
rect 14608 11160 14614 11212
rect 16114 11200 16120 11212
rect 14936 11172 16120 11200
rect 13449 11135 13507 11141
rect 13228 11104 13400 11132
rect 13228 11092 13234 11104
rect 11698 11064 11704 11076
rect 11532 11036 11704 11064
rect 11698 11024 11704 11036
rect 11756 11024 11762 11076
rect 12710 11064 12716 11076
rect 12374 11036 12716 11064
rect 12710 11024 12716 11036
rect 12768 11064 12774 11076
rect 12986 11064 12992 11076
rect 12768 11036 12992 11064
rect 12768 11024 12774 11036
rect 12986 11024 12992 11036
rect 13044 11024 13050 11076
rect 13078 11024 13084 11076
rect 13136 11064 13142 11076
rect 13265 11067 13323 11073
rect 13265 11064 13277 11067
rect 13136 11036 13277 11064
rect 13136 11024 13142 11036
rect 13265 11033 13277 11036
rect 13311 11033 13323 11067
rect 13372 11064 13400 11104
rect 13449 11101 13461 11135
rect 13495 11101 13507 11135
rect 14458 11132 14464 11144
rect 14419 11104 14464 11132
rect 13449 11095 13507 11101
rect 14458 11092 14464 11104
rect 14516 11092 14522 11144
rect 14645 11135 14703 11141
rect 14645 11101 14657 11135
rect 14691 11101 14703 11135
rect 14645 11095 14703 11101
rect 14737 11135 14795 11141
rect 14737 11101 14749 11135
rect 14783 11132 14795 11135
rect 14826 11132 14832 11144
rect 14783 11104 14832 11132
rect 14783 11101 14795 11104
rect 14737 11095 14795 11101
rect 13630 11064 13636 11076
rect 13372 11036 13636 11064
rect 13265 11027 13323 11033
rect 2774 10956 2780 11008
rect 2832 10996 2838 11008
rect 3053 10999 3111 11005
rect 3053 10996 3065 10999
rect 2832 10968 3065 10996
rect 2832 10956 2838 10968
rect 3053 10965 3065 10968
rect 3099 10965 3111 10999
rect 3053 10959 3111 10965
rect 4065 10999 4123 11005
rect 4065 10965 4077 10999
rect 4111 10996 4123 10999
rect 4246 10996 4252 11008
rect 4111 10968 4252 10996
rect 4111 10965 4123 10968
rect 4065 10959 4123 10965
rect 4246 10956 4252 10968
rect 4304 10956 4310 11008
rect 7834 10956 7840 11008
rect 7892 10996 7898 11008
rect 9125 10999 9183 11005
rect 9125 10996 9137 10999
rect 7892 10968 9137 10996
rect 7892 10956 7898 10968
rect 9125 10965 9137 10968
rect 9171 10965 9183 10999
rect 13170 10996 13176 11008
rect 13131 10968 13176 10996
rect 9125 10959 9183 10965
rect 13170 10956 13176 10968
rect 13228 10956 13234 11008
rect 13280 10996 13308 11027
rect 13630 11024 13636 11036
rect 13688 11024 13694 11076
rect 14660 11064 14688 11095
rect 14826 11092 14832 11104
rect 14884 11092 14890 11144
rect 14936 11141 14964 11172
rect 16114 11160 16120 11172
rect 16172 11160 16178 11212
rect 14921 11135 14979 11141
rect 14921 11101 14933 11135
rect 14967 11101 14979 11135
rect 14921 11095 14979 11101
rect 15381 11135 15439 11141
rect 15381 11101 15393 11135
rect 15427 11132 15439 11135
rect 15470 11132 15476 11144
rect 15427 11104 15476 11132
rect 15427 11101 15439 11104
rect 15381 11095 15439 11101
rect 15396 11064 15424 11095
rect 15470 11092 15476 11104
rect 15528 11092 15534 11144
rect 15565 11135 15623 11141
rect 15565 11101 15577 11135
rect 15611 11132 15623 11135
rect 15746 11132 15752 11144
rect 15611 11104 15752 11132
rect 15611 11101 15623 11104
rect 15565 11095 15623 11101
rect 15746 11092 15752 11104
rect 15804 11092 15810 11144
rect 16022 11132 16028 11144
rect 15983 11104 16028 11132
rect 16022 11092 16028 11104
rect 16080 11092 16086 11144
rect 16301 11135 16359 11141
rect 16301 11101 16313 11135
rect 16347 11132 16359 11135
rect 16390 11132 16396 11144
rect 16347 11104 16396 11132
rect 16347 11101 16359 11104
rect 16301 11095 16359 11101
rect 16390 11092 16396 11104
rect 16448 11092 16454 11144
rect 16942 11132 16948 11144
rect 16903 11104 16948 11132
rect 16942 11092 16948 11104
rect 17000 11092 17006 11144
rect 17037 11135 17095 11141
rect 17037 11101 17049 11135
rect 17083 11132 17095 11135
rect 17678 11132 17684 11144
rect 17083 11104 17684 11132
rect 17083 11101 17095 11104
rect 17037 11095 17095 11101
rect 17678 11092 17684 11104
rect 17736 11092 17742 11144
rect 18432 11132 18460 11231
rect 19610 11228 19616 11240
rect 19668 11228 19674 11280
rect 19886 11228 19892 11280
rect 19944 11268 19950 11280
rect 19944 11240 22324 11268
rect 19944 11228 19950 11240
rect 18601 11203 18659 11209
rect 18601 11169 18613 11203
rect 18647 11200 18659 11203
rect 19518 11200 19524 11212
rect 18647 11172 19524 11200
rect 18647 11169 18659 11172
rect 18601 11163 18659 11169
rect 19518 11160 19524 11172
rect 19576 11160 19582 11212
rect 21174 11200 21180 11212
rect 19628 11172 21180 11200
rect 18506 11132 18512 11144
rect 18432 11104 18512 11132
rect 18506 11092 18512 11104
rect 18564 11092 18570 11144
rect 18693 11135 18751 11141
rect 18693 11101 18705 11135
rect 18739 11132 18751 11135
rect 18782 11132 18788 11144
rect 18739 11104 18788 11132
rect 18739 11101 18751 11104
rect 18693 11095 18751 11101
rect 18782 11092 18788 11104
rect 18840 11092 18846 11144
rect 18877 11135 18935 11141
rect 18877 11101 18889 11135
rect 18923 11132 18935 11135
rect 18966 11132 18972 11144
rect 18923 11104 18972 11132
rect 18923 11101 18935 11104
rect 18877 11095 18935 11101
rect 18966 11092 18972 11104
rect 19024 11092 19030 11144
rect 19426 11132 19432 11144
rect 19387 11104 19432 11132
rect 19426 11092 19432 11104
rect 19484 11092 19490 11144
rect 19628 11141 19656 11172
rect 21174 11160 21180 11172
rect 21232 11160 21238 11212
rect 19613 11135 19671 11141
rect 19613 11101 19625 11135
rect 19659 11101 19671 11135
rect 19613 11095 19671 11101
rect 19886 11092 19892 11144
rect 19944 11132 19950 11144
rect 20625 11135 20683 11141
rect 19944 11104 19989 11132
rect 20625 11110 20637 11135
rect 19944 11092 19950 11104
rect 20456 11101 20637 11110
rect 20671 11101 20683 11135
rect 20456 11095 20683 11101
rect 20714 11132 20772 11138
rect 20714 11122 20726 11132
rect 20760 11122 20772 11132
rect 16040 11064 16068 11092
rect 20456 11082 20668 11095
rect 13740 11036 14596 11064
rect 14660 11036 15424 11064
rect 15488 11036 16068 11064
rect 16117 11067 16175 11073
rect 13740 10996 13768 11036
rect 13280 10968 13768 10996
rect 14568 10996 14596 11036
rect 15488 10996 15516 11036
rect 16117 11033 16129 11067
rect 16163 11064 16175 11067
rect 16666 11064 16672 11076
rect 16163 11036 16672 11064
rect 16163 11033 16175 11036
rect 16117 11027 16175 11033
rect 16666 11024 16672 11036
rect 16724 11024 16730 11076
rect 17221 11067 17279 11073
rect 17221 11033 17233 11067
rect 17267 11064 17279 11067
rect 17770 11064 17776 11076
rect 17267 11036 17776 11064
rect 17267 11033 17279 11036
rect 17221 11027 17279 11033
rect 17770 11024 17776 11036
rect 17828 11064 17834 11076
rect 18322 11064 18328 11076
rect 17828 11036 18328 11064
rect 17828 11024 17834 11036
rect 18322 11024 18328 11036
rect 18380 11024 18386 11076
rect 19242 11024 19248 11076
rect 19300 11064 19306 11076
rect 19702 11064 19708 11076
rect 19300 11036 19708 11064
rect 19300 11024 19306 11036
rect 19702 11024 19708 11036
rect 19760 11024 19766 11076
rect 20346 11024 20352 11076
rect 20404 11064 20410 11076
rect 20456 11064 20484 11082
rect 20714 11070 20720 11122
rect 20772 11070 20778 11122
rect 20806 11086 20812 11138
rect 20864 11126 20870 11138
rect 20864 11098 20909 11126
rect 20864 11086 20870 11098
rect 20990 11092 20996 11144
rect 21048 11132 21054 11144
rect 21729 11135 21787 11141
rect 21048 11104 21093 11132
rect 21048 11092 21054 11104
rect 21729 11101 21741 11135
rect 21775 11101 21787 11135
rect 21729 11095 21787 11101
rect 20404 11036 20484 11064
rect 20404 11024 20410 11036
rect 21634 11024 21640 11076
rect 21692 11064 21698 11076
rect 21744 11064 21772 11095
rect 21818 11092 21824 11144
rect 21876 11132 21882 11144
rect 22296 11141 22324 11240
rect 22281 11135 22339 11141
rect 21876 11104 21921 11132
rect 21876 11092 21882 11104
rect 22281 11101 22293 11135
rect 22327 11101 22339 11135
rect 22281 11095 22339 11101
rect 22373 11067 22431 11073
rect 22373 11064 22385 11067
rect 21692 11036 22385 11064
rect 21692 11024 21698 11036
rect 22373 11033 22385 11036
rect 22419 11033 22431 11067
rect 22373 11027 22431 11033
rect 14568 10968 15516 10996
rect 15562 10956 15568 11008
rect 15620 10996 15626 11008
rect 15746 10996 15752 11008
rect 15620 10968 15752 10996
rect 15620 10956 15626 10968
rect 15746 10956 15752 10968
rect 15804 10956 15810 11008
rect 16482 10956 16488 11008
rect 16540 10996 16546 11008
rect 18141 10999 18199 11005
rect 18141 10996 18153 10999
rect 16540 10968 18153 10996
rect 16540 10956 16546 10968
rect 18141 10965 18153 10968
rect 18187 10965 18199 10999
rect 18141 10959 18199 10965
rect 19150 10956 19156 11008
rect 19208 10996 19214 11008
rect 20530 10996 20536 11008
rect 19208 10968 20536 10996
rect 19208 10956 19214 10968
rect 20530 10956 20536 10968
rect 20588 10956 20594 11008
rect 1104 10906 23987 10928
rect 1104 10854 6630 10906
rect 6682 10854 6694 10906
rect 6746 10854 6758 10906
rect 6810 10854 6822 10906
rect 6874 10854 6886 10906
rect 6938 10854 12311 10906
rect 12363 10854 12375 10906
rect 12427 10854 12439 10906
rect 12491 10854 12503 10906
rect 12555 10854 12567 10906
rect 12619 10854 17992 10906
rect 18044 10854 18056 10906
rect 18108 10854 18120 10906
rect 18172 10854 18184 10906
rect 18236 10854 18248 10906
rect 18300 10854 23673 10906
rect 23725 10854 23737 10906
rect 23789 10854 23801 10906
rect 23853 10854 23865 10906
rect 23917 10854 23929 10906
rect 23981 10854 23987 10906
rect 1104 10832 23987 10854
rect 2866 10752 2872 10804
rect 2924 10752 2930 10804
rect 3694 10752 3700 10804
rect 3752 10792 3758 10804
rect 4249 10795 4307 10801
rect 3752 10764 4200 10792
rect 3752 10752 3758 10764
rect 1578 10616 1584 10668
rect 1636 10656 1642 10668
rect 1673 10659 1731 10665
rect 1673 10656 1685 10659
rect 1636 10628 1685 10656
rect 1636 10616 1642 10628
rect 1673 10625 1685 10628
rect 1719 10625 1731 10659
rect 1673 10619 1731 10625
rect 2222 10616 2228 10668
rect 2280 10656 2286 10668
rect 2593 10659 2651 10665
rect 2593 10656 2605 10659
rect 2280 10628 2605 10656
rect 2280 10616 2286 10628
rect 2593 10625 2605 10628
rect 2639 10625 2651 10659
rect 2593 10619 2651 10625
rect 2686 10659 2744 10665
rect 2686 10625 2698 10659
rect 2732 10656 2744 10659
rect 2774 10656 2780 10668
rect 2732 10628 2780 10656
rect 2732 10625 2744 10628
rect 2686 10619 2744 10625
rect 2774 10616 2780 10628
rect 2832 10616 2838 10668
rect 2884 10665 2912 10752
rect 3602 10684 3608 10736
rect 3660 10724 3666 10736
rect 4172 10724 4200 10764
rect 4249 10761 4261 10795
rect 4295 10792 4307 10795
rect 5626 10792 5632 10804
rect 4295 10764 5632 10792
rect 4295 10761 4307 10764
rect 4249 10755 4307 10761
rect 5626 10752 5632 10764
rect 5684 10752 5690 10804
rect 6546 10792 6552 10804
rect 6507 10764 6552 10792
rect 6546 10752 6552 10764
rect 6604 10752 6610 10804
rect 8478 10792 8484 10804
rect 8439 10764 8484 10792
rect 8478 10752 8484 10764
rect 8536 10752 8542 10804
rect 8938 10752 8944 10804
rect 8996 10752 9002 10804
rect 9306 10752 9312 10804
rect 9364 10792 9370 10804
rect 9585 10795 9643 10801
rect 9585 10792 9597 10795
rect 9364 10764 9597 10792
rect 9364 10752 9370 10764
rect 9585 10761 9597 10764
rect 9631 10761 9643 10795
rect 11146 10792 11152 10804
rect 9585 10755 9643 10761
rect 10796 10764 11152 10792
rect 4614 10724 4620 10736
rect 3660 10696 4108 10724
rect 4172 10696 4620 10724
rect 3660 10684 3666 10696
rect 2869 10659 2927 10665
rect 2869 10625 2881 10659
rect 2915 10625 2927 10659
rect 2869 10619 2927 10625
rect 2961 10659 3019 10665
rect 2961 10625 2973 10659
rect 3007 10625 3019 10659
rect 2961 10619 3019 10625
rect 2133 10591 2191 10597
rect 2133 10557 2145 10591
rect 2179 10588 2191 10591
rect 2976 10588 3004 10619
rect 3050 10616 3056 10668
rect 3108 10665 3114 10668
rect 3108 10656 3116 10665
rect 3108 10628 3153 10656
rect 3108 10619 3116 10628
rect 3108 10616 3114 10619
rect 3694 10616 3700 10668
rect 3752 10656 3758 10668
rect 4080 10665 4108 10696
rect 4614 10684 4620 10696
rect 4672 10684 4678 10736
rect 6917 10727 6975 10733
rect 6917 10693 6929 10727
rect 6963 10724 6975 10727
rect 8570 10724 8576 10736
rect 6963 10696 8576 10724
rect 6963 10693 6975 10696
rect 6917 10687 6975 10693
rect 8570 10684 8576 10696
rect 8628 10684 8634 10736
rect 8956 10724 8984 10752
rect 8956 10696 9168 10724
rect 3789 10659 3847 10665
rect 3789 10656 3801 10659
rect 3752 10628 3801 10656
rect 3752 10616 3758 10628
rect 3789 10625 3801 10628
rect 3835 10625 3847 10659
rect 3789 10619 3847 10625
rect 4065 10659 4123 10665
rect 4065 10625 4077 10659
rect 4111 10625 4123 10659
rect 4065 10619 4123 10625
rect 4522 10616 4528 10668
rect 4580 10656 4586 10668
rect 4709 10659 4767 10665
rect 4709 10656 4721 10659
rect 4580 10628 4721 10656
rect 4580 10616 4586 10628
rect 4709 10625 4721 10628
rect 4755 10656 4767 10659
rect 4798 10656 4804 10668
rect 4755 10628 4804 10656
rect 4755 10625 4767 10628
rect 4709 10619 4767 10625
rect 4798 10616 4804 10628
rect 4856 10616 4862 10668
rect 5445 10659 5503 10665
rect 5445 10625 5457 10659
rect 5491 10625 5503 10659
rect 5445 10619 5503 10625
rect 5629 10659 5687 10665
rect 5629 10625 5641 10659
rect 5675 10656 5687 10659
rect 6086 10656 6092 10668
rect 5675 10628 6092 10656
rect 5675 10625 5687 10628
rect 5629 10619 5687 10625
rect 3881 10591 3939 10597
rect 3881 10588 3893 10591
rect 2179 10560 3041 10588
rect 3160 10560 3893 10588
rect 2179 10557 2191 10560
rect 2133 10551 2191 10557
rect 2976 10532 3004 10560
rect 2958 10480 2964 10532
rect 3016 10480 3022 10532
rect 3160 10464 3188 10560
rect 3881 10557 3893 10560
rect 3927 10557 3939 10591
rect 3881 10551 3939 10557
rect 5460 10588 5488 10619
rect 6086 10616 6092 10628
rect 6144 10616 6150 10668
rect 6270 10616 6276 10668
rect 6328 10656 6334 10668
rect 6733 10659 6791 10665
rect 6733 10656 6745 10659
rect 6328 10628 6745 10656
rect 6328 10616 6334 10628
rect 6733 10625 6745 10628
rect 6779 10625 6791 10659
rect 6733 10619 6791 10625
rect 7843 10659 7901 10665
rect 7843 10625 7855 10659
rect 7889 10625 7901 10659
rect 8018 10656 8024 10668
rect 7979 10628 8024 10656
rect 7843 10619 7901 10625
rect 7190 10588 7196 10600
rect 5460 10560 7196 10588
rect 3234 10480 3240 10532
rect 3292 10520 3298 10532
rect 3292 10492 3337 10520
rect 3292 10480 3298 10492
rect 3510 10480 3516 10532
rect 3568 10520 3574 10532
rect 5460 10520 5488 10560
rect 7190 10548 7196 10560
rect 7248 10548 7254 10600
rect 7853 10520 7881 10619
rect 8018 10616 8024 10628
rect 8076 10616 8082 10668
rect 8754 10656 8760 10668
rect 8715 10628 8760 10656
rect 8754 10616 8760 10628
rect 8812 10616 8818 10668
rect 8849 10659 8907 10665
rect 8849 10625 8861 10659
rect 8895 10625 8907 10659
rect 8849 10619 8907 10625
rect 8386 10548 8392 10600
rect 8444 10588 8450 10600
rect 8864 10588 8892 10619
rect 8938 10616 8944 10668
rect 8996 10656 9002 10668
rect 9140 10665 9168 10696
rect 9324 10696 10088 10724
rect 9125 10659 9183 10665
rect 8996 10628 9041 10656
rect 8996 10616 9002 10628
rect 9125 10625 9137 10659
rect 9171 10625 9183 10659
rect 9125 10619 9183 10625
rect 8444 10560 8892 10588
rect 8444 10548 8450 10560
rect 9324 10532 9352 10696
rect 9398 10616 9404 10668
rect 9456 10656 9462 10668
rect 9953 10659 10011 10665
rect 9953 10656 9965 10659
rect 9456 10628 9965 10656
rect 9456 10616 9462 10628
rect 9953 10625 9965 10628
rect 9999 10625 10011 10659
rect 9953 10619 10011 10625
rect 9769 10591 9827 10597
rect 9769 10557 9781 10591
rect 9815 10557 9827 10591
rect 9769 10551 9827 10557
rect 3568 10492 5488 10520
rect 5552 10492 7881 10520
rect 8021 10523 8079 10529
rect 3568 10480 3574 10492
rect 1946 10452 1952 10464
rect 1859 10424 1952 10452
rect 1946 10412 1952 10424
rect 2004 10452 2010 10464
rect 2498 10452 2504 10464
rect 2004 10424 2504 10452
rect 2004 10412 2010 10424
rect 2498 10412 2504 10424
rect 2556 10412 2562 10464
rect 3142 10412 3148 10464
rect 3200 10412 3206 10464
rect 4065 10455 4123 10461
rect 4065 10421 4077 10455
rect 4111 10452 4123 10455
rect 4246 10452 4252 10464
rect 4111 10424 4252 10452
rect 4111 10421 4123 10424
rect 4065 10415 4123 10421
rect 4246 10412 4252 10424
rect 4304 10412 4310 10464
rect 4893 10455 4951 10461
rect 4893 10421 4905 10455
rect 4939 10452 4951 10455
rect 4982 10452 4988 10464
rect 4939 10424 4988 10452
rect 4939 10421 4951 10424
rect 4893 10415 4951 10421
rect 4982 10412 4988 10424
rect 5040 10452 5046 10464
rect 5552 10452 5580 10492
rect 8021 10489 8033 10523
rect 8067 10520 8079 10523
rect 9306 10520 9312 10532
rect 8067 10492 9312 10520
rect 8067 10489 8079 10492
rect 8021 10483 8079 10489
rect 9306 10480 9312 10492
rect 9364 10480 9370 10532
rect 9784 10520 9812 10551
rect 9858 10548 9864 10600
rect 9916 10588 9922 10600
rect 10060 10597 10088 10696
rect 10045 10591 10103 10597
rect 9916 10560 9961 10588
rect 9916 10548 9922 10560
rect 10045 10557 10057 10591
rect 10091 10557 10103 10591
rect 10045 10551 10103 10557
rect 10796 10520 10824 10764
rect 11146 10752 11152 10764
rect 11204 10752 11210 10804
rect 11882 10752 11888 10804
rect 11940 10792 11946 10804
rect 12253 10795 12311 10801
rect 12253 10792 12265 10795
rect 11940 10764 12265 10792
rect 11940 10752 11946 10764
rect 12253 10761 12265 10764
rect 12299 10761 12311 10795
rect 13078 10792 13084 10804
rect 13039 10764 13084 10792
rect 12253 10755 12311 10761
rect 13078 10752 13084 10764
rect 13136 10752 13142 10804
rect 13538 10752 13544 10804
rect 13596 10792 13602 10804
rect 14366 10792 14372 10804
rect 13596 10764 14372 10792
rect 13596 10752 13602 10764
rect 14366 10752 14372 10764
rect 14424 10752 14430 10804
rect 16114 10752 16120 10804
rect 16172 10792 16178 10804
rect 16209 10795 16267 10801
rect 16209 10792 16221 10795
rect 16172 10764 16221 10792
rect 16172 10752 16178 10764
rect 16209 10761 16221 10764
rect 16255 10761 16267 10795
rect 16209 10755 16267 10761
rect 17586 10752 17592 10804
rect 17644 10752 17650 10804
rect 17681 10795 17739 10801
rect 17681 10761 17693 10795
rect 17727 10792 17739 10795
rect 18414 10792 18420 10804
rect 17727 10764 18420 10792
rect 17727 10761 17739 10764
rect 17681 10755 17739 10761
rect 18414 10752 18420 10764
rect 18472 10752 18478 10804
rect 18877 10795 18935 10801
rect 18877 10761 18889 10795
rect 18923 10792 18935 10795
rect 19334 10792 19340 10804
rect 18923 10764 19340 10792
rect 18923 10761 18935 10764
rect 18877 10755 18935 10761
rect 19334 10752 19340 10764
rect 19392 10752 19398 10804
rect 20349 10795 20407 10801
rect 20349 10761 20361 10795
rect 20395 10792 20407 10795
rect 20438 10792 20444 10804
rect 20395 10764 20444 10792
rect 20395 10761 20407 10764
rect 20349 10755 20407 10761
rect 20438 10752 20444 10764
rect 20496 10752 20502 10804
rect 20530 10752 20536 10804
rect 20588 10792 20594 10804
rect 20588 10764 20633 10792
rect 20588 10752 20594 10764
rect 20990 10752 20996 10804
rect 21048 10792 21054 10804
rect 22005 10795 22063 10801
rect 22005 10792 22017 10795
rect 21048 10764 22017 10792
rect 21048 10752 21054 10764
rect 22005 10761 22017 10764
rect 22051 10761 22063 10795
rect 22005 10755 22063 10761
rect 10873 10727 10931 10733
rect 10873 10693 10885 10727
rect 10919 10724 10931 10727
rect 10962 10724 10968 10736
rect 10919 10696 10968 10724
rect 10919 10693 10931 10696
rect 10873 10687 10931 10693
rect 10962 10684 10968 10696
rect 11020 10684 11026 10736
rect 12713 10727 12771 10733
rect 12713 10724 12725 10727
rect 11164 10696 12725 10724
rect 11164 10665 11192 10696
rect 12713 10693 12725 10696
rect 12759 10693 12771 10727
rect 13722 10724 13728 10736
rect 12713 10687 12771 10693
rect 13188 10696 13728 10724
rect 11149 10659 11207 10665
rect 11149 10625 11161 10659
rect 11195 10625 11207 10659
rect 11149 10619 11207 10625
rect 11422 10616 11428 10668
rect 11480 10656 11486 10668
rect 11885 10659 11943 10665
rect 11885 10656 11897 10659
rect 11480 10628 11897 10656
rect 11480 10616 11486 10628
rect 11885 10625 11897 10628
rect 11931 10625 11943 10659
rect 11885 10619 11943 10625
rect 12069 10659 12127 10665
rect 12069 10625 12081 10659
rect 12115 10656 12127 10659
rect 12802 10656 12808 10668
rect 12115 10628 12808 10656
rect 12115 10625 12127 10628
rect 12069 10619 12127 10625
rect 12802 10616 12808 10628
rect 12860 10616 12866 10668
rect 13188 10665 13216 10696
rect 13722 10684 13728 10696
rect 13780 10724 13786 10736
rect 15286 10724 15292 10736
rect 13780 10696 15292 10724
rect 13780 10684 13786 10696
rect 15286 10684 15292 10696
rect 15344 10684 15350 10736
rect 15562 10684 15568 10736
rect 15620 10724 15626 10736
rect 15657 10727 15715 10733
rect 15657 10724 15669 10727
rect 15620 10696 15669 10724
rect 15620 10684 15626 10696
rect 15657 10693 15669 10696
rect 15703 10724 15715 10727
rect 16942 10724 16948 10736
rect 15703 10696 16948 10724
rect 15703 10693 15715 10696
rect 15657 10687 15715 10693
rect 16942 10684 16948 10696
rect 17000 10724 17006 10736
rect 17604 10724 17632 10752
rect 19426 10724 19432 10736
rect 17000 10696 17632 10724
rect 18616 10696 19432 10724
rect 17000 10684 17006 10696
rect 12989 10659 13047 10665
rect 12989 10625 13001 10659
rect 13035 10625 13047 10659
rect 12989 10619 13047 10625
rect 13173 10659 13231 10665
rect 13173 10625 13185 10659
rect 13219 10625 13231 10659
rect 14642 10656 14648 10668
rect 14603 10628 14648 10656
rect 13173 10619 13231 10625
rect 11793 10591 11851 10597
rect 11793 10588 11805 10591
rect 11164 10560 11805 10588
rect 11054 10520 11060 10532
rect 9784 10492 10824 10520
rect 11015 10492 11060 10520
rect 10060 10464 10088 10492
rect 11054 10480 11060 10492
rect 11112 10480 11118 10532
rect 11164 10529 11192 10560
rect 11793 10557 11805 10560
rect 11839 10557 11851 10591
rect 11793 10551 11851 10557
rect 11977 10591 12035 10597
rect 11977 10557 11989 10591
rect 12023 10557 12035 10591
rect 11977 10551 12035 10557
rect 11149 10523 11207 10529
rect 11149 10489 11161 10523
rect 11195 10489 11207 10523
rect 11149 10483 11207 10489
rect 11698 10480 11704 10532
rect 11756 10520 11762 10532
rect 11992 10520 12020 10551
rect 11756 10492 12020 10520
rect 13004 10520 13032 10619
rect 14642 10616 14648 10628
rect 14700 10616 14706 10668
rect 15473 10659 15531 10665
rect 15473 10625 15485 10659
rect 15519 10656 15531 10659
rect 15838 10656 15844 10668
rect 15519 10628 15844 10656
rect 15519 10625 15531 10628
rect 15473 10619 15531 10625
rect 15838 10616 15844 10628
rect 15896 10616 15902 10668
rect 16114 10656 16120 10668
rect 16075 10628 16120 10656
rect 16114 10616 16120 10628
rect 16172 10616 16178 10668
rect 16301 10659 16359 10665
rect 16301 10625 16313 10659
rect 16347 10656 16359 10659
rect 17494 10656 17500 10668
rect 16347 10628 17500 10656
rect 16347 10625 16359 10628
rect 16301 10619 16359 10625
rect 13449 10591 13507 10597
rect 13449 10557 13461 10591
rect 13495 10588 13507 10591
rect 13906 10588 13912 10600
rect 13495 10560 13912 10588
rect 13495 10557 13507 10560
rect 13449 10551 13507 10557
rect 13906 10548 13912 10560
rect 13964 10548 13970 10600
rect 16316 10588 16344 10619
rect 17494 10616 17500 10628
rect 17552 10616 17558 10668
rect 17589 10659 17647 10665
rect 17589 10625 17601 10659
rect 17635 10625 17647 10659
rect 17589 10619 17647 10625
rect 18325 10659 18383 10665
rect 18325 10625 18337 10659
rect 18371 10625 18383 10659
rect 18325 10619 18383 10625
rect 14568 10560 16344 10588
rect 13004 10492 14044 10520
rect 11756 10480 11762 10492
rect 5040 10424 5580 10452
rect 5629 10455 5687 10461
rect 5040 10412 5046 10424
rect 5629 10421 5641 10455
rect 5675 10452 5687 10455
rect 5718 10452 5724 10464
rect 5675 10424 5724 10452
rect 5675 10421 5687 10424
rect 5629 10415 5687 10421
rect 5718 10412 5724 10424
rect 5776 10452 5782 10464
rect 5994 10452 6000 10464
rect 5776 10424 6000 10452
rect 5776 10412 5782 10424
rect 5994 10412 6000 10424
rect 6052 10452 6058 10464
rect 8202 10452 8208 10464
rect 6052 10424 8208 10452
rect 6052 10412 6058 10424
rect 8202 10412 8208 10424
rect 8260 10412 8266 10464
rect 10042 10412 10048 10464
rect 10100 10412 10106 10464
rect 12342 10412 12348 10464
rect 12400 10452 12406 10464
rect 13357 10455 13415 10461
rect 13357 10452 13369 10455
rect 12400 10424 13369 10452
rect 12400 10412 12406 10424
rect 13357 10421 13369 10424
rect 13403 10452 13415 10455
rect 13814 10452 13820 10464
rect 13403 10424 13820 10452
rect 13403 10421 13415 10424
rect 13357 10415 13415 10421
rect 13814 10412 13820 10424
rect 13872 10412 13878 10464
rect 14016 10461 14044 10492
rect 14568 10464 14596 10560
rect 16666 10548 16672 10600
rect 16724 10588 16730 10600
rect 17218 10588 17224 10600
rect 16724 10560 17224 10588
rect 16724 10548 16730 10560
rect 17218 10548 17224 10560
rect 17276 10548 17282 10600
rect 15838 10480 15844 10532
rect 15896 10520 15902 10532
rect 16853 10523 16911 10529
rect 16853 10520 16865 10523
rect 15896 10492 16865 10520
rect 15896 10480 15902 10492
rect 16853 10489 16865 10492
rect 16899 10489 16911 10523
rect 16853 10483 16911 10489
rect 14001 10455 14059 10461
rect 14001 10421 14013 10455
rect 14047 10452 14059 10455
rect 14090 10452 14096 10464
rect 14047 10424 14096 10452
rect 14047 10421 14059 10424
rect 14001 10415 14059 10421
rect 14090 10412 14096 10424
rect 14148 10412 14154 10464
rect 14550 10452 14556 10464
rect 14511 10424 14556 10452
rect 14550 10412 14556 10424
rect 14608 10412 14614 10464
rect 15010 10412 15016 10464
rect 15068 10452 15074 10464
rect 17604 10452 17632 10619
rect 18340 10520 18368 10619
rect 18414 10616 18420 10668
rect 18472 10656 18478 10668
rect 18616 10665 18644 10696
rect 19426 10684 19432 10696
rect 19484 10684 19490 10736
rect 19886 10724 19892 10736
rect 19720 10696 19892 10724
rect 18601 10659 18659 10665
rect 18472 10628 18517 10656
rect 18472 10616 18478 10628
rect 18601 10625 18613 10659
rect 18647 10625 18659 10659
rect 18601 10619 18659 10625
rect 18693 10659 18751 10665
rect 18693 10625 18705 10659
rect 18739 10656 18751 10659
rect 18782 10656 18788 10668
rect 18739 10628 18788 10656
rect 18739 10625 18751 10628
rect 18693 10619 18751 10625
rect 18782 10616 18788 10628
rect 18840 10616 18846 10668
rect 19334 10616 19340 10668
rect 19392 10656 19398 10668
rect 19613 10659 19671 10665
rect 19613 10656 19625 10659
rect 19392 10628 19625 10656
rect 19392 10616 19398 10628
rect 19613 10625 19625 10628
rect 19659 10625 19671 10659
rect 19613 10619 19671 10625
rect 19720 10600 19748 10696
rect 19886 10684 19892 10696
rect 19944 10724 19950 10736
rect 20717 10727 20775 10733
rect 20717 10724 20729 10727
rect 19944 10696 20729 10724
rect 19944 10684 19950 10696
rect 20717 10693 20729 10696
rect 20763 10693 20775 10727
rect 20717 10687 20775 10693
rect 19797 10659 19855 10665
rect 19797 10625 19809 10659
rect 19843 10656 19855 10659
rect 20622 10656 20628 10668
rect 19843 10628 20484 10656
rect 20583 10628 20628 10656
rect 19843 10625 19855 10628
rect 19797 10619 19855 10625
rect 18874 10548 18880 10600
rect 18932 10588 18938 10600
rect 19521 10591 19579 10597
rect 19521 10588 19533 10591
rect 18932 10560 19533 10588
rect 18932 10548 18938 10560
rect 19521 10557 19533 10560
rect 19567 10557 19579 10591
rect 19521 10551 19579 10557
rect 19702 10548 19708 10600
rect 19760 10588 19766 10600
rect 19760 10560 19805 10588
rect 19760 10548 19766 10560
rect 19904 10520 19932 10628
rect 20456 10588 20484 10628
rect 20622 10616 20628 10628
rect 20680 10616 20686 10668
rect 21358 10588 21364 10600
rect 20456 10560 21364 10588
rect 21358 10548 21364 10560
rect 21416 10548 21422 10600
rect 18340 10492 19932 10520
rect 20901 10523 20959 10529
rect 20901 10489 20913 10523
rect 20947 10520 20959 10523
rect 21542 10520 21548 10532
rect 20947 10492 21548 10520
rect 20947 10489 20959 10492
rect 20901 10483 20959 10489
rect 15068 10424 17632 10452
rect 15068 10412 15074 10424
rect 18690 10412 18696 10464
rect 18748 10452 18754 10464
rect 19337 10455 19395 10461
rect 19337 10452 19349 10455
rect 18748 10424 19349 10452
rect 18748 10412 18754 10424
rect 19337 10421 19349 10424
rect 19383 10421 19395 10455
rect 19337 10415 19395 10421
rect 19426 10412 19432 10464
rect 19484 10452 19490 10464
rect 20916 10452 20944 10483
rect 21542 10480 21548 10492
rect 21600 10480 21606 10532
rect 21450 10452 21456 10464
rect 19484 10424 20944 10452
rect 21411 10424 21456 10452
rect 19484 10412 19490 10424
rect 21450 10412 21456 10424
rect 21508 10412 21514 10464
rect 1104 10362 23828 10384
rect 1104 10310 3790 10362
rect 3842 10310 3854 10362
rect 3906 10310 3918 10362
rect 3970 10310 3982 10362
rect 4034 10310 4046 10362
rect 4098 10310 9471 10362
rect 9523 10310 9535 10362
rect 9587 10310 9599 10362
rect 9651 10310 9663 10362
rect 9715 10310 9727 10362
rect 9779 10310 15152 10362
rect 15204 10310 15216 10362
rect 15268 10310 15280 10362
rect 15332 10310 15344 10362
rect 15396 10310 15408 10362
rect 15460 10310 20833 10362
rect 20885 10310 20897 10362
rect 20949 10310 20961 10362
rect 21013 10310 21025 10362
rect 21077 10310 21089 10362
rect 21141 10310 23828 10362
rect 1104 10288 23828 10310
rect 2222 10248 2228 10260
rect 2183 10220 2228 10248
rect 2222 10208 2228 10220
rect 2280 10208 2286 10260
rect 2406 10248 2412 10260
rect 2367 10220 2412 10248
rect 2406 10208 2412 10220
rect 2464 10208 2470 10260
rect 3694 10208 3700 10260
rect 3752 10248 3758 10260
rect 3973 10251 4031 10257
rect 3973 10248 3985 10251
rect 3752 10220 3985 10248
rect 3752 10208 3758 10220
rect 3973 10217 3985 10220
rect 4019 10217 4031 10251
rect 5074 10248 5080 10260
rect 5035 10220 5080 10248
rect 3973 10211 4031 10217
rect 5074 10208 5080 10220
rect 5132 10208 5138 10260
rect 5902 10248 5908 10260
rect 5863 10220 5908 10248
rect 5902 10208 5908 10220
rect 5960 10208 5966 10260
rect 6178 10248 6184 10260
rect 6139 10220 6184 10248
rect 6178 10208 6184 10220
rect 6236 10208 6242 10260
rect 8389 10251 8447 10257
rect 8389 10217 8401 10251
rect 8435 10248 8447 10251
rect 8938 10248 8944 10260
rect 8435 10220 8944 10248
rect 8435 10217 8447 10220
rect 8389 10211 8447 10217
rect 8938 10208 8944 10220
rect 8996 10208 9002 10260
rect 9122 10248 9128 10260
rect 9083 10220 9128 10248
rect 9122 10208 9128 10220
rect 9180 10208 9186 10260
rect 9950 10248 9956 10260
rect 9232 10220 9956 10248
rect 1765 10183 1823 10189
rect 1765 10149 1777 10183
rect 1811 10180 1823 10183
rect 3421 10183 3479 10189
rect 3421 10180 3433 10183
rect 1811 10152 3433 10180
rect 1811 10149 1823 10152
rect 1765 10143 1823 10149
rect 3421 10149 3433 10152
rect 3467 10180 3479 10183
rect 4522 10180 4528 10192
rect 3467 10152 4528 10180
rect 3467 10149 3479 10152
rect 3421 10143 3479 10149
rect 4522 10140 4528 10152
rect 4580 10140 4586 10192
rect 4614 10140 4620 10192
rect 4672 10180 4678 10192
rect 7009 10183 7067 10189
rect 4672 10152 5396 10180
rect 4672 10140 4678 10152
rect 2501 10115 2559 10121
rect 2501 10081 2513 10115
rect 2547 10112 2559 10115
rect 3510 10112 3516 10124
rect 2547 10084 3516 10112
rect 2547 10081 2559 10084
rect 2501 10075 2559 10081
rect 3510 10072 3516 10084
rect 3568 10072 3574 10124
rect 4890 10112 4896 10124
rect 4172 10084 4896 10112
rect 2777 10047 2835 10053
rect 2777 10013 2789 10047
rect 2823 10044 2835 10047
rect 3326 10044 3332 10056
rect 2823 10016 3332 10044
rect 2823 10013 2835 10016
rect 2777 10007 2835 10013
rect 3326 10004 3332 10016
rect 3384 10004 3390 10056
rect 4172 10053 4200 10084
rect 4890 10072 4896 10084
rect 4948 10072 4954 10124
rect 4982 10072 4988 10124
rect 5040 10112 5046 10124
rect 5368 10121 5396 10152
rect 7009 10149 7021 10183
rect 7055 10180 7067 10183
rect 7834 10180 7840 10192
rect 7055 10152 7840 10180
rect 7055 10149 7067 10152
rect 7009 10143 7067 10149
rect 7834 10140 7840 10152
rect 7892 10140 7898 10192
rect 8018 10140 8024 10192
rect 8076 10180 8082 10192
rect 8076 10152 8708 10180
rect 8076 10140 8082 10152
rect 5169 10115 5227 10121
rect 5169 10112 5181 10115
rect 5040 10084 5181 10112
rect 5040 10072 5046 10084
rect 5169 10081 5181 10084
rect 5215 10081 5227 10115
rect 5169 10075 5227 10081
rect 5353 10115 5411 10121
rect 5353 10081 5365 10115
rect 5399 10112 5411 10115
rect 5534 10112 5540 10124
rect 5399 10084 5540 10112
rect 5399 10081 5411 10084
rect 5353 10075 5411 10081
rect 5534 10072 5540 10084
rect 5592 10072 5598 10124
rect 5920 10084 8616 10112
rect 4157 10047 4215 10053
rect 4157 10013 4169 10047
rect 4203 10013 4215 10047
rect 4157 10007 4215 10013
rect 4172 9920 4200 10007
rect 4246 10004 4252 10056
rect 4304 10044 4310 10056
rect 4433 10047 4491 10053
rect 4433 10044 4445 10047
rect 4304 10016 4445 10044
rect 4304 10004 4310 10016
rect 4433 10013 4445 10016
rect 4479 10013 4491 10047
rect 5074 10044 5080 10056
rect 5035 10016 5080 10044
rect 4433 10007 4491 10013
rect 5074 10004 5080 10016
rect 5132 10004 5138 10056
rect 5810 10044 5816 10056
rect 5771 10016 5816 10044
rect 5810 10004 5816 10016
rect 5868 10004 5874 10056
rect 4338 9976 4344 9988
rect 4251 9948 4344 9976
rect 4338 9936 4344 9948
rect 4396 9976 4402 9988
rect 4982 9976 4988 9988
rect 4396 9948 4988 9976
rect 4396 9936 4402 9948
rect 4982 9936 4988 9948
rect 5040 9936 5046 9988
rect 4154 9868 4160 9920
rect 4212 9868 4218 9920
rect 4798 9868 4804 9920
rect 4856 9908 4862 9920
rect 5920 9908 5948 10084
rect 5997 10047 6055 10053
rect 5997 10013 6009 10047
rect 6043 10013 6055 10047
rect 6730 10044 6736 10056
rect 6691 10016 6736 10044
rect 5997 10007 6055 10013
rect 6012 9976 6040 10007
rect 6730 10004 6736 10016
rect 6788 10004 6794 10056
rect 7742 10044 7748 10056
rect 7703 10016 7748 10044
rect 7742 10004 7748 10016
rect 7800 10004 7806 10056
rect 8045 10053 8073 10084
rect 7838 10047 7896 10053
rect 7838 10013 7850 10047
rect 7884 10013 7896 10047
rect 7838 10007 7896 10013
rect 8021 10047 8079 10053
rect 8021 10013 8033 10047
rect 8067 10013 8079 10047
rect 8021 10007 8079 10013
rect 8210 10047 8268 10053
rect 8210 10013 8222 10047
rect 8256 10044 8268 10047
rect 8478 10044 8484 10056
rect 8256 10016 8484 10044
rect 8256 10013 8268 10016
rect 8210 10007 8268 10013
rect 7009 9979 7067 9985
rect 6012 9948 6960 9976
rect 4856 9880 5948 9908
rect 4856 9868 4862 9880
rect 6086 9868 6092 9920
rect 6144 9908 6150 9920
rect 6825 9911 6883 9917
rect 6825 9908 6837 9911
rect 6144 9880 6837 9908
rect 6144 9868 6150 9880
rect 6825 9877 6837 9880
rect 6871 9877 6883 9911
rect 6932 9908 6960 9948
rect 7009 9945 7021 9979
rect 7055 9976 7067 9979
rect 7466 9976 7472 9988
rect 7055 9948 7472 9976
rect 7055 9945 7067 9948
rect 7009 9939 7067 9945
rect 7466 9936 7472 9948
rect 7524 9936 7530 9988
rect 7282 9908 7288 9920
rect 6932 9880 7288 9908
rect 6825 9871 6883 9877
rect 7282 9868 7288 9880
rect 7340 9868 7346 9920
rect 7853 9908 7881 10007
rect 8478 10004 8484 10016
rect 8536 10004 8542 10056
rect 8110 9976 8116 9988
rect 8071 9948 8116 9976
rect 8110 9936 8116 9948
rect 8168 9936 8174 9988
rect 8478 9908 8484 9920
rect 7853 9880 8484 9908
rect 8478 9868 8484 9880
rect 8536 9868 8542 9920
rect 8588 9908 8616 10084
rect 8680 9976 8708 10152
rect 9232 10044 9260 10220
rect 9950 10208 9956 10220
rect 10008 10208 10014 10260
rect 10873 10251 10931 10257
rect 10873 10217 10885 10251
rect 10919 10248 10931 10251
rect 11698 10248 11704 10260
rect 10919 10220 11704 10248
rect 10919 10217 10931 10220
rect 10873 10211 10931 10217
rect 11698 10208 11704 10220
rect 11756 10208 11762 10260
rect 11977 10251 12035 10257
rect 11977 10217 11989 10251
rect 12023 10248 12035 10251
rect 12342 10248 12348 10260
rect 12023 10220 12348 10248
rect 12023 10217 12035 10220
rect 11977 10211 12035 10217
rect 12342 10208 12348 10220
rect 12400 10208 12406 10260
rect 12437 10251 12495 10257
rect 12437 10217 12449 10251
rect 12483 10248 12495 10251
rect 12710 10248 12716 10260
rect 12483 10220 12716 10248
rect 12483 10217 12495 10220
rect 12437 10211 12495 10217
rect 12710 10208 12716 10220
rect 12768 10208 12774 10260
rect 13170 10248 13176 10260
rect 12820 10220 13176 10248
rect 9306 10140 9312 10192
rect 9364 10140 9370 10192
rect 10321 10183 10379 10189
rect 10321 10149 10333 10183
rect 10367 10180 10379 10183
rect 12526 10180 12532 10192
rect 10367 10152 12532 10180
rect 10367 10149 10379 10152
rect 10321 10143 10379 10149
rect 12526 10140 12532 10152
rect 12584 10140 12590 10192
rect 9324 10112 9352 10140
rect 9585 10115 9643 10121
rect 9585 10112 9597 10115
rect 9324 10084 9597 10112
rect 9585 10081 9597 10084
rect 9631 10081 9643 10115
rect 11606 10112 11612 10124
rect 11567 10084 11612 10112
rect 9585 10075 9643 10081
rect 11606 10072 11612 10084
rect 11664 10072 11670 10124
rect 11698 10072 11704 10124
rect 11756 10112 11762 10124
rect 12618 10112 12624 10124
rect 11756 10084 11801 10112
rect 12579 10084 12624 10112
rect 11756 10072 11762 10084
rect 12618 10072 12624 10084
rect 12676 10072 12682 10124
rect 12713 10115 12771 10121
rect 12713 10081 12725 10115
rect 12759 10112 12771 10115
rect 12820 10112 12848 10220
rect 13170 10208 13176 10220
rect 13228 10208 13234 10260
rect 13630 10248 13636 10260
rect 13591 10220 13636 10248
rect 13630 10208 13636 10220
rect 13688 10208 13694 10260
rect 14642 10248 14648 10260
rect 14603 10220 14648 10248
rect 14642 10208 14648 10220
rect 14700 10208 14706 10260
rect 17681 10251 17739 10257
rect 17681 10217 17693 10251
rect 17727 10248 17739 10251
rect 18414 10248 18420 10260
rect 17727 10220 18420 10248
rect 17727 10217 17739 10220
rect 17681 10211 17739 10217
rect 18414 10208 18420 10220
rect 18472 10208 18478 10260
rect 18598 10208 18604 10260
rect 18656 10248 18662 10260
rect 18785 10251 18843 10257
rect 18785 10248 18797 10251
rect 18656 10220 18797 10248
rect 18656 10208 18662 10220
rect 18785 10217 18797 10220
rect 18831 10217 18843 10251
rect 19610 10248 19616 10260
rect 19571 10220 19616 10248
rect 18785 10211 18843 10217
rect 19610 10208 19616 10220
rect 19668 10208 19674 10260
rect 20708 10251 20766 10257
rect 20708 10248 20720 10251
rect 20645 10220 20720 10248
rect 16025 10183 16083 10189
rect 16025 10149 16037 10183
rect 16071 10180 16083 10183
rect 16666 10180 16672 10192
rect 16071 10152 16672 10180
rect 16071 10149 16083 10152
rect 16025 10143 16083 10149
rect 16666 10140 16672 10152
rect 16724 10140 16730 10192
rect 20645 10180 20673 10220
rect 20708 10217 20720 10220
rect 20754 10217 20766 10251
rect 20898 10248 20904 10260
rect 20859 10220 20904 10248
rect 20708 10211 20766 10217
rect 20898 10208 20904 10220
rect 20956 10248 20962 10260
rect 21174 10248 21180 10260
rect 20956 10220 21180 10248
rect 20956 10208 20962 10220
rect 21174 10208 21180 10220
rect 21232 10208 21238 10260
rect 21266 10180 21272 10192
rect 18616 10152 20116 10180
rect 20645 10152 21272 10180
rect 12759 10084 12848 10112
rect 12759 10081 12771 10084
rect 12713 10075 12771 10081
rect 12894 10072 12900 10124
rect 12952 10112 12958 10124
rect 13538 10112 13544 10124
rect 12952 10084 12997 10112
rect 13372 10084 13544 10112
rect 12952 10072 12958 10084
rect 9306 10044 9312 10056
rect 9219 10016 9312 10044
rect 9306 10004 9312 10016
rect 9364 10004 9370 10056
rect 9401 10047 9459 10053
rect 9401 10013 9413 10047
rect 9447 10013 9459 10047
rect 9401 10007 9459 10013
rect 9416 9976 9444 10007
rect 9490 10004 9496 10056
rect 9548 10044 9554 10056
rect 10781 10047 10839 10053
rect 9548 10016 9593 10044
rect 9548 10004 9554 10016
rect 10781 10013 10793 10047
rect 10827 10013 10839 10047
rect 10962 10044 10968 10056
rect 10923 10016 10968 10044
rect 10781 10007 10839 10013
rect 9858 9976 9864 9988
rect 8680 9948 9864 9976
rect 9858 9936 9864 9948
rect 9916 9936 9922 9988
rect 10796 9976 10824 10007
rect 10962 10004 10968 10016
rect 11020 10004 11026 10056
rect 11514 10044 11520 10056
rect 11475 10016 11520 10044
rect 11514 10004 11520 10016
rect 11572 10004 11578 10056
rect 11790 10004 11796 10056
rect 11848 10044 11854 10056
rect 12526 10044 12532 10056
rect 11848 10016 11893 10044
rect 11983 10016 12532 10044
rect 11848 10004 11854 10016
rect 11983 9976 12011 10016
rect 12526 10004 12532 10016
rect 12584 10004 12590 10056
rect 12806 10047 12864 10053
rect 12806 10013 12818 10047
rect 12852 10044 12864 10047
rect 13372 10044 13400 10084
rect 13538 10072 13544 10084
rect 13596 10072 13602 10124
rect 13630 10072 13636 10124
rect 13688 10112 13694 10124
rect 16114 10112 16120 10124
rect 13688 10084 15424 10112
rect 13688 10072 13694 10084
rect 12852 10016 13400 10044
rect 13449 10047 13507 10053
rect 12852 10013 12864 10016
rect 12806 10007 12864 10013
rect 13449 10013 13461 10047
rect 13495 10044 13507 10047
rect 13998 10044 14004 10056
rect 13495 10016 14004 10044
rect 13495 10013 13507 10016
rect 13449 10007 13507 10013
rect 13998 10004 14004 10016
rect 14056 10004 14062 10056
rect 14274 10044 14280 10056
rect 14235 10016 14280 10044
rect 14274 10004 14280 10016
rect 14332 10004 14338 10056
rect 15396 10053 15424 10084
rect 15764 10084 16120 10112
rect 15562 10053 15568 10056
rect 15381 10047 15439 10053
rect 15381 10013 15393 10047
rect 15427 10013 15439 10047
rect 15381 10007 15439 10013
rect 15529 10047 15568 10053
rect 15529 10013 15541 10047
rect 15529 10007 15568 10013
rect 15562 10004 15568 10007
rect 15620 10004 15626 10056
rect 15764 10053 15792 10084
rect 16114 10072 16120 10084
rect 16172 10112 16178 10124
rect 16390 10112 16396 10124
rect 16172 10084 16396 10112
rect 16172 10072 16178 10084
rect 16390 10072 16396 10084
rect 16448 10072 16454 10124
rect 17218 10072 17224 10124
rect 17276 10112 17282 10124
rect 18616 10112 18644 10152
rect 20088 10124 20116 10152
rect 21266 10140 21272 10152
rect 21324 10140 21330 10192
rect 17276 10084 18644 10112
rect 17276 10072 17282 10084
rect 19334 10072 19340 10124
rect 19392 10112 19398 10124
rect 19392 10084 19656 10112
rect 19392 10072 19398 10084
rect 15749 10047 15807 10053
rect 15749 10013 15761 10047
rect 15795 10013 15807 10047
rect 15749 10007 15807 10013
rect 15887 10047 15945 10053
rect 15887 10013 15899 10047
rect 15933 10044 15945 10047
rect 16758 10044 16764 10056
rect 15933 10016 16764 10044
rect 15933 10013 15945 10016
rect 15887 10007 15945 10013
rect 16758 10004 16764 10016
rect 16816 10044 16822 10056
rect 18325 10047 18383 10053
rect 18325 10044 18337 10047
rect 16816 10016 18337 10044
rect 16816 10004 16822 10016
rect 18325 10013 18337 10016
rect 18371 10013 18383 10047
rect 18325 10007 18383 10013
rect 18506 10004 18512 10056
rect 18564 10044 18570 10056
rect 18601 10047 18659 10053
rect 18601 10044 18613 10047
rect 18564 10016 18613 10044
rect 18564 10004 18570 10016
rect 18601 10013 18613 10016
rect 18647 10044 18659 10047
rect 18690 10044 18696 10056
rect 18647 10016 18696 10044
rect 18647 10013 18659 10016
rect 18601 10007 18659 10013
rect 18690 10004 18696 10016
rect 18748 10004 18754 10056
rect 19628 10053 19656 10084
rect 20070 10072 20076 10124
rect 20128 10112 20134 10124
rect 21361 10115 21419 10121
rect 21361 10112 21373 10115
rect 20128 10084 21373 10112
rect 20128 10072 20134 10084
rect 21361 10081 21373 10084
rect 21407 10081 21419 10115
rect 21361 10075 21419 10081
rect 19429 10047 19487 10053
rect 19429 10013 19441 10047
rect 19475 10013 19487 10047
rect 19429 10007 19487 10013
rect 19613 10047 19671 10053
rect 19613 10013 19625 10047
rect 19659 10013 19671 10047
rect 22465 10047 22523 10053
rect 22465 10044 22477 10047
rect 19613 10007 19671 10013
rect 19812 10016 22477 10044
rect 13814 9976 13820 9988
rect 10796 9948 12011 9976
rect 12452 9948 13820 9976
rect 10042 9908 10048 9920
rect 8588 9880 10048 9908
rect 10042 9868 10048 9880
rect 10100 9868 10106 9920
rect 10870 9868 10876 9920
rect 10928 9908 10934 9920
rect 12452 9908 12480 9948
rect 13814 9936 13820 9948
rect 13872 9976 13878 9988
rect 14461 9979 14519 9985
rect 14461 9976 14473 9979
rect 13872 9948 14473 9976
rect 13872 9936 13878 9948
rect 14461 9945 14473 9948
rect 14507 9976 14519 9979
rect 15286 9976 15292 9988
rect 14507 9948 15292 9976
rect 14507 9945 14519 9948
rect 14461 9939 14519 9945
rect 15286 9936 15292 9948
rect 15344 9936 15350 9988
rect 15654 9976 15660 9988
rect 15615 9948 15660 9976
rect 15654 9936 15660 9948
rect 15712 9936 15718 9988
rect 16482 9976 16488 9988
rect 16443 9948 16488 9976
rect 16482 9936 16488 9948
rect 16540 9936 16546 9988
rect 17126 9976 17132 9988
rect 17087 9948 17132 9976
rect 17126 9936 17132 9948
rect 17184 9936 17190 9988
rect 17402 9976 17408 9988
rect 17363 9948 17408 9976
rect 17402 9936 17408 9948
rect 17460 9936 17466 9988
rect 17497 9979 17555 9985
rect 17497 9945 17509 9979
rect 17543 9976 17555 9979
rect 18874 9976 18880 9988
rect 17543 9948 18880 9976
rect 17543 9945 17555 9948
rect 17497 9939 17555 9945
rect 18874 9936 18880 9948
rect 18932 9936 18938 9988
rect 19444 9976 19472 10007
rect 19702 9976 19708 9988
rect 19444 9948 19708 9976
rect 19702 9936 19708 9948
rect 19760 9936 19766 9988
rect 10928 9880 12480 9908
rect 10928 9868 10934 9880
rect 12526 9868 12532 9920
rect 12584 9908 12590 9920
rect 12802 9908 12808 9920
rect 12584 9880 12808 9908
rect 12584 9868 12590 9880
rect 12802 9868 12808 9880
rect 12860 9908 12866 9920
rect 13630 9908 13636 9920
rect 12860 9880 13636 9908
rect 12860 9868 12866 9880
rect 13630 9868 13636 9880
rect 13688 9868 13694 9920
rect 16758 9868 16764 9920
rect 16816 9908 16822 9920
rect 17218 9908 17224 9920
rect 16816 9880 17224 9908
rect 16816 9868 16822 9880
rect 17218 9868 17224 9880
rect 17276 9908 17282 9920
rect 17313 9911 17371 9917
rect 17313 9908 17325 9911
rect 17276 9880 17325 9908
rect 17276 9868 17282 9880
rect 17313 9877 17325 9880
rect 17359 9877 17371 9911
rect 17313 9871 17371 9877
rect 17678 9868 17684 9920
rect 17736 9908 17742 9920
rect 18417 9911 18475 9917
rect 18417 9908 18429 9911
rect 17736 9880 18429 9908
rect 17736 9868 17742 9880
rect 18417 9877 18429 9880
rect 18463 9877 18475 9911
rect 18417 9871 18475 9877
rect 19426 9868 19432 9920
rect 19484 9908 19490 9920
rect 19812 9908 19840 10016
rect 22465 10013 22477 10016
rect 22511 10013 22523 10047
rect 22465 10007 22523 10013
rect 20254 9936 20260 9988
rect 20312 9976 20318 9988
rect 20533 9979 20591 9985
rect 20533 9976 20545 9979
rect 20312 9948 20545 9976
rect 20312 9936 20318 9948
rect 20533 9945 20545 9948
rect 20579 9945 20591 9979
rect 20533 9939 20591 9945
rect 19484 9880 19840 9908
rect 19484 9868 19490 9880
rect 20438 9868 20444 9920
rect 20496 9908 20502 9920
rect 20733 9911 20791 9917
rect 20733 9908 20745 9911
rect 20496 9880 20745 9908
rect 20496 9868 20502 9880
rect 20733 9877 20745 9880
rect 20779 9877 20791 9911
rect 20733 9871 20791 9877
rect 21450 9868 21456 9920
rect 21508 9908 21514 9920
rect 21913 9911 21971 9917
rect 21913 9908 21925 9911
rect 21508 9880 21925 9908
rect 21508 9868 21514 9880
rect 21913 9877 21925 9880
rect 21959 9877 21971 9911
rect 23106 9908 23112 9920
rect 23067 9880 23112 9908
rect 21913 9871 21971 9877
rect 23106 9868 23112 9880
rect 23164 9868 23170 9920
rect 1104 9818 23987 9840
rect 1104 9766 6630 9818
rect 6682 9766 6694 9818
rect 6746 9766 6758 9818
rect 6810 9766 6822 9818
rect 6874 9766 6886 9818
rect 6938 9766 12311 9818
rect 12363 9766 12375 9818
rect 12427 9766 12439 9818
rect 12491 9766 12503 9818
rect 12555 9766 12567 9818
rect 12619 9766 17992 9818
rect 18044 9766 18056 9818
rect 18108 9766 18120 9818
rect 18172 9766 18184 9818
rect 18236 9766 18248 9818
rect 18300 9766 23673 9818
rect 23725 9766 23737 9818
rect 23789 9766 23801 9818
rect 23853 9766 23865 9818
rect 23917 9766 23929 9818
rect 23981 9766 23987 9818
rect 1104 9744 23987 9766
rect 1946 9704 1952 9716
rect 1907 9676 1952 9704
rect 1946 9664 1952 9676
rect 2004 9664 2010 9716
rect 4246 9664 4252 9716
rect 4304 9704 4310 9716
rect 4525 9707 4583 9713
rect 4525 9704 4537 9707
rect 4304 9676 4537 9704
rect 4304 9664 4310 9676
rect 4525 9673 4537 9676
rect 4571 9673 4583 9707
rect 4525 9667 4583 9673
rect 5810 9664 5816 9716
rect 5868 9704 5874 9716
rect 5997 9707 6055 9713
rect 5997 9704 6009 9707
rect 5868 9676 6009 9704
rect 5868 9664 5874 9676
rect 5997 9673 6009 9676
rect 6043 9673 6055 9707
rect 5997 9667 6055 9673
rect 7282 9664 7288 9716
rect 7340 9664 7346 9716
rect 11149 9707 11207 9713
rect 11149 9673 11161 9707
rect 11195 9704 11207 9707
rect 11422 9704 11428 9716
rect 11195 9676 11428 9704
rect 11195 9673 11207 9676
rect 11149 9667 11207 9673
rect 11422 9664 11428 9676
rect 11480 9704 11486 9716
rect 11606 9704 11612 9716
rect 11480 9676 11612 9704
rect 11480 9664 11486 9676
rect 11606 9664 11612 9676
rect 11664 9664 11670 9716
rect 12618 9664 12624 9716
rect 12676 9704 12682 9716
rect 12986 9704 12992 9716
rect 12676 9676 12992 9704
rect 12676 9664 12682 9676
rect 12986 9664 12992 9676
rect 13044 9664 13050 9716
rect 13170 9664 13176 9716
rect 13228 9704 13234 9716
rect 13354 9704 13360 9716
rect 13228 9676 13360 9704
rect 13228 9664 13234 9676
rect 13354 9664 13360 9676
rect 13412 9664 13418 9716
rect 13906 9664 13912 9716
rect 13964 9704 13970 9716
rect 15562 9704 15568 9716
rect 13964 9676 15568 9704
rect 13964 9664 13970 9676
rect 15562 9664 15568 9676
rect 15620 9704 15626 9716
rect 15746 9704 15752 9716
rect 15620 9676 15752 9704
rect 15620 9664 15626 9676
rect 15746 9664 15752 9676
rect 15804 9664 15810 9716
rect 16114 9664 16120 9716
rect 16172 9704 16178 9716
rect 17402 9704 17408 9716
rect 16172 9676 17408 9704
rect 16172 9664 16178 9676
rect 17402 9664 17408 9676
rect 17460 9664 17466 9716
rect 17497 9707 17555 9713
rect 17497 9673 17509 9707
rect 17543 9673 17555 9707
rect 17497 9667 17555 9673
rect 2774 9636 2780 9648
rect 2516 9608 2780 9636
rect 2516 9577 2544 9608
rect 2774 9596 2780 9608
rect 2832 9636 2838 9648
rect 3329 9639 3387 9645
rect 3329 9636 3341 9639
rect 2832 9608 3341 9636
rect 2832 9596 2838 9608
rect 3329 9605 3341 9608
rect 3375 9636 3387 9639
rect 3510 9636 3516 9648
rect 3375 9608 3516 9636
rect 3375 9605 3387 9608
rect 3329 9599 3387 9605
rect 3510 9596 3516 9608
rect 3568 9596 3574 9648
rect 6454 9596 6460 9648
rect 6512 9636 6518 9648
rect 7300 9636 7328 9664
rect 7742 9636 7748 9648
rect 6512 9608 7052 9636
rect 6512 9596 6518 9608
rect 2501 9571 2559 9577
rect 2501 9537 2513 9571
rect 2547 9537 2559 9571
rect 2501 9531 2559 9537
rect 2590 9528 2596 9580
rect 2648 9568 2654 9580
rect 4338 9568 4344 9580
rect 2648 9540 2693 9568
rect 2746 9540 4344 9568
rect 2648 9528 2654 9540
rect 1946 9460 1952 9512
rect 2004 9500 2010 9512
rect 2746 9500 2774 9540
rect 4338 9528 4344 9540
rect 4396 9528 4402 9580
rect 4982 9528 4988 9580
rect 5040 9568 5046 9580
rect 5353 9571 5411 9577
rect 5353 9568 5365 9571
rect 5040 9540 5365 9568
rect 5040 9528 5046 9540
rect 5353 9537 5365 9540
rect 5399 9537 5411 9571
rect 5353 9531 5411 9537
rect 5718 9528 5724 9580
rect 5776 9568 5782 9580
rect 5813 9571 5871 9577
rect 5813 9568 5825 9571
rect 5776 9540 5825 9568
rect 5776 9528 5782 9540
rect 5813 9537 5825 9540
rect 5859 9537 5871 9571
rect 5813 9531 5871 9537
rect 6733 9571 6791 9577
rect 6733 9537 6745 9571
rect 6779 9568 6791 9571
rect 6822 9568 6828 9580
rect 6779 9540 6828 9568
rect 6779 9537 6791 9540
rect 6733 9531 6791 9537
rect 6822 9528 6828 9540
rect 6880 9528 6886 9580
rect 7024 9577 7052 9608
rect 7116 9608 7748 9636
rect 7116 9577 7144 9608
rect 7742 9596 7748 9608
rect 7800 9636 7806 9648
rect 10226 9636 10232 9648
rect 7800 9608 10232 9636
rect 7800 9596 7806 9608
rect 10226 9596 10232 9608
rect 10284 9596 10290 9648
rect 11054 9596 11060 9648
rect 11112 9636 11118 9648
rect 12529 9639 12587 9645
rect 12529 9636 12541 9639
rect 11112 9608 12541 9636
rect 11112 9596 11118 9608
rect 12529 9605 12541 9608
rect 12575 9605 12587 9639
rect 14550 9636 14556 9648
rect 12529 9599 12587 9605
rect 12912 9608 14556 9636
rect 7009 9571 7067 9577
rect 7009 9537 7021 9571
rect 7055 9537 7067 9571
rect 7009 9531 7067 9537
rect 7101 9571 7159 9577
rect 7101 9537 7113 9571
rect 7147 9537 7159 9571
rect 7282 9568 7288 9580
rect 7243 9540 7288 9568
rect 7101 9531 7159 9537
rect 7282 9528 7288 9540
rect 7340 9528 7346 9580
rect 7374 9528 7380 9580
rect 7432 9568 7438 9580
rect 10042 9568 10048 9580
rect 7432 9540 10048 9568
rect 7432 9528 7438 9540
rect 10042 9528 10048 9540
rect 10100 9568 10106 9580
rect 10137 9571 10195 9577
rect 10137 9568 10149 9571
rect 10100 9540 10149 9568
rect 10100 9528 10106 9540
rect 10137 9537 10149 9540
rect 10183 9537 10195 9571
rect 10318 9568 10324 9580
rect 10279 9540 10324 9568
rect 10137 9531 10195 9537
rect 10318 9528 10324 9540
rect 10376 9528 10382 9580
rect 11606 9528 11612 9580
rect 11664 9568 11670 9580
rect 11793 9571 11851 9577
rect 11793 9568 11805 9571
rect 11664 9540 11805 9568
rect 11664 9528 11670 9540
rect 11793 9537 11805 9540
rect 11839 9537 11851 9571
rect 11793 9531 11851 9537
rect 12434 9528 12440 9580
rect 12492 9568 12498 9580
rect 12912 9577 12940 9608
rect 14550 9596 14556 9608
rect 14608 9596 14614 9648
rect 17512 9636 17540 9667
rect 18230 9664 18236 9716
rect 18288 9704 18294 9716
rect 18598 9704 18604 9716
rect 18288 9676 18604 9704
rect 18288 9664 18294 9676
rect 18598 9664 18604 9676
rect 18656 9664 18662 9716
rect 19426 9664 19432 9716
rect 19484 9704 19490 9716
rect 19484 9676 19564 9704
rect 19484 9664 19490 9676
rect 14844 9608 17540 9636
rect 12759 9571 12817 9577
rect 12759 9568 12771 9571
rect 12492 9540 12771 9568
rect 12492 9528 12498 9540
rect 12759 9537 12771 9540
rect 12805 9537 12817 9571
rect 12759 9531 12817 9537
rect 12878 9571 12940 9577
rect 12878 9537 12890 9571
rect 12924 9540 12940 9571
rect 12924 9537 12936 9540
rect 12878 9531 12936 9537
rect 12986 9528 12992 9580
rect 13044 9568 13050 9580
rect 13173 9571 13231 9577
rect 13044 9540 13089 9568
rect 13044 9528 13050 9540
rect 13173 9537 13185 9571
rect 13219 9537 13231 9571
rect 13173 9531 13231 9537
rect 2004 9472 2774 9500
rect 2004 9460 2010 9472
rect 5074 9460 5080 9512
rect 5132 9500 5138 9512
rect 5629 9503 5687 9509
rect 5629 9500 5641 9503
rect 5132 9472 5641 9500
rect 5132 9460 5138 9472
rect 5629 9469 5641 9472
rect 5675 9500 5687 9503
rect 6362 9500 6368 9512
rect 5675 9472 6368 9500
rect 5675 9469 5687 9472
rect 5629 9463 5687 9469
rect 6362 9460 6368 9472
rect 6420 9460 6426 9512
rect 6917 9503 6975 9509
rect 6917 9500 6929 9503
rect 6722 9472 6929 9500
rect 2777 9435 2835 9441
rect 2777 9401 2789 9435
rect 2823 9432 2835 9435
rect 3234 9432 3240 9444
rect 2823 9404 3240 9432
rect 2823 9401 2835 9404
rect 2777 9395 2835 9401
rect 3234 9392 3240 9404
rect 3292 9432 3298 9444
rect 5258 9432 5264 9444
rect 3292 9404 5264 9432
rect 3292 9392 3298 9404
rect 5258 9392 5264 9404
rect 5316 9392 5322 9444
rect 6722 9432 6750 9472
rect 6917 9469 6929 9472
rect 6963 9469 6975 9503
rect 6917 9463 6975 9469
rect 8110 9460 8116 9512
rect 8168 9500 8174 9512
rect 8849 9503 8907 9509
rect 8849 9500 8861 9503
rect 8168 9472 8861 9500
rect 8168 9460 8174 9472
rect 8849 9469 8861 9472
rect 8895 9469 8907 9503
rect 10502 9500 10508 9512
rect 10463 9472 10508 9500
rect 8849 9463 8907 9469
rect 10502 9460 10508 9472
rect 10560 9460 10566 9512
rect 10962 9460 10968 9512
rect 11020 9500 11026 9512
rect 11974 9500 11980 9512
rect 11020 9472 11980 9500
rect 11020 9460 11026 9472
rect 11974 9460 11980 9472
rect 12032 9460 12038 9512
rect 12069 9503 12127 9509
rect 12069 9469 12081 9503
rect 12115 9469 12127 9503
rect 12069 9463 12127 9469
rect 5460 9404 6750 9432
rect 3050 9324 3056 9376
rect 3108 9364 3114 9376
rect 3605 9367 3663 9373
rect 3605 9364 3617 9367
rect 3108 9336 3617 9364
rect 3108 9324 3114 9336
rect 3605 9333 3617 9336
rect 3651 9364 3663 9367
rect 3694 9364 3700 9376
rect 3651 9336 3700 9364
rect 3651 9333 3663 9336
rect 3605 9327 3663 9333
rect 3694 9324 3700 9336
rect 3752 9324 3758 9376
rect 4246 9324 4252 9376
rect 4304 9364 4310 9376
rect 5460 9373 5488 9404
rect 7006 9392 7012 9444
rect 7064 9432 7070 9444
rect 8297 9435 8355 9441
rect 8297 9432 8309 9435
rect 7064 9404 8309 9432
rect 7064 9392 7070 9404
rect 8297 9401 8309 9404
rect 8343 9401 8355 9435
rect 12084 9432 12112 9463
rect 13188 9432 13216 9531
rect 13538 9528 13544 9580
rect 13596 9568 13602 9580
rect 13725 9571 13783 9577
rect 13725 9568 13737 9571
rect 13596 9540 13737 9568
rect 13596 9528 13602 9540
rect 13725 9537 13737 9540
rect 13771 9537 13783 9571
rect 13725 9531 13783 9537
rect 13909 9571 13967 9577
rect 13909 9537 13921 9571
rect 13955 9537 13967 9571
rect 14642 9568 14648 9580
rect 14603 9540 14648 9568
rect 13909 9531 13967 9537
rect 13924 9500 13952 9531
rect 14642 9528 14648 9540
rect 14700 9528 14706 9580
rect 14844 9577 14872 9608
rect 17586 9596 17592 9648
rect 17644 9636 17650 9648
rect 17773 9639 17831 9645
rect 17773 9636 17785 9639
rect 17644 9608 17785 9636
rect 17644 9596 17650 9608
rect 17773 9605 17785 9608
rect 17819 9605 17831 9639
rect 18414 9636 18420 9648
rect 17773 9599 17831 9605
rect 18064 9608 18420 9636
rect 14737 9571 14795 9577
rect 14737 9537 14749 9571
rect 14783 9537 14795 9571
rect 14737 9531 14795 9537
rect 14829 9571 14887 9577
rect 14829 9537 14841 9571
rect 14875 9537 14887 9571
rect 14829 9531 14887 9537
rect 15013 9571 15071 9577
rect 15013 9537 15025 9571
rect 15059 9537 15071 9571
rect 15013 9531 15071 9537
rect 14752 9500 14780 9531
rect 15028 9500 15056 9531
rect 15378 9528 15384 9580
rect 15436 9568 15442 9580
rect 15657 9571 15715 9577
rect 15657 9568 15669 9571
rect 15436 9540 15669 9568
rect 15436 9528 15442 9540
rect 15657 9537 15669 9540
rect 15703 9537 15715 9571
rect 16117 9571 16175 9577
rect 16117 9542 16129 9571
rect 16163 9542 16175 9571
rect 17681 9571 17739 9577
rect 15657 9531 15715 9537
rect 15488 9500 15576 9511
rect 15841 9503 15899 9509
rect 13924 9472 14872 9500
rect 15028 9483 15608 9500
rect 15028 9472 15516 9483
rect 15548 9472 15608 9483
rect 14642 9432 14648 9444
rect 12084 9404 12572 9432
rect 13188 9404 14648 9432
rect 8297 9395 8355 9401
rect 5445 9367 5503 9373
rect 5445 9364 5457 9367
rect 4304 9336 5457 9364
rect 4304 9324 4310 9336
rect 5445 9333 5457 9336
rect 5491 9333 5503 9367
rect 6546 9364 6552 9376
rect 6507 9336 6552 9364
rect 5445 9327 5503 9333
rect 6546 9324 6552 9336
rect 6604 9324 6610 9376
rect 7558 9324 7564 9376
rect 7616 9364 7622 9376
rect 7834 9364 7840 9376
rect 7616 9336 7840 9364
rect 7616 9324 7622 9336
rect 7834 9324 7840 9336
rect 7892 9324 7898 9376
rect 8846 9324 8852 9376
rect 8904 9364 8910 9376
rect 9398 9364 9404 9376
rect 8904 9336 9404 9364
rect 8904 9324 8910 9336
rect 9398 9324 9404 9336
rect 9456 9324 9462 9376
rect 9677 9367 9735 9373
rect 9677 9333 9689 9367
rect 9723 9364 9735 9367
rect 9858 9364 9864 9376
rect 9723 9336 9864 9364
rect 9723 9333 9735 9336
rect 9677 9327 9735 9333
rect 9858 9324 9864 9336
rect 9916 9364 9922 9376
rect 10594 9364 10600 9376
rect 9916 9336 10600 9364
rect 9916 9324 9922 9336
rect 10594 9324 10600 9336
rect 10652 9324 10658 9376
rect 11882 9364 11888 9376
rect 11843 9336 11888 9364
rect 11882 9324 11888 9336
rect 11940 9324 11946 9376
rect 11974 9324 11980 9376
rect 12032 9364 12038 9376
rect 12544 9364 12572 9404
rect 14642 9392 14648 9404
rect 14700 9392 14706 9444
rect 13354 9364 13360 9376
rect 12032 9336 12077 9364
rect 12544 9336 13360 9364
rect 12032 9324 12038 9336
rect 13354 9324 13360 9336
rect 13412 9324 13418 9376
rect 13906 9364 13912 9376
rect 13867 9336 13912 9364
rect 13906 9324 13912 9336
rect 13964 9324 13970 9376
rect 14369 9367 14427 9373
rect 14369 9333 14381 9367
rect 14415 9364 14427 9367
rect 14734 9364 14740 9376
rect 14415 9336 14740 9364
rect 14415 9333 14427 9336
rect 14369 9327 14427 9333
rect 14734 9324 14740 9336
rect 14792 9324 14798 9376
rect 14844 9364 14872 9472
rect 15473 9367 15531 9373
rect 15473 9364 15485 9367
rect 14844 9336 15485 9364
rect 15473 9333 15485 9336
rect 15519 9333 15531 9367
rect 15580 9364 15608 9472
rect 15841 9469 15853 9503
rect 15887 9469 15899 9503
rect 15841 9463 15899 9469
rect 15746 9432 15752 9444
rect 15707 9404 15752 9432
rect 15746 9392 15752 9404
rect 15804 9392 15810 9444
rect 15856 9432 15884 9463
rect 15930 9460 15936 9512
rect 15988 9500 15994 9512
rect 15988 9472 16033 9500
rect 16114 9490 16120 9542
rect 16172 9490 16178 9542
rect 17681 9537 17693 9571
rect 17727 9537 17739 9571
rect 17862 9568 17868 9580
rect 17823 9540 17868 9568
rect 17681 9531 17739 9537
rect 15988 9460 15994 9472
rect 16482 9460 16488 9512
rect 16540 9500 16546 9512
rect 16853 9503 16911 9509
rect 16853 9500 16865 9503
rect 16540 9472 16865 9500
rect 16540 9460 16546 9472
rect 16853 9469 16865 9472
rect 16899 9500 16911 9503
rect 17218 9500 17224 9512
rect 16899 9472 17224 9500
rect 16899 9469 16911 9472
rect 16853 9463 16911 9469
rect 17218 9460 17224 9472
rect 17276 9460 17282 9512
rect 17696 9500 17724 9531
rect 17862 9528 17868 9540
rect 17920 9568 17926 9580
rect 17954 9568 17960 9580
rect 17920 9540 17960 9568
rect 17920 9528 17926 9540
rect 17954 9528 17960 9540
rect 18012 9528 18018 9580
rect 18064 9577 18092 9608
rect 18414 9596 18420 9608
rect 18472 9596 18478 9648
rect 18049 9571 18107 9577
rect 18049 9537 18061 9571
rect 18095 9537 18107 9571
rect 18049 9531 18107 9537
rect 18141 9571 18199 9577
rect 18141 9537 18153 9571
rect 18187 9568 18199 9571
rect 18322 9568 18328 9580
rect 18187 9540 18328 9568
rect 18187 9537 18199 9540
rect 18141 9531 18199 9537
rect 18322 9528 18328 9540
rect 18380 9528 18386 9580
rect 18598 9528 18604 9580
rect 18656 9568 18662 9580
rect 19150 9568 19156 9580
rect 18656 9540 19156 9568
rect 18656 9528 18662 9540
rect 19150 9528 19156 9540
rect 19208 9528 19214 9580
rect 19536 9577 19564 9676
rect 19613 9639 19671 9645
rect 19613 9605 19625 9639
rect 19659 9636 19671 9639
rect 20438 9636 20444 9648
rect 19659 9608 20444 9636
rect 19659 9605 19671 9608
rect 19613 9599 19671 9605
rect 19521 9571 19579 9577
rect 19521 9537 19533 9571
rect 19567 9537 19579 9571
rect 19521 9531 19579 9537
rect 19242 9500 19248 9512
rect 17696 9472 19248 9500
rect 19242 9460 19248 9472
rect 19300 9460 19306 9512
rect 16390 9432 16396 9444
rect 15856 9404 16396 9432
rect 16390 9392 16396 9404
rect 16448 9432 16454 9444
rect 16574 9432 16580 9444
rect 16448 9404 16580 9432
rect 16448 9392 16454 9404
rect 16574 9392 16580 9404
rect 16632 9392 16638 9444
rect 17586 9392 17592 9444
rect 17644 9432 17650 9444
rect 19334 9432 19340 9444
rect 17644 9404 19340 9432
rect 17644 9392 17650 9404
rect 19334 9392 19340 9404
rect 19392 9392 19398 9444
rect 19628 9432 19656 9599
rect 20438 9596 20444 9608
rect 20496 9596 20502 9648
rect 19705 9571 19763 9577
rect 19705 9537 19717 9571
rect 19751 9537 19763 9571
rect 19705 9531 19763 9537
rect 19720 9500 19748 9531
rect 19886 9528 19892 9580
rect 19944 9568 19950 9580
rect 20346 9577 20352 9580
rect 20165 9571 20223 9577
rect 20165 9568 20177 9571
rect 19944 9540 20177 9568
rect 19944 9528 19950 9540
rect 20165 9537 20177 9540
rect 20211 9537 20223 9571
rect 20165 9531 20223 9537
rect 20313 9571 20352 9577
rect 20313 9537 20325 9571
rect 20313 9531 20352 9537
rect 20070 9500 20076 9512
rect 19720 9472 20076 9500
rect 20070 9460 20076 9472
rect 20128 9460 20134 9512
rect 20180 9500 20208 9531
rect 20346 9528 20352 9531
rect 20404 9528 20410 9580
rect 20530 9568 20536 9580
rect 20491 9540 20536 9568
rect 20530 9528 20536 9540
rect 20588 9528 20594 9580
rect 20671 9571 20729 9577
rect 20671 9537 20683 9571
rect 20717 9568 20729 9571
rect 20717 9540 21128 9568
rect 20717 9537 20729 9540
rect 20671 9531 20729 9537
rect 21100 9500 21128 9540
rect 21174 9528 21180 9580
rect 21232 9568 21238 9580
rect 22005 9571 22063 9577
rect 22005 9568 22017 9571
rect 21232 9540 22017 9568
rect 21232 9528 21238 9540
rect 22005 9537 22017 9540
rect 22051 9537 22063 9571
rect 22005 9531 22063 9537
rect 22097 9571 22155 9577
rect 22097 9537 22109 9571
rect 22143 9568 22155 9571
rect 22186 9568 22192 9580
rect 22143 9540 22192 9568
rect 22143 9537 22155 9540
rect 22097 9531 22155 9537
rect 22186 9528 22192 9540
rect 22244 9528 22250 9580
rect 23014 9568 23020 9580
rect 22975 9540 23020 9568
rect 23014 9528 23020 9540
rect 23072 9528 23078 9580
rect 21726 9500 21732 9512
rect 20180 9472 21036 9500
rect 21100 9472 21732 9500
rect 20438 9432 20444 9444
rect 19628 9404 20444 9432
rect 20438 9392 20444 9404
rect 20496 9392 20502 9444
rect 20714 9392 20720 9444
rect 20772 9432 20778 9444
rect 20809 9435 20867 9441
rect 20809 9432 20821 9435
rect 20772 9404 20821 9432
rect 20772 9392 20778 9404
rect 20809 9401 20821 9404
rect 20855 9401 20867 9435
rect 21008 9432 21036 9472
rect 21726 9460 21732 9472
rect 21784 9460 21790 9512
rect 22281 9503 22339 9509
rect 22281 9469 22293 9503
rect 22327 9500 22339 9503
rect 22462 9500 22468 9512
rect 22327 9472 22468 9500
rect 22327 9469 22339 9472
rect 22281 9463 22339 9469
rect 22462 9460 22468 9472
rect 22520 9460 22526 9512
rect 22370 9432 22376 9444
rect 21008 9404 22376 9432
rect 20809 9395 20867 9401
rect 22370 9392 22376 9404
rect 22428 9432 22434 9444
rect 22833 9435 22891 9441
rect 22833 9432 22845 9435
rect 22428 9404 22845 9432
rect 22428 9392 22434 9404
rect 22833 9401 22845 9404
rect 22879 9401 22891 9435
rect 22833 9395 22891 9401
rect 18598 9364 18604 9376
rect 15580 9336 18604 9364
rect 15473 9327 15531 9333
rect 18598 9324 18604 9336
rect 18656 9324 18662 9376
rect 19242 9324 19248 9376
rect 19300 9364 19306 9376
rect 19610 9364 19616 9376
rect 19300 9336 19616 9364
rect 19300 9324 19306 9336
rect 19610 9324 19616 9336
rect 19668 9324 19674 9376
rect 21174 9324 21180 9376
rect 21232 9364 21238 9376
rect 21269 9367 21327 9373
rect 21269 9364 21281 9367
rect 21232 9336 21281 9364
rect 21232 9324 21238 9336
rect 21269 9333 21281 9336
rect 21315 9364 21327 9367
rect 21450 9364 21456 9376
rect 21315 9336 21456 9364
rect 21315 9333 21327 9336
rect 21269 9327 21327 9333
rect 21450 9324 21456 9336
rect 21508 9324 21514 9376
rect 22186 9324 22192 9376
rect 22244 9364 22250 9376
rect 22244 9336 22289 9364
rect 22244 9324 22250 9336
rect 1104 9274 23828 9296
rect 1104 9222 3790 9274
rect 3842 9222 3854 9274
rect 3906 9222 3918 9274
rect 3970 9222 3982 9274
rect 4034 9222 4046 9274
rect 4098 9222 9471 9274
rect 9523 9222 9535 9274
rect 9587 9222 9599 9274
rect 9651 9222 9663 9274
rect 9715 9222 9727 9274
rect 9779 9222 15152 9274
rect 15204 9222 15216 9274
rect 15268 9222 15280 9274
rect 15332 9222 15344 9274
rect 15396 9222 15408 9274
rect 15460 9222 20833 9274
rect 20885 9222 20897 9274
rect 20949 9222 20961 9274
rect 21013 9222 21025 9274
rect 21077 9222 21089 9274
rect 21141 9222 23828 9274
rect 1104 9200 23828 9222
rect 3418 9120 3424 9172
rect 3476 9160 3482 9172
rect 3970 9160 3976 9172
rect 3476 9132 3976 9160
rect 3476 9120 3482 9132
rect 3970 9120 3976 9132
rect 4028 9160 4034 9172
rect 4433 9163 4491 9169
rect 4433 9160 4445 9163
rect 4028 9132 4445 9160
rect 4028 9120 4034 9132
rect 4433 9129 4445 9132
rect 4479 9129 4491 9163
rect 4433 9123 4491 9129
rect 5445 9163 5503 9169
rect 5445 9129 5457 9163
rect 5491 9160 5503 9163
rect 5626 9160 5632 9172
rect 5491 9132 5632 9160
rect 5491 9129 5503 9132
rect 5445 9123 5503 9129
rect 5626 9120 5632 9132
rect 5684 9160 5690 9172
rect 5902 9160 5908 9172
rect 5684 9132 5908 9160
rect 5684 9120 5690 9132
rect 5902 9120 5908 9132
rect 5960 9120 5966 9172
rect 6362 9160 6368 9172
rect 6323 9132 6368 9160
rect 6362 9120 6368 9132
rect 6420 9120 6426 9172
rect 6822 9160 6828 9172
rect 6472 9132 6828 9160
rect 1578 9052 1584 9104
rect 1636 9092 1642 9104
rect 2682 9092 2688 9104
rect 1636 9064 2688 9092
rect 1636 9052 1642 9064
rect 2682 9052 2688 9064
rect 2740 9052 2746 9104
rect 2866 9052 2872 9104
rect 2924 9092 2930 9104
rect 2924 9064 3096 9092
rect 2924 9052 2930 9064
rect 2958 9024 2964 9036
rect 2919 8996 2964 9024
rect 2958 8984 2964 8996
rect 3016 8984 3022 9036
rect 3068 8968 3096 9064
rect 4982 9052 4988 9104
rect 5040 9092 5046 9104
rect 6472 9092 6500 9132
rect 6822 9120 6828 9132
rect 6880 9120 6886 9172
rect 7101 9163 7159 9169
rect 7101 9129 7113 9163
rect 7147 9160 7159 9163
rect 7190 9160 7196 9172
rect 7147 9132 7196 9160
rect 7147 9129 7159 9132
rect 7101 9123 7159 9129
rect 7190 9120 7196 9132
rect 7248 9120 7254 9172
rect 8389 9163 8447 9169
rect 8389 9129 8401 9163
rect 8435 9160 8447 9163
rect 8662 9160 8668 9172
rect 8435 9132 8668 9160
rect 8435 9129 8447 9132
rect 8389 9123 8447 9129
rect 8662 9120 8668 9132
rect 8720 9120 8726 9172
rect 11238 9160 11244 9172
rect 11199 9132 11244 9160
rect 11238 9120 11244 9132
rect 11296 9120 11302 9172
rect 11701 9163 11759 9169
rect 11701 9129 11713 9163
rect 11747 9160 11759 9163
rect 11974 9160 11980 9172
rect 11747 9132 11980 9160
rect 11747 9129 11759 9132
rect 11701 9123 11759 9129
rect 11974 9120 11980 9132
rect 12032 9120 12038 9172
rect 12728 9132 14044 9160
rect 5040 9064 6500 9092
rect 6549 9095 6607 9101
rect 5040 9052 5046 9064
rect 6549 9061 6561 9095
rect 6595 9092 6607 9095
rect 6638 9092 6644 9104
rect 6595 9064 6644 9092
rect 6595 9061 6607 9064
rect 6549 9055 6607 9061
rect 6638 9052 6644 9064
rect 6696 9052 6702 9104
rect 6914 9052 6920 9104
rect 6972 9092 6978 9104
rect 8573 9095 8631 9101
rect 6972 9064 8524 9092
rect 6972 9052 6978 9064
rect 3510 8984 3516 9036
rect 3568 9024 3574 9036
rect 8205 9027 8263 9033
rect 8205 9024 8217 9027
rect 3568 8996 8217 9024
rect 3568 8984 3574 8996
rect 8205 8993 8217 8996
rect 8251 8993 8263 9027
rect 8205 8987 8263 8993
rect 2038 8916 2044 8968
rect 2096 8956 2102 8968
rect 2685 8959 2743 8965
rect 2685 8956 2697 8959
rect 2096 8928 2697 8956
rect 2096 8916 2102 8928
rect 2685 8925 2697 8928
rect 2731 8925 2743 8959
rect 2866 8956 2872 8968
rect 2827 8928 2872 8956
rect 2685 8919 2743 8925
rect 2866 8916 2872 8928
rect 2924 8916 2930 8968
rect 3050 8956 3056 8968
rect 3011 8928 3056 8956
rect 3050 8916 3056 8928
rect 3108 8916 3114 8968
rect 3234 8956 3240 8968
rect 3195 8928 3240 8956
rect 3234 8916 3240 8928
rect 3292 8916 3298 8968
rect 4338 8916 4344 8968
rect 4396 8956 4402 8968
rect 4433 8959 4491 8965
rect 4433 8956 4445 8959
rect 4396 8928 4445 8956
rect 4396 8916 4402 8928
rect 4433 8925 4445 8928
rect 4479 8925 4491 8959
rect 4433 8919 4491 8925
rect 4525 8959 4583 8965
rect 4525 8925 4537 8959
rect 4571 8925 4583 8959
rect 5258 8956 5264 8968
rect 5219 8928 5264 8956
rect 4525 8919 4583 8925
rect 3786 8848 3792 8900
rect 3844 8888 3850 8900
rect 4540 8888 4568 8919
rect 5258 8916 5264 8928
rect 5316 8916 5322 8968
rect 5445 8959 5503 8965
rect 5445 8925 5457 8959
rect 5491 8956 5503 8959
rect 5718 8956 5724 8968
rect 5491 8928 5724 8956
rect 5491 8925 5503 8928
rect 5445 8919 5503 8925
rect 5718 8916 5724 8928
rect 5776 8956 5782 8968
rect 5776 8928 6224 8956
rect 5776 8916 5782 8928
rect 6196 8897 6224 8928
rect 6362 8916 6368 8968
rect 6420 8956 6426 8968
rect 7929 8959 7987 8965
rect 7929 8956 7941 8959
rect 6420 8928 7941 8956
rect 6420 8925 6469 8928
rect 6420 8916 6423 8925
rect 3844 8860 4568 8888
rect 6181 8891 6239 8897
rect 6401 8894 6423 8916
rect 3844 8848 3850 8860
rect 6181 8857 6193 8891
rect 6227 8857 6239 8891
rect 6411 8891 6423 8894
rect 6457 8891 6469 8925
rect 7929 8925 7941 8928
rect 7975 8925 7987 8959
rect 8386 8956 8392 8968
rect 8347 8928 8392 8956
rect 7929 8919 7987 8925
rect 8386 8916 8392 8928
rect 8444 8916 8450 8968
rect 8496 8956 8524 9064
rect 8573 9061 8585 9095
rect 8619 9061 8631 9095
rect 8680 9092 8708 9120
rect 8680 9064 9444 9092
rect 8573 9055 8631 9061
rect 8588 9024 8616 9055
rect 8588 8996 9352 9024
rect 9324 8965 9352 8996
rect 9416 8965 9444 9064
rect 11882 9052 11888 9104
rect 11940 9092 11946 9104
rect 12529 9095 12587 9101
rect 12529 9092 12541 9095
rect 11940 9064 12541 9092
rect 11940 9052 11946 9064
rect 12529 9061 12541 9064
rect 12575 9061 12587 9095
rect 12529 9055 12587 9061
rect 12618 9024 12624 9036
rect 11532 8996 12624 9024
rect 9125 8959 9183 8965
rect 9125 8956 9137 8959
rect 8496 8928 9137 8956
rect 9125 8925 9137 8928
rect 9171 8925 9183 8959
rect 9125 8919 9183 8925
rect 9309 8959 9367 8965
rect 9309 8925 9321 8959
rect 9355 8925 9367 8959
rect 9309 8919 9367 8925
rect 9401 8959 9459 8965
rect 9401 8925 9413 8959
rect 9447 8925 9459 8959
rect 9401 8919 9459 8925
rect 9490 8916 9496 8968
rect 9548 8956 9554 8968
rect 10229 8959 10287 8965
rect 9548 8928 9593 8956
rect 9548 8916 9554 8928
rect 10229 8925 10241 8959
rect 10275 8956 10287 8959
rect 10318 8956 10324 8968
rect 10275 8928 10324 8956
rect 10275 8925 10287 8928
rect 10229 8919 10287 8925
rect 10318 8916 10324 8928
rect 10376 8916 10382 8968
rect 11422 8956 11428 8968
rect 11383 8928 11428 8956
rect 11422 8916 11428 8928
rect 11480 8916 11486 8968
rect 11532 8965 11560 8996
rect 12618 8984 12624 8996
rect 12676 8984 12682 9036
rect 11517 8959 11575 8965
rect 11517 8925 11529 8959
rect 11563 8925 11575 8959
rect 11517 8919 11575 8925
rect 11793 8959 11851 8965
rect 11793 8925 11805 8959
rect 11839 8925 11851 8959
rect 11793 8919 11851 8925
rect 6411 8885 6469 8891
rect 6181 8851 6239 8857
rect 7006 8848 7012 8900
rect 7064 8888 7070 8900
rect 7193 8891 7251 8897
rect 7193 8888 7205 8891
rect 7064 8860 7205 8888
rect 7064 8848 7070 8860
rect 7193 8857 7205 8860
rect 7239 8857 7251 8891
rect 7193 8851 7251 8857
rect 10042 8848 10048 8900
rect 10100 8888 10106 8900
rect 10413 8891 10471 8897
rect 10413 8888 10425 8891
rect 10100 8860 10425 8888
rect 10100 8848 10106 8860
rect 10413 8857 10425 8860
rect 10459 8857 10471 8891
rect 11808 8888 11836 8919
rect 12158 8916 12164 8968
rect 12216 8956 12222 8968
rect 12728 8965 12756 9132
rect 13173 9095 13231 9101
rect 13173 9061 13185 9095
rect 13219 9092 13231 9095
rect 13262 9092 13268 9104
rect 13219 9064 13268 9092
rect 13219 9061 13231 9064
rect 13173 9055 13231 9061
rect 13262 9052 13268 9064
rect 13320 9052 13326 9104
rect 13906 9052 13912 9104
rect 13964 9052 13970 9104
rect 13924 9024 13952 9052
rect 13280 8996 13492 9024
rect 12253 8959 12311 8965
rect 12253 8956 12265 8959
rect 12216 8928 12265 8956
rect 12216 8916 12222 8928
rect 12253 8925 12265 8928
rect 12299 8925 12311 8959
rect 12253 8919 12311 8925
rect 12713 8959 12771 8965
rect 12713 8925 12725 8959
rect 12759 8925 12771 8959
rect 12713 8919 12771 8925
rect 13280 8888 13308 8996
rect 13357 8959 13415 8965
rect 13357 8925 13369 8959
rect 13403 8925 13415 8959
rect 13357 8919 13415 8925
rect 11808 8860 13308 8888
rect 10413 8851 10471 8857
rect 12268 8832 12296 8860
rect 1673 8823 1731 8829
rect 1673 8789 1685 8823
rect 1719 8820 1731 8823
rect 1946 8820 1952 8832
rect 1719 8792 1952 8820
rect 1719 8789 1731 8792
rect 1673 8783 1731 8789
rect 1946 8780 1952 8792
rect 2004 8780 2010 8832
rect 2225 8823 2283 8829
rect 2225 8789 2237 8823
rect 2271 8820 2283 8823
rect 2590 8820 2596 8832
rect 2271 8792 2596 8820
rect 2271 8789 2283 8792
rect 2225 8783 2283 8789
rect 2590 8780 2596 8792
rect 2648 8780 2654 8832
rect 3421 8823 3479 8829
rect 3421 8789 3433 8823
rect 3467 8820 3479 8823
rect 4614 8820 4620 8832
rect 3467 8792 4620 8820
rect 3467 8789 3479 8792
rect 3421 8783 3479 8789
rect 4614 8780 4620 8792
rect 4672 8780 4678 8832
rect 4801 8823 4859 8829
rect 4801 8789 4813 8823
rect 4847 8820 4859 8823
rect 4890 8820 4896 8832
rect 4847 8792 4896 8820
rect 4847 8789 4859 8792
rect 4801 8783 4859 8789
rect 4890 8780 4896 8792
rect 4948 8780 4954 8832
rect 5629 8823 5687 8829
rect 5629 8789 5641 8823
rect 5675 8820 5687 8823
rect 6914 8820 6920 8832
rect 5675 8792 6920 8820
rect 5675 8789 5687 8792
rect 5629 8783 5687 8789
rect 6914 8780 6920 8792
rect 6972 8780 6978 8832
rect 9769 8823 9827 8829
rect 9769 8789 9781 8823
rect 9815 8820 9827 8823
rect 9950 8820 9956 8832
rect 9815 8792 9956 8820
rect 9815 8789 9827 8792
rect 9769 8783 9827 8789
rect 9950 8780 9956 8792
rect 10008 8780 10014 8832
rect 10594 8820 10600 8832
rect 10555 8792 10600 8820
rect 10594 8780 10600 8792
rect 10652 8780 10658 8832
rect 12250 8780 12256 8832
rect 12308 8780 12314 8832
rect 12345 8823 12403 8829
rect 12345 8789 12357 8823
rect 12391 8820 12403 8823
rect 12802 8820 12808 8832
rect 12391 8792 12808 8820
rect 12391 8789 12403 8792
rect 12345 8783 12403 8789
rect 12802 8780 12808 8792
rect 12860 8780 12866 8832
rect 13372 8820 13400 8919
rect 13464 8888 13492 8996
rect 13648 8996 13952 9024
rect 14016 9024 14044 9132
rect 14182 9120 14188 9172
rect 14240 9160 14246 9172
rect 14277 9163 14335 9169
rect 14277 9160 14289 9163
rect 14240 9132 14289 9160
rect 14240 9120 14246 9132
rect 14277 9129 14289 9132
rect 14323 9129 14335 9163
rect 14277 9123 14335 9129
rect 14918 9120 14924 9172
rect 14976 9160 14982 9172
rect 15746 9160 15752 9172
rect 14976 9132 15752 9160
rect 14976 9120 14982 9132
rect 15746 9120 15752 9132
rect 15804 9160 15810 9172
rect 16206 9160 16212 9172
rect 15804 9132 16212 9160
rect 15804 9120 15810 9132
rect 16206 9120 16212 9132
rect 16264 9120 16270 9172
rect 16298 9120 16304 9172
rect 16356 9160 16362 9172
rect 17862 9160 17868 9172
rect 16356 9132 17868 9160
rect 16356 9120 16362 9132
rect 17862 9120 17868 9132
rect 17920 9120 17926 9172
rect 18693 9163 18751 9169
rect 18693 9129 18705 9163
rect 18739 9160 18751 9163
rect 20346 9160 20352 9172
rect 18739 9132 20352 9160
rect 18739 9129 18751 9132
rect 18693 9123 18751 9129
rect 20346 9120 20352 9132
rect 20404 9120 20410 9172
rect 20530 9120 20536 9172
rect 20588 9160 20594 9172
rect 22002 9160 22008 9172
rect 20588 9132 22008 9160
rect 20588 9120 20594 9132
rect 22002 9120 22008 9132
rect 22060 9160 22066 9172
rect 22060 9132 22508 9160
rect 22060 9120 22066 9132
rect 16482 9052 16488 9104
rect 16540 9092 16546 9104
rect 19981 9095 20039 9101
rect 16540 9064 16804 9092
rect 16540 9052 16546 9064
rect 14458 9024 14464 9036
rect 14016 8996 14464 9024
rect 13538 8965 13544 8968
rect 13522 8959 13544 8965
rect 13522 8925 13534 8959
rect 13522 8919 13544 8925
rect 13538 8916 13544 8919
rect 13596 8916 13602 8968
rect 13648 8965 13676 8996
rect 14458 8984 14464 8996
rect 14516 8984 14522 9036
rect 14734 9024 14740 9036
rect 14695 8996 14740 9024
rect 14734 8984 14740 8996
rect 14792 8984 14798 9036
rect 15841 9027 15899 9033
rect 14844 8996 15789 9024
rect 13633 8959 13691 8965
rect 13633 8925 13645 8959
rect 13679 8925 13691 8959
rect 13633 8919 13691 8925
rect 13725 8959 13783 8965
rect 13725 8925 13737 8959
rect 13771 8956 13783 8959
rect 13906 8956 13912 8968
rect 13771 8928 13912 8956
rect 13771 8925 13783 8928
rect 13725 8919 13783 8925
rect 13906 8916 13912 8928
rect 13964 8916 13970 8968
rect 14550 8956 14556 8968
rect 14512 8928 14556 8956
rect 14550 8916 14556 8928
rect 14608 8916 14614 8968
rect 14645 8959 14703 8965
rect 14645 8925 14657 8959
rect 14691 8956 14703 8959
rect 14844 8956 14872 8996
rect 14691 8928 14872 8956
rect 15657 8959 15715 8965
rect 14691 8925 14703 8928
rect 14645 8919 14703 8925
rect 15657 8925 15669 8959
rect 15703 8925 15715 8959
rect 15761 8956 15789 8996
rect 15841 8993 15853 9027
rect 15887 9024 15899 9027
rect 16393 9027 16451 9033
rect 16393 9024 16405 9027
rect 15887 8996 16405 9024
rect 15887 8993 15899 8996
rect 15841 8987 15899 8993
rect 16393 8993 16405 8996
rect 16439 8993 16451 9027
rect 16666 9024 16672 9036
rect 16627 8996 16672 9024
rect 16393 8987 16451 8993
rect 16666 8984 16672 8996
rect 16724 8984 16730 9036
rect 15933 8959 15991 8965
rect 15933 8956 15945 8959
rect 15761 8928 15945 8956
rect 15657 8919 15715 8925
rect 15933 8925 15945 8928
rect 15979 8925 15991 8959
rect 16574 8956 16580 8968
rect 16535 8928 16580 8956
rect 15933 8919 15991 8925
rect 14660 8888 14688 8919
rect 13464 8860 14688 8888
rect 14826 8848 14832 8900
rect 14884 8888 14890 8900
rect 15473 8891 15531 8897
rect 15473 8888 15485 8891
rect 14884 8860 15485 8888
rect 14884 8848 14890 8860
rect 15473 8857 15485 8860
rect 15519 8857 15531 8891
rect 15473 8851 15531 8857
rect 14642 8820 14648 8832
rect 13372 8792 14648 8820
rect 14642 8780 14648 8792
rect 14700 8780 14706 8832
rect 15672 8820 15700 8919
rect 16574 8916 16580 8928
rect 16632 8916 16638 8968
rect 16776 8965 16804 9064
rect 19981 9061 19993 9095
rect 20027 9092 20039 9095
rect 20990 9092 20996 9104
rect 20027 9064 20996 9092
rect 20027 9061 20039 9064
rect 19981 9055 20039 9061
rect 20990 9052 20996 9064
rect 21048 9052 21054 9104
rect 16853 9027 16911 9033
rect 16853 8993 16865 9027
rect 16899 9024 16911 9027
rect 17405 9027 17463 9033
rect 17405 9024 17417 9027
rect 16899 8996 17417 9024
rect 16899 8993 16911 8996
rect 16853 8987 16911 8993
rect 17405 8993 17417 8996
rect 17451 8993 17463 9027
rect 18506 9024 18512 9036
rect 17405 8987 17463 8993
rect 17676 8996 18512 9024
rect 16761 8959 16819 8965
rect 16761 8925 16773 8959
rect 16807 8956 16819 8959
rect 17144 8956 17356 8966
rect 17494 8956 17500 8968
rect 16807 8938 17500 8956
rect 16807 8928 17172 8938
rect 17328 8928 17500 8938
rect 16807 8925 16819 8928
rect 16761 8919 16819 8925
rect 17494 8916 17500 8928
rect 17552 8916 17558 8968
rect 17676 8965 17704 8996
rect 18506 8984 18512 8996
rect 18564 8984 18570 9036
rect 18690 8984 18696 9036
rect 18748 9024 18754 9036
rect 18748 8996 20024 9024
rect 18748 8984 18754 8996
rect 17676 8959 17739 8965
rect 17676 8925 17693 8959
rect 17727 8925 17739 8959
rect 17676 8924 17739 8925
rect 17681 8919 17739 8924
rect 17773 8959 17831 8965
rect 17773 8925 17785 8959
rect 17819 8925 17831 8959
rect 17865 8959 17923 8965
rect 17865 8946 17877 8959
rect 17911 8946 17923 8959
rect 18049 8959 18107 8965
rect 17773 8919 17831 8925
rect 16482 8848 16488 8900
rect 16540 8888 16546 8900
rect 17788 8888 17816 8919
rect 17862 8894 17868 8946
rect 17920 8894 17926 8946
rect 18049 8925 18061 8959
rect 18095 8956 18107 8959
rect 18095 8953 18828 8956
rect 18892 8953 19380 8956
rect 18095 8928 19380 8953
rect 18095 8925 18107 8928
rect 18800 8925 18920 8928
rect 18049 8919 18107 8925
rect 16540 8860 17816 8888
rect 18877 8891 18935 8897
rect 16540 8848 16546 8860
rect 18877 8857 18889 8891
rect 18923 8857 18935 8891
rect 19352 8888 19380 8928
rect 19610 8916 19616 8968
rect 19668 8956 19674 8968
rect 19996 8965 20024 8996
rect 20438 8984 20444 9036
rect 20496 9024 20502 9036
rect 20625 9027 20683 9033
rect 20625 9024 20637 9027
rect 20496 8996 20637 9024
rect 20496 8984 20502 8996
rect 20625 8993 20637 8996
rect 20671 8993 20683 9027
rect 20625 8987 20683 8993
rect 20809 9027 20867 9033
rect 20809 8993 20821 9027
rect 20855 9024 20867 9027
rect 21634 9024 21640 9036
rect 20855 8996 21640 9024
rect 20855 8993 20867 8996
rect 20809 8987 20867 8993
rect 21634 8984 21640 8996
rect 21692 8984 21698 9036
rect 19705 8959 19763 8965
rect 19705 8956 19717 8959
rect 19668 8928 19717 8956
rect 19668 8916 19674 8928
rect 19705 8925 19717 8928
rect 19751 8925 19763 8959
rect 19705 8919 19763 8925
rect 19981 8959 20039 8965
rect 19981 8925 19993 8959
rect 20027 8956 20039 8959
rect 20530 8956 20536 8968
rect 20027 8928 20536 8956
rect 20027 8925 20039 8928
rect 19981 8919 20039 8925
rect 20530 8916 20536 8928
rect 20588 8916 20594 8968
rect 20714 8956 20720 8968
rect 20675 8928 20720 8956
rect 20714 8916 20720 8928
rect 20772 8916 20778 8968
rect 20901 8959 20959 8965
rect 20901 8925 20913 8959
rect 20947 8956 20959 8959
rect 21545 8959 21603 8965
rect 21545 8956 21557 8959
rect 20947 8928 21557 8956
rect 20947 8925 20959 8928
rect 20901 8919 20959 8925
rect 21545 8925 21557 8928
rect 21591 8925 21603 8959
rect 21545 8919 21603 8925
rect 19886 8888 19892 8900
rect 19352 8860 19892 8888
rect 18877 8851 18935 8857
rect 17770 8820 17776 8832
rect 15672 8792 17776 8820
rect 17770 8780 17776 8792
rect 17828 8780 17834 8832
rect 18506 8820 18512 8832
rect 18467 8792 18512 8820
rect 18506 8780 18512 8792
rect 18564 8780 18570 8832
rect 18690 8829 18696 8832
rect 18677 8823 18696 8829
rect 18677 8789 18689 8823
rect 18677 8783 18696 8789
rect 18690 8780 18696 8783
rect 18748 8780 18754 8832
rect 18892 8820 18920 8851
rect 19886 8848 19892 8860
rect 19944 8848 19950 8900
rect 20162 8848 20168 8900
rect 20220 8888 20226 8900
rect 20916 8888 20944 8919
rect 22278 8916 22284 8968
rect 22336 8956 22342 8968
rect 22480 8965 22508 9132
rect 22373 8959 22431 8965
rect 22373 8956 22385 8959
rect 22336 8928 22385 8956
rect 22336 8916 22342 8928
rect 22373 8925 22385 8928
rect 22419 8925 22431 8959
rect 22373 8919 22431 8925
rect 22465 8959 22523 8965
rect 22465 8925 22477 8959
rect 22511 8925 22523 8959
rect 22465 8919 22523 8925
rect 22649 8959 22707 8965
rect 22649 8925 22661 8959
rect 22695 8956 22707 8959
rect 23014 8956 23020 8968
rect 22695 8928 23020 8956
rect 22695 8925 22707 8928
rect 22649 8919 22707 8925
rect 23014 8916 23020 8928
rect 23072 8916 23078 8968
rect 20220 8860 20944 8888
rect 20220 8848 20226 8860
rect 18966 8820 18972 8832
rect 18892 8792 18972 8820
rect 18966 8780 18972 8792
rect 19024 8780 19030 8832
rect 19334 8780 19340 8832
rect 19392 8820 19398 8832
rect 19797 8823 19855 8829
rect 19797 8820 19809 8823
rect 19392 8792 19809 8820
rect 19392 8780 19398 8792
rect 19797 8789 19809 8792
rect 19843 8789 19855 8823
rect 19797 8783 19855 8789
rect 20441 8823 20499 8829
rect 20441 8789 20453 8823
rect 20487 8820 20499 8823
rect 20530 8820 20536 8832
rect 20487 8792 20536 8820
rect 20487 8789 20499 8792
rect 20441 8783 20499 8789
rect 20530 8780 20536 8792
rect 20588 8780 20594 8832
rect 20714 8780 20720 8832
rect 20772 8820 20778 8832
rect 21174 8820 21180 8832
rect 20772 8792 21180 8820
rect 20772 8780 20778 8792
rect 21174 8780 21180 8792
rect 21232 8780 21238 8832
rect 21634 8820 21640 8832
rect 21595 8792 21640 8820
rect 21634 8780 21640 8792
rect 21692 8820 21698 8832
rect 22094 8820 22100 8832
rect 21692 8792 22100 8820
rect 21692 8780 21698 8792
rect 22094 8780 22100 8792
rect 22152 8820 22158 8832
rect 22554 8820 22560 8832
rect 22152 8792 22560 8820
rect 22152 8780 22158 8792
rect 22554 8780 22560 8792
rect 22612 8780 22618 8832
rect 22830 8820 22836 8832
rect 22791 8792 22836 8820
rect 22830 8780 22836 8792
rect 22888 8780 22894 8832
rect 1104 8730 23987 8752
rect 1104 8678 6630 8730
rect 6682 8678 6694 8730
rect 6746 8678 6758 8730
rect 6810 8678 6822 8730
rect 6874 8678 6886 8730
rect 6938 8678 12311 8730
rect 12363 8678 12375 8730
rect 12427 8678 12439 8730
rect 12491 8678 12503 8730
rect 12555 8678 12567 8730
rect 12619 8678 17992 8730
rect 18044 8678 18056 8730
rect 18108 8678 18120 8730
rect 18172 8678 18184 8730
rect 18236 8678 18248 8730
rect 18300 8678 23673 8730
rect 23725 8678 23737 8730
rect 23789 8678 23801 8730
rect 23853 8678 23865 8730
rect 23917 8678 23929 8730
rect 23981 8678 23987 8730
rect 1104 8656 23987 8678
rect 2038 8616 2044 8628
rect 1999 8588 2044 8616
rect 2038 8576 2044 8588
rect 2096 8576 2102 8628
rect 2682 8576 2688 8628
rect 2740 8616 2746 8628
rect 3786 8616 3792 8628
rect 2740 8588 3792 8616
rect 2740 8576 2746 8588
rect 3786 8576 3792 8588
rect 3844 8576 3850 8628
rect 4249 8619 4307 8625
rect 4249 8585 4261 8619
rect 4295 8616 4307 8619
rect 4706 8616 4712 8628
rect 4295 8588 4712 8616
rect 4295 8585 4307 8588
rect 4249 8579 4307 8585
rect 4706 8576 4712 8588
rect 4764 8616 4770 8628
rect 5169 8619 5227 8625
rect 5169 8616 5181 8619
rect 4764 8588 5181 8616
rect 4764 8576 4770 8588
rect 5169 8585 5181 8588
rect 5215 8616 5227 8619
rect 5258 8616 5264 8628
rect 5215 8588 5264 8616
rect 5215 8585 5227 8588
rect 5169 8579 5227 8585
rect 5258 8576 5264 8588
rect 5316 8576 5322 8628
rect 5350 8576 5356 8628
rect 5408 8616 5414 8628
rect 7006 8616 7012 8628
rect 5408 8588 7012 8616
rect 5408 8576 5414 8588
rect 7006 8576 7012 8588
rect 7064 8576 7070 8628
rect 7098 8576 7104 8628
rect 7156 8616 7162 8628
rect 7377 8619 7435 8625
rect 7377 8616 7389 8619
rect 7156 8588 7389 8616
rect 7156 8576 7162 8588
rect 7377 8585 7389 8588
rect 7423 8585 7435 8619
rect 7377 8579 7435 8585
rect 8754 8576 8760 8628
rect 8812 8616 8818 8628
rect 9493 8619 9551 8625
rect 9493 8616 9505 8619
rect 8812 8588 9505 8616
rect 8812 8576 8818 8588
rect 9493 8585 9505 8588
rect 9539 8585 9551 8619
rect 9493 8579 9551 8585
rect 10226 8576 10232 8628
rect 10284 8616 10290 8628
rect 10284 8588 10548 8616
rect 10284 8576 10290 8588
rect 2774 8548 2780 8560
rect 1872 8520 2780 8548
rect 1872 8489 1900 8520
rect 2774 8508 2780 8520
rect 2832 8508 2838 8560
rect 1857 8483 1915 8489
rect 1857 8449 1869 8483
rect 1903 8449 1915 8483
rect 1857 8443 1915 8449
rect 2314 8440 2320 8492
rect 2372 8480 2378 8492
rect 2590 8480 2596 8492
rect 2372 8452 2596 8480
rect 2372 8440 2378 8452
rect 2590 8440 2596 8452
rect 2648 8480 2654 8492
rect 2685 8483 2743 8489
rect 2685 8480 2697 8483
rect 2648 8452 2697 8480
rect 2648 8440 2654 8452
rect 2685 8449 2697 8452
rect 2731 8480 2743 8483
rect 3234 8480 3240 8492
rect 2731 8452 3240 8480
rect 2731 8449 2743 8452
rect 2685 8443 2743 8449
rect 3234 8440 3240 8452
rect 3292 8440 3298 8492
rect 3602 8440 3608 8492
rect 3660 8480 3666 8492
rect 3804 8489 3832 8576
rect 7282 8548 7288 8560
rect 5092 8520 7288 8548
rect 3697 8483 3755 8489
rect 3697 8480 3709 8483
rect 3660 8452 3709 8480
rect 3660 8440 3666 8452
rect 3697 8449 3709 8452
rect 3743 8449 3755 8483
rect 3697 8443 3755 8449
rect 3789 8483 3847 8489
rect 3789 8449 3801 8483
rect 3835 8449 3847 8483
rect 3970 8480 3976 8492
rect 3931 8452 3976 8480
rect 3789 8443 3847 8449
rect 3970 8440 3976 8452
rect 4028 8440 4034 8492
rect 4065 8483 4123 8489
rect 4065 8449 4077 8483
rect 4111 8480 4123 8483
rect 4338 8480 4344 8492
rect 4111 8452 4344 8480
rect 4111 8449 4123 8452
rect 4065 8443 4123 8449
rect 4338 8440 4344 8452
rect 4396 8440 4402 8492
rect 4890 8440 4896 8492
rect 4948 8480 4954 8492
rect 5092 8489 5120 8520
rect 7282 8508 7288 8520
rect 7340 8508 7346 8560
rect 7745 8551 7803 8557
rect 7745 8517 7757 8551
rect 7791 8548 7803 8551
rect 9585 8551 9643 8557
rect 7791 8520 8984 8548
rect 7791 8517 7803 8520
rect 7745 8511 7803 8517
rect 8956 8492 8984 8520
rect 9585 8517 9597 8551
rect 9631 8548 9643 8551
rect 9858 8548 9864 8560
rect 9631 8520 9864 8548
rect 9631 8517 9643 8520
rect 9585 8511 9643 8517
rect 9858 8508 9864 8520
rect 9916 8508 9922 8560
rect 10042 8548 10048 8560
rect 9968 8520 10048 8548
rect 5077 8483 5135 8489
rect 5077 8480 5089 8483
rect 4948 8452 5089 8480
rect 4948 8440 4954 8452
rect 5077 8449 5089 8452
rect 5123 8449 5135 8483
rect 5077 8443 5135 8449
rect 5353 8483 5411 8489
rect 5353 8449 5365 8483
rect 5399 8480 5411 8483
rect 5399 8452 5488 8480
rect 5399 8449 5411 8452
rect 5353 8443 5411 8449
rect 1581 8415 1639 8421
rect 1581 8381 1593 8415
rect 1627 8412 1639 8415
rect 2498 8412 2504 8424
rect 1627 8384 2504 8412
rect 1627 8381 1639 8384
rect 1581 8375 1639 8381
rect 2498 8372 2504 8384
rect 2556 8372 2562 8424
rect 2869 8415 2927 8421
rect 2869 8381 2881 8415
rect 2915 8412 2927 8415
rect 4908 8412 4936 8440
rect 2915 8384 4936 8412
rect 5460 8412 5488 8452
rect 5534 8440 5540 8492
rect 5592 8480 5598 8492
rect 6641 8483 6699 8489
rect 6641 8480 6653 8483
rect 5592 8452 6653 8480
rect 5592 8440 5598 8452
rect 6641 8449 6653 8452
rect 6687 8449 6699 8483
rect 7374 8480 7380 8492
rect 6641 8443 6699 8449
rect 6748 8452 7380 8480
rect 6748 8412 6776 8452
rect 7374 8440 7380 8452
rect 7432 8440 7438 8492
rect 7558 8480 7564 8492
rect 7519 8452 7564 8480
rect 7558 8440 7564 8452
rect 7616 8440 7622 8492
rect 7650 8440 7656 8492
rect 7708 8480 7714 8492
rect 7708 8452 7753 8480
rect 7708 8440 7714 8452
rect 7834 8440 7840 8492
rect 7892 8489 7898 8492
rect 7892 8483 7921 8489
rect 7909 8449 7921 8483
rect 8018 8480 8024 8492
rect 7979 8452 8024 8480
rect 7892 8443 7921 8449
rect 7892 8440 7898 8443
rect 8018 8440 8024 8452
rect 8076 8440 8082 8492
rect 8478 8489 8484 8492
rect 8473 8480 8484 8489
rect 8391 8452 8484 8480
rect 5460 8384 6776 8412
rect 2915 8381 2927 8384
rect 2869 8375 2927 8381
rect 3694 8304 3700 8356
rect 3752 8344 3758 8356
rect 5074 8344 5080 8356
rect 3752 8316 5080 8344
rect 3752 8304 3758 8316
rect 5074 8304 5080 8316
rect 5132 8344 5138 8356
rect 5460 8344 5488 8384
rect 7006 8372 7012 8424
rect 7064 8412 7070 8424
rect 8404 8412 8432 8452
rect 8473 8443 8484 8452
rect 8536 8480 8542 8492
rect 8662 8480 8668 8492
rect 8536 8452 8668 8480
rect 8478 8440 8484 8443
rect 8536 8440 8542 8452
rect 8662 8440 8668 8452
rect 8720 8440 8726 8492
rect 8938 8440 8944 8492
rect 8996 8480 9002 8492
rect 9401 8483 9459 8489
rect 9401 8480 9413 8483
rect 8996 8452 9413 8480
rect 8996 8440 9002 8452
rect 9401 8449 9413 8452
rect 9447 8449 9459 8483
rect 9401 8443 9459 8449
rect 9769 8483 9827 8489
rect 9769 8449 9781 8483
rect 9815 8480 9827 8483
rect 9968 8480 9996 8520
rect 10042 8508 10048 8520
rect 10100 8548 10106 8560
rect 10410 8548 10416 8560
rect 10100 8520 10416 8548
rect 10100 8508 10106 8520
rect 10410 8508 10416 8520
rect 10468 8508 10474 8560
rect 10520 8489 10548 8588
rect 12158 8576 12164 8628
rect 12216 8616 12222 8628
rect 12897 8619 12955 8625
rect 12216 8588 12848 8616
rect 12216 8576 12222 8588
rect 11606 8508 11612 8560
rect 11664 8548 11670 8560
rect 11793 8551 11851 8557
rect 11793 8548 11805 8551
rect 11664 8520 11805 8548
rect 11664 8508 11670 8520
rect 11793 8517 11805 8520
rect 11839 8548 11851 8551
rect 11882 8548 11888 8560
rect 11839 8520 11888 8548
rect 11839 8517 11851 8520
rect 11793 8511 11851 8517
rect 11882 8508 11888 8520
rect 11940 8508 11946 8560
rect 12066 8508 12072 8560
rect 12124 8548 12130 8560
rect 12526 8548 12532 8560
rect 12124 8520 12389 8548
rect 12487 8520 12532 8548
rect 12124 8508 12130 8520
rect 12361 8489 12389 8520
rect 12526 8508 12532 8520
rect 12584 8508 12590 8560
rect 12820 8548 12848 8588
rect 12897 8585 12909 8619
rect 12943 8616 12955 8619
rect 12986 8616 12992 8628
rect 12943 8588 12992 8616
rect 12943 8585 12955 8588
rect 12897 8579 12955 8585
rect 12986 8576 12992 8588
rect 13044 8576 13050 8628
rect 13357 8619 13415 8625
rect 13357 8585 13369 8619
rect 13403 8616 13415 8619
rect 14458 8616 14464 8628
rect 13403 8588 14464 8616
rect 13403 8585 13415 8588
rect 13357 8579 13415 8585
rect 14458 8576 14464 8588
rect 14516 8576 14522 8628
rect 14829 8619 14887 8625
rect 14829 8585 14841 8619
rect 14875 8585 14887 8619
rect 14829 8579 14887 8585
rect 14844 8548 14872 8579
rect 16022 8576 16028 8628
rect 16080 8616 16086 8628
rect 16133 8619 16191 8625
rect 16133 8616 16145 8619
rect 16080 8588 16145 8616
rect 16080 8576 16086 8588
rect 16133 8585 16145 8588
rect 16179 8585 16191 8619
rect 16133 8579 16191 8585
rect 16301 8619 16359 8625
rect 16301 8585 16313 8619
rect 16347 8616 16359 8619
rect 16482 8616 16488 8628
rect 16347 8588 16488 8616
rect 16347 8585 16359 8588
rect 16301 8579 16359 8585
rect 16482 8576 16488 8588
rect 16540 8576 16546 8628
rect 16574 8576 16580 8628
rect 16632 8616 16638 8628
rect 16945 8619 17003 8625
rect 16945 8616 16957 8619
rect 16632 8588 16957 8616
rect 16632 8576 16638 8588
rect 16945 8585 16957 8588
rect 16991 8585 17003 8619
rect 18322 8616 18328 8628
rect 16945 8579 17003 8585
rect 17972 8588 18328 8616
rect 15933 8551 15991 8557
rect 15933 8548 15945 8551
rect 12820 8520 14872 8548
rect 14936 8520 15945 8548
rect 9815 8452 9996 8480
rect 10321 8483 10379 8489
rect 9815 8449 9827 8452
rect 9769 8443 9827 8449
rect 10321 8449 10333 8483
rect 10367 8449 10379 8483
rect 10321 8443 10379 8449
rect 10505 8483 10563 8489
rect 10505 8449 10517 8483
rect 10551 8449 10563 8483
rect 10505 8443 10563 8449
rect 12253 8483 12311 8489
rect 12253 8449 12265 8483
rect 12299 8449 12311 8483
rect 12253 8443 12311 8449
rect 12346 8483 12404 8489
rect 12346 8449 12358 8483
rect 12392 8449 12404 8483
rect 12346 8443 12404 8449
rect 12621 8483 12679 8489
rect 12621 8449 12633 8483
rect 12667 8449 12679 8483
rect 12621 8443 12679 8449
rect 12759 8483 12817 8489
rect 12759 8449 12771 8483
rect 12805 8480 12817 8483
rect 12894 8480 12900 8492
rect 12805 8452 12900 8480
rect 12805 8449 12817 8452
rect 12759 8443 12817 8449
rect 7064 8384 8432 8412
rect 8573 8415 8631 8421
rect 7064 8372 7070 8384
rect 8573 8381 8585 8415
rect 8619 8412 8631 8415
rect 9861 8415 9919 8421
rect 9861 8412 9873 8415
rect 8619 8384 9873 8412
rect 8619 8381 8631 8384
rect 8573 8375 8631 8381
rect 9861 8381 9873 8384
rect 9907 8381 9919 8415
rect 9861 8375 9919 8381
rect 5132 8316 5488 8344
rect 5537 8347 5595 8353
rect 5132 8304 5138 8316
rect 5537 8313 5549 8347
rect 5583 8344 5595 8347
rect 10336 8344 10364 8443
rect 5583 8316 10364 8344
rect 12268 8344 12296 8443
rect 12636 8412 12664 8443
rect 12894 8440 12900 8452
rect 12952 8440 12958 8492
rect 13630 8480 13636 8492
rect 13591 8452 13636 8480
rect 13630 8440 13636 8452
rect 13688 8440 13694 8492
rect 13725 8483 13783 8489
rect 13725 8449 13737 8483
rect 13771 8480 13783 8483
rect 14191 8483 14249 8489
rect 13771 8452 13860 8480
rect 13771 8449 13783 8452
rect 13725 8443 13783 8449
rect 13078 8412 13084 8424
rect 12636 8384 13084 8412
rect 13078 8372 13084 8384
rect 13136 8372 13142 8424
rect 13170 8344 13176 8356
rect 12268 8316 13176 8344
rect 5583 8313 5595 8316
rect 5537 8307 5595 8313
rect 7668 8288 7696 8316
rect 13170 8304 13176 8316
rect 13228 8304 13234 8356
rect 1673 8279 1731 8285
rect 1673 8245 1685 8279
rect 1719 8276 1731 8279
rect 1854 8276 1860 8288
rect 1719 8248 1860 8276
rect 1719 8245 1731 8248
rect 1673 8239 1731 8245
rect 1854 8236 1860 8248
rect 1912 8236 1918 8288
rect 6362 8236 6368 8288
rect 6420 8276 6426 8288
rect 6733 8279 6791 8285
rect 6733 8276 6745 8279
rect 6420 8248 6745 8276
rect 6420 8236 6426 8248
rect 6733 8245 6745 8248
rect 6779 8276 6791 8279
rect 7190 8276 7196 8288
rect 6779 8248 7196 8276
rect 6779 8245 6791 8248
rect 6733 8239 6791 8245
rect 7190 8236 7196 8248
rect 7248 8236 7254 8288
rect 7650 8236 7656 8288
rect 7708 8236 7714 8288
rect 9122 8276 9128 8288
rect 9083 8248 9128 8276
rect 9122 8236 9128 8248
rect 9180 8236 9186 8288
rect 9306 8236 9312 8288
rect 9364 8276 9370 8288
rect 9490 8276 9496 8288
rect 9364 8248 9496 8276
rect 9364 8236 9370 8248
rect 9490 8236 9496 8248
rect 9548 8276 9554 8288
rect 10321 8279 10379 8285
rect 10321 8276 10333 8279
rect 9548 8248 10333 8276
rect 9548 8236 9554 8248
rect 10321 8245 10333 8248
rect 10367 8245 10379 8279
rect 10321 8239 10379 8245
rect 10410 8236 10416 8288
rect 10468 8276 10474 8288
rect 10689 8279 10747 8285
rect 10689 8276 10701 8279
rect 10468 8248 10701 8276
rect 10468 8236 10474 8248
rect 10689 8245 10701 8248
rect 10735 8245 10747 8279
rect 10689 8239 10747 8245
rect 12710 8236 12716 8288
rect 12768 8276 12774 8288
rect 13538 8276 13544 8288
rect 12768 8248 13544 8276
rect 12768 8236 12774 8248
rect 13538 8236 13544 8248
rect 13596 8236 13602 8288
rect 13832 8276 13860 8452
rect 14191 8449 14203 8483
rect 14237 8480 14249 8483
rect 14369 8483 14427 8489
rect 14237 8452 14320 8480
rect 14237 8449 14249 8452
rect 14191 8443 14249 8449
rect 14292 8412 14320 8452
rect 14369 8449 14381 8483
rect 14415 8480 14427 8483
rect 14458 8480 14464 8492
rect 14415 8452 14464 8480
rect 14415 8449 14427 8452
rect 14369 8443 14427 8449
rect 14458 8440 14464 8452
rect 14516 8480 14522 8492
rect 14936 8480 14964 8520
rect 15933 8517 15945 8520
rect 15979 8517 15991 8551
rect 17310 8548 17316 8560
rect 15933 8511 15991 8517
rect 17144 8520 17316 8548
rect 14516 8452 14964 8480
rect 15013 8483 15071 8489
rect 14516 8440 14522 8452
rect 15013 8449 15025 8483
rect 15059 8480 15071 8483
rect 15746 8480 15752 8492
rect 15059 8452 15752 8480
rect 15059 8449 15071 8452
rect 15013 8443 15071 8449
rect 15746 8440 15752 8452
rect 15804 8440 15810 8492
rect 15948 8480 15976 8511
rect 16114 8480 16120 8492
rect 15948 8452 16120 8480
rect 14550 8412 14556 8424
rect 14292 8384 14556 8412
rect 14550 8372 14556 8384
rect 14608 8372 14614 8424
rect 14826 8372 14832 8424
rect 14884 8412 14890 8424
rect 15105 8415 15163 8421
rect 15105 8412 15117 8415
rect 14884 8384 15117 8412
rect 14884 8372 14890 8384
rect 15105 8381 15117 8384
rect 15151 8381 15163 8415
rect 15105 8375 15163 8381
rect 15197 8415 15255 8421
rect 15197 8381 15209 8415
rect 15243 8381 15255 8415
rect 15197 8375 15255 8381
rect 15289 8415 15347 8421
rect 15289 8381 15301 8415
rect 15335 8412 15347 8415
rect 15470 8412 15476 8424
rect 15335 8384 15476 8412
rect 15335 8381 15347 8384
rect 15289 8375 15347 8381
rect 14277 8347 14335 8353
rect 14277 8313 14289 8347
rect 14323 8344 14335 8347
rect 14918 8344 14924 8356
rect 14323 8316 14924 8344
rect 14323 8313 14335 8316
rect 14277 8307 14335 8313
rect 14918 8304 14924 8316
rect 14976 8304 14982 8356
rect 15212 8344 15240 8375
rect 15470 8372 15476 8384
rect 15528 8372 15534 8424
rect 15948 8344 15976 8452
rect 16114 8440 16120 8452
rect 16172 8440 16178 8492
rect 17144 8489 17172 8520
rect 17310 8508 17316 8520
rect 17368 8508 17374 8560
rect 17129 8483 17187 8489
rect 17129 8449 17141 8483
rect 17175 8449 17187 8483
rect 17129 8443 17187 8449
rect 17218 8440 17224 8492
rect 17276 8480 17282 8492
rect 17405 8483 17463 8489
rect 17276 8452 17321 8480
rect 17276 8440 17282 8452
rect 17405 8449 17417 8483
rect 17451 8449 17463 8483
rect 17405 8443 17463 8449
rect 17497 8483 17555 8489
rect 17497 8449 17509 8483
rect 17543 8480 17555 8483
rect 17678 8480 17684 8492
rect 17543 8452 17684 8480
rect 17543 8449 17555 8452
rect 17497 8443 17555 8449
rect 17420 8412 17448 8443
rect 17678 8440 17684 8452
rect 17736 8440 17742 8492
rect 17972 8489 18000 8588
rect 18322 8576 18328 8588
rect 18380 8576 18386 8628
rect 18509 8619 18567 8625
rect 18509 8585 18521 8619
rect 18555 8616 18567 8619
rect 18690 8616 18696 8628
rect 18555 8588 18696 8616
rect 18555 8585 18567 8588
rect 18509 8579 18567 8585
rect 18690 8576 18696 8588
rect 18748 8576 18754 8628
rect 20346 8576 20352 8628
rect 20404 8616 20410 8628
rect 20533 8619 20591 8625
rect 20533 8616 20545 8619
rect 20404 8588 20545 8616
rect 20404 8576 20410 8588
rect 20533 8585 20545 8588
rect 20579 8585 20591 8619
rect 20533 8579 20591 8585
rect 20622 8576 20628 8628
rect 20680 8616 20686 8628
rect 22002 8616 22008 8628
rect 20680 8588 22008 8616
rect 20680 8576 20686 8588
rect 22002 8576 22008 8588
rect 22060 8576 22066 8628
rect 22097 8619 22155 8625
rect 22097 8585 22109 8619
rect 22143 8616 22155 8619
rect 22278 8616 22284 8628
rect 22143 8588 22284 8616
rect 22143 8585 22155 8588
rect 22097 8579 22155 8585
rect 22278 8576 22284 8588
rect 22336 8576 22342 8628
rect 22462 8616 22468 8628
rect 22423 8588 22468 8616
rect 22462 8576 22468 8588
rect 22520 8576 22526 8628
rect 23014 8576 23020 8628
rect 23072 8616 23078 8628
rect 23109 8619 23167 8625
rect 23109 8616 23121 8619
rect 23072 8588 23121 8616
rect 23072 8576 23078 8588
rect 23109 8585 23121 8588
rect 23155 8585 23167 8619
rect 23109 8579 23167 8585
rect 18414 8548 18420 8560
rect 18064 8520 18420 8548
rect 18064 8489 18092 8520
rect 18414 8508 18420 8520
rect 18472 8508 18478 8560
rect 22830 8548 22836 8560
rect 19812 8520 22836 8548
rect 17957 8483 18015 8489
rect 17957 8449 17969 8483
rect 18003 8449 18015 8483
rect 17957 8443 18015 8449
rect 18049 8483 18107 8489
rect 18049 8449 18061 8483
rect 18095 8449 18107 8483
rect 18230 8480 18236 8492
rect 18191 8452 18236 8480
rect 18049 8443 18107 8449
rect 18230 8440 18236 8452
rect 18288 8440 18294 8492
rect 18325 8483 18383 8489
rect 18325 8449 18337 8483
rect 18371 8480 18383 8483
rect 18782 8480 18788 8492
rect 18371 8452 18788 8480
rect 18371 8449 18383 8452
rect 18325 8443 18383 8449
rect 18782 8440 18788 8452
rect 18840 8440 18846 8492
rect 19518 8440 19524 8492
rect 19576 8480 19582 8492
rect 19812 8489 19840 8520
rect 22830 8508 22836 8520
rect 22888 8508 22894 8560
rect 19705 8483 19763 8489
rect 19705 8480 19717 8483
rect 19576 8452 19717 8480
rect 19576 8440 19582 8452
rect 19705 8449 19717 8452
rect 19751 8449 19763 8483
rect 19705 8443 19763 8449
rect 19797 8483 19855 8489
rect 19797 8449 19809 8483
rect 19843 8449 19855 8483
rect 19797 8443 19855 8449
rect 19886 8440 19892 8492
rect 19944 8480 19950 8492
rect 19944 8452 19989 8480
rect 19944 8440 19950 8452
rect 20070 8440 20076 8492
rect 20128 8480 20134 8492
rect 20714 8480 20720 8492
rect 20128 8452 20173 8480
rect 20675 8452 20720 8480
rect 20128 8440 20134 8452
rect 20714 8440 20720 8452
rect 20772 8440 20778 8492
rect 20809 8483 20867 8489
rect 20809 8449 20821 8483
rect 20855 8449 20867 8483
rect 20990 8480 20996 8492
rect 20951 8452 20996 8480
rect 20809 8443 20867 8449
rect 18414 8412 18420 8424
rect 17420 8384 18420 8412
rect 18414 8372 18420 8384
rect 18472 8372 18478 8424
rect 18966 8412 18972 8424
rect 18524 8384 18972 8412
rect 15212 8316 15976 8344
rect 17218 8304 17224 8356
rect 17276 8344 17282 8356
rect 18230 8344 18236 8356
rect 17276 8316 18236 8344
rect 17276 8304 17282 8316
rect 18230 8304 18236 8316
rect 18288 8304 18294 8356
rect 14734 8276 14740 8288
rect 13832 8248 14740 8276
rect 14734 8236 14740 8248
rect 14792 8236 14798 8288
rect 16117 8279 16175 8285
rect 16117 8245 16129 8279
rect 16163 8276 16175 8279
rect 16298 8276 16304 8288
rect 16163 8248 16304 8276
rect 16163 8245 16175 8248
rect 16117 8239 16175 8245
rect 16298 8236 16304 8248
rect 16356 8236 16362 8288
rect 18046 8236 18052 8288
rect 18104 8276 18110 8288
rect 18524 8276 18552 8384
rect 18966 8372 18972 8384
rect 19024 8412 19030 8424
rect 19024 8384 20484 8412
rect 19024 8372 19030 8384
rect 20456 8294 20484 8384
rect 20622 8372 20628 8424
rect 20680 8412 20686 8424
rect 20824 8412 20852 8443
rect 20990 8440 20996 8452
rect 21048 8440 21054 8492
rect 21085 8483 21143 8489
rect 21085 8449 21097 8483
rect 21131 8480 21143 8483
rect 21634 8480 21640 8492
rect 21131 8452 21640 8480
rect 21131 8449 21143 8452
rect 21085 8443 21143 8449
rect 21634 8440 21640 8452
rect 21692 8440 21698 8492
rect 21726 8440 21732 8492
rect 21784 8480 21790 8492
rect 22005 8483 22063 8489
rect 22005 8480 22017 8483
rect 21784 8452 22017 8480
rect 21784 8440 21790 8452
rect 22005 8449 22017 8452
rect 22051 8449 22063 8483
rect 22005 8443 22063 8449
rect 22281 8483 22339 8489
rect 22281 8449 22293 8483
rect 22327 8480 22339 8483
rect 22370 8480 22376 8492
rect 22327 8452 22376 8480
rect 22327 8449 22339 8452
rect 22281 8443 22339 8449
rect 22370 8440 22376 8452
rect 22428 8440 22434 8492
rect 22925 8483 22983 8489
rect 22925 8449 22937 8483
rect 22971 8449 22983 8483
rect 22925 8443 22983 8449
rect 20680 8384 20852 8412
rect 20680 8372 20686 8384
rect 21358 8372 21364 8424
rect 21416 8412 21422 8424
rect 22940 8412 22968 8443
rect 21416 8384 22968 8412
rect 21416 8372 21422 8384
rect 20806 8304 20812 8356
rect 20864 8344 20870 8356
rect 20864 8316 21956 8344
rect 20864 8304 20870 8316
rect 18104 8248 18552 8276
rect 18104 8236 18110 8248
rect 19334 8236 19340 8288
rect 19392 8276 19398 8288
rect 19429 8279 19487 8285
rect 19429 8276 19441 8279
rect 19392 8248 19441 8276
rect 19392 8236 19398 8248
rect 19429 8245 19441 8248
rect 19475 8245 19487 8279
rect 20456 8276 20576 8294
rect 21082 8276 21088 8288
rect 20456 8266 21088 8276
rect 20548 8248 21088 8266
rect 19429 8239 19487 8245
rect 21082 8236 21088 8248
rect 21140 8236 21146 8288
rect 21928 8276 21956 8316
rect 22002 8304 22008 8356
rect 22060 8344 22066 8356
rect 22186 8344 22192 8356
rect 22060 8316 22192 8344
rect 22060 8304 22066 8316
rect 22186 8304 22192 8316
rect 22244 8304 22250 8356
rect 22554 8276 22560 8288
rect 21928 8248 22560 8276
rect 22554 8236 22560 8248
rect 22612 8276 22618 8288
rect 23014 8276 23020 8288
rect 22612 8248 23020 8276
rect 22612 8236 22618 8248
rect 23014 8236 23020 8248
rect 23072 8236 23078 8288
rect 1104 8186 23828 8208
rect 1104 8134 3790 8186
rect 3842 8134 3854 8186
rect 3906 8134 3918 8186
rect 3970 8134 3982 8186
rect 4034 8134 4046 8186
rect 4098 8134 9471 8186
rect 9523 8134 9535 8186
rect 9587 8134 9599 8186
rect 9651 8134 9663 8186
rect 9715 8134 9727 8186
rect 9779 8134 15152 8186
rect 15204 8134 15216 8186
rect 15268 8134 15280 8186
rect 15332 8134 15344 8186
rect 15396 8134 15408 8186
rect 15460 8134 20833 8186
rect 20885 8134 20897 8186
rect 20949 8134 20961 8186
rect 21013 8134 21025 8186
rect 21077 8134 21089 8186
rect 21141 8134 23828 8186
rect 1104 8112 23828 8134
rect 1765 8075 1823 8081
rect 1765 8041 1777 8075
rect 1811 8072 1823 8075
rect 1946 8072 1952 8084
rect 1811 8044 1952 8072
rect 1811 8041 1823 8044
rect 1765 8035 1823 8041
rect 1946 8032 1952 8044
rect 2004 8032 2010 8084
rect 2685 8075 2743 8081
rect 2685 8041 2697 8075
rect 2731 8072 2743 8075
rect 2866 8072 2872 8084
rect 2731 8044 2872 8072
rect 2731 8041 2743 8044
rect 2685 8035 2743 8041
rect 2866 8032 2872 8044
rect 2924 8032 2930 8084
rect 3329 8075 3387 8081
rect 3329 8041 3341 8075
rect 3375 8072 3387 8075
rect 3510 8072 3516 8084
rect 3375 8044 3516 8072
rect 3375 8041 3387 8044
rect 3329 8035 3387 8041
rect 3510 8032 3516 8044
rect 3568 8032 3574 8084
rect 4249 8075 4307 8081
rect 4249 8041 4261 8075
rect 4295 8072 4307 8075
rect 4338 8072 4344 8084
rect 4295 8044 4344 8072
rect 4295 8041 4307 8044
rect 4249 8035 4307 8041
rect 4338 8032 4344 8044
rect 4396 8032 4402 8084
rect 5077 8075 5135 8081
rect 5077 8041 5089 8075
rect 5123 8072 5135 8075
rect 5166 8072 5172 8084
rect 5123 8044 5172 8072
rect 5123 8041 5135 8044
rect 5077 8035 5135 8041
rect 5166 8032 5172 8044
rect 5224 8032 5230 8084
rect 6454 8032 6460 8084
rect 6512 8072 6518 8084
rect 7285 8075 7343 8081
rect 7285 8072 7297 8075
rect 6512 8044 7297 8072
rect 6512 8032 6518 8044
rect 7285 8041 7297 8044
rect 7331 8041 7343 8075
rect 7285 8035 7343 8041
rect 2774 8004 2780 8016
rect 2424 7976 2780 8004
rect 2314 7877 2320 7880
rect 2299 7871 2320 7877
rect 2299 7837 2311 7871
rect 2299 7831 2320 7837
rect 2314 7828 2320 7831
rect 2372 7828 2378 7880
rect 2424 7877 2452 7976
rect 2774 7964 2780 7976
rect 2832 7964 2838 8016
rect 4706 8004 4712 8016
rect 4667 7976 4712 8004
rect 4706 7964 4712 7976
rect 4764 7964 4770 8016
rect 5261 8007 5319 8013
rect 5261 7973 5273 8007
rect 5307 8004 5319 8007
rect 6270 8004 6276 8016
rect 5307 7976 6276 8004
rect 5307 7973 5319 7976
rect 5261 7967 5319 7973
rect 6270 7964 6276 7976
rect 6328 8004 6334 8016
rect 7300 8004 7328 8035
rect 7558 8032 7564 8084
rect 7616 8072 7622 8084
rect 7745 8075 7803 8081
rect 7745 8072 7757 8075
rect 7616 8044 7757 8072
rect 7616 8032 7622 8044
rect 7745 8041 7757 8044
rect 7791 8041 7803 8075
rect 7745 8035 7803 8041
rect 9677 8075 9735 8081
rect 9677 8041 9689 8075
rect 9723 8072 9735 8075
rect 9858 8072 9864 8084
rect 9723 8044 9864 8072
rect 9723 8041 9735 8044
rect 9677 8035 9735 8041
rect 9858 8032 9864 8044
rect 9916 8032 9922 8084
rect 10778 8032 10784 8084
rect 10836 8072 10842 8084
rect 10873 8075 10931 8081
rect 10873 8072 10885 8075
rect 10836 8044 10885 8072
rect 10836 8032 10842 8044
rect 10873 8041 10885 8044
rect 10919 8041 10931 8075
rect 10873 8035 10931 8041
rect 12897 8075 12955 8081
rect 12897 8041 12909 8075
rect 12943 8072 12955 8075
rect 13354 8072 13360 8084
rect 12943 8044 13360 8072
rect 12943 8041 12955 8044
rect 12897 8035 12955 8041
rect 13354 8032 13360 8044
rect 13412 8032 13418 8084
rect 14642 8072 14648 8084
rect 14603 8044 14648 8072
rect 14642 8032 14648 8044
rect 14700 8032 14706 8084
rect 15746 8072 15752 8084
rect 15707 8044 15752 8072
rect 15746 8032 15752 8044
rect 15804 8072 15810 8084
rect 16482 8072 16488 8084
rect 15804 8044 16488 8072
rect 15804 8032 15810 8044
rect 16482 8032 16488 8044
rect 16540 8072 16546 8084
rect 16945 8075 17003 8081
rect 16945 8072 16957 8075
rect 16540 8044 16957 8072
rect 16540 8032 16546 8044
rect 16945 8041 16957 8044
rect 16991 8041 17003 8075
rect 17770 8072 17776 8084
rect 17731 8044 17776 8072
rect 16945 8035 17003 8041
rect 17770 8032 17776 8044
rect 17828 8032 17834 8084
rect 18782 8032 18788 8084
rect 18840 8072 18846 8084
rect 19429 8075 19487 8081
rect 19429 8072 19441 8075
rect 18840 8044 19441 8072
rect 18840 8032 18846 8044
rect 19429 8041 19441 8044
rect 19475 8041 19487 8075
rect 19429 8035 19487 8041
rect 19797 8075 19855 8081
rect 19797 8041 19809 8075
rect 19843 8072 19855 8075
rect 19886 8072 19892 8084
rect 19843 8044 19892 8072
rect 19843 8041 19855 8044
rect 19797 8035 19855 8041
rect 19886 8032 19892 8044
rect 19944 8032 19950 8084
rect 20254 8072 20260 8084
rect 20215 8044 20260 8072
rect 20254 8032 20260 8044
rect 20312 8032 20318 8084
rect 10229 8007 10287 8013
rect 6328 7976 6868 8004
rect 7300 7976 8248 8004
rect 6328 7964 6334 7976
rect 3421 7939 3479 7945
rect 3421 7936 3433 7939
rect 2516 7908 3433 7936
rect 2516 7880 2544 7908
rect 3421 7905 3433 7908
rect 3467 7905 3479 7939
rect 3421 7899 3479 7905
rect 4246 7896 4252 7948
rect 4304 7936 4310 7948
rect 5626 7936 5632 7948
rect 4304 7908 5632 7936
rect 4304 7896 4310 7908
rect 5626 7896 5632 7908
rect 5684 7936 5690 7948
rect 6362 7936 6368 7948
rect 5684 7908 6368 7936
rect 5684 7896 5690 7908
rect 2409 7871 2467 7877
rect 2409 7837 2421 7871
rect 2455 7837 2467 7871
rect 2409 7831 2467 7837
rect 2498 7828 2504 7880
rect 2556 7868 2562 7880
rect 2556 7840 2601 7868
rect 2556 7828 2562 7840
rect 2682 7828 2688 7880
rect 2740 7868 2746 7880
rect 3145 7871 3203 7877
rect 3145 7868 3157 7871
rect 2740 7840 3157 7868
rect 2740 7828 2746 7840
rect 3145 7837 3157 7840
rect 3191 7837 3203 7871
rect 3145 7831 3203 7837
rect 3237 7871 3295 7877
rect 3237 7837 3249 7871
rect 3283 7868 3295 7871
rect 3510 7868 3516 7880
rect 3283 7840 3516 7868
rect 3283 7837 3295 7840
rect 3237 7831 3295 7837
rect 3510 7828 3516 7840
rect 3568 7828 3574 7880
rect 5994 7868 6000 7880
rect 5092 7840 6000 7868
rect 5092 7809 5120 7840
rect 5994 7828 6000 7840
rect 6052 7828 6058 7880
rect 6288 7877 6316 7908
rect 6362 7896 6368 7908
rect 6420 7896 6426 7948
rect 6546 7936 6552 7948
rect 6507 7908 6552 7936
rect 6546 7896 6552 7908
rect 6604 7896 6610 7948
rect 6840 7936 6868 7976
rect 6840 7908 7880 7936
rect 6273 7871 6331 7877
rect 6273 7837 6285 7871
rect 6319 7837 6331 7871
rect 6454 7868 6460 7880
rect 6415 7840 6460 7868
rect 6273 7831 6331 7837
rect 6454 7828 6460 7840
rect 6512 7828 6518 7880
rect 7190 7868 7196 7880
rect 7151 7840 7196 7868
rect 7190 7828 7196 7840
rect 7248 7828 7254 7880
rect 7469 7871 7527 7877
rect 7469 7868 7481 7871
rect 7300 7840 7481 7868
rect 5077 7803 5135 7809
rect 5077 7769 5089 7803
rect 5123 7769 5135 7803
rect 5077 7763 5135 7769
rect 5626 7760 5632 7812
rect 5684 7800 5690 7812
rect 7300 7800 7328 7840
rect 7469 7837 7481 7840
rect 7515 7837 7527 7871
rect 7469 7831 7527 7837
rect 7561 7871 7619 7877
rect 7561 7837 7573 7871
rect 7607 7868 7619 7871
rect 7650 7868 7656 7880
rect 7607 7840 7656 7868
rect 7607 7837 7619 7840
rect 7561 7831 7619 7837
rect 7650 7828 7656 7840
rect 7708 7828 7714 7880
rect 7745 7871 7803 7877
rect 7745 7837 7757 7871
rect 7791 7837 7803 7871
rect 7852 7868 7880 7908
rect 8220 7880 8248 7976
rect 10229 7973 10241 8007
rect 10275 8004 10287 8007
rect 11146 8004 11152 8016
rect 10275 7976 11152 8004
rect 10275 7973 10287 7976
rect 10229 7967 10287 7973
rect 11146 7964 11152 7976
rect 11204 7964 11210 8016
rect 11514 7964 11520 8016
rect 11572 8004 11578 8016
rect 16022 8004 16028 8016
rect 11572 7976 16028 8004
rect 11572 7964 11578 7976
rect 16022 7964 16028 7976
rect 16080 8004 16086 8016
rect 16209 8007 16267 8013
rect 16080 7976 16160 8004
rect 16080 7964 16086 7976
rect 10410 7936 10416 7948
rect 9324 7908 10416 7936
rect 7926 7868 7932 7880
rect 7852 7840 7932 7868
rect 7745 7831 7803 7837
rect 5684 7772 7328 7800
rect 7760 7800 7788 7831
rect 7926 7828 7932 7840
rect 7984 7828 7990 7880
rect 8202 7868 8208 7880
rect 8115 7840 8208 7868
rect 8202 7828 8208 7840
rect 8260 7828 8266 7880
rect 8386 7868 8392 7880
rect 8347 7840 8392 7868
rect 8386 7828 8392 7840
rect 8444 7868 8450 7880
rect 9324 7877 9352 7908
rect 10410 7896 10416 7908
rect 10468 7896 10474 7948
rect 12069 7939 12127 7945
rect 12069 7905 12081 7939
rect 12115 7936 12127 7939
rect 12158 7936 12164 7948
rect 12115 7908 12164 7936
rect 12115 7905 12127 7908
rect 12069 7899 12127 7905
rect 12158 7896 12164 7908
rect 12216 7936 12222 7948
rect 12894 7936 12900 7948
rect 12216 7908 12900 7936
rect 12216 7896 12222 7908
rect 12894 7896 12900 7908
rect 12952 7936 12958 7948
rect 14550 7936 14556 7948
rect 12952 7908 14556 7936
rect 12952 7896 12958 7908
rect 14550 7896 14556 7908
rect 14608 7896 14614 7948
rect 15102 7936 15108 7948
rect 14844 7908 15108 7936
rect 9125 7871 9183 7877
rect 9125 7868 9137 7871
rect 8444 7840 9137 7868
rect 8444 7828 8450 7840
rect 9125 7837 9137 7840
rect 9171 7837 9183 7871
rect 9125 7831 9183 7837
rect 9309 7871 9367 7877
rect 9309 7837 9321 7871
rect 9355 7837 9367 7871
rect 9309 7831 9367 7837
rect 9401 7871 9459 7877
rect 9401 7837 9413 7871
rect 9447 7837 9459 7871
rect 9401 7831 9459 7837
rect 9493 7871 9551 7877
rect 9493 7837 9505 7871
rect 9539 7868 9551 7871
rect 10042 7868 10048 7880
rect 9539 7840 10048 7868
rect 9539 7837 9551 7840
rect 9493 7831 9551 7837
rect 8754 7800 8760 7812
rect 7760 7772 8760 7800
rect 5684 7760 5690 7772
rect 8754 7760 8760 7772
rect 8812 7760 8818 7812
rect 9416 7800 9444 7831
rect 10042 7828 10048 7840
rect 10100 7828 10106 7880
rect 10594 7828 10600 7880
rect 10652 7868 10658 7880
rect 10689 7871 10747 7877
rect 10689 7868 10701 7871
rect 10652 7840 10701 7868
rect 10652 7828 10658 7840
rect 10689 7837 10701 7840
rect 10735 7837 10747 7871
rect 10689 7831 10747 7837
rect 11609 7871 11667 7877
rect 11609 7837 11621 7871
rect 11655 7868 11667 7871
rect 11790 7868 11796 7880
rect 11655 7840 11796 7868
rect 11655 7837 11667 7840
rect 11609 7831 11667 7837
rect 11790 7828 11796 7840
rect 11848 7828 11854 7880
rect 11882 7828 11888 7880
rect 11940 7868 11946 7880
rect 13081 7871 13139 7877
rect 11940 7840 11985 7868
rect 11940 7828 11946 7840
rect 13081 7837 13093 7871
rect 13127 7837 13139 7871
rect 13081 7831 13139 7837
rect 13173 7871 13231 7877
rect 13173 7837 13185 7871
rect 13219 7837 13231 7871
rect 13354 7868 13360 7880
rect 13315 7840 13360 7868
rect 13173 7831 13231 7837
rect 11698 7800 11704 7812
rect 9416 7772 9536 7800
rect 11659 7772 11704 7800
rect 6089 7735 6147 7741
rect 6089 7701 6101 7735
rect 6135 7732 6147 7735
rect 7282 7732 7288 7744
rect 6135 7704 7288 7732
rect 6135 7701 6147 7704
rect 6089 7695 6147 7701
rect 7282 7692 7288 7704
rect 7340 7692 7346 7744
rect 7650 7692 7656 7744
rect 7708 7732 7714 7744
rect 8297 7735 8355 7741
rect 8297 7732 8309 7735
rect 7708 7704 8309 7732
rect 7708 7692 7714 7704
rect 8297 7701 8309 7704
rect 8343 7732 8355 7735
rect 9508 7732 9536 7772
rect 11698 7760 11704 7772
rect 11756 7760 11762 7812
rect 9582 7732 9588 7744
rect 8343 7704 9588 7732
rect 8343 7701 8355 7704
rect 8297 7695 8355 7701
rect 9582 7692 9588 7704
rect 9640 7692 9646 7744
rect 13096 7732 13124 7831
rect 13188 7800 13216 7831
rect 13354 7828 13360 7840
rect 13412 7828 13418 7880
rect 13446 7828 13452 7880
rect 13504 7868 13510 7880
rect 14844 7877 14872 7908
rect 15102 7896 15108 7908
rect 15160 7896 15166 7948
rect 14829 7871 14887 7877
rect 13504 7840 13549 7868
rect 13504 7828 13510 7840
rect 14829 7837 14841 7871
rect 14875 7837 14887 7871
rect 14829 7831 14887 7837
rect 14918 7828 14924 7880
rect 14976 7868 14982 7880
rect 15289 7871 15347 7877
rect 14976 7840 15021 7868
rect 14976 7828 14982 7840
rect 15289 7837 15301 7871
rect 15335 7868 15347 7871
rect 15335 7840 15884 7868
rect 15335 7837 15347 7840
rect 15289 7831 15347 7837
rect 13188 7772 14136 7800
rect 14108 7744 14136 7772
rect 14366 7760 14372 7812
rect 14424 7800 14430 7812
rect 14734 7800 14740 7812
rect 14424 7772 14740 7800
rect 14424 7760 14430 7772
rect 14734 7760 14740 7772
rect 14792 7800 14798 7812
rect 15013 7803 15071 7809
rect 15013 7800 15025 7803
rect 14792 7772 15025 7800
rect 14792 7760 14798 7772
rect 15013 7769 15025 7772
rect 15059 7769 15071 7803
rect 15013 7763 15071 7769
rect 15151 7803 15209 7809
rect 15151 7769 15163 7803
rect 15197 7800 15209 7803
rect 15378 7800 15384 7812
rect 15197 7772 15384 7800
rect 15197 7769 15209 7772
rect 15151 7763 15209 7769
rect 15378 7760 15384 7772
rect 15436 7800 15442 7812
rect 15654 7800 15660 7812
rect 15436 7772 15660 7800
rect 15436 7760 15442 7772
rect 15654 7760 15660 7772
rect 15712 7760 15718 7812
rect 15856 7800 15884 7840
rect 15930 7828 15936 7880
rect 15988 7868 15994 7880
rect 16132 7877 16160 7976
rect 16209 7973 16221 8007
rect 16255 7973 16267 8007
rect 16850 8004 16856 8016
rect 16811 7976 16856 8004
rect 16209 7967 16267 7973
rect 16224 7918 16252 7967
rect 16850 7964 16856 7976
rect 16908 7964 16914 8016
rect 22278 8004 22284 8016
rect 17880 7976 22284 8004
rect 16761 7939 16819 7945
rect 16085 7871 16160 7877
rect 15988 7840 16033 7868
rect 15988 7828 15994 7840
rect 16085 7837 16097 7871
rect 16131 7840 16160 7871
rect 16206 7866 16212 7918
rect 16264 7866 16270 7918
rect 16761 7905 16773 7939
rect 16807 7936 16819 7939
rect 16942 7936 16948 7948
rect 16807 7908 16948 7936
rect 16807 7905 16819 7908
rect 16761 7899 16819 7905
rect 16942 7896 16948 7908
rect 17000 7896 17006 7948
rect 16131 7837 16143 7840
rect 16085 7831 16143 7837
rect 16298 7828 16304 7880
rect 16356 7868 16362 7880
rect 16356 7840 16401 7868
rect 16356 7828 16362 7840
rect 16850 7828 16856 7880
rect 16908 7868 16914 7880
rect 17037 7871 17095 7877
rect 17037 7868 17049 7871
rect 16908 7840 17049 7868
rect 16908 7828 16914 7840
rect 17037 7837 17049 7840
rect 17083 7837 17095 7871
rect 17037 7831 17095 7837
rect 16206 7800 16212 7812
rect 15856 7772 16212 7800
rect 16206 7760 16212 7772
rect 16264 7800 16270 7812
rect 17880 7800 17908 7976
rect 22278 7964 22284 7976
rect 22336 7964 22342 8016
rect 19334 7936 19340 7948
rect 18248 7908 19340 7936
rect 17957 7871 18015 7877
rect 17957 7837 17969 7871
rect 18003 7837 18015 7871
rect 17957 7831 18015 7837
rect 16264 7772 17908 7800
rect 16264 7760 16270 7772
rect 13998 7732 14004 7744
rect 13096 7704 14004 7732
rect 13998 7692 14004 7704
rect 14056 7692 14062 7744
rect 14090 7692 14096 7744
rect 14148 7732 14154 7744
rect 14918 7732 14924 7744
rect 14148 7704 14924 7732
rect 14148 7692 14154 7704
rect 14918 7692 14924 7704
rect 14976 7732 14982 7744
rect 16666 7732 16672 7744
rect 14976 7704 16672 7732
rect 14976 7692 14982 7704
rect 16666 7692 16672 7704
rect 16724 7732 16730 7744
rect 17678 7732 17684 7744
rect 16724 7704 17684 7732
rect 16724 7692 16730 7704
rect 17678 7692 17684 7704
rect 17736 7692 17742 7744
rect 17972 7732 18000 7831
rect 18046 7828 18052 7880
rect 18104 7868 18110 7880
rect 18248 7877 18276 7908
rect 19334 7896 19340 7908
rect 19392 7896 19398 7948
rect 20717 7939 20775 7945
rect 20717 7905 20729 7939
rect 20763 7936 20775 7939
rect 21269 7939 21327 7945
rect 21269 7936 21281 7939
rect 20763 7908 21281 7936
rect 20763 7905 20775 7908
rect 20717 7899 20775 7905
rect 21269 7905 21281 7908
rect 21315 7905 21327 7939
rect 21269 7899 21327 7905
rect 18233 7871 18291 7877
rect 18104 7840 18149 7868
rect 18104 7828 18110 7840
rect 18233 7837 18245 7871
rect 18279 7837 18291 7871
rect 18233 7831 18291 7837
rect 18325 7871 18383 7877
rect 18325 7837 18337 7871
rect 18371 7837 18383 7871
rect 18325 7831 18383 7837
rect 18340 7800 18368 7831
rect 18414 7828 18420 7880
rect 18472 7868 18478 7880
rect 19429 7871 19487 7877
rect 19429 7868 19441 7871
rect 18472 7840 19441 7868
rect 18472 7828 18478 7840
rect 19429 7837 19441 7840
rect 19475 7837 19487 7871
rect 19429 7831 19487 7837
rect 19613 7871 19671 7877
rect 19613 7837 19625 7871
rect 19659 7868 19671 7871
rect 20162 7868 20168 7880
rect 19659 7840 20168 7868
rect 19659 7837 19671 7840
rect 19613 7831 19671 7837
rect 20162 7828 20168 7840
rect 20220 7828 20226 7880
rect 20441 7871 20499 7877
rect 20441 7837 20453 7871
rect 20487 7837 20499 7871
rect 20441 7831 20499 7837
rect 18598 7800 18604 7812
rect 18340 7772 18604 7800
rect 18598 7760 18604 7772
rect 18656 7760 18662 7812
rect 20456 7800 20484 7831
rect 20530 7828 20536 7880
rect 20588 7868 20594 7880
rect 20809 7871 20867 7877
rect 20588 7840 20633 7868
rect 20588 7828 20594 7840
rect 20809 7837 20821 7871
rect 20855 7837 20867 7871
rect 20809 7831 20867 7837
rect 20714 7800 20720 7812
rect 20456 7772 20720 7800
rect 20714 7760 20720 7772
rect 20772 7760 20778 7812
rect 18322 7732 18328 7744
rect 17972 7704 18328 7732
rect 18322 7692 18328 7704
rect 18380 7692 18386 7744
rect 18877 7735 18935 7741
rect 18877 7701 18889 7735
rect 18923 7732 18935 7735
rect 19334 7732 19340 7744
rect 18923 7704 19340 7732
rect 18923 7701 18935 7704
rect 18877 7695 18935 7701
rect 19334 7692 19340 7704
rect 19392 7692 19398 7744
rect 20346 7692 20352 7744
rect 20404 7732 20410 7744
rect 20824 7732 20852 7831
rect 21358 7828 21364 7880
rect 21416 7868 21422 7880
rect 21453 7871 21511 7877
rect 21453 7868 21465 7871
rect 21416 7840 21465 7868
rect 21416 7828 21422 7840
rect 21453 7837 21465 7840
rect 21499 7837 21511 7871
rect 21726 7868 21732 7880
rect 21687 7840 21732 7868
rect 21453 7831 21511 7837
rect 21726 7828 21732 7840
rect 21784 7828 21790 7880
rect 22094 7760 22100 7812
rect 22152 7800 22158 7812
rect 22741 7803 22799 7809
rect 22741 7800 22753 7803
rect 22152 7772 22753 7800
rect 22152 7760 22158 7772
rect 22741 7769 22753 7772
rect 22787 7769 22799 7803
rect 22741 7763 22799 7769
rect 21634 7732 21640 7744
rect 20404 7704 20852 7732
rect 21595 7704 21640 7732
rect 20404 7692 20410 7704
rect 21634 7692 21640 7704
rect 21692 7692 21698 7744
rect 22186 7692 22192 7744
rect 22244 7732 22250 7744
rect 22281 7735 22339 7741
rect 22281 7732 22293 7735
rect 22244 7704 22293 7732
rect 22244 7692 22250 7704
rect 22281 7701 22293 7704
rect 22327 7732 22339 7735
rect 23014 7732 23020 7744
rect 22327 7704 23020 7732
rect 22327 7701 22339 7704
rect 22281 7695 22339 7701
rect 23014 7692 23020 7704
rect 23072 7692 23078 7744
rect 1104 7642 23987 7664
rect 1104 7590 6630 7642
rect 6682 7590 6694 7642
rect 6746 7590 6758 7642
rect 6810 7590 6822 7642
rect 6874 7590 6886 7642
rect 6938 7590 12311 7642
rect 12363 7590 12375 7642
rect 12427 7590 12439 7642
rect 12491 7590 12503 7642
rect 12555 7590 12567 7642
rect 12619 7590 17992 7642
rect 18044 7590 18056 7642
rect 18108 7590 18120 7642
rect 18172 7590 18184 7642
rect 18236 7590 18248 7642
rect 18300 7590 23673 7642
rect 23725 7590 23737 7642
rect 23789 7590 23801 7642
rect 23853 7590 23865 7642
rect 23917 7590 23929 7642
rect 23981 7590 23987 7642
rect 1104 7568 23987 7590
rect 2961 7531 3019 7537
rect 2961 7497 2973 7531
rect 3007 7528 3019 7531
rect 3142 7528 3148 7540
rect 3007 7500 3148 7528
rect 3007 7497 3019 7500
rect 2961 7491 3019 7497
rect 3142 7488 3148 7500
rect 3200 7488 3206 7540
rect 3234 7488 3240 7540
rect 3292 7528 3298 7540
rect 4985 7531 5043 7537
rect 3292 7500 4660 7528
rect 3292 7488 3298 7500
rect 2130 7420 2136 7472
rect 2188 7460 2194 7472
rect 2501 7463 2559 7469
rect 2501 7460 2513 7463
rect 2188 7432 2513 7460
rect 2188 7420 2194 7432
rect 2501 7429 2513 7432
rect 2547 7460 2559 7463
rect 2682 7460 2688 7472
rect 2547 7432 2688 7460
rect 2547 7429 2559 7432
rect 2501 7423 2559 7429
rect 2682 7420 2688 7432
rect 2740 7460 2746 7472
rect 4632 7469 4660 7500
rect 4985 7497 4997 7531
rect 5031 7528 5043 7531
rect 5534 7528 5540 7540
rect 5031 7500 5540 7528
rect 5031 7497 5043 7500
rect 4985 7491 5043 7497
rect 5534 7488 5540 7500
rect 5592 7488 5598 7540
rect 8110 7528 8116 7540
rect 5644 7500 8116 7528
rect 3605 7463 3663 7469
rect 3605 7460 3617 7463
rect 2740 7432 3617 7460
rect 2740 7420 2746 7432
rect 3605 7429 3617 7432
rect 3651 7429 3663 7463
rect 3605 7423 3663 7429
rect 4617 7463 4675 7469
rect 4617 7429 4629 7463
rect 4663 7460 4675 7463
rect 5644 7460 5672 7500
rect 8110 7488 8116 7500
rect 8168 7488 8174 7540
rect 8294 7488 8300 7540
rect 8352 7528 8358 7540
rect 8849 7531 8907 7537
rect 8849 7528 8861 7531
rect 8352 7500 8861 7528
rect 8352 7488 8358 7500
rect 8849 7497 8861 7500
rect 8895 7497 8907 7531
rect 8849 7491 8907 7497
rect 9306 7488 9312 7540
rect 9364 7488 9370 7540
rect 11698 7528 11704 7540
rect 10888 7500 11704 7528
rect 4663 7432 5672 7460
rect 4663 7429 4675 7432
rect 4617 7423 4675 7429
rect 6362 7420 6368 7472
rect 6420 7460 6426 7472
rect 6420 7432 7880 7460
rect 6420 7420 6426 7432
rect 2041 7395 2099 7401
rect 2041 7361 2053 7395
rect 2087 7392 2099 7395
rect 2406 7392 2412 7404
rect 2087 7364 2412 7392
rect 2087 7361 2099 7364
rect 2041 7355 2099 7361
rect 2406 7352 2412 7364
rect 2464 7352 2470 7404
rect 2774 7352 2780 7404
rect 2832 7392 2838 7404
rect 3421 7395 3479 7401
rect 2832 7364 2877 7392
rect 2832 7352 2838 7364
rect 3421 7361 3433 7395
rect 3467 7392 3479 7395
rect 3510 7392 3516 7404
rect 3467 7364 3516 7392
rect 3467 7361 3479 7364
rect 3421 7355 3479 7361
rect 3510 7352 3516 7364
rect 3568 7352 3574 7404
rect 4798 7392 4804 7404
rect 4759 7364 4804 7392
rect 4798 7352 4804 7364
rect 4856 7392 4862 7404
rect 5350 7392 5356 7404
rect 4856 7364 5356 7392
rect 4856 7352 4862 7364
rect 5350 7352 5356 7364
rect 5408 7352 5414 7404
rect 5534 7352 5540 7404
rect 5592 7392 5598 7404
rect 5718 7392 5724 7404
rect 5592 7364 5724 7392
rect 5592 7352 5598 7364
rect 5718 7352 5724 7364
rect 5776 7352 5782 7404
rect 5810 7352 5816 7404
rect 5868 7392 5874 7404
rect 7285 7395 7343 7401
rect 5868 7364 6500 7392
rect 5868 7352 5874 7364
rect 1854 7284 1860 7336
rect 1912 7324 1918 7336
rect 2685 7327 2743 7333
rect 2685 7324 2697 7327
rect 1912 7296 2697 7324
rect 1912 7284 1918 7296
rect 2685 7293 2697 7296
rect 2731 7293 2743 7327
rect 2685 7287 2743 7293
rect 2700 7256 2728 7287
rect 2866 7284 2872 7336
rect 2924 7324 2930 7336
rect 3050 7324 3056 7336
rect 2924 7296 3056 7324
rect 2924 7284 2930 7296
rect 3050 7284 3056 7296
rect 3108 7324 3114 7336
rect 5828 7324 5856 7352
rect 3108 7296 5856 7324
rect 5997 7327 6055 7333
rect 3108 7284 3114 7296
rect 5997 7293 6009 7327
rect 6043 7324 6055 7327
rect 6086 7324 6092 7336
rect 6043 7296 6092 7324
rect 6043 7293 6055 7296
rect 5997 7287 6055 7293
rect 6012 7256 6040 7287
rect 6086 7284 6092 7296
rect 6144 7324 6150 7336
rect 6362 7324 6368 7336
rect 6144 7296 6368 7324
rect 6144 7284 6150 7296
rect 6362 7284 6368 7296
rect 6420 7284 6426 7336
rect 2700 7228 6040 7256
rect 6472 7256 6500 7364
rect 7285 7361 7297 7395
rect 7331 7392 7343 7395
rect 7466 7392 7472 7404
rect 7331 7364 7472 7392
rect 7331 7361 7343 7364
rect 7285 7355 7343 7361
rect 7466 7352 7472 7364
rect 7524 7352 7530 7404
rect 7852 7401 7880 7432
rect 7926 7420 7932 7472
rect 7984 7420 7990 7472
rect 8662 7420 8668 7472
rect 8720 7460 8726 7472
rect 9324 7460 9352 7488
rect 10888 7469 10916 7500
rect 11698 7488 11704 7500
rect 11756 7488 11762 7540
rect 12253 7531 12311 7537
rect 12253 7497 12265 7531
rect 12299 7528 12311 7531
rect 12897 7531 12955 7537
rect 12897 7528 12909 7531
rect 12299 7500 12909 7528
rect 12299 7497 12311 7500
rect 12253 7491 12311 7497
rect 12897 7497 12909 7500
rect 12943 7497 12955 7531
rect 12897 7491 12955 7497
rect 12986 7488 12992 7540
rect 13044 7528 13050 7540
rect 13044 7500 13089 7528
rect 13044 7488 13050 7500
rect 13998 7488 14004 7540
rect 14056 7528 14062 7540
rect 15289 7531 15347 7537
rect 15289 7528 15301 7531
rect 14056 7500 15301 7528
rect 14056 7488 14062 7500
rect 15289 7497 15301 7500
rect 15335 7497 15347 7531
rect 15289 7491 15347 7497
rect 15470 7488 15476 7540
rect 15528 7528 15534 7540
rect 17405 7531 17463 7537
rect 15528 7500 15792 7528
rect 15528 7488 15534 7500
rect 10873 7463 10931 7469
rect 8720 7432 10272 7460
rect 8720 7420 8726 7432
rect 7837 7395 7895 7401
rect 7837 7361 7849 7395
rect 7883 7361 7895 7395
rect 7944 7392 7972 7420
rect 9033 7395 9091 7401
rect 9033 7392 9045 7395
rect 7944 7364 9045 7392
rect 7837 7355 7895 7361
rect 9033 7361 9045 7364
rect 9079 7361 9091 7395
rect 9306 7392 9312 7404
rect 9267 7364 9312 7392
rect 9033 7355 9091 7361
rect 7006 7333 7012 7336
rect 6997 7327 7012 7333
rect 6997 7293 7009 7327
rect 6997 7287 7012 7293
rect 7006 7284 7012 7287
rect 7064 7284 7070 7336
rect 7374 7284 7380 7336
rect 7432 7284 7438 7336
rect 7745 7327 7803 7333
rect 7745 7293 7757 7327
rect 7791 7293 7803 7327
rect 7745 7287 7803 7293
rect 7760 7256 7788 7287
rect 6472 7228 7788 7256
rect 7852 7256 7880 7355
rect 9306 7352 9312 7364
rect 9364 7352 9370 7404
rect 9582 7352 9588 7404
rect 9640 7392 9646 7404
rect 10244 7401 10272 7432
rect 10873 7429 10885 7463
rect 10919 7429 10931 7463
rect 10873 7423 10931 7429
rect 11238 7420 11244 7472
rect 11296 7460 11302 7472
rect 11974 7460 11980 7472
rect 11296 7432 11980 7460
rect 11296 7420 11302 7432
rect 11974 7420 11980 7432
rect 12032 7420 12038 7472
rect 12713 7463 12771 7469
rect 12713 7429 12725 7463
rect 12759 7460 12771 7463
rect 13354 7460 13360 7472
rect 12759 7432 13360 7460
rect 12759 7429 12771 7432
rect 12713 7423 12771 7429
rect 13354 7420 13360 7432
rect 13412 7420 13418 7472
rect 13538 7420 13544 7472
rect 13596 7460 13602 7472
rect 14829 7463 14887 7469
rect 13596 7432 14412 7460
rect 13596 7420 13602 7432
rect 14384 7404 14412 7432
rect 14829 7429 14841 7463
rect 14875 7460 14887 7463
rect 15378 7460 15384 7472
rect 14875 7432 15384 7460
rect 14875 7429 14887 7432
rect 14829 7423 14887 7429
rect 15378 7420 15384 7432
rect 15436 7420 15442 7472
rect 9953 7395 10011 7401
rect 9953 7392 9965 7395
rect 9640 7364 9965 7392
rect 9640 7352 9646 7364
rect 9953 7361 9965 7364
rect 9999 7361 10011 7395
rect 9953 7355 10011 7361
rect 10137 7395 10195 7401
rect 10137 7361 10149 7395
rect 10183 7361 10195 7395
rect 10137 7355 10195 7361
rect 10229 7395 10287 7401
rect 10229 7361 10241 7395
rect 10275 7361 10287 7395
rect 11146 7392 11152 7404
rect 11107 7364 11152 7392
rect 10229 7355 10287 7361
rect 7926 7284 7932 7336
rect 7984 7324 7990 7336
rect 9125 7327 9183 7333
rect 9125 7324 9137 7327
rect 7984 7296 9137 7324
rect 7984 7284 7990 7296
rect 9125 7293 9137 7296
rect 9171 7293 9183 7327
rect 9125 7287 9183 7293
rect 10152 7256 10180 7355
rect 11146 7352 11152 7364
rect 11204 7352 11210 7404
rect 11701 7395 11759 7401
rect 11701 7361 11713 7395
rect 11747 7361 11759 7395
rect 11701 7355 11759 7361
rect 11885 7395 11943 7401
rect 11885 7361 11897 7395
rect 11931 7361 11943 7395
rect 11885 7355 11943 7361
rect 12069 7395 12127 7401
rect 12069 7361 12081 7395
rect 12115 7392 12127 7395
rect 12158 7392 12164 7404
rect 12115 7364 12164 7392
rect 12115 7361 12127 7364
rect 12069 7355 12127 7361
rect 10410 7284 10416 7336
rect 10468 7324 10474 7336
rect 11716 7324 11744 7355
rect 10468 7296 11744 7324
rect 11900 7324 11928 7355
rect 12158 7352 12164 7364
rect 12216 7352 12222 7404
rect 12894 7352 12900 7404
rect 12952 7392 12958 7404
rect 13081 7395 13139 7401
rect 13081 7392 13093 7395
rect 12952 7364 13093 7392
rect 12952 7352 12958 7364
rect 13081 7361 13093 7364
rect 13127 7392 13139 7395
rect 13722 7392 13728 7404
rect 13127 7364 13728 7392
rect 13127 7361 13139 7364
rect 13081 7355 13139 7361
rect 13722 7352 13728 7364
rect 13780 7352 13786 7404
rect 14182 7392 14188 7404
rect 14143 7364 14188 7392
rect 14182 7352 14188 7364
rect 14240 7352 14246 7404
rect 14366 7392 14372 7404
rect 14327 7364 14372 7392
rect 14366 7352 14372 7364
rect 14424 7352 14430 7404
rect 14461 7395 14519 7401
rect 14461 7361 14473 7395
rect 14507 7361 14519 7395
rect 14461 7355 14519 7361
rect 12710 7324 12716 7336
rect 11900 7296 12716 7324
rect 10468 7284 10474 7296
rect 7852 7228 10180 7256
rect 11716 7256 11744 7296
rect 12710 7284 12716 7296
rect 12768 7284 12774 7336
rect 14476 7324 14504 7355
rect 14550 7352 14556 7404
rect 14608 7392 14614 7404
rect 14608 7364 14653 7392
rect 14608 7352 14614 7364
rect 14734 7352 14740 7404
rect 14792 7392 14798 7404
rect 15764 7401 15792 7500
rect 16224 7500 17356 7528
rect 15749 7395 15807 7401
rect 14792 7364 15608 7392
rect 14792 7352 14798 7364
rect 15010 7324 15016 7336
rect 14476 7296 15016 7324
rect 15010 7284 15016 7296
rect 15068 7284 15074 7336
rect 15102 7284 15108 7336
rect 15160 7324 15166 7336
rect 15580 7333 15608 7364
rect 15749 7361 15761 7395
rect 15795 7361 15807 7395
rect 15749 7355 15807 7361
rect 15473 7327 15531 7333
rect 15473 7324 15485 7327
rect 15160 7296 15485 7324
rect 15160 7284 15166 7296
rect 15473 7293 15485 7296
rect 15519 7293 15531 7327
rect 15473 7287 15531 7293
rect 15565 7327 15623 7333
rect 15565 7293 15577 7327
rect 15611 7293 15623 7327
rect 15565 7287 15623 7293
rect 12066 7256 12072 7268
rect 11716 7228 12072 7256
rect 1857 7191 1915 7197
rect 1857 7157 1869 7191
rect 1903 7188 1915 7191
rect 2038 7188 2044 7200
rect 1903 7160 2044 7188
rect 1903 7157 1915 7160
rect 1857 7151 1915 7157
rect 2038 7148 2044 7160
rect 2096 7148 2102 7200
rect 2498 7188 2504 7200
rect 2459 7160 2504 7188
rect 2498 7148 2504 7160
rect 2556 7148 2562 7200
rect 3694 7188 3700 7200
rect 3655 7160 3700 7188
rect 3694 7148 3700 7160
rect 3752 7148 3758 7200
rect 4522 7148 4528 7200
rect 4580 7188 4586 7200
rect 5074 7188 5080 7200
rect 4580 7160 5080 7188
rect 4580 7148 4586 7160
rect 5074 7148 5080 7160
rect 5132 7148 5138 7200
rect 5902 7148 5908 7200
rect 5960 7188 5966 7200
rect 7760 7188 7788 7228
rect 12066 7216 12072 7228
rect 12124 7216 12130 7268
rect 13265 7259 13323 7265
rect 13265 7225 13277 7259
rect 13311 7256 13323 7259
rect 13630 7256 13636 7268
rect 13311 7228 13636 7256
rect 13311 7225 13323 7228
rect 13265 7219 13323 7225
rect 13630 7216 13636 7228
rect 13688 7216 13694 7268
rect 15488 7256 15516 7287
rect 15654 7284 15660 7336
rect 15712 7324 15718 7336
rect 16224 7324 16252 7500
rect 16482 7420 16488 7472
rect 16540 7460 16546 7472
rect 17328 7460 17356 7500
rect 17405 7497 17417 7531
rect 17451 7528 17463 7531
rect 17862 7528 17868 7540
rect 17451 7500 17868 7528
rect 17451 7497 17463 7500
rect 17405 7491 17463 7497
rect 17862 7488 17868 7500
rect 17920 7488 17926 7540
rect 18064 7500 19564 7528
rect 18064 7460 18092 7500
rect 16540 7432 16988 7460
rect 17328 7432 18092 7460
rect 16540 7420 16546 7432
rect 16666 7352 16672 7404
rect 16724 7392 16730 7404
rect 16960 7401 16988 7432
rect 18138 7420 18144 7472
rect 18196 7460 18202 7472
rect 18598 7460 18604 7472
rect 18196 7432 18604 7460
rect 18196 7420 18202 7432
rect 18598 7420 18604 7432
rect 18656 7460 18662 7472
rect 18782 7460 18788 7472
rect 18656 7432 18788 7460
rect 18656 7420 18662 7432
rect 18782 7420 18788 7432
rect 18840 7420 18846 7472
rect 19536 7460 19564 7500
rect 19610 7488 19616 7540
rect 19668 7528 19674 7540
rect 20165 7531 20223 7537
rect 20165 7528 20177 7531
rect 19668 7500 20177 7528
rect 19668 7488 19674 7500
rect 20165 7497 20177 7500
rect 20211 7528 20223 7531
rect 21634 7528 21640 7540
rect 20211 7500 21640 7528
rect 20211 7497 20223 7500
rect 20165 7491 20223 7497
rect 21634 7488 21640 7500
rect 21692 7488 21698 7540
rect 21910 7488 21916 7540
rect 21968 7528 21974 7540
rect 22005 7531 22063 7537
rect 22005 7528 22017 7531
rect 21968 7500 22017 7528
rect 21968 7488 21974 7500
rect 22005 7497 22017 7500
rect 22051 7497 22063 7531
rect 23014 7528 23020 7540
rect 22975 7500 23020 7528
rect 22005 7491 22063 7497
rect 23014 7488 23020 7500
rect 23072 7488 23078 7540
rect 19536 7432 19748 7460
rect 16853 7395 16911 7401
rect 16853 7392 16865 7395
rect 16724 7364 16865 7392
rect 16724 7352 16730 7364
rect 16853 7361 16865 7364
rect 16899 7361 16911 7395
rect 16853 7355 16911 7361
rect 16945 7395 17003 7401
rect 16945 7361 16957 7395
rect 16991 7361 17003 7395
rect 16945 7355 17003 7361
rect 17129 7395 17187 7401
rect 17129 7361 17141 7395
rect 17175 7361 17187 7395
rect 17129 7355 17187 7361
rect 15712 7296 16252 7324
rect 15712 7284 15718 7296
rect 16390 7284 16396 7336
rect 16448 7324 16454 7336
rect 17144 7324 17172 7355
rect 17218 7352 17224 7404
rect 17276 7392 17282 7404
rect 17865 7395 17923 7401
rect 17276 7364 17321 7392
rect 17276 7352 17282 7364
rect 17865 7361 17877 7395
rect 17911 7361 17923 7395
rect 17865 7355 17923 7361
rect 17770 7324 17776 7336
rect 16448 7296 17776 7324
rect 16448 7284 16454 7296
rect 17770 7284 17776 7296
rect 17828 7284 17834 7336
rect 17880 7324 17908 7355
rect 17954 7352 17960 7404
rect 18012 7392 18018 7404
rect 18049 7395 18107 7401
rect 18049 7392 18061 7395
rect 18012 7364 18061 7392
rect 18012 7352 18018 7364
rect 18049 7361 18061 7364
rect 18095 7392 18107 7395
rect 18966 7392 18972 7404
rect 18095 7364 18828 7392
rect 18927 7364 18972 7392
rect 18095 7361 18107 7364
rect 18049 7355 18107 7361
rect 18800 7336 18828 7364
rect 18966 7352 18972 7364
rect 19024 7352 19030 7404
rect 19334 7352 19340 7404
rect 19392 7392 19398 7404
rect 19610 7392 19616 7404
rect 19392 7364 19616 7392
rect 19392 7352 19398 7364
rect 19610 7352 19616 7364
rect 19668 7352 19674 7404
rect 19720 7401 19748 7432
rect 19794 7420 19800 7472
rect 19852 7460 19858 7472
rect 20993 7463 21051 7469
rect 19852 7432 19897 7460
rect 19852 7420 19858 7432
rect 20993 7429 21005 7463
rect 21039 7460 21051 7463
rect 21266 7460 21272 7472
rect 21039 7432 21272 7460
rect 21039 7429 21051 7432
rect 20993 7423 21051 7429
rect 21266 7420 21272 7432
rect 21324 7420 21330 7472
rect 19705 7395 19763 7401
rect 19705 7361 19717 7395
rect 19751 7361 19763 7395
rect 19978 7392 19984 7404
rect 19939 7364 19984 7392
rect 19705 7355 19763 7361
rect 18138 7324 18144 7336
rect 17880 7296 18144 7324
rect 18138 7284 18144 7296
rect 18196 7284 18202 7336
rect 18230 7284 18236 7336
rect 18288 7324 18294 7336
rect 18325 7327 18383 7333
rect 18325 7324 18337 7327
rect 18288 7296 18337 7324
rect 18288 7284 18294 7296
rect 18325 7293 18337 7296
rect 18371 7293 18383 7327
rect 18325 7287 18383 7293
rect 18782 7284 18788 7336
rect 18840 7284 18846 7336
rect 15838 7256 15844 7268
rect 15488 7228 15844 7256
rect 15838 7216 15844 7228
rect 15896 7216 15902 7268
rect 16298 7216 16304 7268
rect 16356 7256 16362 7268
rect 18877 7259 18935 7265
rect 18877 7256 18889 7259
rect 16356 7228 18889 7256
rect 16356 7216 16362 7228
rect 18877 7225 18889 7228
rect 18923 7256 18935 7259
rect 19426 7256 19432 7268
rect 18923 7228 19432 7256
rect 18923 7225 18935 7228
rect 18877 7219 18935 7225
rect 19426 7216 19432 7228
rect 19484 7216 19490 7268
rect 19720 7256 19748 7355
rect 19978 7352 19984 7364
rect 20036 7392 20042 7404
rect 20625 7395 20683 7401
rect 20625 7392 20637 7395
rect 20036 7364 20637 7392
rect 20036 7352 20042 7364
rect 20625 7361 20637 7364
rect 20671 7361 20683 7395
rect 20806 7392 20812 7404
rect 20767 7364 20812 7392
rect 20625 7355 20683 7361
rect 20806 7352 20812 7364
rect 20864 7352 20870 7404
rect 21726 7352 21732 7404
rect 21784 7392 21790 7404
rect 22189 7395 22247 7401
rect 22189 7392 22201 7395
rect 21784 7364 22201 7392
rect 21784 7352 21790 7364
rect 22189 7361 22201 7364
rect 22235 7361 22247 7395
rect 22189 7355 22247 7361
rect 22278 7352 22284 7404
rect 22336 7392 22342 7404
rect 22465 7395 22523 7401
rect 22336 7364 22381 7392
rect 22336 7352 22342 7364
rect 22465 7361 22477 7395
rect 22511 7361 22523 7395
rect 22465 7355 22523 7361
rect 21266 7256 21272 7268
rect 19720 7228 21272 7256
rect 21266 7216 21272 7228
rect 21324 7256 21330 7268
rect 21542 7256 21548 7268
rect 21324 7228 21548 7256
rect 21324 7216 21330 7228
rect 21542 7216 21548 7228
rect 21600 7216 21606 7268
rect 8294 7188 8300 7200
rect 5960 7160 6005 7188
rect 7760 7160 8300 7188
rect 5960 7148 5966 7160
rect 8294 7148 8300 7160
rect 8352 7148 8358 7200
rect 9122 7188 9128 7200
rect 9083 7160 9128 7188
rect 9122 7148 9128 7160
rect 9180 7148 9186 7200
rect 9769 7191 9827 7197
rect 9769 7157 9781 7191
rect 9815 7188 9827 7191
rect 9858 7188 9864 7200
rect 9815 7160 9864 7188
rect 9815 7157 9827 7160
rect 9769 7151 9827 7157
rect 9858 7148 9864 7160
rect 9916 7148 9922 7200
rect 12084 7188 12112 7216
rect 14182 7188 14188 7200
rect 12084 7160 14188 7188
rect 14182 7148 14188 7160
rect 14240 7148 14246 7200
rect 15930 7148 15936 7200
rect 15988 7188 15994 7200
rect 17494 7188 17500 7200
rect 15988 7160 17500 7188
rect 15988 7148 15994 7160
rect 17494 7148 17500 7160
rect 17552 7188 17558 7200
rect 18233 7191 18291 7197
rect 18233 7188 18245 7191
rect 17552 7160 18245 7188
rect 17552 7148 17558 7160
rect 18233 7157 18245 7160
rect 18279 7188 18291 7191
rect 18690 7188 18696 7200
rect 18279 7160 18696 7188
rect 18279 7157 18291 7160
rect 18233 7151 18291 7157
rect 18690 7148 18696 7160
rect 18748 7148 18754 7200
rect 18966 7148 18972 7200
rect 19024 7188 19030 7200
rect 22480 7188 22508 7355
rect 22554 7352 22560 7404
rect 22612 7392 22618 7404
rect 22612 7364 22657 7392
rect 22612 7352 22618 7364
rect 19024 7160 22508 7188
rect 19024 7148 19030 7160
rect 1104 7098 23828 7120
rect 1104 7046 3790 7098
rect 3842 7046 3854 7098
rect 3906 7046 3918 7098
rect 3970 7046 3982 7098
rect 4034 7046 4046 7098
rect 4098 7046 9471 7098
rect 9523 7046 9535 7098
rect 9587 7046 9599 7098
rect 9651 7046 9663 7098
rect 9715 7046 9727 7098
rect 9779 7046 15152 7098
rect 15204 7046 15216 7098
rect 15268 7046 15280 7098
rect 15332 7046 15344 7098
rect 15396 7046 15408 7098
rect 15460 7046 20833 7098
rect 20885 7046 20897 7098
rect 20949 7046 20961 7098
rect 21013 7046 21025 7098
rect 21077 7046 21089 7098
rect 21141 7046 23828 7098
rect 1104 7024 23828 7046
rect 1762 6944 1768 6996
rect 1820 6984 1826 6996
rect 2225 6987 2283 6993
rect 2225 6984 2237 6987
rect 1820 6956 2237 6984
rect 1820 6944 1826 6956
rect 2225 6953 2237 6956
rect 2271 6984 2283 6987
rect 3510 6984 3516 6996
rect 2271 6956 3516 6984
rect 2271 6953 2283 6956
rect 2225 6947 2283 6953
rect 3510 6944 3516 6956
rect 3568 6944 3574 6996
rect 3694 6944 3700 6996
rect 3752 6984 3758 6996
rect 5074 6984 5080 6996
rect 3752 6956 5080 6984
rect 3752 6944 3758 6956
rect 2409 6919 2467 6925
rect 2409 6885 2421 6919
rect 2455 6916 2467 6919
rect 2866 6916 2872 6928
rect 2455 6888 2872 6916
rect 2455 6885 2467 6888
rect 2409 6879 2467 6885
rect 2866 6876 2872 6888
rect 2924 6876 2930 6928
rect 2961 6783 3019 6789
rect 2961 6749 2973 6783
rect 3007 6780 3019 6783
rect 3326 6780 3332 6792
rect 3007 6752 3332 6780
rect 3007 6749 3019 6752
rect 2961 6743 3019 6749
rect 3326 6740 3332 6752
rect 3384 6740 3390 6792
rect 3973 6783 4031 6789
rect 3973 6749 3985 6783
rect 4019 6749 4031 6783
rect 3973 6743 4031 6749
rect 4157 6783 4215 6789
rect 4157 6749 4169 6783
rect 4203 6780 4215 6783
rect 4264 6780 4292 6956
rect 5074 6944 5080 6956
rect 5132 6984 5138 6996
rect 5258 6984 5264 6996
rect 5132 6956 5264 6984
rect 5132 6944 5138 6956
rect 5258 6944 5264 6956
rect 5316 6944 5322 6996
rect 6454 6944 6460 6996
rect 6512 6984 6518 6996
rect 6641 6987 6699 6993
rect 6641 6984 6653 6987
rect 6512 6956 6653 6984
rect 6512 6944 6518 6956
rect 6641 6953 6653 6956
rect 6687 6953 6699 6987
rect 10594 6984 10600 6996
rect 6641 6947 6699 6953
rect 7668 6956 7972 6984
rect 10555 6956 10600 6984
rect 4890 6876 4896 6928
rect 4948 6916 4954 6928
rect 4948 6888 5212 6916
rect 4948 6876 4954 6888
rect 5076 6851 5134 6857
rect 5076 6848 5088 6851
rect 4540 6820 5088 6848
rect 4540 6792 4568 6820
rect 5076 6817 5088 6820
rect 5122 6817 5134 6851
rect 5184 6848 5212 6888
rect 5994 6876 6000 6928
rect 6052 6916 6058 6928
rect 6052 6888 6776 6916
rect 6052 6876 6058 6888
rect 5184 6820 5304 6848
rect 5076 6811 5134 6817
rect 4522 6780 4528 6792
rect 4203 6752 4292 6780
rect 4483 6752 4528 6780
rect 4203 6749 4215 6752
rect 4157 6743 4215 6749
rect 2041 6715 2099 6721
rect 2041 6681 2053 6715
rect 2087 6712 2099 6715
rect 2130 6712 2136 6724
rect 2087 6684 2136 6712
rect 2087 6681 2099 6684
rect 2041 6675 2099 6681
rect 2130 6672 2136 6684
rect 2188 6672 2194 6724
rect 3418 6712 3424 6724
rect 2240 6684 3424 6712
rect 2240 6656 2268 6684
rect 3418 6672 3424 6684
rect 3476 6672 3482 6724
rect 3988 6712 4016 6743
rect 4522 6740 4528 6752
rect 4580 6740 4586 6792
rect 5276 6789 5304 6820
rect 5350 6808 5356 6860
rect 5408 6848 5414 6860
rect 5408 6820 5453 6848
rect 5408 6808 5414 6820
rect 5902 6808 5908 6860
rect 5960 6848 5966 6860
rect 6365 6851 6423 6857
rect 6365 6848 6377 6851
rect 5960 6820 6377 6848
rect 5960 6808 5966 6820
rect 6365 6817 6377 6820
rect 6411 6817 6423 6851
rect 6748 6848 6776 6888
rect 7668 6848 7696 6956
rect 7742 6876 7748 6928
rect 7800 6876 7806 6928
rect 6748 6820 7696 6848
rect 7760 6848 7788 6876
rect 7944 6857 7972 6956
rect 10594 6944 10600 6956
rect 10652 6944 10658 6996
rect 11146 6984 11152 6996
rect 11107 6956 11152 6984
rect 11146 6944 11152 6956
rect 11204 6944 11210 6996
rect 12986 6944 12992 6996
rect 13044 6984 13050 6996
rect 13173 6987 13231 6993
rect 13173 6984 13185 6987
rect 13044 6956 13185 6984
rect 13044 6944 13050 6956
rect 13173 6953 13185 6956
rect 13219 6953 13231 6987
rect 14918 6984 14924 6996
rect 14879 6956 14924 6984
rect 13173 6947 13231 6953
rect 14918 6944 14924 6956
rect 14976 6944 14982 6996
rect 15381 6987 15439 6993
rect 15381 6953 15393 6987
rect 15427 6984 15439 6987
rect 15470 6984 15476 6996
rect 15427 6956 15476 6984
rect 15427 6953 15439 6956
rect 15381 6947 15439 6953
rect 15470 6944 15476 6956
rect 15528 6944 15534 6996
rect 15565 6987 15623 6993
rect 15565 6953 15577 6987
rect 15611 6984 15623 6987
rect 16298 6984 16304 6996
rect 15611 6956 16304 6984
rect 15611 6953 15623 6956
rect 15565 6947 15623 6953
rect 16298 6944 16304 6956
rect 16356 6984 16362 6996
rect 17586 6984 17592 6996
rect 16356 6956 16528 6984
rect 16356 6944 16362 6956
rect 8478 6876 8484 6928
rect 8536 6916 8542 6928
rect 8938 6916 8944 6928
rect 8536 6888 8944 6916
rect 8536 6876 8542 6888
rect 8938 6876 8944 6888
rect 8996 6916 9002 6928
rect 9490 6916 9496 6928
rect 8996 6888 9496 6916
rect 8996 6876 9002 6888
rect 9490 6876 9496 6888
rect 9548 6876 9554 6928
rect 11974 6876 11980 6928
rect 12032 6916 12038 6928
rect 15930 6916 15936 6928
rect 12032 6888 15936 6916
rect 12032 6876 12038 6888
rect 15930 6876 15936 6888
rect 15988 6916 15994 6928
rect 16390 6916 16396 6928
rect 15988 6888 16396 6916
rect 15988 6876 15994 6888
rect 16390 6876 16396 6888
rect 16448 6876 16454 6928
rect 16500 6925 16528 6956
rect 16592 6956 17592 6984
rect 16485 6919 16543 6925
rect 16485 6885 16497 6919
rect 16531 6885 16543 6919
rect 16485 6879 16543 6885
rect 7837 6851 7895 6857
rect 7837 6848 7849 6851
rect 7760 6820 7849 6848
rect 6365 6811 6423 6817
rect 7837 6817 7849 6820
rect 7883 6817 7895 6851
rect 7837 6811 7895 6817
rect 7929 6851 7987 6857
rect 7929 6817 7941 6851
rect 7975 6817 7987 6851
rect 7929 6811 7987 6817
rect 8021 6851 8079 6857
rect 8021 6817 8033 6851
rect 8067 6848 8079 6851
rect 8202 6848 8208 6860
rect 8067 6820 8208 6848
rect 8067 6817 8079 6820
rect 8021 6811 8079 6817
rect 8202 6808 8208 6820
rect 8260 6808 8266 6860
rect 8386 6808 8392 6860
rect 8444 6848 8450 6860
rect 9585 6851 9643 6857
rect 9585 6848 9597 6851
rect 8444 6820 9597 6848
rect 8444 6808 8450 6820
rect 9585 6817 9597 6820
rect 9631 6817 9643 6851
rect 9585 6811 9643 6817
rect 10873 6851 10931 6857
rect 10873 6817 10885 6851
rect 10919 6848 10931 6851
rect 11238 6848 11244 6860
rect 10919 6820 11244 6848
rect 10919 6817 10931 6820
rect 10873 6811 10931 6817
rect 11238 6808 11244 6820
rect 11296 6808 11302 6860
rect 13538 6848 13544 6860
rect 11348 6820 13544 6848
rect 5169 6783 5227 6789
rect 5169 6749 5181 6783
rect 5215 6749 5227 6783
rect 5169 6743 5227 6749
rect 5260 6783 5318 6789
rect 5260 6749 5272 6783
rect 5306 6749 5318 6783
rect 5260 6743 5318 6749
rect 6457 6783 6515 6789
rect 6457 6749 6469 6783
rect 6503 6780 6515 6783
rect 7098 6780 7104 6792
rect 6503 6752 7104 6780
rect 6503 6749 6515 6752
rect 6457 6743 6515 6749
rect 4338 6712 4344 6724
rect 3988 6684 4344 6712
rect 4338 6672 4344 6684
rect 4396 6672 4402 6724
rect 4433 6715 4491 6721
rect 4433 6681 4445 6715
rect 4479 6712 4491 6715
rect 4798 6712 4804 6724
rect 4479 6684 4804 6712
rect 4479 6681 4491 6684
rect 4433 6675 4491 6681
rect 4798 6672 4804 6684
rect 4856 6672 4862 6724
rect 5184 6712 5212 6743
rect 7098 6740 7104 6752
rect 7156 6740 7162 6792
rect 7466 6740 7472 6792
rect 7524 6780 7530 6792
rect 7745 6783 7803 6789
rect 7745 6780 7757 6783
rect 7524 6752 7757 6780
rect 7524 6740 7530 6752
rect 7745 6749 7757 6752
rect 7791 6749 7803 6783
rect 7745 6743 7803 6749
rect 8110 6740 8116 6792
rect 8168 6780 8174 6792
rect 9309 6783 9367 6789
rect 9309 6780 9321 6783
rect 8168 6752 9321 6780
rect 8168 6740 8174 6752
rect 9309 6749 9321 6752
rect 9355 6749 9367 6783
rect 9309 6743 9367 6749
rect 9401 6783 9459 6789
rect 9401 6749 9413 6783
rect 9447 6749 9459 6783
rect 9401 6743 9459 6749
rect 5994 6712 6000 6724
rect 5092 6684 5212 6712
rect 5955 6684 6000 6712
rect 5092 6656 5120 6684
rect 5994 6672 6000 6684
rect 6052 6672 6058 6724
rect 7190 6672 7196 6724
rect 7248 6712 7254 6724
rect 9416 6712 9444 6743
rect 9490 6740 9496 6792
rect 9548 6780 9554 6792
rect 10965 6783 11023 6789
rect 10965 6780 10977 6783
rect 9548 6752 9593 6780
rect 10060 6752 10977 6780
rect 9548 6740 9554 6752
rect 7248 6684 9444 6712
rect 7248 6672 7254 6684
rect 2222 6644 2228 6656
rect 2183 6616 2228 6644
rect 2222 6604 2228 6616
rect 2280 6604 2286 6656
rect 2682 6604 2688 6656
rect 2740 6644 2746 6656
rect 3145 6647 3203 6653
rect 3145 6644 3157 6647
rect 2740 6616 3157 6644
rect 2740 6604 2746 6616
rect 3145 6613 3157 6616
rect 3191 6613 3203 6647
rect 3145 6607 3203 6613
rect 5074 6604 5080 6656
rect 5132 6604 5138 6656
rect 5537 6647 5595 6653
rect 5537 6613 5549 6647
rect 5583 6644 5595 6647
rect 7006 6644 7012 6656
rect 5583 6616 7012 6644
rect 5583 6613 5595 6616
rect 5537 6607 5595 6613
rect 7006 6604 7012 6616
rect 7064 6604 7070 6656
rect 7101 6647 7159 6653
rect 7101 6613 7113 6647
rect 7147 6644 7159 6647
rect 7374 6644 7380 6656
rect 7147 6616 7380 6644
rect 7147 6613 7159 6616
rect 7101 6607 7159 6613
rect 7374 6604 7380 6616
rect 7432 6604 7438 6656
rect 7466 6604 7472 6656
rect 7524 6644 7530 6656
rect 8018 6644 8024 6656
rect 7524 6616 8024 6644
rect 7524 6604 7530 6616
rect 8018 6604 8024 6616
rect 8076 6604 8082 6656
rect 8202 6644 8208 6656
rect 8163 6616 8208 6644
rect 8202 6604 8208 6616
rect 8260 6604 8266 6656
rect 8570 6604 8576 6656
rect 8628 6644 8634 6656
rect 9125 6647 9183 6653
rect 9125 6644 9137 6647
rect 8628 6616 9137 6644
rect 8628 6604 8634 6616
rect 9125 6613 9137 6616
rect 9171 6613 9183 6647
rect 9125 6607 9183 6613
rect 9398 6604 9404 6656
rect 9456 6644 9462 6656
rect 10060 6644 10088 6752
rect 10965 6749 10977 6752
rect 11011 6780 11023 6783
rect 11348 6780 11376 6820
rect 11698 6780 11704 6792
rect 11011 6752 11376 6780
rect 11659 6752 11704 6780
rect 11011 6749 11023 6752
rect 10965 6743 11023 6749
rect 11698 6740 11704 6752
rect 11756 6740 11762 6792
rect 12544 6789 12572 6820
rect 13538 6808 13544 6820
rect 13596 6848 13602 6860
rect 13814 6848 13820 6860
rect 13596 6820 13820 6848
rect 13596 6808 13602 6820
rect 13814 6808 13820 6820
rect 13872 6808 13878 6860
rect 13906 6808 13912 6860
rect 13964 6848 13970 6860
rect 14369 6851 14427 6857
rect 14369 6848 14381 6851
rect 13964 6820 14381 6848
rect 13964 6808 13970 6820
rect 14369 6817 14381 6820
rect 14415 6848 14427 6851
rect 16592 6848 16620 6956
rect 17586 6944 17592 6956
rect 17644 6944 17650 6996
rect 17770 6944 17776 6996
rect 17828 6984 17834 6996
rect 20438 6984 20444 6996
rect 17828 6956 20444 6984
rect 17828 6944 17834 6956
rect 20438 6944 20444 6956
rect 20496 6984 20502 6996
rect 20496 6956 21404 6984
rect 20496 6944 20502 6956
rect 17494 6876 17500 6928
rect 17552 6876 17558 6928
rect 18230 6876 18236 6928
rect 18288 6916 18294 6928
rect 18601 6919 18659 6925
rect 18601 6916 18613 6919
rect 18288 6888 18613 6916
rect 18288 6876 18294 6888
rect 18601 6885 18613 6888
rect 18647 6916 18659 6919
rect 18966 6916 18972 6928
rect 18647 6888 18972 6916
rect 18647 6885 18659 6888
rect 18601 6879 18659 6885
rect 18966 6876 18972 6888
rect 19024 6876 19030 6928
rect 20180 6888 20484 6916
rect 14415 6820 16620 6848
rect 17512 6848 17540 6876
rect 17957 6851 18015 6857
rect 17512 6820 17632 6848
rect 14415 6817 14427 6820
rect 14369 6811 14427 6817
rect 12529 6783 12587 6789
rect 12529 6749 12541 6783
rect 12575 6780 12587 6783
rect 13078 6780 13084 6792
rect 12575 6752 12609 6780
rect 13039 6752 13084 6780
rect 12575 6749 12587 6752
rect 12529 6743 12587 6749
rect 13078 6740 13084 6752
rect 13136 6740 13142 6792
rect 13170 6740 13176 6792
rect 13228 6780 13234 6792
rect 13265 6783 13323 6789
rect 13265 6780 13277 6783
rect 13228 6752 13277 6780
rect 13228 6740 13234 6752
rect 13265 6749 13277 6752
rect 13311 6749 13323 6783
rect 13265 6743 13323 6749
rect 14182 6740 14188 6792
rect 14240 6780 14246 6792
rect 16209 6783 16267 6789
rect 16209 6780 16221 6783
rect 14240 6752 16221 6780
rect 14240 6740 14246 6752
rect 16209 6749 16221 6752
rect 16255 6749 16267 6783
rect 16209 6743 16267 6749
rect 16393 6783 16451 6789
rect 16393 6749 16405 6783
rect 16439 6749 16451 6783
rect 16574 6780 16580 6792
rect 16535 6752 16580 6780
rect 16393 6743 16451 6749
rect 10505 6715 10563 6721
rect 10505 6681 10517 6715
rect 10551 6712 10563 6715
rect 11054 6712 11060 6724
rect 10551 6684 11060 6712
rect 10551 6681 10563 6684
rect 10505 6675 10563 6681
rect 11054 6672 11060 6684
rect 11112 6672 11118 6724
rect 12437 6715 12495 6721
rect 12437 6681 12449 6715
rect 12483 6712 12495 6715
rect 13096 6712 13124 6740
rect 12483 6684 13124 6712
rect 15749 6715 15807 6721
rect 12483 6681 12495 6684
rect 12437 6675 12495 6681
rect 15749 6681 15761 6715
rect 15795 6712 15807 6715
rect 15930 6712 15936 6724
rect 15795 6684 15936 6712
rect 15795 6681 15807 6684
rect 15749 6675 15807 6681
rect 15930 6672 15936 6684
rect 15988 6672 15994 6724
rect 9456 6616 10088 6644
rect 9456 6604 9462 6616
rect 10226 6604 10232 6656
rect 10284 6644 10290 6656
rect 11422 6644 11428 6656
rect 10284 6616 11428 6644
rect 10284 6604 10290 6616
rect 11422 6604 11428 6616
rect 11480 6644 11486 6656
rect 11701 6647 11759 6653
rect 11701 6644 11713 6647
rect 11480 6616 11713 6644
rect 11480 6604 11486 6616
rect 11701 6613 11713 6616
rect 11747 6613 11759 6647
rect 11701 6607 11759 6613
rect 14366 6604 14372 6656
rect 14424 6644 14430 6656
rect 15549 6647 15607 6653
rect 15549 6644 15561 6647
rect 14424 6616 15561 6644
rect 14424 6604 14430 6616
rect 15549 6613 15561 6616
rect 15595 6644 15607 6647
rect 16408 6644 16436 6743
rect 16574 6740 16580 6752
rect 16632 6740 16638 6792
rect 16669 6783 16727 6789
rect 16669 6749 16681 6783
rect 16715 6780 16727 6783
rect 16850 6780 16856 6792
rect 16715 6752 16856 6780
rect 16715 6749 16727 6752
rect 16669 6743 16727 6749
rect 16850 6740 16856 6752
rect 16908 6740 16914 6792
rect 17310 6780 17316 6792
rect 17271 6752 17316 6780
rect 17310 6740 17316 6752
rect 17368 6740 17374 6792
rect 17402 6740 17408 6792
rect 17460 6777 17466 6792
rect 17604 6789 17632 6820
rect 17957 6817 17969 6851
rect 18003 6848 18015 6851
rect 18874 6848 18880 6860
rect 18003 6820 18880 6848
rect 18003 6817 18015 6820
rect 17957 6811 18015 6817
rect 18874 6808 18880 6820
rect 18932 6808 18938 6860
rect 19794 6848 19800 6860
rect 18984 6820 19800 6848
rect 17497 6783 17555 6789
rect 17497 6777 17509 6783
rect 17460 6749 17509 6777
rect 17543 6749 17555 6783
rect 17460 6740 17466 6749
rect 17497 6743 17555 6749
rect 17589 6783 17647 6789
rect 17589 6749 17601 6783
rect 17635 6749 17647 6783
rect 17589 6743 17647 6749
rect 17678 6740 17684 6792
rect 17736 6780 17742 6792
rect 18230 6780 18236 6792
rect 17736 6752 18236 6780
rect 17736 6740 17742 6752
rect 18230 6740 18236 6752
rect 18288 6740 18294 6792
rect 18414 6780 18420 6792
rect 18375 6752 18420 6780
rect 18414 6740 18420 6752
rect 18472 6740 18478 6792
rect 18509 6783 18567 6789
rect 18509 6749 18521 6783
rect 18555 6780 18567 6783
rect 18690 6780 18696 6792
rect 18555 6752 18696 6780
rect 18555 6749 18567 6752
rect 18509 6743 18567 6749
rect 18690 6740 18696 6752
rect 18748 6740 18754 6792
rect 18984 6780 19012 6820
rect 19794 6808 19800 6820
rect 19852 6808 19858 6860
rect 20180 6848 20208 6888
rect 20346 6848 20352 6860
rect 19996 6820 20208 6848
rect 20307 6820 20352 6848
rect 18800 6752 19012 6780
rect 16592 6712 16620 6740
rect 17034 6712 17040 6724
rect 16592 6684 17040 6712
rect 17034 6672 17040 6684
rect 17092 6672 17098 6724
rect 17328 6712 17356 6740
rect 18800 6712 18828 6752
rect 19334 6740 19340 6792
rect 19392 6780 19398 6792
rect 19705 6783 19763 6789
rect 19705 6780 19717 6783
rect 19392 6752 19717 6780
rect 19392 6740 19398 6752
rect 19705 6749 19717 6752
rect 19751 6749 19763 6783
rect 19886 6780 19892 6792
rect 19847 6752 19892 6780
rect 19705 6743 19763 6749
rect 19886 6740 19892 6752
rect 19944 6740 19950 6792
rect 19996 6789 20024 6820
rect 20346 6808 20352 6820
rect 20404 6808 20410 6860
rect 20456 6848 20484 6888
rect 21266 6876 21272 6928
rect 21324 6876 21330 6928
rect 20530 6848 20536 6860
rect 20456 6820 20536 6848
rect 20530 6808 20536 6820
rect 20588 6808 20594 6860
rect 20714 6808 20720 6860
rect 20772 6848 20778 6860
rect 20809 6851 20867 6857
rect 20809 6848 20821 6851
rect 20772 6820 20821 6848
rect 20772 6808 20778 6820
rect 20809 6817 20821 6820
rect 20855 6817 20867 6851
rect 21284 6848 21312 6876
rect 20809 6811 20867 6817
rect 21100 6820 21312 6848
rect 21376 6848 21404 6956
rect 22005 6919 22063 6925
rect 22005 6885 22017 6919
rect 22051 6885 22063 6919
rect 22005 6879 22063 6885
rect 22020 6848 22048 6879
rect 21376 6820 22048 6848
rect 19981 6783 20039 6789
rect 19981 6749 19993 6783
rect 20027 6749 20039 6783
rect 19981 6743 20039 6749
rect 20070 6740 20076 6792
rect 20128 6780 20134 6792
rect 20622 6780 20628 6792
rect 20128 6752 20628 6780
rect 20128 6740 20134 6752
rect 20622 6740 20628 6752
rect 20680 6740 20686 6792
rect 21100 6789 21128 6820
rect 21085 6783 21143 6789
rect 21085 6749 21097 6783
rect 21131 6749 21143 6783
rect 21085 6743 21143 6749
rect 21177 6783 21235 6789
rect 21177 6749 21189 6783
rect 21223 6749 21235 6783
rect 21177 6743 21235 6749
rect 21269 6783 21327 6789
rect 21269 6749 21281 6783
rect 21315 6749 21327 6783
rect 21450 6780 21456 6792
rect 21411 6752 21456 6780
rect 21269 6743 21327 6749
rect 17328 6684 18828 6712
rect 18874 6672 18880 6724
rect 18932 6712 18938 6724
rect 18932 6684 18977 6712
rect 18932 6672 18938 6684
rect 19794 6672 19800 6724
rect 19852 6712 19858 6724
rect 21192 6712 21220 6743
rect 19852 6684 21220 6712
rect 21284 6712 21312 6743
rect 21450 6740 21456 6752
rect 21508 6740 21514 6792
rect 22189 6783 22247 6789
rect 22189 6780 22201 6783
rect 22066 6752 22201 6780
rect 22066 6712 22094 6752
rect 22189 6749 22201 6752
rect 22235 6749 22247 6783
rect 22189 6743 22247 6749
rect 21284 6684 22094 6712
rect 19852 6672 19858 6684
rect 15595 6616 16436 6644
rect 16853 6647 16911 6653
rect 15595 6613 15607 6616
rect 15549 6607 15607 6613
rect 16853 6613 16865 6647
rect 16899 6644 16911 6647
rect 18414 6644 18420 6656
rect 16899 6616 18420 6644
rect 16899 6613 16911 6616
rect 16853 6607 16911 6613
rect 18414 6604 18420 6616
rect 18472 6604 18478 6656
rect 18782 6644 18788 6656
rect 18743 6616 18788 6644
rect 18782 6604 18788 6616
rect 18840 6604 18846 6656
rect 19334 6604 19340 6656
rect 19392 6644 19398 6656
rect 19702 6644 19708 6656
rect 19392 6616 19708 6644
rect 19392 6604 19398 6616
rect 19702 6604 19708 6616
rect 19760 6644 19766 6656
rect 21284 6644 21312 6684
rect 19760 6616 21312 6644
rect 19760 6604 19766 6616
rect 1104 6554 23987 6576
rect 1104 6502 6630 6554
rect 6682 6502 6694 6554
rect 6746 6502 6758 6554
rect 6810 6502 6822 6554
rect 6874 6502 6886 6554
rect 6938 6502 12311 6554
rect 12363 6502 12375 6554
rect 12427 6502 12439 6554
rect 12491 6502 12503 6554
rect 12555 6502 12567 6554
rect 12619 6502 17992 6554
rect 18044 6502 18056 6554
rect 18108 6502 18120 6554
rect 18172 6502 18184 6554
rect 18236 6502 18248 6554
rect 18300 6502 23673 6554
rect 23725 6502 23737 6554
rect 23789 6502 23801 6554
rect 23853 6502 23865 6554
rect 23917 6502 23929 6554
rect 23981 6502 23987 6554
rect 1104 6480 23987 6502
rect 3418 6400 3424 6452
rect 3476 6440 3482 6452
rect 4249 6443 4307 6449
rect 4249 6440 4261 6443
rect 3476 6412 4261 6440
rect 3476 6400 3482 6412
rect 4249 6409 4261 6412
rect 4295 6409 4307 6443
rect 4249 6403 4307 6409
rect 4338 6400 4344 6452
rect 4396 6440 4402 6452
rect 4890 6440 4896 6452
rect 4396 6412 4896 6440
rect 4396 6400 4402 6412
rect 4890 6400 4896 6412
rect 4948 6400 4954 6452
rect 5166 6440 5172 6452
rect 5127 6412 5172 6440
rect 5166 6400 5172 6412
rect 5224 6400 5230 6452
rect 5261 6443 5319 6449
rect 5261 6409 5273 6443
rect 5307 6440 5319 6443
rect 5626 6440 5632 6452
rect 5307 6412 5632 6440
rect 5307 6409 5319 6412
rect 5261 6403 5319 6409
rect 5626 6400 5632 6412
rect 5684 6400 5690 6452
rect 6546 6440 6552 6452
rect 6380 6412 6552 6440
rect 1854 6372 1860 6384
rect 1688 6344 1860 6372
rect 1688 6313 1716 6344
rect 1854 6332 1860 6344
rect 1912 6332 1918 6384
rect 2130 6332 2136 6384
rect 2188 6372 2194 6384
rect 2188 6344 2774 6372
rect 2188 6332 2194 6344
rect 1673 6307 1731 6313
rect 1673 6273 1685 6307
rect 1719 6273 1731 6307
rect 1673 6267 1731 6273
rect 1762 6264 1768 6316
rect 1820 6304 1826 6316
rect 1820 6276 1865 6304
rect 1820 6264 1826 6276
rect 1946 6264 1952 6316
rect 2004 6304 2010 6316
rect 2593 6307 2651 6313
rect 2004 6276 2049 6304
rect 2004 6264 2010 6276
rect 2593 6273 2605 6307
rect 2639 6273 2651 6307
rect 2746 6304 2774 6344
rect 3602 6332 3608 6384
rect 3660 6372 3666 6384
rect 3789 6375 3847 6381
rect 3789 6372 3801 6375
rect 3660 6344 3801 6372
rect 3660 6332 3666 6344
rect 3789 6341 3801 6344
rect 3835 6372 3847 6375
rect 4522 6372 4528 6384
rect 3835 6344 4528 6372
rect 3835 6341 3847 6344
rect 3789 6335 3847 6341
rect 4522 6332 4528 6344
rect 4580 6372 4586 6384
rect 4985 6375 5043 6381
rect 4985 6372 4997 6375
rect 4580 6344 4997 6372
rect 4580 6332 4586 6344
rect 4985 6341 4997 6344
rect 5031 6341 5043 6375
rect 6380 6372 6408 6412
rect 6546 6400 6552 6412
rect 6604 6440 6610 6452
rect 7190 6440 7196 6452
rect 6604 6412 6960 6440
rect 7151 6412 7196 6440
rect 6604 6400 6610 6412
rect 4985 6335 5043 6341
rect 5092 6344 6408 6372
rect 2869 6307 2927 6313
rect 2869 6304 2881 6307
rect 2746 6276 2881 6304
rect 2593 6267 2651 6273
rect 2869 6273 2881 6276
rect 2915 6273 2927 6307
rect 2869 6267 2927 6273
rect 3237 6307 3295 6313
rect 3237 6273 3249 6307
rect 3283 6304 3295 6307
rect 5092 6304 5120 6344
rect 6454 6332 6460 6384
rect 6512 6372 6518 6384
rect 6932 6381 6960 6412
rect 7190 6400 7196 6412
rect 7248 6400 7254 6452
rect 7929 6443 7987 6449
rect 7929 6409 7941 6443
rect 7975 6440 7987 6443
rect 9030 6440 9036 6452
rect 7975 6412 8616 6440
rect 8991 6412 9036 6440
rect 7975 6409 7987 6412
rect 7929 6403 7987 6409
rect 6825 6375 6883 6381
rect 6825 6372 6837 6375
rect 6512 6344 6837 6372
rect 6512 6332 6518 6344
rect 6825 6341 6837 6344
rect 6871 6341 6883 6375
rect 6825 6335 6883 6341
rect 6917 6375 6975 6381
rect 6917 6341 6929 6375
rect 6963 6341 6975 6375
rect 6917 6335 6975 6341
rect 3283 6276 5120 6304
rect 5353 6307 5411 6313
rect 3283 6273 3295 6276
rect 3237 6267 3295 6273
rect 5353 6273 5365 6307
rect 5399 6304 5411 6307
rect 5810 6304 5816 6316
rect 5399 6276 5816 6304
rect 5399 6273 5411 6276
rect 5353 6267 5411 6273
rect 1578 6196 1584 6248
rect 1636 6236 1642 6248
rect 1857 6239 1915 6245
rect 1857 6236 1869 6239
rect 1636 6208 1869 6236
rect 1636 6196 1642 6208
rect 1857 6205 1869 6208
rect 1903 6205 1915 6239
rect 1857 6199 1915 6205
rect 2038 6196 2044 6248
rect 2096 6236 2102 6248
rect 2608 6236 2636 6267
rect 5810 6264 5816 6276
rect 5868 6264 5874 6316
rect 6549 6307 6607 6313
rect 6549 6273 6561 6307
rect 6595 6273 6607 6307
rect 6549 6267 6607 6273
rect 2096 6208 2636 6236
rect 2096 6196 2102 6208
rect 2608 6168 2636 6208
rect 3053 6239 3111 6245
rect 3053 6205 3065 6239
rect 3099 6236 3111 6239
rect 4246 6236 4252 6248
rect 3099 6208 4252 6236
rect 3099 6205 3111 6208
rect 3053 6199 3111 6205
rect 4246 6196 4252 6208
rect 4304 6196 4310 6248
rect 3694 6168 3700 6180
rect 2608 6140 3700 6168
rect 3694 6128 3700 6140
rect 3752 6128 3758 6180
rect 3786 6128 3792 6180
rect 3844 6168 3850 6180
rect 3844 6140 3889 6168
rect 3844 6128 3850 6140
rect 4890 6128 4896 6180
rect 4948 6168 4954 6180
rect 5537 6171 5595 6177
rect 5537 6168 5549 6171
rect 4948 6140 5549 6168
rect 4948 6128 4954 6140
rect 5537 6137 5549 6140
rect 5583 6137 5595 6171
rect 6564 6168 6592 6267
rect 6638 6264 6644 6316
rect 6696 6304 6702 6316
rect 7098 6313 7104 6316
rect 7055 6307 7104 6313
rect 7055 6304 7067 6307
rect 6696 6276 6741 6304
rect 7011 6276 7067 6304
rect 6696 6264 6702 6276
rect 7055 6273 7067 6276
rect 7101 6273 7104 6307
rect 7055 6267 7104 6273
rect 7098 6264 7104 6267
rect 7156 6304 7162 6316
rect 7558 6304 7564 6316
rect 7156 6276 7564 6304
rect 7156 6264 7162 6276
rect 7558 6264 7564 6276
rect 7616 6304 7622 6316
rect 8018 6304 8024 6316
rect 7616 6276 8024 6304
rect 7616 6264 7622 6276
rect 8018 6264 8024 6276
rect 8076 6264 8082 6316
rect 6730 6196 6736 6248
rect 6788 6236 6794 6248
rect 8128 6236 8156 6412
rect 8478 6372 8484 6384
rect 8404 6344 8484 6372
rect 8404 6313 8432 6344
rect 8478 6332 8484 6344
rect 8536 6332 8542 6384
rect 8588 6372 8616 6412
rect 9030 6400 9036 6412
rect 9088 6400 9094 6452
rect 9306 6400 9312 6452
rect 9364 6440 9370 6452
rect 9493 6443 9551 6449
rect 9493 6440 9505 6443
rect 9364 6412 9505 6440
rect 9364 6400 9370 6412
rect 9493 6409 9505 6412
rect 9539 6409 9551 6443
rect 11149 6443 11207 6449
rect 9493 6403 9551 6409
rect 9646 6412 11100 6440
rect 9646 6372 9674 6412
rect 8588 6344 9674 6372
rect 11072 6372 11100 6412
rect 11149 6409 11161 6443
rect 11195 6440 11207 6443
rect 11790 6440 11796 6452
rect 11195 6412 11796 6440
rect 11195 6409 11207 6412
rect 11149 6403 11207 6409
rect 11790 6400 11796 6412
rect 11848 6400 11854 6452
rect 16206 6440 16212 6452
rect 16167 6412 16212 6440
rect 16206 6400 16212 6412
rect 16264 6400 16270 6452
rect 17037 6443 17095 6449
rect 17037 6409 17049 6443
rect 17083 6440 17095 6443
rect 18138 6440 18144 6452
rect 17083 6412 18144 6440
rect 17083 6409 17095 6412
rect 17037 6403 17095 6409
rect 11698 6372 11704 6384
rect 11072 6344 11704 6372
rect 11698 6332 11704 6344
rect 11756 6332 11762 6384
rect 12713 6375 12771 6381
rect 12713 6341 12725 6375
rect 12759 6372 12771 6375
rect 12894 6372 12900 6384
rect 12759 6344 12900 6372
rect 12759 6341 12771 6344
rect 12713 6335 12771 6341
rect 12894 6332 12900 6344
rect 12952 6332 12958 6384
rect 13906 6372 13912 6384
rect 13867 6344 13912 6372
rect 13906 6332 13912 6344
rect 13964 6332 13970 6384
rect 15746 6372 15752 6384
rect 14660 6344 15752 6372
rect 8389 6307 8447 6313
rect 8389 6273 8401 6307
rect 8435 6273 8447 6307
rect 8570 6304 8576 6316
rect 8531 6276 8576 6304
rect 8389 6267 8447 6273
rect 8570 6264 8576 6276
rect 8628 6264 8634 6316
rect 8665 6307 8723 6313
rect 8665 6282 8677 6307
rect 8711 6282 8723 6307
rect 6788 6208 8156 6236
rect 8662 6230 8668 6282
rect 8720 6230 8726 6282
rect 8754 6264 8760 6316
rect 8812 6304 8818 6316
rect 9677 6307 9735 6313
rect 8812 6276 8905 6304
rect 8812 6264 8818 6276
rect 9677 6273 9689 6307
rect 9723 6304 9735 6307
rect 10134 6304 10140 6316
rect 9723 6276 10140 6304
rect 9723 6273 9735 6276
rect 9677 6267 9735 6273
rect 10134 6264 10140 6276
rect 10192 6264 10198 6316
rect 10689 6307 10747 6313
rect 10689 6304 10701 6307
rect 10428 6276 10701 6304
rect 6788 6196 6794 6208
rect 8772 6168 8800 6264
rect 9953 6239 10011 6245
rect 9953 6205 9965 6239
rect 9999 6236 10011 6239
rect 10226 6236 10232 6248
rect 9999 6208 10232 6236
rect 9999 6205 10011 6208
rect 9953 6199 10011 6205
rect 10226 6196 10232 6208
rect 10284 6196 10290 6248
rect 6564 6140 8800 6168
rect 9861 6171 9919 6177
rect 5537 6131 5595 6137
rect 9861 6137 9873 6171
rect 9907 6168 9919 6171
rect 10042 6168 10048 6180
rect 9907 6140 10048 6168
rect 9907 6137 9919 6140
rect 9861 6131 9919 6137
rect 10042 6128 10048 6140
rect 10100 6128 10106 6180
rect 10428 6168 10456 6276
rect 10689 6273 10701 6276
rect 10735 6273 10747 6307
rect 10689 6267 10747 6273
rect 10870 6264 10876 6316
rect 10928 6304 10934 6316
rect 11977 6307 12035 6313
rect 10928 6276 10973 6304
rect 10928 6264 10934 6276
rect 11977 6273 11989 6307
rect 12023 6304 12035 6307
rect 12434 6304 12440 6316
rect 12023 6276 12440 6304
rect 12023 6273 12035 6276
rect 11977 6267 12035 6273
rect 12434 6264 12440 6276
rect 12492 6304 12498 6316
rect 14660 6313 14688 6344
rect 15746 6332 15752 6344
rect 15804 6332 15810 6384
rect 15838 6332 15844 6384
rect 15896 6372 15902 6384
rect 17052 6372 17080 6403
rect 18138 6400 18144 6412
rect 18196 6400 18202 6452
rect 19518 6400 19524 6452
rect 19576 6440 19582 6452
rect 19797 6443 19855 6449
rect 19797 6440 19809 6443
rect 19576 6412 19809 6440
rect 19576 6400 19582 6412
rect 19797 6409 19809 6412
rect 19843 6409 19855 6443
rect 19797 6403 19855 6409
rect 20530 6400 20536 6452
rect 20588 6440 20594 6452
rect 21269 6443 21327 6449
rect 21269 6440 21281 6443
rect 20588 6412 21281 6440
rect 20588 6400 20594 6412
rect 21269 6409 21281 6412
rect 21315 6440 21327 6443
rect 21818 6440 21824 6452
rect 21315 6412 21824 6440
rect 21315 6409 21327 6412
rect 21269 6403 21327 6409
rect 21818 6400 21824 6412
rect 21876 6400 21882 6452
rect 15896 6344 17080 6372
rect 15896 6332 15902 6344
rect 17678 6332 17684 6384
rect 17736 6372 17742 6384
rect 19334 6372 19340 6384
rect 17736 6344 18276 6372
rect 19295 6344 19340 6372
rect 17736 6332 17742 6344
rect 13173 6307 13231 6313
rect 13173 6304 13185 6307
rect 12492 6276 13185 6304
rect 12492 6264 12498 6276
rect 13173 6273 13185 6276
rect 13219 6273 13231 6307
rect 13173 6267 13231 6273
rect 14461 6307 14519 6313
rect 14461 6273 14473 6307
rect 14507 6273 14519 6307
rect 14461 6267 14519 6273
rect 14645 6307 14703 6313
rect 14645 6273 14657 6307
rect 14691 6273 14703 6307
rect 14645 6267 14703 6273
rect 15381 6307 15439 6313
rect 15381 6273 15393 6307
rect 15427 6304 15439 6307
rect 15470 6304 15476 6316
rect 15427 6276 15476 6304
rect 15427 6273 15439 6276
rect 15381 6267 15439 6273
rect 10502 6196 10508 6248
rect 10560 6236 10566 6248
rect 10781 6239 10839 6245
rect 10781 6236 10793 6239
rect 10560 6208 10793 6236
rect 10560 6196 10566 6208
rect 10781 6205 10793 6208
rect 10827 6205 10839 6239
rect 10781 6199 10839 6205
rect 10965 6239 11023 6245
rect 10965 6205 10977 6239
rect 11011 6236 11023 6239
rect 11054 6236 11060 6248
rect 11011 6208 11060 6236
rect 11011 6205 11023 6208
rect 10965 6199 11023 6205
rect 11054 6196 11060 6208
rect 11112 6196 11118 6248
rect 12345 6239 12403 6245
rect 12345 6236 12357 6239
rect 11151 6208 12357 6236
rect 11151 6168 11179 6208
rect 12345 6205 12357 6208
rect 12391 6236 12403 6239
rect 13078 6236 13084 6248
rect 12391 6208 13084 6236
rect 12391 6205 12403 6208
rect 12345 6199 12403 6205
rect 13078 6196 13084 6208
rect 13136 6196 13142 6248
rect 13538 6236 13544 6248
rect 13499 6208 13544 6236
rect 13538 6196 13544 6208
rect 13596 6196 13602 6248
rect 13630 6196 13636 6248
rect 13688 6236 13694 6248
rect 14476 6236 14504 6267
rect 15470 6264 15476 6276
rect 15528 6264 15534 6316
rect 16114 6304 16120 6316
rect 16075 6276 16120 6304
rect 16114 6264 16120 6276
rect 16172 6264 16178 6316
rect 16298 6304 16304 6316
rect 16259 6276 16304 6304
rect 16298 6264 16304 6276
rect 16356 6264 16362 6316
rect 16390 6264 16396 6316
rect 16448 6304 16454 6316
rect 16853 6307 16911 6313
rect 16853 6304 16865 6307
rect 16448 6276 16865 6304
rect 16448 6264 16454 6276
rect 16853 6273 16865 6276
rect 16899 6273 16911 6307
rect 16853 6267 16911 6273
rect 17037 6307 17095 6313
rect 17037 6273 17049 6307
rect 17083 6304 17095 6307
rect 17310 6304 17316 6316
rect 17083 6276 17316 6304
rect 17083 6273 17095 6276
rect 17037 6267 17095 6273
rect 17052 6236 17080 6267
rect 17310 6264 17316 6276
rect 17368 6264 17374 6316
rect 17770 6264 17776 6316
rect 17828 6304 17834 6316
rect 18248 6313 18276 6344
rect 19334 6332 19340 6344
rect 19392 6332 19398 6384
rect 20548 6372 20576 6400
rect 20180 6344 20576 6372
rect 18141 6307 18199 6313
rect 18141 6304 18153 6307
rect 17828 6276 18153 6304
rect 17828 6264 17834 6276
rect 18141 6273 18153 6276
rect 18187 6273 18199 6307
rect 18141 6267 18199 6273
rect 18233 6307 18291 6313
rect 18233 6273 18245 6307
rect 18279 6304 18291 6307
rect 18782 6304 18788 6316
rect 18279 6276 18788 6304
rect 18279 6273 18291 6276
rect 18233 6267 18291 6273
rect 18782 6264 18788 6276
rect 18840 6264 18846 6316
rect 18966 6304 18972 6316
rect 18927 6276 18972 6304
rect 18966 6264 18972 6276
rect 19024 6264 19030 6316
rect 19150 6264 19156 6316
rect 19208 6304 19214 6316
rect 20180 6313 20208 6344
rect 19245 6307 19303 6313
rect 19245 6304 19257 6307
rect 19208 6276 19257 6304
rect 19208 6264 19214 6276
rect 19245 6273 19257 6276
rect 19291 6273 19303 6307
rect 19245 6267 19303 6273
rect 20073 6307 20131 6313
rect 20073 6273 20085 6307
rect 20119 6273 20131 6307
rect 20073 6267 20131 6273
rect 20165 6307 20223 6313
rect 20165 6273 20177 6307
rect 20211 6273 20223 6307
rect 20165 6267 20223 6273
rect 18046 6236 18052 6248
rect 13688 6208 14504 6236
rect 14844 6208 17080 6236
rect 18007 6208 18052 6236
rect 13688 6196 13694 6208
rect 10428 6140 11179 6168
rect 11882 6128 11888 6180
rect 11940 6168 11946 6180
rect 12115 6171 12173 6177
rect 12115 6168 12127 6171
rect 11940 6140 12127 6168
rect 11940 6128 11946 6140
rect 12115 6137 12127 6140
rect 12161 6137 12173 6171
rect 12115 6131 12173 6137
rect 12253 6171 12311 6177
rect 12253 6137 12265 6171
rect 12299 6168 12311 6171
rect 12894 6168 12900 6180
rect 12299 6140 12900 6168
rect 12299 6137 12311 6140
rect 12253 6131 12311 6137
rect 12894 6128 12900 6140
rect 12952 6128 12958 6180
rect 14844 6177 14872 6208
rect 18046 6196 18052 6208
rect 18104 6196 18110 6248
rect 18325 6239 18383 6245
rect 18325 6205 18337 6239
rect 18371 6205 18383 6239
rect 18325 6199 18383 6205
rect 14829 6171 14887 6177
rect 14829 6137 14841 6171
rect 14875 6137 14887 6171
rect 14829 6131 14887 6137
rect 14918 6128 14924 6180
rect 14976 6168 14982 6180
rect 17954 6168 17960 6180
rect 14976 6140 17960 6168
rect 14976 6128 14982 6140
rect 17954 6128 17960 6140
rect 18012 6128 18018 6180
rect 18138 6128 18144 6180
rect 18196 6168 18202 6180
rect 18340 6168 18368 6199
rect 19978 6196 19984 6248
rect 20036 6236 20042 6248
rect 20088 6236 20116 6267
rect 20254 6264 20260 6316
rect 20312 6304 20318 6316
rect 20453 6307 20511 6313
rect 20312 6276 20357 6304
rect 20312 6264 20318 6276
rect 20453 6273 20465 6307
rect 20499 6304 20511 6307
rect 20499 6276 20576 6304
rect 20499 6273 20511 6276
rect 20453 6267 20511 6273
rect 20548 6236 20576 6276
rect 20714 6264 20720 6316
rect 20772 6304 20778 6316
rect 21085 6307 21143 6313
rect 21085 6304 21097 6307
rect 20772 6276 21097 6304
rect 20772 6264 20778 6276
rect 21085 6273 21097 6276
rect 21131 6273 21143 6307
rect 21085 6267 21143 6273
rect 20036 6208 20116 6236
rect 20456 6208 20576 6236
rect 20901 6239 20959 6245
rect 20036 6196 20042 6208
rect 20456 6180 20484 6208
rect 20901 6205 20913 6239
rect 20947 6236 20959 6239
rect 21174 6236 21180 6248
rect 20947 6208 21180 6236
rect 20947 6205 20959 6208
rect 20901 6199 20959 6205
rect 21174 6196 21180 6208
rect 21232 6196 21238 6248
rect 19886 6168 19892 6180
rect 18196 6140 18368 6168
rect 18432 6140 19892 6168
rect 18196 6128 18202 6140
rect 2038 6060 2044 6112
rect 2096 6100 2102 6112
rect 2133 6103 2191 6109
rect 2133 6100 2145 6103
rect 2096 6072 2145 6100
rect 2096 6060 2102 6072
rect 2133 6069 2145 6072
rect 2179 6069 2191 6103
rect 2133 6063 2191 6069
rect 4525 6103 4583 6109
rect 4525 6069 4537 6103
rect 4571 6100 4583 6103
rect 5442 6100 5448 6112
rect 4571 6072 5448 6100
rect 4571 6069 4583 6072
rect 4525 6063 4583 6069
rect 5442 6060 5448 6072
rect 5500 6060 5506 6112
rect 8018 6060 8024 6112
rect 8076 6100 8082 6112
rect 10686 6100 10692 6112
rect 8076 6072 10692 6100
rect 8076 6060 8082 6072
rect 10686 6060 10692 6072
rect 10744 6060 10750 6112
rect 12802 6060 12808 6112
rect 12860 6100 12866 6112
rect 13311 6103 13369 6109
rect 13311 6100 13323 6103
rect 12860 6072 13323 6100
rect 12860 6060 12866 6072
rect 13311 6069 13323 6072
rect 13357 6069 13369 6103
rect 13311 6063 13369 6069
rect 13446 6060 13452 6112
rect 13504 6100 13510 6112
rect 14642 6100 14648 6112
rect 13504 6072 13549 6100
rect 14603 6072 14648 6100
rect 13504 6060 13510 6072
rect 14642 6060 14648 6072
rect 14700 6060 14706 6112
rect 15565 6103 15623 6109
rect 15565 6069 15577 6103
rect 15611 6100 15623 6103
rect 16114 6100 16120 6112
rect 15611 6072 16120 6100
rect 15611 6069 15623 6072
rect 15565 6063 15623 6069
rect 16114 6060 16120 6072
rect 16172 6100 16178 6112
rect 18432 6100 18460 6140
rect 19886 6128 19892 6140
rect 19944 6168 19950 6180
rect 20254 6168 20260 6180
rect 19944 6140 20260 6168
rect 19944 6128 19950 6140
rect 20254 6128 20260 6140
rect 20312 6128 20318 6180
rect 20438 6128 20444 6180
rect 20496 6128 20502 6180
rect 16172 6072 18460 6100
rect 18509 6103 18567 6109
rect 16172 6060 16178 6072
rect 18509 6069 18521 6103
rect 18555 6100 18567 6103
rect 18690 6100 18696 6112
rect 18555 6072 18696 6100
rect 18555 6069 18567 6072
rect 18509 6063 18567 6069
rect 18690 6060 18696 6072
rect 18748 6060 18754 6112
rect 19334 6060 19340 6112
rect 19392 6100 19398 6112
rect 19610 6100 19616 6112
rect 19392 6072 19616 6100
rect 19392 6060 19398 6072
rect 19610 6060 19616 6072
rect 19668 6060 19674 6112
rect 22094 6060 22100 6112
rect 22152 6100 22158 6112
rect 22152 6072 22197 6100
rect 22152 6060 22158 6072
rect 1104 6010 23828 6032
rect 1104 5958 3790 6010
rect 3842 5958 3854 6010
rect 3906 5958 3918 6010
rect 3970 5958 3982 6010
rect 4034 5958 4046 6010
rect 4098 5958 9471 6010
rect 9523 5958 9535 6010
rect 9587 5958 9599 6010
rect 9651 5958 9663 6010
rect 9715 5958 9727 6010
rect 9779 5958 15152 6010
rect 15204 5958 15216 6010
rect 15268 5958 15280 6010
rect 15332 5958 15344 6010
rect 15396 5958 15408 6010
rect 15460 5958 20833 6010
rect 20885 5958 20897 6010
rect 20949 5958 20961 6010
rect 21013 5958 21025 6010
rect 21077 5958 21089 6010
rect 21141 5958 23828 6010
rect 1104 5936 23828 5958
rect 4065 5899 4123 5905
rect 4065 5865 4077 5899
rect 4111 5896 4123 5899
rect 5166 5896 5172 5908
rect 4111 5868 5172 5896
rect 4111 5865 4123 5868
rect 4065 5859 4123 5865
rect 5166 5856 5172 5868
rect 5224 5856 5230 5908
rect 7837 5899 7895 5905
rect 7837 5865 7849 5899
rect 7883 5896 7895 5899
rect 8110 5896 8116 5908
rect 7883 5868 8116 5896
rect 7883 5865 7895 5868
rect 7837 5859 7895 5865
rect 8110 5856 8116 5868
rect 8168 5856 8174 5908
rect 8570 5856 8576 5908
rect 8628 5896 8634 5908
rect 9125 5899 9183 5905
rect 9125 5896 9137 5899
rect 8628 5868 9137 5896
rect 8628 5856 8634 5868
rect 9125 5865 9137 5868
rect 9171 5865 9183 5899
rect 9125 5859 9183 5865
rect 10229 5899 10287 5905
rect 10229 5865 10241 5899
rect 10275 5896 10287 5899
rect 11238 5896 11244 5908
rect 10275 5868 11244 5896
rect 10275 5865 10287 5868
rect 10229 5859 10287 5865
rect 1486 5788 1492 5840
rect 1544 5828 1550 5840
rect 2317 5831 2375 5837
rect 2317 5828 2329 5831
rect 1544 5800 2329 5828
rect 1544 5788 1550 5800
rect 2317 5797 2329 5800
rect 2363 5797 2375 5831
rect 7466 5828 7472 5840
rect 2317 5791 2375 5797
rect 6104 5800 7472 5828
rect 1578 5720 1584 5772
rect 1636 5760 1642 5772
rect 2682 5760 2688 5772
rect 1636 5732 2452 5760
rect 1636 5720 1642 5732
rect 1946 5692 1952 5704
rect 1859 5664 1952 5692
rect 1946 5652 1952 5664
rect 2004 5652 2010 5704
rect 2133 5695 2191 5701
rect 2133 5661 2145 5695
rect 2179 5661 2191 5695
rect 2133 5655 2191 5661
rect 1964 5556 1992 5652
rect 2148 5624 2176 5655
rect 2222 5652 2228 5704
rect 2280 5692 2286 5704
rect 2424 5701 2452 5732
rect 2516 5732 2688 5760
rect 2409 5695 2467 5701
rect 2280 5664 2325 5692
rect 2280 5652 2286 5664
rect 2409 5661 2421 5695
rect 2455 5661 2467 5695
rect 2409 5655 2467 5661
rect 2314 5624 2320 5636
rect 2148 5596 2320 5624
rect 2314 5584 2320 5596
rect 2372 5584 2378 5636
rect 2516 5624 2544 5732
rect 2682 5720 2688 5732
rect 2740 5760 2746 5772
rect 2740 5732 4016 5760
rect 2740 5720 2746 5732
rect 3053 5695 3111 5701
rect 3053 5692 3065 5695
rect 2424 5596 2544 5624
rect 2608 5664 3065 5692
rect 2222 5556 2228 5568
rect 1964 5528 2228 5556
rect 2222 5516 2228 5528
rect 2280 5556 2286 5568
rect 2424 5556 2452 5596
rect 2280 5528 2452 5556
rect 2280 5516 2286 5528
rect 2498 5516 2504 5568
rect 2556 5556 2562 5568
rect 2608 5565 2636 5664
rect 3053 5661 3065 5664
rect 3099 5661 3111 5695
rect 3053 5655 3111 5661
rect 3237 5695 3295 5701
rect 3237 5661 3249 5695
rect 3283 5692 3295 5695
rect 3602 5692 3608 5704
rect 3283 5664 3608 5692
rect 3283 5661 3295 5664
rect 3237 5655 3295 5661
rect 3602 5652 3608 5664
rect 3660 5652 3666 5704
rect 3988 5701 4016 5732
rect 4614 5720 4620 5772
rect 4672 5760 4678 5772
rect 4672 5732 5120 5760
rect 4672 5720 4678 5732
rect 5092 5704 5120 5732
rect 6104 5704 6132 5800
rect 7466 5788 7472 5800
rect 7524 5788 7530 5840
rect 9766 5788 9772 5840
rect 9824 5828 9830 5840
rect 10042 5828 10048 5840
rect 9824 5800 10048 5828
rect 9824 5788 9830 5800
rect 10042 5788 10048 5800
rect 10100 5788 10106 5840
rect 10410 5828 10416 5840
rect 10371 5800 10416 5828
rect 10410 5788 10416 5800
rect 10468 5788 10474 5840
rect 11164 5837 11192 5868
rect 11238 5856 11244 5868
rect 11296 5856 11302 5908
rect 11514 5856 11520 5908
rect 11572 5896 11578 5908
rect 12253 5899 12311 5905
rect 12253 5896 12265 5899
rect 11572 5868 12265 5896
rect 11572 5856 11578 5868
rect 12253 5865 12265 5868
rect 12299 5896 12311 5899
rect 12802 5896 12808 5908
rect 12299 5868 12808 5896
rect 12299 5865 12311 5868
rect 12253 5859 12311 5865
rect 12802 5856 12808 5868
rect 12860 5856 12866 5908
rect 12894 5856 12900 5908
rect 12952 5896 12958 5908
rect 13354 5896 13360 5908
rect 12952 5868 13360 5896
rect 12952 5856 12958 5868
rect 13354 5856 13360 5868
rect 13412 5856 13418 5908
rect 13906 5856 13912 5908
rect 13964 5896 13970 5908
rect 14277 5899 14335 5905
rect 14277 5896 14289 5899
rect 13964 5868 14289 5896
rect 13964 5856 13970 5868
rect 14277 5865 14289 5868
rect 14323 5865 14335 5899
rect 14277 5859 14335 5865
rect 14645 5899 14703 5905
rect 14645 5865 14657 5899
rect 14691 5896 14703 5899
rect 14826 5896 14832 5908
rect 14691 5868 14832 5896
rect 14691 5865 14703 5868
rect 14645 5859 14703 5865
rect 14826 5856 14832 5868
rect 14884 5856 14890 5908
rect 16669 5899 16727 5905
rect 16669 5865 16681 5899
rect 16715 5896 16727 5899
rect 16758 5896 16764 5908
rect 16715 5868 16764 5896
rect 16715 5865 16727 5868
rect 16669 5859 16727 5865
rect 16758 5856 16764 5868
rect 16816 5856 16822 5908
rect 18233 5899 18291 5905
rect 18233 5865 18245 5899
rect 18279 5896 18291 5899
rect 18322 5896 18328 5908
rect 18279 5868 18328 5896
rect 18279 5865 18291 5868
rect 18233 5859 18291 5865
rect 18322 5856 18328 5868
rect 18380 5856 18386 5908
rect 18414 5856 18420 5908
rect 18472 5896 18478 5908
rect 18472 5868 18552 5896
rect 18472 5856 18478 5868
rect 11149 5831 11207 5837
rect 11149 5797 11161 5831
rect 11195 5828 11207 5831
rect 11195 5800 11229 5828
rect 11195 5797 11207 5800
rect 11149 5791 11207 5797
rect 12986 5788 12992 5840
rect 13044 5828 13050 5840
rect 13449 5831 13507 5837
rect 13449 5828 13461 5831
rect 13044 5800 13461 5828
rect 13044 5788 13050 5800
rect 13449 5797 13461 5800
rect 13495 5797 13507 5831
rect 13449 5791 13507 5797
rect 16025 5831 16083 5837
rect 16025 5797 16037 5831
rect 16071 5828 16083 5831
rect 17218 5828 17224 5840
rect 16071 5800 17224 5828
rect 16071 5797 16083 5800
rect 16025 5791 16083 5797
rect 17218 5788 17224 5800
rect 17276 5788 17282 5840
rect 18524 5837 18552 5868
rect 19610 5856 19616 5908
rect 19668 5896 19674 5908
rect 20438 5896 20444 5908
rect 19668 5868 20444 5896
rect 19668 5856 19674 5868
rect 20438 5856 20444 5868
rect 20496 5856 20502 5908
rect 20533 5899 20591 5905
rect 20533 5865 20545 5899
rect 20579 5896 20591 5899
rect 20622 5896 20628 5908
rect 20579 5868 20628 5896
rect 20579 5865 20591 5868
rect 20533 5859 20591 5865
rect 20622 5856 20628 5868
rect 20680 5856 20686 5908
rect 18509 5831 18567 5837
rect 18509 5797 18521 5831
rect 18555 5797 18567 5831
rect 18966 5828 18972 5840
rect 18509 5791 18567 5797
rect 18616 5800 18972 5828
rect 8202 5760 8208 5772
rect 7392 5732 8208 5760
rect 3973 5695 4031 5701
rect 3973 5661 3985 5695
rect 4019 5661 4031 5695
rect 4890 5692 4896 5704
rect 4851 5664 4896 5692
rect 3973 5655 4031 5661
rect 4890 5652 4896 5664
rect 4948 5652 4954 5704
rect 5074 5692 5080 5704
rect 4987 5664 5080 5692
rect 5074 5652 5080 5664
rect 5132 5652 5138 5704
rect 5442 5692 5448 5704
rect 5403 5664 5448 5692
rect 5442 5652 5448 5664
rect 5500 5652 5506 5704
rect 6086 5692 6092 5704
rect 6047 5664 6092 5692
rect 6086 5652 6092 5664
rect 6144 5652 6150 5704
rect 6270 5692 6276 5704
rect 6231 5664 6276 5692
rect 6270 5652 6276 5664
rect 6328 5692 6334 5704
rect 6638 5692 6644 5704
rect 6328 5664 6644 5692
rect 6328 5652 6334 5664
rect 6638 5652 6644 5664
rect 6696 5652 6702 5704
rect 7282 5692 7288 5704
rect 7243 5664 7288 5692
rect 7282 5652 7288 5664
rect 7340 5652 7346 5704
rect 7392 5701 7420 5732
rect 8202 5720 8208 5732
rect 8260 5760 8266 5772
rect 8260 5732 9352 5760
rect 8260 5720 8266 5732
rect 7377 5695 7435 5701
rect 7377 5661 7389 5695
rect 7423 5661 7435 5695
rect 7558 5692 7564 5704
rect 7519 5664 7564 5692
rect 7377 5655 7435 5661
rect 7558 5652 7564 5664
rect 7616 5652 7622 5704
rect 7650 5652 7656 5704
rect 7708 5692 7714 5704
rect 7708 5664 7753 5692
rect 7708 5652 7714 5664
rect 8294 5652 8300 5704
rect 8352 5692 8358 5704
rect 8570 5692 8576 5704
rect 8352 5664 8576 5692
rect 8352 5652 8358 5664
rect 8570 5652 8576 5664
rect 8628 5652 8634 5704
rect 9324 5701 9352 5732
rect 13078 5720 13084 5772
rect 13136 5760 13142 5772
rect 14369 5763 14427 5769
rect 14369 5760 14381 5763
rect 13136 5732 14381 5760
rect 13136 5720 13142 5732
rect 14369 5729 14381 5732
rect 14415 5729 14427 5763
rect 14369 5723 14427 5729
rect 15010 5720 15016 5772
rect 15068 5760 15074 5772
rect 15749 5763 15807 5769
rect 15749 5760 15761 5763
rect 15068 5732 15761 5760
rect 15068 5720 15074 5732
rect 15749 5729 15761 5732
rect 15795 5760 15807 5763
rect 15838 5760 15844 5772
rect 15795 5732 15844 5760
rect 15795 5729 15807 5732
rect 15749 5723 15807 5729
rect 15838 5720 15844 5732
rect 15896 5720 15902 5772
rect 18616 5760 18644 5800
rect 18966 5788 18972 5800
rect 19024 5788 19030 5840
rect 19334 5788 19340 5840
rect 19392 5828 19398 5840
rect 21177 5831 21235 5837
rect 21177 5828 21189 5831
rect 19392 5800 21189 5828
rect 19392 5788 19398 5800
rect 21177 5797 21189 5800
rect 21223 5797 21235 5831
rect 21177 5791 21235 5797
rect 18524 5732 18644 5760
rect 9309 5695 9367 5701
rect 9309 5661 9321 5695
rect 9355 5661 9367 5695
rect 9490 5692 9496 5704
rect 9451 5664 9496 5692
rect 9309 5655 9367 5661
rect 9490 5652 9496 5664
rect 9548 5652 9554 5704
rect 9585 5695 9643 5701
rect 9585 5661 9597 5695
rect 9631 5692 9643 5695
rect 9858 5692 9864 5704
rect 9631 5664 9864 5692
rect 9631 5661 9643 5664
rect 9585 5655 9643 5661
rect 9858 5652 9864 5664
rect 9916 5652 9922 5704
rect 10042 5692 10048 5704
rect 10003 5664 10048 5692
rect 10042 5652 10048 5664
rect 10100 5652 10106 5704
rect 10229 5695 10287 5701
rect 10229 5661 10241 5695
rect 10275 5692 10287 5695
rect 10778 5692 10784 5704
rect 10275 5664 10784 5692
rect 10275 5661 10287 5664
rect 10229 5655 10287 5661
rect 10778 5652 10784 5664
rect 10836 5652 10842 5704
rect 10962 5652 10968 5704
rect 11020 5692 11026 5704
rect 11057 5695 11115 5701
rect 11057 5692 11069 5695
rect 11020 5664 11069 5692
rect 11020 5652 11026 5664
rect 11057 5661 11069 5664
rect 11103 5661 11115 5695
rect 11057 5655 11115 5661
rect 11241 5695 11299 5701
rect 11241 5661 11253 5695
rect 11287 5661 11299 5695
rect 11241 5655 11299 5661
rect 11333 5695 11391 5701
rect 11333 5661 11345 5695
rect 11379 5692 11391 5695
rect 11422 5692 11428 5704
rect 11379 5664 11428 5692
rect 11379 5661 11391 5664
rect 11333 5655 11391 5661
rect 6549 5627 6607 5633
rect 6549 5593 6561 5627
rect 6595 5624 6607 5627
rect 8202 5624 8208 5636
rect 6595 5596 8208 5624
rect 6595 5593 6607 5596
rect 6549 5587 6607 5593
rect 8202 5584 8208 5596
rect 8260 5584 8266 5636
rect 10796 5624 10824 5652
rect 11256 5624 11284 5655
rect 11422 5652 11428 5664
rect 11480 5652 11486 5704
rect 11609 5695 11667 5701
rect 11609 5661 11621 5695
rect 11655 5692 11667 5695
rect 13541 5695 13599 5701
rect 11655 5664 12434 5692
rect 11655 5661 11667 5664
rect 11609 5655 11667 5661
rect 12406 5636 12434 5664
rect 13541 5661 13553 5695
rect 13587 5692 13599 5695
rect 13630 5692 13636 5704
rect 13587 5664 13636 5692
rect 13587 5661 13599 5664
rect 13541 5655 13599 5661
rect 13630 5652 13636 5664
rect 13688 5652 13694 5704
rect 13725 5695 13783 5701
rect 13725 5661 13737 5695
rect 13771 5661 13783 5695
rect 13725 5655 13783 5661
rect 10796 5596 11284 5624
rect 11882 5584 11888 5636
rect 11940 5624 11946 5636
rect 12161 5627 12219 5633
rect 12161 5624 12173 5627
rect 11940 5596 12173 5624
rect 11940 5584 11946 5596
rect 12161 5593 12173 5596
rect 12207 5593 12219 5627
rect 12406 5596 12440 5636
rect 12161 5587 12219 5593
rect 12434 5584 12440 5596
rect 12492 5624 12498 5636
rect 13740 5624 13768 5655
rect 13814 5652 13820 5704
rect 13872 5692 13878 5704
rect 14277 5695 14335 5701
rect 14277 5692 14289 5695
rect 13872 5664 14289 5692
rect 13872 5652 13878 5664
rect 14277 5661 14289 5664
rect 14323 5661 14335 5695
rect 14277 5655 14335 5661
rect 15657 5695 15715 5701
rect 15657 5661 15669 5695
rect 15703 5661 15715 5695
rect 16482 5692 16488 5704
rect 16443 5664 16488 5692
rect 15657 5655 15715 5661
rect 14642 5624 14648 5636
rect 12492 5596 14648 5624
rect 12492 5584 12498 5596
rect 14642 5584 14648 5596
rect 14700 5584 14706 5636
rect 2593 5559 2651 5565
rect 2593 5556 2605 5559
rect 2556 5528 2605 5556
rect 2556 5516 2562 5528
rect 2593 5525 2605 5528
rect 2639 5525 2651 5559
rect 2593 5519 2651 5525
rect 3145 5559 3203 5565
rect 3145 5525 3157 5559
rect 3191 5556 3203 5559
rect 4246 5556 4252 5568
rect 3191 5528 4252 5556
rect 3191 5525 3203 5528
rect 3145 5519 3203 5525
rect 4246 5516 4252 5528
rect 4304 5516 4310 5568
rect 4430 5516 4436 5568
rect 4488 5556 4494 5568
rect 6730 5556 6736 5568
rect 4488 5528 6736 5556
rect 4488 5516 4494 5528
rect 6730 5516 6736 5528
rect 6788 5516 6794 5568
rect 8294 5516 8300 5568
rect 8352 5556 8358 5568
rect 8481 5559 8539 5565
rect 8481 5556 8493 5559
rect 8352 5528 8493 5556
rect 8352 5516 8358 5528
rect 8481 5525 8493 5528
rect 8527 5556 8539 5559
rect 9306 5556 9312 5568
rect 8527 5528 9312 5556
rect 8527 5525 8539 5528
rect 8481 5519 8539 5525
rect 9306 5516 9312 5528
rect 9364 5516 9370 5568
rect 13170 5516 13176 5568
rect 13228 5556 13234 5568
rect 15672 5556 15700 5655
rect 16482 5652 16488 5664
rect 16540 5652 16546 5704
rect 16666 5692 16672 5704
rect 16627 5664 16672 5692
rect 16666 5652 16672 5664
rect 16724 5652 16730 5704
rect 16942 5652 16948 5704
rect 17000 5692 17006 5704
rect 17313 5695 17371 5701
rect 17313 5692 17325 5695
rect 17000 5664 17325 5692
rect 17000 5652 17006 5664
rect 17313 5661 17325 5664
rect 17359 5661 17371 5695
rect 17313 5655 17371 5661
rect 18322 5652 18328 5704
rect 18380 5692 18386 5704
rect 18417 5695 18475 5701
rect 18417 5692 18429 5695
rect 18380 5664 18429 5692
rect 18380 5652 18386 5664
rect 18417 5661 18429 5664
rect 18463 5661 18475 5695
rect 18524 5692 18552 5732
rect 18690 5720 18696 5772
rect 18748 5760 18754 5772
rect 18748 5732 18793 5760
rect 18748 5720 18754 5732
rect 19150 5720 19156 5772
rect 19208 5760 19214 5772
rect 19208 5732 20392 5760
rect 19208 5720 19214 5732
rect 20364 5701 20392 5732
rect 18601 5695 18659 5701
rect 18601 5692 18613 5695
rect 18524 5664 18613 5692
rect 18417 5655 18475 5661
rect 18601 5661 18613 5664
rect 18647 5661 18659 5695
rect 18601 5655 18659 5661
rect 18877 5695 18935 5701
rect 18877 5661 18889 5695
rect 18923 5692 18935 5695
rect 20349 5695 20407 5701
rect 18923 5664 19748 5692
rect 18923 5661 18935 5664
rect 18877 5655 18935 5661
rect 16684 5624 16712 5652
rect 17589 5627 17647 5633
rect 17589 5624 17601 5627
rect 16684 5596 17601 5624
rect 17589 5593 17601 5596
rect 17635 5593 17647 5627
rect 17589 5587 17647 5593
rect 18690 5584 18696 5636
rect 18748 5624 18754 5636
rect 18748 5596 19334 5624
rect 18748 5584 18754 5596
rect 19306 5568 19334 5596
rect 19426 5584 19432 5636
rect 19484 5624 19490 5636
rect 19521 5627 19579 5633
rect 19521 5624 19533 5627
rect 19484 5596 19533 5624
rect 19484 5584 19490 5596
rect 19521 5593 19533 5596
rect 19567 5593 19579 5627
rect 19521 5587 19579 5593
rect 19306 5556 19340 5568
rect 13228 5528 15700 5556
rect 19247 5528 19340 5556
rect 13228 5516 13234 5528
rect 19334 5516 19340 5528
rect 19392 5556 19398 5568
rect 19613 5559 19671 5565
rect 19613 5556 19625 5559
rect 19392 5528 19625 5556
rect 19392 5516 19398 5528
rect 19613 5525 19625 5528
rect 19659 5525 19671 5559
rect 19720 5556 19748 5664
rect 20349 5661 20361 5695
rect 20395 5661 20407 5695
rect 20349 5655 20407 5661
rect 20717 5695 20775 5701
rect 20717 5661 20729 5695
rect 20763 5661 20775 5695
rect 20717 5655 20775 5661
rect 20530 5584 20536 5636
rect 20588 5624 20594 5636
rect 20732 5624 20760 5655
rect 20588 5596 20760 5624
rect 20588 5584 20594 5596
rect 20625 5559 20683 5565
rect 20625 5556 20637 5559
rect 19720 5528 20637 5556
rect 19613 5519 19671 5525
rect 20625 5525 20637 5528
rect 20671 5525 20683 5559
rect 20625 5519 20683 5525
rect 1104 5466 23987 5488
rect 1104 5414 6630 5466
rect 6682 5414 6694 5466
rect 6746 5414 6758 5466
rect 6810 5414 6822 5466
rect 6874 5414 6886 5466
rect 6938 5414 12311 5466
rect 12363 5414 12375 5466
rect 12427 5414 12439 5466
rect 12491 5414 12503 5466
rect 12555 5414 12567 5466
rect 12619 5414 17992 5466
rect 18044 5414 18056 5466
rect 18108 5414 18120 5466
rect 18172 5414 18184 5466
rect 18236 5414 18248 5466
rect 18300 5414 23673 5466
rect 23725 5414 23737 5466
rect 23789 5414 23801 5466
rect 23853 5414 23865 5466
rect 23917 5414 23929 5466
rect 23981 5414 23987 5466
rect 1104 5392 23987 5414
rect 2774 5352 2780 5364
rect 1964 5324 2780 5352
rect 1964 5225 1992 5324
rect 2774 5312 2780 5324
rect 2832 5312 2838 5364
rect 3418 5352 3424 5364
rect 3379 5324 3424 5352
rect 3418 5312 3424 5324
rect 3476 5312 3482 5364
rect 3510 5312 3516 5364
rect 3568 5352 3574 5364
rect 5169 5355 5227 5361
rect 3568 5324 4844 5352
rect 3568 5312 3574 5324
rect 2130 5244 2136 5296
rect 2188 5284 2194 5296
rect 2501 5287 2559 5293
rect 2188 5256 2360 5284
rect 2188 5244 2194 5256
rect 1949 5219 2007 5225
rect 1949 5185 1961 5219
rect 1995 5185 2007 5219
rect 1949 5179 2007 5185
rect 2041 5219 2099 5225
rect 2041 5185 2053 5219
rect 2087 5185 2099 5219
rect 2222 5216 2228 5228
rect 2183 5188 2228 5216
rect 2041 5179 2099 5185
rect 2056 5148 2084 5179
rect 2222 5176 2228 5188
rect 2280 5176 2286 5228
rect 2332 5225 2360 5256
rect 2501 5253 2513 5287
rect 2547 5284 2559 5287
rect 2547 5256 4752 5284
rect 2547 5253 2559 5256
rect 2501 5247 2559 5253
rect 4724 5228 4752 5256
rect 2317 5219 2375 5225
rect 2317 5185 2329 5219
rect 2363 5185 2375 5219
rect 2317 5179 2375 5185
rect 3237 5219 3295 5225
rect 3237 5185 3249 5219
rect 3283 5216 3295 5219
rect 3326 5216 3332 5228
rect 3283 5188 3332 5216
rect 3283 5185 3295 5188
rect 3237 5179 3295 5185
rect 3326 5176 3332 5188
rect 3384 5176 3390 5228
rect 4706 5216 4712 5228
rect 4619 5188 4712 5216
rect 4706 5176 4712 5188
rect 4764 5176 4770 5228
rect 4816 5216 4844 5324
rect 5169 5321 5181 5355
rect 5215 5352 5227 5355
rect 6270 5352 6276 5364
rect 5215 5324 6276 5352
rect 5215 5321 5227 5324
rect 5169 5315 5227 5321
rect 6270 5312 6276 5324
rect 6328 5312 6334 5364
rect 7745 5355 7803 5361
rect 7745 5321 7757 5355
rect 7791 5352 7803 5355
rect 8662 5352 8668 5364
rect 7791 5324 8668 5352
rect 7791 5321 7803 5324
rect 7745 5315 7803 5321
rect 8662 5312 8668 5324
rect 8720 5312 8726 5364
rect 8846 5352 8852 5364
rect 8807 5324 8852 5352
rect 8846 5312 8852 5324
rect 8904 5312 8910 5364
rect 11057 5355 11115 5361
rect 11057 5321 11069 5355
rect 11103 5352 11115 5355
rect 11882 5352 11888 5364
rect 11103 5324 11888 5352
rect 11103 5321 11115 5324
rect 11057 5315 11115 5321
rect 11882 5312 11888 5324
rect 11940 5312 11946 5364
rect 13630 5312 13636 5364
rect 13688 5352 13694 5364
rect 15013 5355 15071 5361
rect 13688 5324 14688 5352
rect 13688 5312 13694 5324
rect 5626 5244 5632 5296
rect 5684 5284 5690 5296
rect 5721 5287 5779 5293
rect 5721 5284 5733 5287
rect 5684 5256 5733 5284
rect 5684 5244 5690 5256
rect 5721 5253 5733 5256
rect 5767 5253 5779 5287
rect 5721 5247 5779 5253
rect 4893 5219 4951 5225
rect 4893 5216 4905 5219
rect 4816 5188 4905 5216
rect 4893 5185 4905 5188
rect 4939 5185 4951 5219
rect 4893 5179 4951 5185
rect 4982 5176 4988 5228
rect 5040 5216 5046 5228
rect 5813 5219 5871 5225
rect 5040 5188 5085 5216
rect 5040 5176 5046 5188
rect 5813 5185 5825 5219
rect 5859 5185 5871 5219
rect 6288 5216 6316 5312
rect 6546 5244 6552 5296
rect 6604 5284 6610 5296
rect 7469 5287 7527 5293
rect 7469 5284 7481 5287
rect 6604 5256 7481 5284
rect 6604 5244 6610 5256
rect 7469 5253 7481 5256
rect 7515 5253 7527 5287
rect 7469 5247 7527 5253
rect 7834 5244 7840 5296
rect 7892 5284 7898 5296
rect 8110 5284 8116 5296
rect 7892 5256 8116 5284
rect 7892 5244 7898 5256
rect 8110 5244 8116 5256
rect 8168 5284 8174 5296
rect 9677 5287 9735 5293
rect 9677 5284 9689 5287
rect 8168 5256 9689 5284
rect 8168 5244 8174 5256
rect 9677 5253 9689 5256
rect 9723 5284 9735 5287
rect 10134 5284 10140 5296
rect 9723 5256 10140 5284
rect 9723 5253 9735 5256
rect 9677 5247 9735 5253
rect 10134 5244 10140 5256
rect 10192 5244 10198 5296
rect 10502 5244 10508 5296
rect 10560 5284 10566 5296
rect 10689 5287 10747 5293
rect 10689 5284 10701 5287
rect 10560 5256 10701 5284
rect 10560 5244 10566 5256
rect 10689 5253 10701 5256
rect 10735 5253 10747 5287
rect 10689 5247 10747 5253
rect 10905 5287 10963 5293
rect 10905 5253 10917 5287
rect 10951 5284 10963 5287
rect 11330 5284 11336 5296
rect 10951 5256 11336 5284
rect 10951 5253 10963 5256
rect 10905 5247 10963 5253
rect 11330 5244 11336 5256
rect 11388 5244 11394 5296
rect 11440 5256 12112 5284
rect 7193 5219 7251 5225
rect 7193 5216 7205 5219
rect 6288 5188 7205 5216
rect 5813 5179 5871 5185
rect 7193 5185 7205 5188
rect 7239 5185 7251 5219
rect 7374 5216 7380 5228
rect 7335 5188 7380 5216
rect 7193 5179 7251 5185
rect 2056 5120 2360 5148
rect 2332 5092 2360 5120
rect 2774 5108 2780 5160
rect 2832 5148 2838 5160
rect 3605 5151 3663 5157
rect 3605 5148 3617 5151
rect 2832 5120 3617 5148
rect 2832 5108 2838 5120
rect 3605 5117 3617 5120
rect 3651 5117 3663 5151
rect 3605 5111 3663 5117
rect 3694 5108 3700 5160
rect 3752 5148 3758 5160
rect 4801 5151 4859 5157
rect 4801 5148 4813 5151
rect 3752 5120 4813 5148
rect 3752 5108 3758 5120
rect 4801 5117 4813 5120
rect 4847 5148 4859 5151
rect 5534 5148 5540 5160
rect 4847 5120 5540 5148
rect 4847 5117 4859 5120
rect 4801 5111 4859 5117
rect 5534 5108 5540 5120
rect 5592 5108 5598 5160
rect 2314 5040 2320 5092
rect 2372 5080 2378 5092
rect 4065 5083 4123 5089
rect 4065 5080 4077 5083
rect 2372 5052 4077 5080
rect 2372 5040 2378 5052
rect 3160 5021 3188 5052
rect 4065 5049 4077 5052
rect 4111 5080 4123 5083
rect 5828 5080 5856 5179
rect 7374 5176 7380 5188
rect 7432 5176 7438 5228
rect 7561 5219 7619 5225
rect 7561 5185 7573 5219
rect 7607 5216 7619 5219
rect 7607 5188 8432 5216
rect 7607 5185 7619 5188
rect 7561 5179 7619 5185
rect 4111 5052 5856 5080
rect 4111 5049 4123 5052
rect 4065 5043 4123 5049
rect 5994 5040 6000 5092
rect 6052 5080 6058 5092
rect 8018 5080 8024 5092
rect 6052 5052 8024 5080
rect 6052 5040 6058 5052
rect 8018 5040 8024 5052
rect 8076 5040 8082 5092
rect 8404 5080 8432 5188
rect 8846 5176 8852 5228
rect 8904 5216 8910 5228
rect 9861 5219 9919 5225
rect 9861 5216 9873 5219
rect 8904 5188 9873 5216
rect 8904 5176 8910 5188
rect 9861 5185 9873 5188
rect 9907 5185 9919 5219
rect 9861 5179 9919 5185
rect 10778 5176 10784 5228
rect 10836 5216 10842 5228
rect 11440 5216 11468 5256
rect 11790 5216 11796 5228
rect 10836 5188 11468 5216
rect 11751 5188 11796 5216
rect 10836 5176 10842 5188
rect 11790 5176 11796 5188
rect 11848 5176 11854 5228
rect 11885 5219 11943 5225
rect 11885 5185 11897 5219
rect 11931 5216 11943 5219
rect 11974 5216 11980 5228
rect 11931 5188 11980 5216
rect 11931 5185 11943 5188
rect 11885 5179 11943 5185
rect 11974 5176 11980 5188
rect 12032 5176 12038 5228
rect 12084 5225 12112 5256
rect 12250 5244 12256 5296
rect 12308 5284 12314 5296
rect 12308 5256 13124 5284
rect 12308 5244 12314 5256
rect 12069 5219 12127 5225
rect 12069 5185 12081 5219
rect 12115 5216 12127 5219
rect 12710 5216 12716 5228
rect 12115 5188 12716 5216
rect 12115 5185 12127 5188
rect 12069 5179 12127 5185
rect 12710 5176 12716 5188
rect 12768 5176 12774 5228
rect 13096 5225 13124 5256
rect 13354 5244 13360 5296
rect 13412 5284 13418 5296
rect 13412 5256 13860 5284
rect 13412 5244 13418 5256
rect 13832 5228 13860 5256
rect 12805 5219 12863 5225
rect 12805 5185 12817 5219
rect 12851 5185 12863 5219
rect 12805 5179 12863 5185
rect 13081 5219 13139 5225
rect 13081 5185 13093 5219
rect 13127 5216 13139 5219
rect 13814 5216 13820 5228
rect 13127 5188 13676 5216
rect 13727 5188 13820 5216
rect 13127 5185 13139 5188
rect 13081 5179 13139 5185
rect 8478 5108 8484 5160
rect 8536 5148 8542 5160
rect 8573 5151 8631 5157
rect 8573 5148 8585 5151
rect 8536 5120 8585 5148
rect 8536 5108 8542 5120
rect 8573 5117 8585 5120
rect 8619 5117 8631 5151
rect 8754 5148 8760 5160
rect 8715 5120 8760 5148
rect 8573 5111 8631 5117
rect 8754 5108 8760 5120
rect 8812 5108 8818 5160
rect 9214 5108 9220 5160
rect 9272 5148 9278 5160
rect 10045 5151 10103 5157
rect 10045 5148 10057 5151
rect 9272 5120 10057 5148
rect 9272 5108 9278 5120
rect 10045 5117 10057 5120
rect 10091 5117 10103 5151
rect 10045 5111 10103 5117
rect 11514 5108 11520 5160
rect 11572 5148 11578 5160
rect 12820 5148 12848 5179
rect 13354 5148 13360 5160
rect 11572 5120 13360 5148
rect 11572 5108 11578 5120
rect 13354 5108 13360 5120
rect 13412 5108 13418 5160
rect 13541 5151 13599 5157
rect 13541 5117 13553 5151
rect 13587 5117 13599 5151
rect 13648 5148 13676 5188
rect 13814 5176 13820 5188
rect 13872 5176 13878 5228
rect 13906 5176 13912 5228
rect 13964 5216 13970 5228
rect 14660 5225 14688 5324
rect 15013 5321 15025 5355
rect 15059 5352 15071 5355
rect 15470 5352 15476 5364
rect 15059 5324 15476 5352
rect 15059 5321 15071 5324
rect 15013 5315 15071 5321
rect 15470 5312 15476 5324
rect 15528 5312 15534 5364
rect 15838 5312 15844 5364
rect 15896 5352 15902 5364
rect 16117 5355 16175 5361
rect 16117 5352 16129 5355
rect 15896 5324 16129 5352
rect 15896 5312 15902 5324
rect 16117 5321 16129 5324
rect 16163 5352 16175 5355
rect 16390 5352 16396 5364
rect 16163 5324 16396 5352
rect 16163 5321 16175 5324
rect 16117 5315 16175 5321
rect 16390 5312 16396 5324
rect 16448 5312 16454 5364
rect 16945 5355 17003 5361
rect 16945 5321 16957 5355
rect 16991 5352 17003 5355
rect 17126 5352 17132 5364
rect 16991 5324 17132 5352
rect 16991 5321 17003 5324
rect 16945 5315 17003 5321
rect 17126 5312 17132 5324
rect 17184 5312 17190 5364
rect 18414 5312 18420 5364
rect 18472 5352 18478 5364
rect 18785 5355 18843 5361
rect 18785 5352 18797 5355
rect 18472 5324 18797 5352
rect 18472 5312 18478 5324
rect 18785 5321 18797 5324
rect 18831 5321 18843 5355
rect 18785 5315 18843 5321
rect 18966 5312 18972 5364
rect 19024 5352 19030 5364
rect 19429 5355 19487 5361
rect 19429 5352 19441 5355
rect 19024 5324 19441 5352
rect 19024 5312 19030 5324
rect 19429 5321 19441 5324
rect 19475 5321 19487 5355
rect 19429 5315 19487 5321
rect 20441 5355 20499 5361
rect 20441 5321 20453 5355
rect 20487 5352 20499 5355
rect 20622 5352 20628 5364
rect 20487 5324 20628 5352
rect 20487 5321 20499 5324
rect 20441 5315 20499 5321
rect 14734 5244 14740 5296
rect 14792 5284 14798 5296
rect 15562 5284 15568 5296
rect 14792 5256 15568 5284
rect 14792 5244 14798 5256
rect 15562 5244 15568 5256
rect 15620 5244 15626 5296
rect 16574 5244 16580 5296
rect 16632 5284 16638 5296
rect 16632 5256 17080 5284
rect 16632 5244 16638 5256
rect 14645 5219 14703 5225
rect 13964 5188 14009 5216
rect 13964 5176 13970 5188
rect 14645 5185 14657 5219
rect 14691 5185 14703 5219
rect 14645 5179 14703 5185
rect 14829 5219 14887 5225
rect 14829 5185 14841 5219
rect 14875 5216 14887 5219
rect 16482 5216 16488 5228
rect 14875 5188 16488 5216
rect 14875 5185 14887 5188
rect 14829 5179 14887 5185
rect 16482 5176 16488 5188
rect 16540 5176 16546 5228
rect 13924 5148 13952 5176
rect 13648 5120 13952 5148
rect 14093 5151 14151 5157
rect 13541 5111 13599 5117
rect 14093 5117 14105 5151
rect 14139 5148 14151 5151
rect 16684 5148 16712 5256
rect 16850 5216 16856 5228
rect 16811 5188 16856 5216
rect 16850 5176 16856 5188
rect 16908 5176 16914 5228
rect 17052 5225 17080 5256
rect 17037 5219 17095 5225
rect 17037 5185 17049 5219
rect 17083 5185 17095 5219
rect 17144 5216 17172 5312
rect 20456 5284 20484 5315
rect 20622 5312 20628 5324
rect 20680 5312 20686 5364
rect 19904 5256 20484 5284
rect 18325 5219 18383 5225
rect 18325 5216 18337 5219
rect 17144 5188 18337 5216
rect 17037 5179 17095 5185
rect 18325 5185 18337 5188
rect 18371 5185 18383 5219
rect 18598 5216 18604 5228
rect 18559 5188 18604 5216
rect 18325 5179 18383 5185
rect 18598 5176 18604 5188
rect 18656 5176 18662 5228
rect 19610 5216 19616 5228
rect 19571 5188 19616 5216
rect 19610 5176 19616 5188
rect 19668 5176 19674 5228
rect 19904 5225 19932 5256
rect 19889 5219 19947 5225
rect 19889 5185 19901 5219
rect 19935 5185 19947 5219
rect 20346 5216 20352 5228
rect 20307 5188 20352 5216
rect 19889 5179 19947 5185
rect 20346 5176 20352 5188
rect 20404 5176 20410 5228
rect 20533 5219 20591 5225
rect 20533 5185 20545 5219
rect 20579 5216 20591 5219
rect 20714 5216 20720 5228
rect 20579 5188 20720 5216
rect 20579 5185 20591 5188
rect 20533 5179 20591 5185
rect 14139 5120 16712 5148
rect 14139 5117 14151 5120
rect 14093 5111 14151 5117
rect 9030 5080 9036 5092
rect 8404 5052 9036 5080
rect 9030 5040 9036 5052
rect 9088 5080 9094 5092
rect 9490 5080 9496 5092
rect 9088 5052 9496 5080
rect 9088 5040 9094 5052
rect 9490 5040 9496 5052
rect 9548 5040 9554 5092
rect 11238 5040 11244 5092
rect 11296 5080 11302 5092
rect 11977 5083 12035 5089
rect 11977 5080 11989 5083
rect 11296 5052 11989 5080
rect 11296 5040 11302 5052
rect 11977 5049 11989 5052
rect 12023 5080 12035 5083
rect 12342 5080 12348 5092
rect 12023 5052 12348 5080
rect 12023 5049 12035 5052
rect 11977 5043 12035 5049
rect 12342 5040 12348 5052
rect 12400 5040 12406 5092
rect 12805 5083 12863 5089
rect 12805 5049 12817 5083
rect 12851 5080 12863 5083
rect 13170 5080 13176 5092
rect 12851 5052 13176 5080
rect 12851 5049 12863 5052
rect 12805 5043 12863 5049
rect 13170 5040 13176 5052
rect 13228 5040 13234 5092
rect 13556 5080 13584 5111
rect 19426 5108 19432 5160
rect 19484 5148 19490 5160
rect 20548 5148 20576 5179
rect 20714 5176 20720 5188
rect 20772 5176 20778 5228
rect 19484 5120 20576 5148
rect 19484 5108 19490 5120
rect 13556 5052 14688 5080
rect 14660 5024 14688 5052
rect 17126 5040 17132 5092
rect 17184 5080 17190 5092
rect 18417 5083 18475 5089
rect 18417 5080 18429 5083
rect 17184 5052 18429 5080
rect 17184 5040 17190 5052
rect 18417 5049 18429 5052
rect 18463 5080 18475 5083
rect 18690 5080 18696 5092
rect 18463 5052 18696 5080
rect 18463 5049 18475 5052
rect 18417 5043 18475 5049
rect 18690 5040 18696 5052
rect 18748 5040 18754 5092
rect 20346 5040 20352 5092
rect 20404 5080 20410 5092
rect 21174 5080 21180 5092
rect 20404 5052 21180 5080
rect 20404 5040 20410 5052
rect 21174 5040 21180 5052
rect 21232 5040 21238 5092
rect 3145 5015 3203 5021
rect 3145 4981 3157 5015
rect 3191 5012 3203 5015
rect 3191 4984 3225 5012
rect 3191 4981 3203 4984
rect 3145 4975 3203 4981
rect 6270 4972 6276 5024
rect 6328 5012 6334 5024
rect 6641 5015 6699 5021
rect 6641 5012 6653 5015
rect 6328 4984 6653 5012
rect 6328 4972 6334 4984
rect 6641 4981 6653 4984
rect 6687 5012 6699 5015
rect 7282 5012 7288 5024
rect 6687 4984 7288 5012
rect 6687 4981 6699 4984
rect 6641 4975 6699 4981
rect 7282 4972 7288 4984
rect 7340 4972 7346 5024
rect 9214 5012 9220 5024
rect 9175 4984 9220 5012
rect 9214 4972 9220 4984
rect 9272 4972 9278 5024
rect 10870 5012 10876 5024
rect 10831 4984 10876 5012
rect 10870 4972 10876 4984
rect 10928 4972 10934 5024
rect 13630 5012 13636 5024
rect 13591 4984 13636 5012
rect 13630 4972 13636 4984
rect 13688 4972 13694 5024
rect 14642 5012 14648 5024
rect 14603 4984 14648 5012
rect 14642 4972 14648 4984
rect 14700 4972 14706 5024
rect 15562 4972 15568 5024
rect 15620 5012 15626 5024
rect 17497 5015 17555 5021
rect 17497 5012 17509 5015
rect 15620 4984 17509 5012
rect 15620 4972 15626 4984
rect 17497 4981 17509 4984
rect 17543 4981 17555 5015
rect 17497 4975 17555 4981
rect 19797 5015 19855 5021
rect 19797 4981 19809 5015
rect 19843 5012 19855 5015
rect 20530 5012 20536 5024
rect 19843 4984 20536 5012
rect 19843 4981 19855 4984
rect 19797 4975 19855 4981
rect 20530 4972 20536 4984
rect 20588 4972 20594 5024
rect 1104 4922 23828 4944
rect 1104 4870 3790 4922
rect 3842 4870 3854 4922
rect 3906 4870 3918 4922
rect 3970 4870 3982 4922
rect 4034 4870 4046 4922
rect 4098 4870 9471 4922
rect 9523 4870 9535 4922
rect 9587 4870 9599 4922
rect 9651 4870 9663 4922
rect 9715 4870 9727 4922
rect 9779 4870 15152 4922
rect 15204 4870 15216 4922
rect 15268 4870 15280 4922
rect 15332 4870 15344 4922
rect 15396 4870 15408 4922
rect 15460 4870 20833 4922
rect 20885 4870 20897 4922
rect 20949 4870 20961 4922
rect 21013 4870 21025 4922
rect 21077 4870 21089 4922
rect 21141 4870 23828 4922
rect 1104 4848 23828 4870
rect 1670 4808 1676 4820
rect 1583 4780 1676 4808
rect 1670 4768 1676 4780
rect 1728 4808 1734 4820
rect 2314 4808 2320 4820
rect 1728 4780 2320 4808
rect 1728 4768 1734 4780
rect 2314 4768 2320 4780
rect 2372 4768 2378 4820
rect 2498 4808 2504 4820
rect 2459 4780 2504 4808
rect 2498 4768 2504 4780
rect 2556 4768 2562 4820
rect 4062 4808 4068 4820
rect 4023 4780 4068 4808
rect 4062 4768 4068 4780
rect 4120 4768 4126 4820
rect 7377 4811 7435 4817
rect 7377 4777 7389 4811
rect 7423 4808 7435 4811
rect 7926 4808 7932 4820
rect 7423 4780 7932 4808
rect 7423 4777 7435 4780
rect 7377 4771 7435 4777
rect 7926 4768 7932 4780
rect 7984 4768 7990 4820
rect 8018 4768 8024 4820
rect 8076 4808 8082 4820
rect 8386 4808 8392 4820
rect 8076 4780 8121 4808
rect 8347 4780 8392 4808
rect 8076 4768 8082 4780
rect 8386 4768 8392 4780
rect 8444 4768 8450 4820
rect 11514 4808 11520 4820
rect 11475 4780 11520 4808
rect 11514 4768 11520 4780
rect 11572 4768 11578 4820
rect 12250 4808 12256 4820
rect 12211 4780 12256 4808
rect 12250 4768 12256 4780
rect 12308 4768 12314 4820
rect 12342 4768 12348 4820
rect 12400 4808 12406 4820
rect 13173 4811 13231 4817
rect 13173 4808 13185 4811
rect 12400 4780 13185 4808
rect 12400 4768 12406 4780
rect 13173 4777 13185 4780
rect 13219 4777 13231 4811
rect 13173 4771 13231 4777
rect 14369 4811 14427 4817
rect 14369 4777 14381 4811
rect 14415 4808 14427 4811
rect 15562 4808 15568 4820
rect 14415 4780 15568 4808
rect 14415 4777 14427 4780
rect 14369 4771 14427 4777
rect 15562 4768 15568 4780
rect 15620 4768 15626 4820
rect 15657 4811 15715 4817
rect 15657 4777 15669 4811
rect 15703 4777 15715 4811
rect 15657 4771 15715 4777
rect 15841 4811 15899 4817
rect 15841 4777 15853 4811
rect 15887 4808 15899 4811
rect 16850 4808 16856 4820
rect 15887 4780 16856 4808
rect 15887 4777 15899 4780
rect 15841 4771 15899 4777
rect 2685 4743 2743 4749
rect 2685 4709 2697 4743
rect 2731 4740 2743 4743
rect 3234 4740 3240 4752
rect 2731 4712 3240 4740
rect 2731 4709 2743 4712
rect 2685 4703 2743 4709
rect 3234 4700 3240 4712
rect 3292 4700 3298 4752
rect 3418 4700 3424 4752
rect 3476 4740 3482 4752
rect 3476 4712 4568 4740
rect 3476 4700 3482 4712
rect 4246 4672 4252 4684
rect 2148 4644 3280 4672
rect 4207 4644 4252 4672
rect 2038 4564 2044 4616
rect 2096 4604 2102 4616
rect 2148 4613 2176 4644
rect 2133 4607 2191 4613
rect 2133 4604 2145 4607
rect 2096 4576 2145 4604
rect 2096 4564 2102 4576
rect 2133 4573 2145 4576
rect 2179 4573 2191 4607
rect 2133 4567 2191 4573
rect 2501 4607 2559 4613
rect 2501 4573 2513 4607
rect 2547 4604 2559 4607
rect 2774 4604 2780 4616
rect 2547 4576 2780 4604
rect 2547 4573 2559 4576
rect 2501 4567 2559 4573
rect 2774 4564 2780 4576
rect 2832 4564 2838 4616
rect 3252 4613 3280 4644
rect 4246 4632 4252 4644
rect 4304 4632 4310 4684
rect 3237 4607 3295 4613
rect 3237 4573 3249 4607
rect 3283 4573 3295 4607
rect 3237 4567 3295 4573
rect 3421 4607 3479 4613
rect 3421 4573 3433 4607
rect 3467 4604 3479 4607
rect 3602 4604 3608 4616
rect 3467 4576 3608 4604
rect 3467 4573 3479 4576
rect 3421 4567 3479 4573
rect 3602 4564 3608 4576
rect 3660 4564 3666 4616
rect 4062 4564 4068 4616
rect 4120 4604 4126 4616
rect 4341 4607 4399 4613
rect 4341 4604 4353 4607
rect 4120 4576 4353 4604
rect 4120 4564 4126 4576
rect 4341 4573 4353 4576
rect 4387 4573 4399 4607
rect 4540 4604 4568 4712
rect 4706 4700 4712 4752
rect 4764 4740 4770 4752
rect 5350 4740 5356 4752
rect 4764 4712 5356 4740
rect 4764 4700 4770 4712
rect 5350 4700 5356 4712
rect 5408 4700 5414 4752
rect 5534 4700 5540 4752
rect 5592 4740 5598 4752
rect 6086 4740 6092 4752
rect 5592 4712 6092 4740
rect 5592 4700 5598 4712
rect 6086 4700 6092 4712
rect 6144 4740 6150 4752
rect 6144 4712 6776 4740
rect 6144 4700 6150 4712
rect 4617 4675 4675 4681
rect 4617 4641 4629 4675
rect 4663 4672 4675 4675
rect 5813 4675 5871 4681
rect 5813 4672 5825 4675
rect 4663 4644 5825 4672
rect 4663 4641 4675 4644
rect 4617 4635 4675 4641
rect 5813 4641 5825 4644
rect 5859 4641 5871 4675
rect 5813 4635 5871 4641
rect 5166 4604 5172 4616
rect 4540 4576 5028 4604
rect 5127 4576 5172 4604
rect 4341 4567 4399 4573
rect 3329 4539 3387 4545
rect 3329 4505 3341 4539
rect 3375 4536 3387 4539
rect 4522 4536 4528 4548
rect 3375 4508 4528 4536
rect 3375 4505 3387 4508
rect 3329 4499 3387 4505
rect 4522 4496 4528 4508
rect 4580 4496 4586 4548
rect 4614 4496 4620 4548
rect 4672 4536 4678 4548
rect 4709 4539 4767 4545
rect 4709 4536 4721 4539
rect 4672 4508 4721 4536
rect 4672 4496 4678 4508
rect 4709 4505 4721 4508
rect 4755 4505 4767 4539
rect 5000 4536 5028 4576
rect 5166 4564 5172 4576
rect 5224 4564 5230 4616
rect 5537 4607 5595 4613
rect 5537 4573 5549 4607
rect 5583 4573 5595 4607
rect 5537 4567 5595 4573
rect 5629 4607 5687 4613
rect 5629 4573 5641 4607
rect 5675 4604 5687 4607
rect 6546 4604 6552 4616
rect 5675 4576 6552 4604
rect 5675 4573 5687 4576
rect 5629 4567 5687 4573
rect 5552 4536 5580 4567
rect 6546 4564 6552 4576
rect 6604 4564 6610 4616
rect 6748 4613 6776 4712
rect 6914 4700 6920 4752
rect 6972 4740 6978 4752
rect 9858 4740 9864 4752
rect 6972 4712 9864 4740
rect 6972 4700 6978 4712
rect 7024 4613 7052 4712
rect 9858 4700 9864 4712
rect 9916 4700 9922 4752
rect 10042 4700 10048 4752
rect 10100 4740 10106 4752
rect 10321 4743 10379 4749
rect 10321 4740 10333 4743
rect 10100 4712 10333 4740
rect 10100 4700 10106 4712
rect 10321 4709 10333 4712
rect 10367 4740 10379 4743
rect 10594 4740 10600 4752
rect 10367 4712 10600 4740
rect 10367 4709 10379 4712
rect 10321 4703 10379 4709
rect 10594 4700 10600 4712
rect 10652 4700 10658 4752
rect 11054 4700 11060 4752
rect 11112 4740 11118 4752
rect 11112 4712 11284 4740
rect 11112 4700 11118 4712
rect 7190 4632 7196 4684
rect 7248 4672 7254 4684
rect 7929 4675 7987 4681
rect 7929 4672 7941 4675
rect 7248 4644 7941 4672
rect 7248 4632 7254 4644
rect 7929 4641 7941 4644
rect 7975 4672 7987 4675
rect 9585 4675 9643 4681
rect 7975 4644 9536 4672
rect 7975 4641 7987 4644
rect 7929 4635 7987 4641
rect 6733 4607 6791 4613
rect 6733 4573 6745 4607
rect 6779 4573 6791 4607
rect 6733 4567 6791 4573
rect 6917 4607 6975 4613
rect 6917 4573 6929 4607
rect 6963 4573 6975 4607
rect 6917 4567 6975 4573
rect 7009 4607 7067 4613
rect 7009 4573 7021 4607
rect 7055 4573 7067 4607
rect 7009 4567 7067 4573
rect 7101 4607 7159 4613
rect 7101 4573 7113 4607
rect 7147 4604 7159 4607
rect 7466 4604 7472 4616
rect 7147 4576 7472 4604
rect 7147 4573 7159 4576
rect 7101 4567 7159 4573
rect 5000 4508 5580 4536
rect 6932 4536 6960 4567
rect 7466 4564 7472 4576
rect 7524 4564 7530 4616
rect 8110 4564 8116 4616
rect 8168 4604 8174 4616
rect 9140 4613 9168 4644
rect 8205 4607 8263 4613
rect 8205 4604 8217 4607
rect 8168 4576 8217 4604
rect 8168 4564 8174 4576
rect 8205 4573 8217 4576
rect 8251 4573 8263 4607
rect 8205 4567 8263 4573
rect 9125 4607 9183 4613
rect 9125 4573 9137 4607
rect 9171 4573 9183 4607
rect 9125 4567 9183 4573
rect 9217 4607 9275 4613
rect 9217 4573 9229 4607
rect 9263 4604 9275 4607
rect 9306 4604 9312 4616
rect 9263 4576 9312 4604
rect 9263 4573 9275 4576
rect 9217 4567 9275 4573
rect 9306 4564 9312 4576
rect 9364 4564 9370 4616
rect 9401 4607 9459 4613
rect 9401 4573 9413 4607
rect 9447 4573 9459 4607
rect 9508 4604 9536 4644
rect 9585 4641 9597 4675
rect 9631 4672 9643 4675
rect 9631 4644 11179 4672
rect 9631 4641 9643 4644
rect 9585 4635 9643 4641
rect 10045 4607 10103 4613
rect 10045 4604 10057 4607
rect 9508 4576 10057 4604
rect 9401 4567 9459 4573
rect 10045 4573 10057 4576
rect 10091 4604 10103 4607
rect 10226 4604 10232 4616
rect 10091 4576 10232 4604
rect 10091 4573 10103 4576
rect 10045 4567 10103 4573
rect 7190 4536 7196 4548
rect 6932 4508 7196 4536
rect 4709 4499 4767 4505
rect 3234 4428 3240 4480
rect 3292 4468 3298 4480
rect 5258 4468 5264 4480
rect 3292 4440 5264 4468
rect 3292 4428 3298 4440
rect 5258 4428 5264 4440
rect 5316 4428 5322 4480
rect 5350 4428 5356 4480
rect 5408 4468 5414 4480
rect 5552 4468 5580 4508
rect 7190 4496 7196 4508
rect 7248 4496 7254 4548
rect 7282 4496 7288 4548
rect 7340 4536 7346 4548
rect 9416 4536 9444 4567
rect 10226 4564 10232 4576
rect 10284 4564 10290 4616
rect 10870 4604 10876 4616
rect 10831 4576 10876 4604
rect 10870 4564 10876 4576
rect 10928 4564 10934 4616
rect 11151 4610 11179 4644
rect 11256 4613 11284 4712
rect 11882 4700 11888 4752
rect 11940 4740 11946 4752
rect 12437 4743 12495 4749
rect 12437 4740 12449 4743
rect 11940 4712 12449 4740
rect 11940 4700 11946 4712
rect 12437 4709 12449 4712
rect 12483 4709 12495 4743
rect 12437 4703 12495 4709
rect 13541 4743 13599 4749
rect 13541 4709 13553 4743
rect 13587 4709 13599 4743
rect 13541 4703 13599 4709
rect 12066 4632 12072 4684
rect 12124 4672 12130 4684
rect 12345 4675 12403 4681
rect 12345 4672 12357 4675
rect 12124 4644 12357 4672
rect 12124 4632 12130 4644
rect 12345 4641 12357 4644
rect 12391 4641 12403 4675
rect 12345 4635 12403 4641
rect 12710 4632 12716 4684
rect 12768 4672 12774 4684
rect 13265 4675 13323 4681
rect 13265 4672 13277 4675
rect 12768 4644 13277 4672
rect 12768 4632 12774 4644
rect 13265 4641 13277 4644
rect 13311 4641 13323 4675
rect 13265 4635 13323 4641
rect 11036 4604 11094 4610
rect 11036 4570 11048 4604
rect 11082 4570 11094 4604
rect 11036 4564 11094 4570
rect 11136 4604 11194 4610
rect 11136 4570 11148 4604
rect 11182 4570 11194 4604
rect 11136 4564 11194 4570
rect 11241 4607 11299 4613
rect 11241 4573 11253 4607
rect 11287 4573 11299 4607
rect 11241 4567 11299 4573
rect 11882 4564 11888 4616
rect 11940 4604 11946 4616
rect 11977 4607 12035 4613
rect 11977 4604 11989 4607
rect 11940 4576 11989 4604
rect 11940 4564 11946 4576
rect 11977 4573 11989 4576
rect 12023 4573 12035 4607
rect 11977 4567 12035 4573
rect 12161 4607 12219 4613
rect 12161 4573 12173 4607
rect 12207 4573 12219 4607
rect 12161 4567 12219 4573
rect 7340 4508 9444 4536
rect 7340 4496 7346 4508
rect 7834 4468 7840 4480
rect 5408 4440 5453 4468
rect 5552 4440 7840 4468
rect 5408 4428 5414 4440
rect 7834 4428 7840 4440
rect 7892 4428 7898 4480
rect 9416 4468 9444 4508
rect 9490 4496 9496 4548
rect 9548 4536 9554 4548
rect 10137 4539 10195 4545
rect 10137 4536 10149 4539
rect 9548 4508 10149 4536
rect 9548 4496 9554 4508
rect 10137 4505 10149 4508
rect 10183 4505 10195 4539
rect 10318 4536 10324 4548
rect 10279 4508 10324 4536
rect 10137 4499 10195 4505
rect 10318 4496 10324 4508
rect 10376 4496 10382 4548
rect 10502 4496 10508 4548
rect 10560 4536 10566 4548
rect 11051 4536 11079 4564
rect 11151 4536 11179 4564
rect 11330 4536 11336 4548
rect 10560 4508 11100 4536
rect 11151 4508 11336 4536
rect 10560 4496 10566 4508
rect 10336 4468 10364 4496
rect 9416 4440 10364 4468
rect 11072 4468 11100 4508
rect 11330 4496 11336 4508
rect 11388 4496 11394 4548
rect 12176 4536 12204 4567
rect 12250 4564 12256 4616
rect 12308 4604 12314 4616
rect 13173 4607 13231 4613
rect 13173 4604 13185 4607
rect 12308 4576 13185 4604
rect 12308 4564 12314 4576
rect 13173 4573 13185 4576
rect 13219 4573 13231 4607
rect 13173 4567 13231 4573
rect 13556 4536 13584 4703
rect 13814 4632 13820 4684
rect 13872 4672 13878 4684
rect 14507 4675 14565 4681
rect 14507 4672 14519 4675
rect 13872 4644 14519 4672
rect 13872 4632 13878 4644
rect 14507 4641 14519 4644
rect 14553 4641 14565 4675
rect 14918 4672 14924 4684
rect 14831 4644 14924 4672
rect 14507 4635 14565 4641
rect 14918 4632 14924 4644
rect 14976 4672 14982 4684
rect 15672 4672 15700 4771
rect 16850 4768 16856 4780
rect 16908 4768 16914 4820
rect 18233 4811 18291 4817
rect 18233 4777 18245 4811
rect 18279 4808 18291 4811
rect 18322 4808 18328 4820
rect 18279 4780 18328 4808
rect 18279 4777 18291 4780
rect 18233 4771 18291 4777
rect 18322 4768 18328 4780
rect 18380 4808 18386 4820
rect 19521 4811 19579 4817
rect 19521 4808 19533 4811
rect 18380 4780 19533 4808
rect 18380 4768 18386 4780
rect 19521 4777 19533 4780
rect 19567 4808 19579 4811
rect 22094 4808 22100 4820
rect 19567 4780 22100 4808
rect 19567 4777 19579 4780
rect 19521 4771 19579 4777
rect 22094 4768 22100 4780
rect 22152 4768 22158 4820
rect 16390 4740 16396 4752
rect 16351 4712 16396 4740
rect 16390 4700 16396 4712
rect 16448 4740 16454 4752
rect 16945 4743 17003 4749
rect 16945 4740 16957 4743
rect 16448 4712 16957 4740
rect 16448 4700 16454 4712
rect 16945 4709 16957 4712
rect 16991 4740 17003 4743
rect 17126 4740 17132 4752
rect 16991 4712 17132 4740
rect 16991 4709 17003 4712
rect 16945 4703 17003 4709
rect 17126 4700 17132 4712
rect 17184 4700 17190 4752
rect 17681 4743 17739 4749
rect 17681 4709 17693 4743
rect 17727 4740 17739 4743
rect 18506 4740 18512 4752
rect 17727 4712 18512 4740
rect 17727 4709 17739 4712
rect 17681 4703 17739 4709
rect 18506 4700 18512 4712
rect 18564 4700 18570 4752
rect 14976 4644 15700 4672
rect 14976 4632 14982 4644
rect 17586 4632 17592 4684
rect 17644 4672 17650 4684
rect 18693 4675 18751 4681
rect 18693 4672 18705 4675
rect 17644 4644 18705 4672
rect 17644 4632 17650 4644
rect 18693 4641 18705 4644
rect 18739 4641 18751 4675
rect 18693 4635 18751 4641
rect 13906 4564 13912 4616
rect 13964 4604 13970 4616
rect 14645 4607 14703 4613
rect 14645 4604 14657 4607
rect 13964 4576 14657 4604
rect 13964 4564 13970 4576
rect 14645 4573 14657 4576
rect 14691 4573 14703 4607
rect 20346 4604 20352 4616
rect 14645 4567 14703 4573
rect 14936 4576 20352 4604
rect 14936 4536 14964 4576
rect 20346 4564 20352 4576
rect 20404 4564 20410 4616
rect 12176 4508 13584 4536
rect 14568 4508 14964 4536
rect 14568 4480 14596 4508
rect 15010 4496 15016 4548
rect 15068 4536 15074 4548
rect 15068 4508 15113 4536
rect 15068 4496 15074 4508
rect 15194 4496 15200 4548
rect 15252 4536 15258 4548
rect 15473 4539 15531 4545
rect 15473 4536 15485 4539
rect 15252 4508 15485 4536
rect 15252 4496 15258 4508
rect 15473 4505 15485 4508
rect 15519 4536 15531 4539
rect 16482 4536 16488 4548
rect 15519 4508 16488 4536
rect 15519 4505 15531 4508
rect 15473 4499 15531 4505
rect 16482 4496 16488 4508
rect 16540 4496 16546 4548
rect 11882 4468 11888 4480
rect 11072 4440 11888 4468
rect 11882 4428 11888 4440
rect 11940 4428 11946 4480
rect 12713 4471 12771 4477
rect 12713 4437 12725 4471
rect 12759 4468 12771 4471
rect 14550 4468 14556 4480
rect 12759 4440 14556 4468
rect 12759 4437 12771 4440
rect 12713 4431 12771 4437
rect 14550 4428 14556 4440
rect 14608 4428 14614 4480
rect 15028 4468 15056 4496
rect 15673 4471 15731 4477
rect 15673 4468 15685 4471
rect 15028 4440 15685 4468
rect 15673 4437 15685 4440
rect 15719 4437 15731 4471
rect 15673 4431 15731 4437
rect 1104 4378 23987 4400
rect 1104 4326 6630 4378
rect 6682 4326 6694 4378
rect 6746 4326 6758 4378
rect 6810 4326 6822 4378
rect 6874 4326 6886 4378
rect 6938 4326 12311 4378
rect 12363 4326 12375 4378
rect 12427 4326 12439 4378
rect 12491 4326 12503 4378
rect 12555 4326 12567 4378
rect 12619 4326 17992 4378
rect 18044 4326 18056 4378
rect 18108 4326 18120 4378
rect 18172 4326 18184 4378
rect 18236 4326 18248 4378
rect 18300 4326 23673 4378
rect 23725 4326 23737 4378
rect 23789 4326 23801 4378
rect 23853 4326 23865 4378
rect 23917 4326 23929 4378
rect 23981 4326 23987 4378
rect 1104 4304 23987 4326
rect 1670 4264 1676 4276
rect 1631 4236 1676 4264
rect 1670 4224 1676 4236
rect 1728 4264 1734 4276
rect 2133 4267 2191 4273
rect 2133 4264 2145 4267
rect 1728 4236 2145 4264
rect 1728 4224 1734 4236
rect 2133 4233 2145 4236
rect 2179 4233 2191 4267
rect 2133 4227 2191 4233
rect 4062 4224 4068 4276
rect 4120 4264 4126 4276
rect 4249 4267 4307 4273
rect 4249 4264 4261 4267
rect 4120 4236 4261 4264
rect 4120 4224 4126 4236
rect 4249 4233 4261 4236
rect 4295 4233 4307 4267
rect 4249 4227 4307 4233
rect 4341 4267 4399 4273
rect 4341 4233 4353 4267
rect 4387 4264 4399 4267
rect 4706 4264 4712 4276
rect 4387 4236 4712 4264
rect 4387 4233 4399 4236
rect 4341 4227 4399 4233
rect 4706 4224 4712 4236
rect 4764 4224 4770 4276
rect 5258 4224 5264 4276
rect 5316 4264 5322 4276
rect 7190 4264 7196 4276
rect 5316 4236 7098 4264
rect 7151 4236 7196 4264
rect 5316 4224 5322 4236
rect 4985 4199 5043 4205
rect 4985 4196 4997 4199
rect 4264 4168 4997 4196
rect 2038 4088 2044 4140
rect 2096 4128 2102 4140
rect 2685 4131 2743 4137
rect 2685 4128 2697 4131
rect 2096 4100 2697 4128
rect 2096 4088 2102 4100
rect 2685 4097 2697 4100
rect 2731 4097 2743 4131
rect 2866 4128 2872 4140
rect 2827 4100 2872 4128
rect 2685 4091 2743 4097
rect 2866 4088 2872 4100
rect 2924 4088 2930 4140
rect 3329 4131 3387 4137
rect 3329 4097 3341 4131
rect 3375 4128 3387 4131
rect 3418 4128 3424 4140
rect 3375 4100 3424 4128
rect 3375 4097 3387 4100
rect 3329 4091 3387 4097
rect 3418 4088 3424 4100
rect 3476 4088 3482 4140
rect 3513 4131 3571 4137
rect 3513 4097 3525 4131
rect 3559 4128 3571 4131
rect 4264 4128 4292 4168
rect 4985 4165 4997 4168
rect 5031 4196 5043 4199
rect 5166 4196 5172 4208
rect 5031 4168 5172 4196
rect 5031 4165 5043 4168
rect 4985 4159 5043 4165
rect 5166 4156 5172 4168
rect 5224 4156 5230 4208
rect 6917 4199 6975 4205
rect 6917 4196 6929 4199
rect 6564 4168 6929 4196
rect 3559 4100 4292 4128
rect 3559 4097 3571 4100
rect 3513 4091 3571 4097
rect 4338 4088 4344 4140
rect 4396 4128 4402 4140
rect 4433 4131 4491 4137
rect 4433 4128 4445 4131
rect 4396 4100 4445 4128
rect 4396 4088 4402 4100
rect 4433 4097 4445 4100
rect 4479 4128 4491 4131
rect 4890 4128 4896 4140
rect 4479 4100 4896 4128
rect 4479 4097 4491 4100
rect 4433 4091 4491 4097
rect 4890 4088 4896 4100
rect 4948 4088 4954 4140
rect 5074 4128 5080 4140
rect 5035 4100 5080 4128
rect 5074 4088 5080 4100
rect 5132 4088 5138 4140
rect 5721 4131 5779 4137
rect 5721 4097 5733 4131
rect 5767 4128 5779 4131
rect 6564 4128 6592 4168
rect 6917 4165 6929 4168
rect 6963 4165 6975 4199
rect 7070 4196 7098 4236
rect 7190 4224 7196 4236
rect 7248 4224 7254 4276
rect 10410 4224 10416 4276
rect 10468 4264 10474 4276
rect 13005 4267 13063 4273
rect 13005 4264 13017 4267
rect 10468 4236 13017 4264
rect 10468 4224 10474 4236
rect 8478 4196 8484 4208
rect 7070 4168 8484 4196
rect 6917 4159 6975 4165
rect 8478 4156 8484 4168
rect 8536 4156 8542 4208
rect 8956 4168 9260 4196
rect 5767 4100 6592 4128
rect 6707 4131 6765 4137
rect 5767 4097 5779 4100
rect 5721 4091 5779 4097
rect 6707 4097 6719 4131
rect 6753 4128 6765 4131
rect 6753 4097 6776 4128
rect 6707 4091 6776 4097
rect 2777 4063 2835 4069
rect 2777 4029 2789 4063
rect 2823 4060 2835 4063
rect 3973 4063 4031 4069
rect 3973 4060 3985 4063
rect 2823 4032 3985 4060
rect 2823 4029 2835 4032
rect 2777 4023 2835 4029
rect 3973 4029 3985 4032
rect 4019 4060 4031 4063
rect 5736 4060 5764 4091
rect 5994 4060 6000 4072
rect 4019 4032 5764 4060
rect 5955 4032 6000 4060
rect 4019 4029 4031 4032
rect 3973 4023 4031 4029
rect 5994 4020 6000 4032
rect 6052 4020 6058 4072
rect 6546 4060 6552 4072
rect 6507 4032 6552 4060
rect 6546 4020 6552 4032
rect 6604 4020 6610 4072
rect 6748 4060 6776 4091
rect 6822 4088 6828 4140
rect 6880 4128 6886 4140
rect 7009 4131 7067 4137
rect 6880 4100 6925 4128
rect 6880 4088 6886 4100
rect 7009 4097 7021 4131
rect 7055 4128 7067 4131
rect 7653 4131 7711 4137
rect 7653 4128 7665 4131
rect 7055 4100 7665 4128
rect 7055 4097 7067 4100
rect 7009 4091 7067 4097
rect 7653 4097 7665 4100
rect 7699 4097 7711 4131
rect 7834 4128 7840 4140
rect 7795 4100 7840 4128
rect 7653 4091 7711 4097
rect 7834 4088 7840 4100
rect 7892 4088 7898 4140
rect 8021 4131 8079 4137
rect 8021 4097 8033 4131
rect 8067 4097 8079 4131
rect 8021 4091 8079 4097
rect 8113 4131 8171 4137
rect 8113 4097 8125 4131
rect 8159 4097 8171 4131
rect 8113 4091 8171 4097
rect 6914 4060 6920 4072
rect 6748 4032 6920 4060
rect 6914 4020 6920 4032
rect 6972 4020 6978 4072
rect 7098 4020 7104 4072
rect 7156 4060 7162 4072
rect 8036 4060 8064 4091
rect 7156 4032 8064 4060
rect 8128 4060 8156 4091
rect 8202 4088 8208 4140
rect 8260 4128 8266 4140
rect 8956 4128 8984 4168
rect 9122 4128 9128 4140
rect 8260 4100 8984 4128
rect 9083 4100 9128 4128
rect 8260 4088 8266 4100
rect 9122 4088 9128 4100
rect 9180 4088 9186 4140
rect 9232 4128 9260 4168
rect 11330 4156 11336 4208
rect 11388 4196 11394 4208
rect 11388 4168 12020 4196
rect 11388 4156 11394 4168
rect 9401 4131 9459 4137
rect 9401 4128 9413 4131
rect 9232 4100 9413 4128
rect 9401 4097 9413 4100
rect 9447 4097 9459 4131
rect 9950 4128 9956 4140
rect 9911 4100 9956 4128
rect 9401 4091 9459 4097
rect 9950 4088 9956 4100
rect 10008 4088 10014 4140
rect 10137 4131 10195 4137
rect 10137 4097 10149 4131
rect 10183 4097 10195 4131
rect 10137 4091 10195 4097
rect 8294 4060 8300 4072
rect 8128 4032 8300 4060
rect 7156 4020 7162 4032
rect 8294 4020 8300 4032
rect 8352 4060 8358 4072
rect 8570 4060 8576 4072
rect 8352 4032 8576 4060
rect 8352 4020 8358 4032
rect 8570 4020 8576 4032
rect 8628 4020 8634 4072
rect 9214 4020 9220 4072
rect 9272 4060 9278 4072
rect 10152 4060 10180 4091
rect 10870 4088 10876 4140
rect 10928 4128 10934 4140
rect 11514 4128 11520 4140
rect 10928 4100 11520 4128
rect 10928 4088 10934 4100
rect 11514 4088 11520 4100
rect 11572 4128 11578 4140
rect 11701 4131 11759 4137
rect 11701 4128 11713 4131
rect 11572 4100 11713 4128
rect 11572 4088 11578 4100
rect 11701 4097 11713 4100
rect 11747 4097 11759 4131
rect 11882 4128 11888 4140
rect 11843 4100 11888 4128
rect 11701 4091 11759 4097
rect 11882 4088 11888 4100
rect 11940 4088 11946 4140
rect 11992 4137 12020 4168
rect 12084 4137 12112 4236
rect 13005 4233 13017 4236
rect 13051 4233 13063 4267
rect 15194 4264 15200 4276
rect 15155 4236 15200 4264
rect 13005 4227 13063 4233
rect 15194 4224 15200 4236
rect 15252 4224 15258 4276
rect 17126 4264 17132 4276
rect 17087 4236 17132 4264
rect 17126 4224 17132 4236
rect 17184 4264 17190 4276
rect 18877 4267 18935 4273
rect 18877 4264 18889 4267
rect 17184 4236 18889 4264
rect 17184 4224 17190 4236
rect 18877 4233 18889 4236
rect 18923 4233 18935 4267
rect 18877 4227 18935 4233
rect 12434 4156 12440 4208
rect 12492 4196 12498 4208
rect 12805 4199 12863 4205
rect 12805 4196 12817 4199
rect 12492 4168 12817 4196
rect 12492 4156 12498 4168
rect 12805 4165 12817 4168
rect 12851 4165 12863 4199
rect 15933 4199 15991 4205
rect 12805 4159 12863 4165
rect 13464 4168 13860 4196
rect 11977 4131 12035 4137
rect 11977 4097 11989 4131
rect 12023 4097 12035 4131
rect 11977 4091 12035 4097
rect 12069 4131 12127 4137
rect 12069 4097 12081 4131
rect 12115 4097 12127 4131
rect 13464 4128 13492 4168
rect 12069 4091 12127 4097
rect 12176 4100 13492 4128
rect 9272 4032 10180 4060
rect 9272 4020 9278 4032
rect 10226 4020 10232 4072
rect 10284 4060 10290 4072
rect 10505 4063 10563 4069
rect 10505 4060 10517 4063
rect 10284 4032 10517 4060
rect 10284 4020 10290 4032
rect 10505 4029 10517 4032
rect 10551 4060 10563 4063
rect 11238 4060 11244 4072
rect 10551 4032 11244 4060
rect 10551 4029 10563 4032
rect 10505 4023 10563 4029
rect 11238 4020 11244 4032
rect 11296 4020 11302 4072
rect 11422 4020 11428 4072
rect 11480 4060 11486 4072
rect 11790 4060 11796 4072
rect 11480 4032 11796 4060
rect 11480 4020 11486 4032
rect 11790 4020 11796 4032
rect 11848 4060 11854 4072
rect 12176 4060 12204 4100
rect 13538 4088 13544 4140
rect 13596 4128 13602 4140
rect 13725 4131 13783 4137
rect 13725 4128 13737 4131
rect 13596 4100 13737 4128
rect 13596 4088 13602 4100
rect 13725 4097 13737 4100
rect 13771 4097 13783 4131
rect 13832 4128 13860 4168
rect 15933 4165 15945 4199
rect 15979 4196 15991 4199
rect 16666 4196 16672 4208
rect 15979 4168 16672 4196
rect 15979 4165 15991 4168
rect 15933 4159 15991 4165
rect 16666 4156 16672 4168
rect 16724 4156 16730 4208
rect 14369 4131 14427 4137
rect 14369 4128 14381 4131
rect 13832 4100 14381 4128
rect 13725 4091 13783 4097
rect 14369 4097 14381 4100
rect 14415 4128 14427 4131
rect 15289 4131 15347 4137
rect 15289 4128 15301 4131
rect 14415 4100 15301 4128
rect 14415 4097 14427 4100
rect 14369 4091 14427 4097
rect 15289 4097 15301 4100
rect 15335 4128 15347 4131
rect 15746 4128 15752 4140
rect 15335 4100 15752 4128
rect 15335 4097 15347 4100
rect 15289 4091 15347 4097
rect 15746 4088 15752 4100
rect 15804 4088 15810 4140
rect 11848 4032 12204 4060
rect 12345 4063 12403 4069
rect 11848 4020 11854 4032
rect 12345 4029 12357 4063
rect 12391 4060 12403 4063
rect 13630 4060 13636 4072
rect 12391 4032 13636 4060
rect 12391 4029 12403 4032
rect 12345 4023 12403 4029
rect 13630 4020 13636 4032
rect 13688 4020 13694 4072
rect 4154 3952 4160 4004
rect 4212 3992 4218 4004
rect 4706 3992 4712 4004
rect 4212 3964 4712 3992
rect 4212 3952 4218 3964
rect 4706 3952 4712 3964
rect 4764 3952 4770 4004
rect 5537 3995 5595 4001
rect 5537 3961 5549 3995
rect 5583 3992 5595 3995
rect 6086 3992 6092 4004
rect 5583 3964 6092 3992
rect 5583 3961 5595 3964
rect 5537 3955 5595 3961
rect 6086 3952 6092 3964
rect 6144 3952 6150 4004
rect 10134 3952 10140 4004
rect 10192 3992 10198 4004
rect 10318 3992 10324 4004
rect 10192 3964 10324 3992
rect 10192 3952 10198 3964
rect 10318 3952 10324 3964
rect 10376 3992 10382 4004
rect 10873 3995 10931 4001
rect 10873 3992 10885 3995
rect 10376 3964 10885 3992
rect 10376 3952 10382 3964
rect 10873 3961 10885 3964
rect 10919 3992 10931 3995
rect 12158 3992 12164 4004
rect 10919 3964 12164 3992
rect 10919 3961 10931 3964
rect 10873 3955 10931 3961
rect 12158 3952 12164 3964
rect 12216 3952 12222 4004
rect 13173 3995 13231 4001
rect 13173 3961 13185 3995
rect 13219 3992 13231 3995
rect 13446 3992 13452 4004
rect 13219 3964 13452 3992
rect 13219 3961 13231 3964
rect 13173 3955 13231 3961
rect 13446 3952 13452 3964
rect 13504 3952 13510 4004
rect 3421 3927 3479 3933
rect 3421 3893 3433 3927
rect 3467 3924 3479 3927
rect 5626 3924 5632 3936
rect 3467 3896 5632 3924
rect 3467 3893 3479 3896
rect 3421 3887 3479 3893
rect 5626 3884 5632 3896
rect 5684 3924 5690 3936
rect 5905 3927 5963 3933
rect 5905 3924 5917 3927
rect 5684 3896 5917 3924
rect 5684 3884 5690 3896
rect 5905 3893 5917 3896
rect 5951 3924 5963 3927
rect 7466 3924 7472 3936
rect 5951 3896 7472 3924
rect 5951 3893 5963 3896
rect 5905 3887 5963 3893
rect 7466 3884 7472 3896
rect 7524 3884 7530 3936
rect 11330 3884 11336 3936
rect 11388 3924 11394 3936
rect 11514 3924 11520 3936
rect 11388 3896 11520 3924
rect 11388 3884 11394 3896
rect 11514 3884 11520 3896
rect 11572 3924 11578 3936
rect 12250 3924 12256 3936
rect 11572 3896 12256 3924
rect 11572 3884 11578 3896
rect 12250 3884 12256 3896
rect 12308 3924 12314 3936
rect 12989 3927 13047 3933
rect 12989 3924 13001 3927
rect 12308 3896 13001 3924
rect 12308 3884 12314 3896
rect 12989 3893 13001 3896
rect 13035 3893 13047 3927
rect 12989 3887 13047 3893
rect 1104 3834 23828 3856
rect 1104 3782 3790 3834
rect 3842 3782 3854 3834
rect 3906 3782 3918 3834
rect 3970 3782 3982 3834
rect 4034 3782 4046 3834
rect 4098 3782 9471 3834
rect 9523 3782 9535 3834
rect 9587 3782 9599 3834
rect 9651 3782 9663 3834
rect 9715 3782 9727 3834
rect 9779 3782 15152 3834
rect 15204 3782 15216 3834
rect 15268 3782 15280 3834
rect 15332 3782 15344 3834
rect 15396 3782 15408 3834
rect 15460 3782 20833 3834
rect 20885 3782 20897 3834
rect 20949 3782 20961 3834
rect 21013 3782 21025 3834
rect 21077 3782 21089 3834
rect 21141 3782 23828 3834
rect 1104 3760 23828 3782
rect 4154 3720 4160 3732
rect 1964 3692 4160 3720
rect 1964 3525 1992 3692
rect 4154 3680 4160 3692
rect 4212 3680 4218 3732
rect 4246 3680 4252 3732
rect 4304 3720 4310 3732
rect 4433 3723 4491 3729
rect 4433 3720 4445 3723
rect 4304 3692 4445 3720
rect 4304 3680 4310 3692
rect 4433 3689 4445 3692
rect 4479 3689 4491 3723
rect 4433 3683 4491 3689
rect 4522 3680 4528 3732
rect 4580 3720 4586 3732
rect 4580 3692 4625 3720
rect 4580 3680 4586 3692
rect 4706 3680 4712 3732
rect 4764 3720 4770 3732
rect 6362 3720 6368 3732
rect 4764 3692 6368 3720
rect 4764 3680 4770 3692
rect 6362 3680 6368 3692
rect 6420 3680 6426 3732
rect 6454 3680 6460 3732
rect 6512 3720 6518 3732
rect 6641 3723 6699 3729
rect 6641 3720 6653 3723
rect 6512 3692 6653 3720
rect 6512 3680 6518 3692
rect 6641 3689 6653 3692
rect 6687 3689 6699 3723
rect 6641 3683 6699 3689
rect 8481 3723 8539 3729
rect 8481 3689 8493 3723
rect 8527 3720 8539 3723
rect 8754 3720 8760 3732
rect 8527 3692 8760 3720
rect 8527 3689 8539 3692
rect 8481 3683 8539 3689
rect 8754 3680 8760 3692
rect 8812 3680 8818 3732
rect 9769 3723 9827 3729
rect 9769 3689 9781 3723
rect 9815 3720 9827 3723
rect 10870 3720 10876 3732
rect 9815 3692 10876 3720
rect 9815 3689 9827 3692
rect 9769 3683 9827 3689
rect 10870 3680 10876 3692
rect 10928 3680 10934 3732
rect 11054 3680 11060 3732
rect 11112 3720 11118 3732
rect 11241 3723 11299 3729
rect 11241 3720 11253 3723
rect 11112 3692 11253 3720
rect 11112 3680 11118 3692
rect 11241 3689 11253 3692
rect 11287 3720 11299 3723
rect 11790 3720 11796 3732
rect 11287 3692 11796 3720
rect 11287 3689 11299 3692
rect 11241 3683 11299 3689
rect 11790 3680 11796 3692
rect 11848 3680 11854 3732
rect 11882 3680 11888 3732
rect 11940 3720 11946 3732
rect 12342 3720 12348 3732
rect 11940 3692 12348 3720
rect 11940 3680 11946 3692
rect 12342 3680 12348 3692
rect 12400 3680 12406 3732
rect 12437 3723 12495 3729
rect 12437 3689 12449 3723
rect 12483 3720 12495 3723
rect 12710 3720 12716 3732
rect 12483 3692 12716 3720
rect 12483 3689 12495 3692
rect 12437 3683 12495 3689
rect 12710 3680 12716 3692
rect 12768 3680 12774 3732
rect 12989 3723 13047 3729
rect 12989 3689 13001 3723
rect 13035 3720 13047 3723
rect 13538 3720 13544 3732
rect 13035 3692 13544 3720
rect 13035 3689 13047 3692
rect 12989 3683 13047 3689
rect 13538 3680 13544 3692
rect 13596 3720 13602 3732
rect 16025 3723 16083 3729
rect 16025 3720 16037 3723
rect 13596 3692 16037 3720
rect 13596 3680 13602 3692
rect 16025 3689 16037 3692
rect 16071 3689 16083 3723
rect 16025 3683 16083 3689
rect 16666 3680 16672 3732
rect 16724 3720 16730 3732
rect 16761 3723 16819 3729
rect 16761 3720 16773 3723
rect 16724 3692 16773 3720
rect 16724 3680 16730 3692
rect 16761 3689 16773 3692
rect 16807 3689 16819 3723
rect 16761 3683 16819 3689
rect 2133 3655 2191 3661
rect 2133 3621 2145 3655
rect 2179 3652 2191 3655
rect 4341 3655 4399 3661
rect 4341 3652 4353 3655
rect 2179 3624 4353 3652
rect 2179 3621 2191 3624
rect 2133 3615 2191 3621
rect 4341 3621 4353 3624
rect 4387 3621 4399 3655
rect 4341 3615 4399 3621
rect 4890 3612 4896 3664
rect 4948 3652 4954 3664
rect 4948 3624 4993 3652
rect 4948 3612 4954 3624
rect 5350 3612 5356 3664
rect 5408 3652 5414 3664
rect 7101 3655 7159 3661
rect 7101 3652 7113 3655
rect 5408 3624 5948 3652
rect 5408 3612 5414 3624
rect 3142 3584 3148 3596
rect 2608 3556 3148 3584
rect 2608 3525 2636 3556
rect 3142 3544 3148 3556
rect 3200 3544 3206 3596
rect 1949 3519 2007 3525
rect 1949 3485 1961 3519
rect 1995 3485 2007 3519
rect 1949 3479 2007 3485
rect 2133 3519 2191 3525
rect 2133 3485 2145 3519
rect 2179 3485 2191 3519
rect 2133 3479 2191 3485
rect 2593 3519 2651 3525
rect 2593 3485 2605 3519
rect 2639 3485 2651 3519
rect 2593 3479 2651 3485
rect 2777 3519 2835 3525
rect 2777 3485 2789 3519
rect 2823 3516 2835 3519
rect 3418 3516 3424 3528
rect 2823 3488 3280 3516
rect 3379 3488 3424 3516
rect 2823 3485 2835 3488
rect 2777 3479 2835 3485
rect 2148 3448 2176 3479
rect 2866 3448 2872 3460
rect 2148 3420 2872 3448
rect 2866 3408 2872 3420
rect 2924 3408 2930 3460
rect 3252 3448 3280 3488
rect 3418 3476 3424 3488
rect 3476 3476 3482 3528
rect 4157 3519 4215 3525
rect 4157 3485 4169 3519
rect 4203 3516 4215 3519
rect 4430 3516 4436 3528
rect 4203 3488 4436 3516
rect 4203 3485 4215 3488
rect 4157 3479 4215 3485
rect 4430 3476 4436 3488
rect 4488 3476 4494 3528
rect 4614 3516 4620 3528
rect 4575 3488 4620 3516
rect 4614 3476 4620 3488
rect 4672 3476 4678 3528
rect 5537 3519 5595 3525
rect 5537 3485 5549 3519
rect 5583 3485 5595 3519
rect 5920 3516 5948 3624
rect 6012 3624 7113 3652
rect 6012 3593 6040 3624
rect 7101 3621 7113 3624
rect 7147 3621 7159 3655
rect 7101 3615 7159 3621
rect 7742 3612 7748 3664
rect 7800 3652 7806 3664
rect 10318 3652 10324 3664
rect 7800 3624 10324 3652
rect 7800 3612 7806 3624
rect 10318 3612 10324 3624
rect 10376 3612 10382 3664
rect 10781 3655 10839 3661
rect 10781 3621 10793 3655
rect 10827 3652 10839 3655
rect 15010 3652 15016 3664
rect 10827 3624 15016 3652
rect 10827 3621 10839 3624
rect 10781 3615 10839 3621
rect 15010 3612 15016 3624
rect 15068 3612 15074 3664
rect 5997 3587 6055 3593
rect 5997 3553 6009 3587
rect 6043 3553 6055 3587
rect 5997 3547 6055 3553
rect 6086 3544 6092 3596
rect 6144 3584 6150 3596
rect 6822 3584 6828 3596
rect 6144 3556 6189 3584
rect 6380 3556 6828 3584
rect 6144 3544 6150 3556
rect 6380 3525 6408 3556
rect 6822 3544 6828 3556
rect 6880 3584 6886 3596
rect 8846 3584 8852 3596
rect 6880 3556 8852 3584
rect 6880 3544 6886 3556
rect 7484 3528 7512 3556
rect 8846 3544 8852 3556
rect 8904 3544 8910 3596
rect 9214 3544 9220 3596
rect 9272 3584 9278 3596
rect 9493 3587 9551 3593
rect 9493 3584 9505 3587
rect 9272 3556 9505 3584
rect 9272 3544 9278 3556
rect 9493 3553 9505 3556
rect 9539 3553 9551 3587
rect 9493 3547 9551 3553
rect 9585 3587 9643 3593
rect 9585 3553 9597 3587
rect 9631 3584 9643 3587
rect 10134 3584 10140 3596
rect 9631 3556 10140 3584
rect 9631 3553 9643 3556
rect 9585 3547 9643 3553
rect 10134 3544 10140 3556
rect 10192 3544 10198 3596
rect 10686 3584 10692 3596
rect 10336 3556 10692 3584
rect 6365 3519 6423 3525
rect 6365 3516 6377 3519
rect 5920 3488 6377 3516
rect 5537 3479 5595 3485
rect 6365 3485 6377 3488
rect 6411 3485 6423 3519
rect 6365 3479 6423 3485
rect 5552 3448 5580 3479
rect 6454 3476 6460 3528
rect 6512 3516 6518 3528
rect 7098 3516 7104 3528
rect 6512 3488 7104 3516
rect 6512 3476 6518 3488
rect 7098 3476 7104 3488
rect 7156 3476 7162 3528
rect 7282 3516 7288 3528
rect 7243 3488 7288 3516
rect 7282 3476 7288 3488
rect 7340 3476 7346 3528
rect 7466 3476 7472 3528
rect 7524 3516 7530 3528
rect 7653 3519 7711 3525
rect 7524 3488 7617 3516
rect 7524 3476 7530 3488
rect 7653 3485 7665 3519
rect 7699 3516 7711 3519
rect 7834 3516 7840 3528
rect 7699 3488 7840 3516
rect 7699 3485 7711 3488
rect 7653 3479 7711 3485
rect 7834 3476 7840 3488
rect 7892 3516 7898 3528
rect 8113 3519 8171 3525
rect 8113 3516 8125 3519
rect 7892 3488 8125 3516
rect 7892 3476 7898 3488
rect 8113 3485 8125 3488
rect 8159 3485 8171 3519
rect 8113 3479 8171 3485
rect 8202 3476 8208 3528
rect 8260 3516 8266 3528
rect 9122 3516 9128 3528
rect 8260 3488 8432 3516
rect 9083 3488 9128 3516
rect 8260 3476 8266 3488
rect 7377 3451 7435 3457
rect 3252 3420 4660 3448
rect 5552 3420 5764 3448
rect 2682 3380 2688 3392
rect 2643 3352 2688 3380
rect 2682 3340 2688 3352
rect 2740 3340 2746 3392
rect 3234 3380 3240 3392
rect 3195 3352 3240 3380
rect 3234 3340 3240 3352
rect 3292 3340 3298 3392
rect 4632 3380 4660 3420
rect 5534 3380 5540 3392
rect 4632 3352 5540 3380
rect 5534 3340 5540 3352
rect 5592 3340 5598 3392
rect 5736 3380 5764 3420
rect 7377 3417 7389 3451
rect 7423 3448 7435 3451
rect 7742 3448 7748 3460
rect 7423 3420 7748 3448
rect 7423 3417 7435 3420
rect 7377 3411 7435 3417
rect 7742 3408 7748 3420
rect 7800 3408 7806 3460
rect 8294 3448 8300 3460
rect 8255 3420 8300 3448
rect 8294 3408 8300 3420
rect 8352 3408 8358 3460
rect 8404 3448 8432 3488
rect 9122 3476 9128 3488
rect 9180 3476 9186 3528
rect 10226 3516 10232 3528
rect 10187 3488 10232 3516
rect 10226 3476 10232 3488
rect 10284 3476 10290 3528
rect 10336 3525 10364 3556
rect 10686 3544 10692 3556
rect 10744 3544 10750 3596
rect 11606 3544 11612 3596
rect 11664 3584 11670 3596
rect 12069 3587 12127 3593
rect 12069 3584 12081 3587
rect 11664 3556 12081 3584
rect 11664 3544 11670 3556
rect 12069 3553 12081 3556
rect 12115 3553 12127 3587
rect 12250 3584 12256 3596
rect 12211 3556 12256 3584
rect 12069 3547 12127 3553
rect 10321 3519 10379 3525
rect 10321 3485 10333 3519
rect 10367 3485 10379 3519
rect 10321 3479 10379 3485
rect 10505 3519 10563 3525
rect 10505 3485 10517 3519
rect 10551 3485 10563 3519
rect 10505 3479 10563 3485
rect 9217 3451 9275 3457
rect 9217 3448 9229 3451
rect 8404 3420 9229 3448
rect 9217 3417 9229 3420
rect 9263 3417 9275 3451
rect 9950 3448 9956 3460
rect 9217 3411 9275 3417
rect 9416 3420 9956 3448
rect 8570 3380 8576 3392
rect 5736 3352 8576 3380
rect 8570 3340 8576 3352
rect 8628 3340 8634 3392
rect 9416 3389 9444 3420
rect 9950 3408 9956 3420
rect 10008 3408 10014 3460
rect 10520 3448 10548 3479
rect 10594 3476 10600 3528
rect 10652 3516 10658 3528
rect 11241 3519 11299 3525
rect 10652 3488 10697 3516
rect 10652 3476 10658 3488
rect 11241 3485 11253 3519
rect 11287 3485 11299 3519
rect 11422 3516 11428 3528
rect 11383 3488 11428 3516
rect 11241 3479 11299 3485
rect 11256 3448 11284 3479
rect 11422 3476 11428 3488
rect 11480 3476 11486 3528
rect 11514 3476 11520 3528
rect 11572 3516 11578 3528
rect 11882 3516 11888 3528
rect 11572 3488 11888 3516
rect 11572 3476 11578 3488
rect 11882 3476 11888 3488
rect 11940 3516 11946 3528
rect 11977 3519 12035 3525
rect 11977 3516 11989 3519
rect 11940 3488 11989 3516
rect 11940 3476 11946 3488
rect 11977 3485 11989 3488
rect 12023 3485 12035 3519
rect 11977 3479 12035 3485
rect 12084 3448 12112 3547
rect 12250 3544 12256 3556
rect 12308 3544 12314 3596
rect 12161 3519 12219 3525
rect 12161 3485 12173 3519
rect 12207 3516 12219 3519
rect 12342 3516 12348 3528
rect 12207 3488 12348 3516
rect 12207 3485 12219 3488
rect 12161 3479 12219 3485
rect 12342 3476 12348 3488
rect 12400 3476 12406 3528
rect 13541 3519 13599 3525
rect 13541 3485 13553 3519
rect 13587 3516 13599 3519
rect 13906 3516 13912 3528
rect 13587 3488 13912 3516
rect 13587 3485 13599 3488
rect 13541 3479 13599 3485
rect 13906 3476 13912 3488
rect 13964 3516 13970 3528
rect 15013 3519 15071 3525
rect 15013 3516 15025 3519
rect 13964 3488 15025 3516
rect 13964 3476 13970 3488
rect 15013 3485 15025 3488
rect 15059 3516 15071 3519
rect 15746 3516 15752 3528
rect 15059 3488 15752 3516
rect 15059 3485 15071 3488
rect 15013 3479 15071 3485
rect 15746 3476 15752 3488
rect 15804 3476 15810 3528
rect 23293 3519 23351 3525
rect 23293 3485 23305 3519
rect 23339 3516 23351 3519
rect 23382 3516 23388 3528
rect 23339 3488 23388 3516
rect 23339 3485 23351 3488
rect 23293 3479 23351 3485
rect 23382 3476 23388 3488
rect 23440 3476 23446 3528
rect 14277 3451 14335 3457
rect 14277 3448 14289 3451
rect 10520 3420 12020 3448
rect 12084 3420 14289 3448
rect 11992 3392 12020 3420
rect 14277 3417 14289 3420
rect 14323 3448 14335 3451
rect 14366 3448 14372 3460
rect 14323 3420 14372 3448
rect 14323 3417 14335 3420
rect 14277 3411 14335 3417
rect 14366 3408 14372 3420
rect 14424 3448 14430 3460
rect 15473 3451 15531 3457
rect 15473 3448 15485 3451
rect 14424 3420 15485 3448
rect 14424 3408 14430 3420
rect 15473 3417 15485 3420
rect 15519 3417 15531 3451
rect 17954 3448 17960 3460
rect 17915 3420 17960 3448
rect 15473 3411 15531 3417
rect 17954 3408 17960 3420
rect 18012 3408 18018 3460
rect 9401 3383 9459 3389
rect 9401 3349 9413 3383
rect 9447 3349 9459 3383
rect 9401 3343 9459 3349
rect 11974 3340 11980 3392
rect 12032 3340 12038 3392
rect 17310 3380 17316 3392
rect 17271 3352 17316 3380
rect 17310 3340 17316 3352
rect 17368 3340 17374 3392
rect 1104 3290 23987 3312
rect 1104 3238 6630 3290
rect 6682 3238 6694 3290
rect 6746 3238 6758 3290
rect 6810 3238 6822 3290
rect 6874 3238 6886 3290
rect 6938 3238 12311 3290
rect 12363 3238 12375 3290
rect 12427 3238 12439 3290
rect 12491 3238 12503 3290
rect 12555 3238 12567 3290
rect 12619 3238 17992 3290
rect 18044 3238 18056 3290
rect 18108 3238 18120 3290
rect 18172 3238 18184 3290
rect 18236 3238 18248 3290
rect 18300 3238 23673 3290
rect 23725 3238 23737 3290
rect 23789 3238 23801 3290
rect 23853 3238 23865 3290
rect 23917 3238 23929 3290
rect 23981 3238 23987 3290
rect 1104 3216 23987 3238
rect 1670 3176 1676 3188
rect 1631 3148 1676 3176
rect 1670 3136 1676 3148
rect 1728 3136 1734 3188
rect 4890 3136 4896 3188
rect 4948 3176 4954 3188
rect 7101 3179 7159 3185
rect 7101 3176 7113 3179
rect 4948 3148 7113 3176
rect 4948 3136 4954 3148
rect 7101 3145 7113 3148
rect 7147 3145 7159 3179
rect 7101 3139 7159 3145
rect 7374 3136 7380 3188
rect 7432 3176 7438 3188
rect 7745 3179 7803 3185
rect 7745 3176 7757 3179
rect 7432 3148 7757 3176
rect 7432 3136 7438 3148
rect 7745 3145 7757 3148
rect 7791 3145 7803 3179
rect 7745 3139 7803 3145
rect 8205 3179 8263 3185
rect 8205 3145 8217 3179
rect 8251 3176 8263 3179
rect 9122 3176 9128 3188
rect 8251 3148 9128 3176
rect 8251 3145 8263 3148
rect 8205 3139 8263 3145
rect 9122 3136 9128 3148
rect 9180 3136 9186 3188
rect 11057 3179 11115 3185
rect 11057 3145 11069 3179
rect 11103 3176 11115 3179
rect 11514 3176 11520 3188
rect 11103 3148 11520 3176
rect 11103 3145 11115 3148
rect 11057 3139 11115 3145
rect 11514 3136 11520 3148
rect 11572 3136 11578 3188
rect 11790 3136 11796 3188
rect 11848 3176 11854 3188
rect 11901 3179 11959 3185
rect 11901 3176 11913 3179
rect 11848 3148 11913 3176
rect 11848 3136 11854 3148
rect 11901 3145 11913 3148
rect 11947 3145 11959 3179
rect 12066 3176 12072 3188
rect 12027 3148 12072 3176
rect 11901 3139 11959 3145
rect 12066 3136 12072 3148
rect 12124 3136 12130 3188
rect 13906 3176 13912 3188
rect 13867 3148 13912 3176
rect 13906 3136 13912 3148
rect 13964 3136 13970 3188
rect 14366 3176 14372 3188
rect 14327 3148 14372 3176
rect 14366 3136 14372 3148
rect 14424 3136 14430 3188
rect 17402 3176 17408 3188
rect 17363 3148 17408 3176
rect 17402 3136 17408 3148
rect 17460 3136 17466 3188
rect 7926 3108 7932 3120
rect 4816 3080 7932 3108
rect 2498 3040 2504 3052
rect 2459 3012 2504 3040
rect 2498 3000 2504 3012
rect 2556 3000 2562 3052
rect 4816 3049 4844 3080
rect 7926 3068 7932 3080
rect 7984 3068 7990 3120
rect 8478 3068 8484 3120
rect 8536 3108 8542 3120
rect 8573 3111 8631 3117
rect 8573 3108 8585 3111
rect 8536 3080 8585 3108
rect 8536 3068 8542 3080
rect 8573 3077 8585 3080
rect 8619 3108 8631 3111
rect 8938 3108 8944 3120
rect 8619 3080 8944 3108
rect 8619 3077 8631 3080
rect 8573 3071 8631 3077
rect 8938 3068 8944 3080
rect 8996 3068 9002 3120
rect 9214 3068 9220 3120
rect 9272 3108 9278 3120
rect 10410 3108 10416 3120
rect 9272 3080 9674 3108
rect 10371 3080 10416 3108
rect 9272 3068 9278 3080
rect 4801 3043 4859 3049
rect 4801 3009 4813 3043
rect 4847 3009 4859 3043
rect 4801 3003 4859 3009
rect 5537 3043 5595 3049
rect 5537 3009 5549 3043
rect 5583 3040 5595 3043
rect 5626 3040 5632 3052
rect 5583 3012 5632 3040
rect 5583 3009 5595 3012
rect 5537 3003 5595 3009
rect 5626 3000 5632 3012
rect 5684 3000 5690 3052
rect 5721 3043 5779 3049
rect 5721 3009 5733 3043
rect 5767 3040 5779 3043
rect 5902 3040 5908 3052
rect 5767 3012 5908 3040
rect 5767 3009 5779 3012
rect 5721 3003 5779 3009
rect 5902 3000 5908 3012
rect 5960 3000 5966 3052
rect 7282 3040 7288 3052
rect 6472 3012 7288 3040
rect 4157 2975 4215 2981
rect 4157 2941 4169 2975
rect 4203 2972 4215 2975
rect 6472 2972 6500 3012
rect 7282 3000 7288 3012
rect 7340 3000 7346 3052
rect 8294 3000 8300 3052
rect 8352 3040 8358 3052
rect 8389 3043 8447 3049
rect 8389 3040 8401 3043
rect 8352 3012 8401 3040
rect 8352 3000 8358 3012
rect 8389 3009 8401 3012
rect 8435 3009 8447 3043
rect 8389 3003 8447 3009
rect 8665 3043 8723 3049
rect 8665 3009 8677 3043
rect 8711 3009 8723 3043
rect 8665 3003 8723 3009
rect 7374 2972 7380 2984
rect 4203 2944 6500 2972
rect 6564 2944 7380 2972
rect 4203 2941 4215 2944
rect 4157 2935 4215 2941
rect 3513 2907 3571 2913
rect 3513 2873 3525 2907
rect 3559 2904 3571 2907
rect 6454 2904 6460 2916
rect 3559 2876 6460 2904
rect 3559 2873 3571 2876
rect 3513 2867 3571 2873
rect 6454 2864 6460 2876
rect 6512 2864 6518 2916
rect 2130 2796 2136 2848
rect 2188 2836 2194 2848
rect 2317 2839 2375 2845
rect 2317 2836 2329 2839
rect 2188 2808 2329 2836
rect 2188 2796 2194 2808
rect 2317 2805 2329 2808
rect 2363 2805 2375 2839
rect 2317 2799 2375 2805
rect 4522 2796 4528 2848
rect 4580 2836 4586 2848
rect 5261 2839 5319 2845
rect 5261 2836 5273 2839
rect 4580 2808 5273 2836
rect 4580 2796 4586 2808
rect 5261 2805 5273 2808
rect 5307 2805 5319 2839
rect 5261 2799 5319 2805
rect 5537 2839 5595 2845
rect 5537 2805 5549 2839
rect 5583 2836 5595 2839
rect 6564 2836 6592 2944
rect 7374 2932 7380 2944
rect 7432 2972 7438 2984
rect 7469 2975 7527 2981
rect 7469 2972 7481 2975
rect 7432 2944 7481 2972
rect 7432 2932 7438 2944
rect 7469 2941 7481 2944
rect 7515 2941 7527 2975
rect 7469 2935 7527 2941
rect 7561 2975 7619 2981
rect 7561 2941 7573 2975
rect 7607 2972 7619 2975
rect 8478 2972 8484 2984
rect 7607 2944 8484 2972
rect 7607 2941 7619 2944
rect 7561 2935 7619 2941
rect 8478 2932 8484 2944
rect 8536 2932 8542 2984
rect 8680 2972 8708 3003
rect 8846 3000 8852 3052
rect 8904 3040 8910 3052
rect 9125 3043 9183 3049
rect 9125 3040 9137 3043
rect 8904 3012 9137 3040
rect 8904 3000 8910 3012
rect 9125 3009 9137 3012
rect 9171 3009 9183 3043
rect 9306 3040 9312 3052
rect 9267 3012 9312 3040
rect 9125 3003 9183 3009
rect 9306 3000 9312 3012
rect 9364 3000 9370 3052
rect 9493 2975 9551 2981
rect 9493 2972 9505 2975
rect 8680 2944 9505 2972
rect 9493 2941 9505 2944
rect 9539 2941 9551 2975
rect 9646 2972 9674 3080
rect 10410 3068 10416 3080
rect 10468 3068 10474 3120
rect 11698 3108 11704 3120
rect 11659 3080 11704 3108
rect 11698 3068 11704 3080
rect 11756 3068 11762 3120
rect 12158 3068 12164 3120
rect 12216 3108 12222 3120
rect 14921 3111 14979 3117
rect 14921 3108 14933 3111
rect 12216 3080 14933 3108
rect 12216 3068 12222 3080
rect 14921 3077 14933 3080
rect 14967 3077 14979 3111
rect 14921 3071 14979 3077
rect 10957 3052 11015 3055
rect 10318 3040 10324 3052
rect 10279 3012 10324 3040
rect 10318 3000 10324 3012
rect 10376 3000 10382 3052
rect 10505 3043 10563 3049
rect 10505 3009 10517 3043
rect 10551 3040 10563 3043
rect 10957 3040 10968 3052
rect 10551 3012 10968 3040
rect 10551 3009 10563 3012
rect 10957 3009 10968 3012
rect 10505 3003 10563 3009
rect 10962 3000 10968 3009
rect 11020 3000 11026 3052
rect 9646 2944 13216 2972
rect 9493 2935 9551 2941
rect 6638 2864 6644 2916
rect 6696 2904 6702 2916
rect 6696 2876 6741 2904
rect 6696 2864 6702 2876
rect 9858 2864 9864 2916
rect 9916 2904 9922 2916
rect 13188 2913 13216 2944
rect 12529 2907 12587 2913
rect 12529 2904 12541 2907
rect 9916 2876 12541 2904
rect 9916 2864 9922 2876
rect 12529 2873 12541 2876
rect 12575 2873 12587 2907
rect 12529 2867 12587 2873
rect 13173 2907 13231 2913
rect 13173 2873 13185 2907
rect 13219 2873 13231 2907
rect 13173 2867 13231 2873
rect 5583 2808 6592 2836
rect 5583 2805 5595 2808
rect 5537 2799 5595 2805
rect 11330 2796 11336 2848
rect 11388 2836 11394 2848
rect 11885 2839 11943 2845
rect 11885 2836 11897 2839
rect 11388 2808 11897 2836
rect 11388 2796 11394 2808
rect 11885 2805 11897 2808
rect 11931 2805 11943 2839
rect 11885 2799 11943 2805
rect 15654 2796 15660 2848
rect 15712 2836 15718 2848
rect 15749 2839 15807 2845
rect 15749 2836 15761 2839
rect 15712 2808 15761 2836
rect 15712 2796 15718 2808
rect 15749 2805 15761 2808
rect 15795 2805 15807 2839
rect 16850 2836 16856 2848
rect 16811 2808 16856 2836
rect 15749 2799 15807 2805
rect 16850 2796 16856 2808
rect 16908 2796 16914 2848
rect 18322 2836 18328 2848
rect 18283 2808 18328 2836
rect 18322 2796 18328 2808
rect 18380 2796 18386 2848
rect 20714 2796 20720 2848
rect 20772 2836 20778 2848
rect 20901 2839 20959 2845
rect 20901 2836 20913 2839
rect 20772 2808 20913 2836
rect 20772 2796 20778 2808
rect 20901 2805 20913 2808
rect 20947 2805 20959 2839
rect 20901 2799 20959 2805
rect 22738 2796 22744 2848
rect 22796 2836 22802 2848
rect 22833 2839 22891 2845
rect 22833 2836 22845 2839
rect 22796 2808 22845 2836
rect 22796 2796 22802 2808
rect 22833 2805 22845 2808
rect 22879 2805 22891 2839
rect 22833 2799 22891 2805
rect 1104 2746 23828 2768
rect 1104 2694 3790 2746
rect 3842 2694 3854 2746
rect 3906 2694 3918 2746
rect 3970 2694 3982 2746
rect 4034 2694 4046 2746
rect 4098 2694 9471 2746
rect 9523 2694 9535 2746
rect 9587 2694 9599 2746
rect 9651 2694 9663 2746
rect 9715 2694 9727 2746
rect 9779 2694 15152 2746
rect 15204 2694 15216 2746
rect 15268 2694 15280 2746
rect 15332 2694 15344 2746
rect 15396 2694 15408 2746
rect 15460 2694 20833 2746
rect 20885 2694 20897 2746
rect 20949 2694 20961 2746
rect 21013 2694 21025 2746
rect 21077 2694 21089 2746
rect 21141 2694 23828 2746
rect 1104 2672 23828 2694
rect 7834 2632 7840 2644
rect 7795 2604 7840 2632
rect 7834 2592 7840 2604
rect 7892 2592 7898 2644
rect 8478 2592 8484 2644
rect 8536 2632 8542 2644
rect 9125 2635 9183 2641
rect 9125 2632 9137 2635
rect 8536 2604 9137 2632
rect 8536 2592 8542 2604
rect 9125 2601 9137 2604
rect 9171 2601 9183 2635
rect 11793 2635 11851 2641
rect 9125 2595 9183 2601
rect 9232 2604 11284 2632
rect 5074 2564 5080 2576
rect 4987 2536 5080 2564
rect 1854 2428 1860 2440
rect 1815 2400 1860 2428
rect 1854 2388 1860 2400
rect 1912 2388 1918 2440
rect 2685 2431 2743 2437
rect 2685 2397 2697 2431
rect 2731 2428 2743 2431
rect 3234 2428 3240 2440
rect 2731 2400 3240 2428
rect 2731 2397 2743 2400
rect 2685 2391 2743 2397
rect 3234 2388 3240 2400
rect 3292 2388 3298 2440
rect 3418 2428 3424 2440
rect 3379 2400 3424 2428
rect 3418 2388 3424 2400
rect 3476 2388 3482 2440
rect 4246 2428 4252 2440
rect 4207 2400 4252 2428
rect 4246 2388 4252 2400
rect 4304 2388 4310 2440
rect 5000 2437 5028 2536
rect 5074 2524 5080 2536
rect 5132 2564 5138 2576
rect 9232 2564 9260 2604
rect 5132 2536 9260 2564
rect 10505 2567 10563 2573
rect 5132 2524 5138 2536
rect 10505 2533 10517 2567
rect 10551 2564 10563 2567
rect 11146 2564 11152 2576
rect 10551 2536 11152 2564
rect 10551 2533 10563 2536
rect 10505 2527 10563 2533
rect 11146 2524 11152 2536
rect 11204 2524 11210 2576
rect 11256 2564 11284 2604
rect 11793 2601 11805 2635
rect 11839 2632 11851 2635
rect 11974 2632 11980 2644
rect 11839 2604 11980 2632
rect 11839 2601 11851 2604
rect 11793 2595 11851 2601
rect 11974 2592 11980 2604
rect 12032 2592 12038 2644
rect 16850 2632 16856 2644
rect 12406 2604 16856 2632
rect 12406 2564 12434 2604
rect 16850 2592 16856 2604
rect 16908 2592 16914 2644
rect 17310 2564 17316 2576
rect 11256 2536 12434 2564
rect 16224 2536 17316 2564
rect 8294 2496 8300 2508
rect 5736 2468 8300 2496
rect 5736 2437 5764 2468
rect 8294 2456 8300 2468
rect 8352 2456 8358 2508
rect 8938 2456 8944 2508
rect 8996 2496 9002 2508
rect 9493 2499 9551 2505
rect 9493 2496 9505 2499
rect 8996 2468 9505 2496
rect 8996 2456 9002 2468
rect 9493 2465 9505 2468
rect 9539 2465 9551 2499
rect 9493 2459 9551 2465
rect 4985 2431 5043 2437
rect 4985 2397 4997 2431
rect 5031 2397 5043 2431
rect 4985 2391 5043 2397
rect 5721 2431 5779 2437
rect 5721 2397 5733 2431
rect 5767 2397 5779 2431
rect 5721 2391 5779 2397
rect 5810 2388 5816 2440
rect 5868 2428 5874 2440
rect 6825 2431 6883 2437
rect 6825 2428 6837 2431
rect 5868 2400 6837 2428
rect 5868 2388 5874 2400
rect 6825 2397 6837 2400
rect 6871 2397 6883 2431
rect 7374 2428 7380 2440
rect 7335 2400 7380 2428
rect 6825 2391 6883 2397
rect 1486 2252 1492 2304
rect 1544 2292 1550 2304
rect 1673 2295 1731 2301
rect 1673 2292 1685 2295
rect 1544 2264 1685 2292
rect 1544 2252 1550 2264
rect 1673 2261 1685 2264
rect 1719 2261 1731 2295
rect 1673 2255 1731 2261
rect 2501 2295 2559 2301
rect 2501 2261 2513 2295
rect 2547 2292 2559 2295
rect 2774 2292 2780 2304
rect 2547 2264 2780 2292
rect 2547 2261 2559 2264
rect 2501 2255 2559 2261
rect 2774 2252 2780 2264
rect 2832 2252 2838 2304
rect 3237 2295 3295 2301
rect 3237 2261 3249 2295
rect 3283 2292 3295 2295
rect 3418 2292 3424 2304
rect 3283 2264 3424 2292
rect 3283 2261 3295 2264
rect 3237 2255 3295 2261
rect 3418 2252 3424 2264
rect 3476 2252 3482 2304
rect 4062 2292 4068 2304
rect 4023 2264 4068 2292
rect 4062 2252 4068 2264
rect 4120 2252 4126 2304
rect 4706 2252 4712 2304
rect 4764 2292 4770 2304
rect 4801 2295 4859 2301
rect 4801 2292 4813 2295
rect 4764 2264 4813 2292
rect 4764 2252 4770 2264
rect 4801 2261 4813 2264
rect 4847 2261 4859 2295
rect 4801 2255 4859 2261
rect 5350 2252 5356 2304
rect 5408 2292 5414 2304
rect 5537 2295 5595 2301
rect 5537 2292 5549 2295
rect 5408 2264 5549 2292
rect 5408 2252 5414 2264
rect 5537 2261 5549 2264
rect 5583 2261 5595 2295
rect 5537 2255 5595 2261
rect 5994 2252 6000 2304
rect 6052 2292 6058 2304
rect 6641 2295 6699 2301
rect 6641 2292 6653 2295
rect 6052 2264 6653 2292
rect 6052 2252 6058 2264
rect 6641 2261 6653 2264
rect 6687 2261 6699 2295
rect 6840 2292 6868 2391
rect 7374 2388 7380 2400
rect 7432 2388 7438 2440
rect 7466 2388 7472 2440
rect 7524 2428 7530 2440
rect 7650 2428 7656 2440
rect 7524 2400 7569 2428
rect 7611 2400 7656 2428
rect 7524 2388 7530 2400
rect 7650 2388 7656 2400
rect 7708 2388 7714 2440
rect 8573 2431 8631 2437
rect 8573 2397 8585 2431
rect 8619 2397 8631 2431
rect 8573 2391 8631 2397
rect 8588 2360 8616 2391
rect 9030 2388 9036 2440
rect 9088 2428 9094 2440
rect 9309 2431 9367 2437
rect 9309 2428 9321 2431
rect 9088 2400 9321 2428
rect 9088 2388 9094 2400
rect 9309 2397 9321 2400
rect 9355 2397 9367 2431
rect 9309 2391 9367 2397
rect 11149 2431 11207 2437
rect 11149 2397 11161 2431
rect 11195 2397 11207 2431
rect 11149 2391 11207 2397
rect 10502 2360 10508 2372
rect 8588 2332 10508 2360
rect 10502 2320 10508 2332
rect 10560 2320 10566 2372
rect 11164 2360 11192 2391
rect 11606 2388 11612 2440
rect 11664 2428 11670 2440
rect 11701 2431 11759 2437
rect 11701 2428 11713 2431
rect 11664 2400 11713 2428
rect 11664 2388 11670 2400
rect 11701 2397 11713 2400
rect 11747 2397 11759 2431
rect 11882 2428 11888 2440
rect 11843 2400 11888 2428
rect 11701 2391 11759 2397
rect 11882 2388 11888 2400
rect 11940 2388 11946 2440
rect 12529 2431 12587 2437
rect 12529 2397 12541 2431
rect 12575 2428 12587 2431
rect 12710 2428 12716 2440
rect 12575 2400 12716 2428
rect 12575 2397 12587 2400
rect 12529 2391 12587 2397
rect 12710 2388 12716 2400
rect 12768 2388 12774 2440
rect 13078 2388 13084 2440
rect 13136 2428 13142 2440
rect 13173 2431 13231 2437
rect 13173 2428 13185 2431
rect 13136 2400 13185 2428
rect 13136 2388 13142 2400
rect 13173 2397 13185 2400
rect 13219 2397 13231 2431
rect 13173 2391 13231 2397
rect 13722 2388 13728 2440
rect 13780 2428 13786 2440
rect 14277 2431 14335 2437
rect 14277 2428 14289 2431
rect 13780 2400 14289 2428
rect 13780 2388 13786 2400
rect 14277 2397 14289 2400
rect 14323 2397 14335 2431
rect 14277 2391 14335 2397
rect 14366 2388 14372 2440
rect 14424 2428 14430 2440
rect 14921 2431 14979 2437
rect 14921 2428 14933 2431
rect 14424 2400 14933 2428
rect 14424 2388 14430 2400
rect 14921 2397 14933 2400
rect 14967 2397 14979 2431
rect 14921 2391 14979 2397
rect 15010 2388 15016 2440
rect 15068 2428 15074 2440
rect 15565 2431 15623 2437
rect 15565 2428 15577 2431
rect 15068 2400 15577 2428
rect 15068 2388 15074 2400
rect 15565 2397 15577 2400
rect 15611 2397 15623 2431
rect 15565 2391 15623 2397
rect 11790 2360 11796 2372
rect 11164 2332 11796 2360
rect 11790 2320 11796 2332
rect 11848 2320 11854 2372
rect 16224 2369 16252 2536
rect 17310 2524 17316 2536
rect 17368 2524 17374 2576
rect 16298 2388 16304 2440
rect 16356 2428 16362 2440
rect 16853 2431 16911 2437
rect 16853 2428 16865 2431
rect 16356 2400 16865 2428
rect 16356 2388 16362 2400
rect 16853 2397 16865 2400
rect 16899 2397 16911 2431
rect 16853 2391 16911 2397
rect 16942 2388 16948 2440
rect 17000 2428 17006 2440
rect 17497 2431 17555 2437
rect 17497 2428 17509 2431
rect 17000 2400 17509 2428
rect 17000 2388 17006 2400
rect 17497 2397 17509 2400
rect 17543 2397 17555 2431
rect 17497 2391 17555 2397
rect 17586 2388 17592 2440
rect 17644 2428 17650 2440
rect 18141 2431 18199 2437
rect 18141 2428 18153 2431
rect 17644 2400 18153 2428
rect 17644 2388 17650 2400
rect 18141 2397 18153 2400
rect 18187 2397 18199 2431
rect 18141 2391 18199 2397
rect 18874 2388 18880 2440
rect 18932 2428 18938 2440
rect 19429 2431 19487 2437
rect 19429 2428 19441 2431
rect 18932 2400 19441 2428
rect 18932 2388 18938 2400
rect 19429 2397 19441 2400
rect 19475 2397 19487 2431
rect 19429 2391 19487 2397
rect 19518 2388 19524 2440
rect 19576 2428 19582 2440
rect 20073 2431 20131 2437
rect 20073 2428 20085 2431
rect 19576 2400 20085 2428
rect 19576 2388 19582 2400
rect 20073 2397 20085 2400
rect 20119 2397 20131 2431
rect 20073 2391 20131 2397
rect 20162 2388 20168 2440
rect 20220 2428 20226 2440
rect 20717 2431 20775 2437
rect 20717 2428 20729 2431
rect 20220 2400 20729 2428
rect 20220 2388 20226 2400
rect 20717 2397 20729 2400
rect 20763 2397 20775 2431
rect 20717 2391 20775 2397
rect 21450 2388 21456 2440
rect 21508 2428 21514 2440
rect 22005 2431 22063 2437
rect 22005 2428 22017 2431
rect 21508 2400 22017 2428
rect 21508 2388 21514 2400
rect 22005 2397 22017 2400
rect 22051 2397 22063 2431
rect 22005 2391 22063 2397
rect 22094 2388 22100 2440
rect 22152 2428 22158 2440
rect 22649 2431 22707 2437
rect 22649 2428 22661 2431
rect 22152 2400 22661 2428
rect 22152 2388 22158 2400
rect 22649 2397 22661 2400
rect 22695 2397 22707 2431
rect 22649 2391 22707 2397
rect 16209 2363 16267 2369
rect 16209 2360 16221 2363
rect 12406 2332 16221 2360
rect 12406 2292 12434 2332
rect 16209 2329 16221 2332
rect 16255 2329 16267 2363
rect 16209 2323 16267 2329
rect 16390 2320 16396 2372
rect 16448 2360 16454 2372
rect 18785 2363 18843 2369
rect 18785 2360 18797 2363
rect 16448 2332 18797 2360
rect 16448 2320 16454 2332
rect 18785 2329 18797 2332
rect 18831 2329 18843 2363
rect 18785 2323 18843 2329
rect 6840 2264 12434 2292
rect 6641 2255 6699 2261
rect 1104 2202 23987 2224
rect 1104 2150 6630 2202
rect 6682 2150 6694 2202
rect 6746 2150 6758 2202
rect 6810 2150 6822 2202
rect 6874 2150 6886 2202
rect 6938 2150 12311 2202
rect 12363 2150 12375 2202
rect 12427 2150 12439 2202
rect 12491 2150 12503 2202
rect 12555 2150 12567 2202
rect 12619 2150 17992 2202
rect 18044 2150 18056 2202
rect 18108 2150 18120 2202
rect 18172 2150 18184 2202
rect 18236 2150 18248 2202
rect 18300 2150 23673 2202
rect 23725 2150 23737 2202
rect 23789 2150 23801 2202
rect 23853 2150 23865 2202
rect 23917 2150 23929 2202
rect 23981 2150 23987 2202
rect 1104 2128 23987 2150
rect 8202 2048 8208 2100
rect 8260 2088 8266 2100
rect 16390 2088 16396 2100
rect 8260 2060 16396 2088
rect 8260 2048 8266 2060
rect 16390 2048 16396 2060
rect 16448 2048 16454 2100
<< via1 >>
rect 3790 22278 3842 22330
rect 3854 22278 3906 22330
rect 3918 22278 3970 22330
rect 3982 22278 4034 22330
rect 4046 22278 4098 22330
rect 9471 22278 9523 22330
rect 9535 22278 9587 22330
rect 9599 22278 9651 22330
rect 9663 22278 9715 22330
rect 9727 22278 9779 22330
rect 15152 22278 15204 22330
rect 15216 22278 15268 22330
rect 15280 22278 15332 22330
rect 15344 22278 15396 22330
rect 15408 22278 15460 22330
rect 20833 22278 20885 22330
rect 20897 22278 20949 22330
rect 20961 22278 21013 22330
rect 21025 22278 21077 22330
rect 21089 22278 21141 22330
rect 9772 22015 9824 22024
rect 9772 21981 9781 22015
rect 9781 21981 9815 22015
rect 9815 21981 9824 22015
rect 9772 21972 9824 21981
rect 12440 21972 12492 22024
rect 13084 22015 13136 22024
rect 7472 21904 7524 21956
rect 10140 21904 10192 21956
rect 11336 21904 11388 21956
rect 7564 21836 7616 21888
rect 11428 21836 11480 21888
rect 13084 21981 13093 22015
rect 13093 21981 13127 22015
rect 13127 21981 13136 22015
rect 13084 21972 13136 21981
rect 17408 21972 17460 22024
rect 22376 21972 22428 22024
rect 14372 21904 14424 21956
rect 13544 21836 13596 21888
rect 13728 21879 13780 21888
rect 13728 21845 13737 21879
rect 13737 21845 13771 21879
rect 13771 21845 13780 21879
rect 14556 21904 14608 21956
rect 14648 21879 14700 21888
rect 13728 21836 13780 21845
rect 14648 21845 14657 21879
rect 14657 21845 14691 21879
rect 14691 21845 14700 21879
rect 14648 21836 14700 21845
rect 17500 21879 17552 21888
rect 17500 21845 17509 21879
rect 17509 21845 17543 21879
rect 17543 21845 17552 21879
rect 17500 21836 17552 21845
rect 6630 21734 6682 21786
rect 6694 21734 6746 21786
rect 6758 21734 6810 21786
rect 6822 21734 6874 21786
rect 6886 21734 6938 21786
rect 12311 21734 12363 21786
rect 12375 21734 12427 21786
rect 12439 21734 12491 21786
rect 12503 21734 12555 21786
rect 12567 21734 12619 21786
rect 17992 21734 18044 21786
rect 18056 21734 18108 21786
rect 18120 21734 18172 21786
rect 18184 21734 18236 21786
rect 18248 21734 18300 21786
rect 23673 21734 23725 21786
rect 23737 21734 23789 21786
rect 23801 21734 23853 21786
rect 23865 21734 23917 21786
rect 23929 21734 23981 21786
rect 9312 21496 9364 21548
rect 11244 21496 11296 21548
rect 14648 21539 14700 21548
rect 14648 21505 14657 21539
rect 14657 21505 14691 21539
rect 14691 21505 14700 21539
rect 14648 21496 14700 21505
rect 9772 21471 9824 21480
rect 9772 21437 9781 21471
rect 9781 21437 9815 21471
rect 9815 21437 9824 21471
rect 9772 21428 9824 21437
rect 13084 21471 13136 21480
rect 13084 21437 13093 21471
rect 13093 21437 13127 21471
rect 13127 21437 13136 21471
rect 13084 21428 13136 21437
rect 14188 21471 14240 21480
rect 11060 21360 11112 21412
rect 7104 21292 7156 21344
rect 11520 21292 11572 21344
rect 11796 21292 11848 21344
rect 13360 21360 13412 21412
rect 14188 21437 14197 21471
rect 14197 21437 14231 21471
rect 14231 21437 14240 21471
rect 14188 21428 14240 21437
rect 17500 21360 17552 21412
rect 13452 21292 13504 21344
rect 3790 21190 3842 21242
rect 3854 21190 3906 21242
rect 3918 21190 3970 21242
rect 3982 21190 4034 21242
rect 4046 21190 4098 21242
rect 9471 21190 9523 21242
rect 9535 21190 9587 21242
rect 9599 21190 9651 21242
rect 9663 21190 9715 21242
rect 9727 21190 9779 21242
rect 15152 21190 15204 21242
rect 15216 21190 15268 21242
rect 15280 21190 15332 21242
rect 15344 21190 15396 21242
rect 15408 21190 15460 21242
rect 20833 21190 20885 21242
rect 20897 21190 20949 21242
rect 20961 21190 21013 21242
rect 21025 21190 21077 21242
rect 21089 21190 21141 21242
rect 2504 21088 2556 21140
rect 7104 21088 7156 21140
rect 9864 21088 9916 21140
rect 11152 21088 11204 21140
rect 11796 21088 11848 21140
rect 9312 21020 9364 21072
rect 13452 20995 13504 21004
rect 13452 20961 13461 20995
rect 13461 20961 13495 20995
rect 13495 20961 13504 20995
rect 13452 20952 13504 20961
rect 5540 20884 5592 20936
rect 13360 20927 13412 20936
rect 13360 20893 13369 20927
rect 13369 20893 13403 20927
rect 13403 20893 13412 20927
rect 13360 20884 13412 20893
rect 6184 20816 6236 20868
rect 7656 20816 7708 20868
rect 8944 20816 8996 20868
rect 4896 20791 4948 20800
rect 4896 20757 4905 20791
rect 4905 20757 4939 20791
rect 4939 20757 4948 20791
rect 4896 20748 4948 20757
rect 8116 20791 8168 20800
rect 8116 20757 8125 20791
rect 8125 20757 8159 20791
rect 8159 20757 8168 20791
rect 8116 20748 8168 20757
rect 6630 20646 6682 20698
rect 6694 20646 6746 20698
rect 6758 20646 6810 20698
rect 6822 20646 6874 20698
rect 6886 20646 6938 20698
rect 12311 20646 12363 20698
rect 12375 20646 12427 20698
rect 12439 20646 12491 20698
rect 12503 20646 12555 20698
rect 12567 20646 12619 20698
rect 17992 20646 18044 20698
rect 18056 20646 18108 20698
rect 18120 20646 18172 20698
rect 18184 20646 18236 20698
rect 18248 20646 18300 20698
rect 23673 20646 23725 20698
rect 23737 20646 23789 20698
rect 23801 20646 23853 20698
rect 23865 20646 23917 20698
rect 23929 20646 23981 20698
rect 14188 20544 14240 20596
rect 12716 20476 12768 20528
rect 4896 20408 4948 20460
rect 5540 20408 5592 20460
rect 7288 20408 7340 20460
rect 11152 20451 11204 20460
rect 11152 20417 11161 20451
rect 11161 20417 11195 20451
rect 11195 20417 11204 20451
rect 11152 20408 11204 20417
rect 14372 20476 14424 20528
rect 13728 20408 13780 20460
rect 4436 20204 4488 20256
rect 8116 20204 8168 20256
rect 10416 20204 10468 20256
rect 11244 20204 11296 20256
rect 3790 20102 3842 20154
rect 3854 20102 3906 20154
rect 3918 20102 3970 20154
rect 3982 20102 4034 20154
rect 4046 20102 4098 20154
rect 9471 20102 9523 20154
rect 9535 20102 9587 20154
rect 9599 20102 9651 20154
rect 9663 20102 9715 20154
rect 9727 20102 9779 20154
rect 15152 20102 15204 20154
rect 15216 20102 15268 20154
rect 15280 20102 15332 20154
rect 15344 20102 15396 20154
rect 15408 20102 15460 20154
rect 20833 20102 20885 20154
rect 20897 20102 20949 20154
rect 20961 20102 21013 20154
rect 21025 20102 21077 20154
rect 21089 20102 21141 20154
rect 11152 19907 11204 19916
rect 11152 19873 11161 19907
rect 11161 19873 11195 19907
rect 11195 19873 11204 19907
rect 11152 19864 11204 19873
rect 5540 19796 5592 19848
rect 8300 19796 8352 19848
rect 11704 19796 11756 19848
rect 4252 19771 4304 19780
rect 4252 19737 4286 19771
rect 4286 19737 4304 19771
rect 4252 19728 4304 19737
rect 2136 19660 2188 19712
rect 6368 19660 6420 19712
rect 8208 19660 8260 19712
rect 10784 19660 10836 19712
rect 18328 19728 18380 19780
rect 10968 19660 11020 19712
rect 11612 19703 11664 19712
rect 11612 19669 11621 19703
rect 11621 19669 11655 19703
rect 11655 19669 11664 19703
rect 11612 19660 11664 19669
rect 6630 19558 6682 19610
rect 6694 19558 6746 19610
rect 6758 19558 6810 19610
rect 6822 19558 6874 19610
rect 6886 19558 6938 19610
rect 12311 19558 12363 19610
rect 12375 19558 12427 19610
rect 12439 19558 12491 19610
rect 12503 19558 12555 19610
rect 12567 19558 12619 19610
rect 17992 19558 18044 19610
rect 18056 19558 18108 19610
rect 18120 19558 18172 19610
rect 18184 19558 18236 19610
rect 18248 19558 18300 19610
rect 23673 19558 23725 19610
rect 23737 19558 23789 19610
rect 23801 19558 23853 19610
rect 23865 19558 23917 19610
rect 23929 19558 23981 19610
rect 3700 19499 3752 19508
rect 3700 19465 3709 19499
rect 3709 19465 3743 19499
rect 3743 19465 3752 19499
rect 3700 19456 3752 19465
rect 7104 19499 7156 19508
rect 7104 19465 7113 19499
rect 7113 19465 7147 19499
rect 7147 19465 7156 19499
rect 7104 19456 7156 19465
rect 5908 19388 5960 19440
rect 5540 19320 5592 19372
rect 8944 19159 8996 19168
rect 8944 19125 8953 19159
rect 8953 19125 8987 19159
rect 8987 19125 8996 19159
rect 8944 19116 8996 19125
rect 3790 19014 3842 19066
rect 3854 19014 3906 19066
rect 3918 19014 3970 19066
rect 3982 19014 4034 19066
rect 4046 19014 4098 19066
rect 9471 19014 9523 19066
rect 9535 19014 9587 19066
rect 9599 19014 9651 19066
rect 9663 19014 9715 19066
rect 9727 19014 9779 19066
rect 15152 19014 15204 19066
rect 15216 19014 15268 19066
rect 15280 19014 15332 19066
rect 15344 19014 15396 19066
rect 15408 19014 15460 19066
rect 20833 19014 20885 19066
rect 20897 19014 20949 19066
rect 20961 19014 21013 19066
rect 21025 19014 21077 19066
rect 21089 19014 21141 19066
rect 4252 18912 4304 18964
rect 18328 18912 18380 18964
rect 2320 18751 2372 18760
rect 2320 18717 2329 18751
rect 2329 18717 2363 18751
rect 2363 18717 2372 18751
rect 2320 18708 2372 18717
rect 5540 18708 5592 18760
rect 11704 18819 11756 18828
rect 11704 18785 11713 18819
rect 11713 18785 11747 18819
rect 11747 18785 11756 18819
rect 11704 18776 11756 18785
rect 8300 18708 8352 18760
rect 8392 18708 8444 18760
rect 18420 18751 18472 18760
rect 6092 18683 6144 18692
rect 6092 18649 6110 18683
rect 6110 18649 6144 18683
rect 6092 18640 6144 18649
rect 5080 18572 5132 18624
rect 8024 18572 8076 18624
rect 11704 18572 11756 18624
rect 18420 18717 18429 18751
rect 18429 18717 18463 18751
rect 18463 18717 18472 18751
rect 18420 18708 18472 18717
rect 13452 18572 13504 18624
rect 6630 18470 6682 18522
rect 6694 18470 6746 18522
rect 6758 18470 6810 18522
rect 6822 18470 6874 18522
rect 6886 18470 6938 18522
rect 12311 18470 12363 18522
rect 12375 18470 12427 18522
rect 12439 18470 12491 18522
rect 12503 18470 12555 18522
rect 12567 18470 12619 18522
rect 17992 18470 18044 18522
rect 18056 18470 18108 18522
rect 18120 18470 18172 18522
rect 18184 18470 18236 18522
rect 18248 18470 18300 18522
rect 23673 18470 23725 18522
rect 23737 18470 23789 18522
rect 23801 18470 23853 18522
rect 23865 18470 23917 18522
rect 23929 18470 23981 18522
rect 4344 18232 4396 18284
rect 7380 18275 7432 18284
rect 7380 18241 7414 18275
rect 7414 18241 7432 18275
rect 7380 18232 7432 18241
rect 8300 18232 8352 18284
rect 9312 18232 9364 18284
rect 12072 18232 12124 18284
rect 7104 18207 7156 18216
rect 3516 18071 3568 18080
rect 3516 18037 3525 18071
rect 3525 18037 3559 18071
rect 3559 18037 3568 18071
rect 3516 18028 3568 18037
rect 4620 18028 4672 18080
rect 7104 18173 7113 18207
rect 7113 18173 7147 18207
rect 7147 18173 7156 18207
rect 7104 18164 7156 18173
rect 11888 18096 11940 18148
rect 9128 18028 9180 18080
rect 11796 18071 11848 18080
rect 11796 18037 11805 18071
rect 11805 18037 11839 18071
rect 11839 18037 11848 18071
rect 11796 18028 11848 18037
rect 3790 17926 3842 17978
rect 3854 17926 3906 17978
rect 3918 17926 3970 17978
rect 3982 17926 4034 17978
rect 4046 17926 4098 17978
rect 9471 17926 9523 17978
rect 9535 17926 9587 17978
rect 9599 17926 9651 17978
rect 9663 17926 9715 17978
rect 9727 17926 9779 17978
rect 15152 17926 15204 17978
rect 15216 17926 15268 17978
rect 15280 17926 15332 17978
rect 15344 17926 15396 17978
rect 15408 17926 15460 17978
rect 20833 17926 20885 17978
rect 20897 17926 20949 17978
rect 20961 17926 21013 17978
rect 21025 17926 21077 17978
rect 21089 17926 21141 17978
rect 5540 17867 5592 17876
rect 5540 17833 5549 17867
rect 5549 17833 5583 17867
rect 5583 17833 5592 17867
rect 5540 17824 5592 17833
rect 8116 17824 8168 17876
rect 4620 17620 4672 17672
rect 7472 17663 7524 17672
rect 7472 17629 7481 17663
rect 7481 17629 7515 17663
rect 7515 17629 7524 17663
rect 7472 17620 7524 17629
rect 9312 17620 9364 17672
rect 11152 17620 11204 17672
rect 2504 17552 2556 17604
rect 7012 17595 7064 17604
rect 7012 17561 7021 17595
rect 7021 17561 7055 17595
rect 7055 17561 7064 17595
rect 7012 17552 7064 17561
rect 11796 17552 11848 17604
rect 12992 17552 13044 17604
rect 3424 17527 3476 17536
rect 3424 17493 3433 17527
rect 3433 17493 3467 17527
rect 3467 17493 3476 17527
rect 3424 17484 3476 17493
rect 6000 17484 6052 17536
rect 10876 17484 10928 17536
rect 16028 17484 16080 17536
rect 6630 17382 6682 17434
rect 6694 17382 6746 17434
rect 6758 17382 6810 17434
rect 6822 17382 6874 17434
rect 6886 17382 6938 17434
rect 12311 17382 12363 17434
rect 12375 17382 12427 17434
rect 12439 17382 12491 17434
rect 12503 17382 12555 17434
rect 12567 17382 12619 17434
rect 17992 17382 18044 17434
rect 18056 17382 18108 17434
rect 18120 17382 18172 17434
rect 18184 17382 18236 17434
rect 18248 17382 18300 17434
rect 23673 17382 23725 17434
rect 23737 17382 23789 17434
rect 23801 17382 23853 17434
rect 23865 17382 23917 17434
rect 23929 17382 23981 17434
rect 11796 17280 11848 17332
rect 14004 17280 14056 17332
rect 3240 17187 3292 17196
rect 4620 17212 4672 17264
rect 3240 17153 3258 17187
rect 3258 17153 3292 17187
rect 3240 17144 3292 17153
rect 4252 17187 4304 17196
rect 4252 17153 4286 17187
rect 4286 17153 4304 17187
rect 4252 17144 4304 17153
rect 7104 17144 7156 17196
rect 7748 17144 7800 17196
rect 9312 17144 9364 17196
rect 11796 17144 11848 17196
rect 13084 17008 13136 17060
rect 2228 16940 2280 16992
rect 5356 16983 5408 16992
rect 5356 16949 5365 16983
rect 5365 16949 5399 16983
rect 5399 16949 5408 16983
rect 5356 16940 5408 16949
rect 8484 16940 8536 16992
rect 11796 16983 11848 16992
rect 11796 16949 11805 16983
rect 11805 16949 11839 16983
rect 11839 16949 11848 16983
rect 11796 16940 11848 16949
rect 3790 16838 3842 16890
rect 3854 16838 3906 16890
rect 3918 16838 3970 16890
rect 3982 16838 4034 16890
rect 4046 16838 4098 16890
rect 9471 16838 9523 16890
rect 9535 16838 9587 16890
rect 9599 16838 9651 16890
rect 9663 16838 9715 16890
rect 9727 16838 9779 16890
rect 15152 16838 15204 16890
rect 15216 16838 15268 16890
rect 15280 16838 15332 16890
rect 15344 16838 15396 16890
rect 15408 16838 15460 16890
rect 20833 16838 20885 16890
rect 20897 16838 20949 16890
rect 20961 16838 21013 16890
rect 21025 16838 21077 16890
rect 21089 16838 21141 16890
rect 2504 16779 2556 16788
rect 2504 16745 2513 16779
rect 2513 16745 2547 16779
rect 2547 16745 2556 16779
rect 2504 16736 2556 16745
rect 2228 16668 2280 16720
rect 5540 16736 5592 16788
rect 4620 16643 4672 16652
rect 4620 16609 4629 16643
rect 4629 16609 4663 16643
rect 4663 16609 4672 16643
rect 4620 16600 4672 16609
rect 8300 16643 8352 16652
rect 8300 16609 8309 16643
rect 8309 16609 8343 16643
rect 8343 16609 8352 16643
rect 8300 16600 8352 16609
rect 9312 16600 9364 16652
rect 2504 16532 2556 16584
rect 3056 16532 3108 16584
rect 3516 16532 3568 16584
rect 16580 16532 16632 16584
rect 3700 16464 3752 16516
rect 4712 16396 4764 16448
rect 7472 16464 7524 16516
rect 7932 16464 7984 16516
rect 7840 16396 7892 16448
rect 9312 16396 9364 16448
rect 11980 16396 12032 16448
rect 6630 16294 6682 16346
rect 6694 16294 6746 16346
rect 6758 16294 6810 16346
rect 6822 16294 6874 16346
rect 6886 16294 6938 16346
rect 12311 16294 12363 16346
rect 12375 16294 12427 16346
rect 12439 16294 12491 16346
rect 12503 16294 12555 16346
rect 12567 16294 12619 16346
rect 17992 16294 18044 16346
rect 18056 16294 18108 16346
rect 18120 16294 18172 16346
rect 18184 16294 18236 16346
rect 18248 16294 18300 16346
rect 23673 16294 23725 16346
rect 23737 16294 23789 16346
rect 23801 16294 23853 16346
rect 23865 16294 23917 16346
rect 23929 16294 23981 16346
rect 2320 16192 2372 16244
rect 4620 16192 4672 16244
rect 5908 16235 5960 16244
rect 5908 16201 5917 16235
rect 5917 16201 5951 16235
rect 5951 16201 5960 16235
rect 5908 16192 5960 16201
rect 7012 16192 7064 16244
rect 8300 16235 8352 16244
rect 8300 16201 8309 16235
rect 8309 16201 8343 16235
rect 8343 16201 8352 16235
rect 8300 16192 8352 16201
rect 8944 16124 8996 16176
rect 1584 16056 1636 16108
rect 3700 16056 3752 16108
rect 4160 15988 4212 16040
rect 2964 15920 3016 15972
rect 5172 16099 5224 16108
rect 5172 16065 5181 16099
rect 5181 16065 5215 16099
rect 5215 16065 5224 16099
rect 5172 16056 5224 16065
rect 5724 16056 5776 16108
rect 6000 16099 6052 16108
rect 6000 16065 6009 16099
rect 6009 16065 6043 16099
rect 6043 16065 6052 16099
rect 6000 16056 6052 16065
rect 7104 16099 7156 16108
rect 7104 16065 7113 16099
rect 7113 16065 7147 16099
rect 7147 16065 7156 16099
rect 7380 16099 7432 16108
rect 7104 16056 7156 16065
rect 7380 16065 7389 16099
rect 7389 16065 7423 16099
rect 7423 16065 7432 16099
rect 7380 16056 7432 16065
rect 8116 16056 8168 16108
rect 12808 16056 12860 16108
rect 7196 15988 7248 16040
rect 11060 15988 11112 16040
rect 5816 15920 5868 15972
rect 7564 15920 7616 15972
rect 4804 15895 4856 15904
rect 4804 15861 4813 15895
rect 4813 15861 4847 15895
rect 4847 15861 4856 15895
rect 4804 15852 4856 15861
rect 6552 15852 6604 15904
rect 9312 15852 9364 15904
rect 11060 15895 11112 15904
rect 11060 15861 11069 15895
rect 11069 15861 11103 15895
rect 11103 15861 11112 15895
rect 11060 15852 11112 15861
rect 11796 15852 11848 15904
rect 14188 15895 14240 15904
rect 14188 15861 14197 15895
rect 14197 15861 14231 15895
rect 14231 15861 14240 15895
rect 14188 15852 14240 15861
rect 3790 15750 3842 15802
rect 3854 15750 3906 15802
rect 3918 15750 3970 15802
rect 3982 15750 4034 15802
rect 4046 15750 4098 15802
rect 9471 15750 9523 15802
rect 9535 15750 9587 15802
rect 9599 15750 9651 15802
rect 9663 15750 9715 15802
rect 9727 15750 9779 15802
rect 15152 15750 15204 15802
rect 15216 15750 15268 15802
rect 15280 15750 15332 15802
rect 15344 15750 15396 15802
rect 15408 15750 15460 15802
rect 20833 15750 20885 15802
rect 20897 15750 20949 15802
rect 20961 15750 21013 15802
rect 21025 15750 21077 15802
rect 21089 15750 21141 15802
rect 1584 15691 1636 15700
rect 1584 15657 1593 15691
rect 1593 15657 1627 15691
rect 1627 15657 1636 15691
rect 1584 15648 1636 15657
rect 2504 15691 2556 15700
rect 2504 15657 2513 15691
rect 2513 15657 2547 15691
rect 2547 15657 2556 15691
rect 2504 15648 2556 15657
rect 4712 15648 4764 15700
rect 7104 15648 7156 15700
rect 8392 15691 8444 15700
rect 8392 15657 8401 15691
rect 8401 15657 8435 15691
rect 8435 15657 8444 15691
rect 8392 15648 8444 15657
rect 12808 15691 12860 15700
rect 12808 15657 12817 15691
rect 12817 15657 12851 15691
rect 12851 15657 12860 15691
rect 12808 15648 12860 15657
rect 16580 15691 16632 15700
rect 16580 15657 16589 15691
rect 16589 15657 16623 15691
rect 16623 15657 16632 15691
rect 16580 15648 16632 15657
rect 5448 15580 5500 15632
rect 7380 15580 7432 15632
rect 1952 15512 2004 15564
rect 3424 15512 3476 15564
rect 7196 15555 7248 15564
rect 7196 15521 7205 15555
rect 7205 15521 7239 15555
rect 7239 15521 7248 15555
rect 7196 15512 7248 15521
rect 8024 15512 8076 15564
rect 9220 15512 9272 15564
rect 11152 15555 11204 15564
rect 11152 15521 11161 15555
rect 11161 15521 11195 15555
rect 11195 15521 11204 15555
rect 11152 15512 11204 15521
rect 1860 15444 1912 15496
rect 3056 15444 3108 15496
rect 4528 15444 4580 15496
rect 4620 15444 4672 15496
rect 4160 15376 4212 15428
rect 4804 15376 4856 15428
rect 5264 15376 5316 15428
rect 6276 15444 6328 15496
rect 7564 15444 7616 15496
rect 9128 15487 9180 15496
rect 9128 15453 9137 15487
rect 9137 15453 9171 15487
rect 9171 15453 9180 15487
rect 9128 15444 9180 15453
rect 9404 15444 9456 15496
rect 11060 15444 11112 15496
rect 11428 15512 11480 15564
rect 12256 15512 12308 15564
rect 11980 15487 12032 15496
rect 11980 15453 11989 15487
rect 11989 15453 12023 15487
rect 12023 15453 12032 15487
rect 11980 15444 12032 15453
rect 12808 15444 12860 15496
rect 13084 15487 13136 15496
rect 13084 15453 13093 15487
rect 13093 15453 13127 15487
rect 13127 15453 13136 15487
rect 13268 15487 13320 15496
rect 13084 15444 13136 15453
rect 13268 15453 13277 15487
rect 13277 15453 13311 15487
rect 13311 15453 13320 15487
rect 13268 15444 13320 15453
rect 13636 15512 13688 15564
rect 14188 15512 14240 15564
rect 13912 15444 13964 15496
rect 14556 15487 14608 15496
rect 14556 15453 14565 15487
rect 14565 15453 14599 15487
rect 14599 15453 14608 15487
rect 14556 15444 14608 15453
rect 15292 15444 15344 15496
rect 7472 15376 7524 15428
rect 8300 15376 8352 15428
rect 9864 15376 9916 15428
rect 2504 15308 2556 15360
rect 2872 15351 2924 15360
rect 2872 15317 2881 15351
rect 2881 15317 2915 15351
rect 2915 15317 2924 15351
rect 2872 15308 2924 15317
rect 3976 15351 4028 15360
rect 3976 15317 3985 15351
rect 3985 15317 4019 15351
rect 4019 15317 4028 15351
rect 3976 15308 4028 15317
rect 4988 15308 5040 15360
rect 5448 15308 5500 15360
rect 5908 15351 5960 15360
rect 5908 15317 5917 15351
rect 5917 15317 5951 15351
rect 5951 15317 5960 15351
rect 5908 15308 5960 15317
rect 8024 15351 8076 15360
rect 8024 15317 8033 15351
rect 8033 15317 8067 15351
rect 8067 15317 8076 15351
rect 8024 15308 8076 15317
rect 10692 15308 10744 15360
rect 11152 15308 11204 15360
rect 19064 15376 19116 15428
rect 16948 15351 17000 15360
rect 16948 15317 16957 15351
rect 16957 15317 16991 15351
rect 16991 15317 17000 15351
rect 16948 15308 17000 15317
rect 17040 15351 17092 15360
rect 17040 15317 17049 15351
rect 17049 15317 17083 15351
rect 17083 15317 17092 15351
rect 17040 15308 17092 15317
rect 18696 15308 18748 15360
rect 6630 15206 6682 15258
rect 6694 15206 6746 15258
rect 6758 15206 6810 15258
rect 6822 15206 6874 15258
rect 6886 15206 6938 15258
rect 12311 15206 12363 15258
rect 12375 15206 12427 15258
rect 12439 15206 12491 15258
rect 12503 15206 12555 15258
rect 12567 15206 12619 15258
rect 17992 15206 18044 15258
rect 18056 15206 18108 15258
rect 18120 15206 18172 15258
rect 18184 15206 18236 15258
rect 18248 15206 18300 15258
rect 23673 15206 23725 15258
rect 23737 15206 23789 15258
rect 23801 15206 23853 15258
rect 23865 15206 23917 15258
rect 23929 15206 23981 15258
rect 2504 15079 2556 15088
rect 2504 15045 2513 15079
rect 2513 15045 2547 15079
rect 2547 15045 2556 15079
rect 2504 15036 2556 15045
rect 4252 15104 4304 15156
rect 4344 15147 4396 15156
rect 4344 15113 4353 15147
rect 4353 15113 4387 15147
rect 4387 15113 4396 15147
rect 4344 15104 4396 15113
rect 4528 15104 4580 15156
rect 1860 14968 1912 15020
rect 2596 14968 2648 15020
rect 5172 15036 5224 15088
rect 5540 15104 5592 15156
rect 7748 15104 7800 15156
rect 11612 15104 11664 15156
rect 13268 15104 13320 15156
rect 14556 15147 14608 15156
rect 14556 15113 14565 15147
rect 14565 15113 14599 15147
rect 14599 15113 14608 15147
rect 14556 15104 14608 15113
rect 15292 15147 15344 15156
rect 15292 15113 15301 15147
rect 15301 15113 15335 15147
rect 15335 15113 15344 15147
rect 15292 15104 15344 15113
rect 3148 14968 3200 15020
rect 3516 15011 3568 15020
rect 3516 14977 3525 15011
rect 3525 14977 3559 15011
rect 3559 14977 3568 15011
rect 3516 14968 3568 14977
rect 2044 14943 2096 14952
rect 2044 14909 2053 14943
rect 2053 14909 2087 14943
rect 2087 14909 2096 14943
rect 2044 14900 2096 14909
rect 2688 14900 2740 14952
rect 3700 15011 3752 15020
rect 3700 14977 3709 15011
rect 3709 14977 3743 15011
rect 3743 14977 3752 15011
rect 4528 15011 4580 15020
rect 3700 14968 3752 14977
rect 4528 14977 4537 15011
rect 4537 14977 4571 15011
rect 4571 14977 4580 15011
rect 4528 14968 4580 14977
rect 4620 15011 4672 15020
rect 4620 14977 4629 15011
rect 4629 14977 4663 15011
rect 4663 14977 4672 15011
rect 4620 14968 4672 14977
rect 4804 14968 4856 15020
rect 5448 14968 5500 15020
rect 6644 15079 6696 15088
rect 6644 15045 6653 15079
rect 6653 15045 6687 15079
rect 6687 15045 6696 15079
rect 6644 15036 6696 15045
rect 8300 15079 8352 15088
rect 8300 15045 8309 15079
rect 8309 15045 8343 15079
rect 8343 15045 8352 15079
rect 8300 15036 8352 15045
rect 10784 15079 10836 15088
rect 10784 15045 10793 15079
rect 10793 15045 10827 15079
rect 10827 15045 10836 15079
rect 10784 15036 10836 15045
rect 3976 14900 4028 14952
rect 8024 14968 8076 15020
rect 8392 14968 8444 15020
rect 8484 15011 8536 15020
rect 8484 14977 8493 15011
rect 8493 14977 8527 15011
rect 8527 14977 8536 15011
rect 8484 14968 8536 14977
rect 9312 14968 9364 15020
rect 11520 14968 11572 15020
rect 13084 15036 13136 15088
rect 14096 15036 14148 15088
rect 15476 15079 15528 15088
rect 12808 15011 12860 15020
rect 12808 14977 12817 15011
rect 12817 14977 12851 15011
rect 12851 14977 12860 15011
rect 12808 14968 12860 14977
rect 13820 15011 13872 15020
rect 13820 14977 13829 15011
rect 13829 14977 13863 15011
rect 13863 14977 13872 15011
rect 13820 14968 13872 14977
rect 11060 14943 11112 14952
rect 11060 14909 11069 14943
rect 11069 14909 11103 14943
rect 11103 14909 11112 14943
rect 11060 14900 11112 14909
rect 2504 14832 2556 14884
rect 3148 14832 3200 14884
rect 3332 14832 3384 14884
rect 8852 14832 8904 14884
rect 9404 14832 9456 14884
rect 11244 14832 11296 14884
rect 11428 14832 11480 14884
rect 14280 14968 14332 15020
rect 15476 15045 15485 15079
rect 15485 15045 15519 15079
rect 15519 15045 15528 15079
rect 15476 15036 15528 15045
rect 16764 15036 16816 15088
rect 19248 15104 19300 15156
rect 16212 14968 16264 15020
rect 16580 14968 16632 15020
rect 17132 15011 17184 15020
rect 17132 14977 17141 15011
rect 17141 14977 17175 15011
rect 17175 14977 17184 15011
rect 17132 14968 17184 14977
rect 18696 15011 18748 15020
rect 18696 14977 18705 15011
rect 18705 14977 18739 15011
rect 18739 14977 18748 15011
rect 18696 14968 18748 14977
rect 18604 14900 18656 14952
rect 14188 14832 14240 14884
rect 14556 14832 14608 14884
rect 15844 14875 15896 14884
rect 1860 14807 1912 14816
rect 1860 14773 1869 14807
rect 1869 14773 1903 14807
rect 1903 14773 1912 14807
rect 1860 14764 1912 14773
rect 1952 14764 2004 14816
rect 2872 14807 2924 14816
rect 2872 14773 2881 14807
rect 2881 14773 2915 14807
rect 2915 14773 2924 14807
rect 2872 14764 2924 14773
rect 3700 14764 3752 14816
rect 5356 14807 5408 14816
rect 5356 14773 5365 14807
rect 5365 14773 5399 14807
rect 5399 14773 5408 14807
rect 5356 14764 5408 14773
rect 6460 14764 6512 14816
rect 7012 14764 7064 14816
rect 8944 14764 8996 14816
rect 9220 14807 9272 14816
rect 9220 14773 9229 14807
rect 9229 14773 9263 14807
rect 9263 14773 9272 14807
rect 9220 14764 9272 14773
rect 10508 14807 10560 14816
rect 10508 14773 10517 14807
rect 10517 14773 10551 14807
rect 10551 14773 10560 14807
rect 10508 14764 10560 14773
rect 10784 14764 10836 14816
rect 12348 14764 12400 14816
rect 13544 14764 13596 14816
rect 14372 14764 14424 14816
rect 15844 14841 15853 14875
rect 15853 14841 15887 14875
rect 15887 14841 15896 14875
rect 15844 14832 15896 14841
rect 17040 14832 17092 14884
rect 19616 14968 19668 15020
rect 18328 14807 18380 14816
rect 18328 14773 18337 14807
rect 18337 14773 18371 14807
rect 18371 14773 18380 14807
rect 18328 14764 18380 14773
rect 3790 14662 3842 14714
rect 3854 14662 3906 14714
rect 3918 14662 3970 14714
rect 3982 14662 4034 14714
rect 4046 14662 4098 14714
rect 9471 14662 9523 14714
rect 9535 14662 9587 14714
rect 9599 14662 9651 14714
rect 9663 14662 9715 14714
rect 9727 14662 9779 14714
rect 15152 14662 15204 14714
rect 15216 14662 15268 14714
rect 15280 14662 15332 14714
rect 15344 14662 15396 14714
rect 15408 14662 15460 14714
rect 20833 14662 20885 14714
rect 20897 14662 20949 14714
rect 20961 14662 21013 14714
rect 21025 14662 21077 14714
rect 21089 14662 21141 14714
rect 1768 14560 1820 14612
rect 2136 14603 2188 14612
rect 2136 14569 2145 14603
rect 2145 14569 2179 14603
rect 2179 14569 2188 14603
rect 2136 14560 2188 14569
rect 2596 14603 2648 14612
rect 2596 14569 2605 14603
rect 2605 14569 2639 14603
rect 2639 14569 2648 14603
rect 2596 14560 2648 14569
rect 2688 14560 2740 14612
rect 3148 14560 3200 14612
rect 4160 14560 4212 14612
rect 1584 14424 1636 14476
rect 3700 14424 3752 14476
rect 3976 14492 4028 14544
rect 5632 14560 5684 14612
rect 6368 14560 6420 14612
rect 6828 14560 6880 14612
rect 4344 14492 4396 14544
rect 4988 14492 5040 14544
rect 5264 14492 5316 14544
rect 8024 14560 8076 14612
rect 10784 14603 10836 14612
rect 10784 14569 10793 14603
rect 10793 14569 10827 14603
rect 10827 14569 10836 14603
rect 10784 14560 10836 14569
rect 5724 14467 5776 14476
rect 2872 14356 2924 14408
rect 5448 14399 5500 14408
rect 2412 14288 2464 14340
rect 2964 14331 3016 14340
rect 2964 14297 2973 14331
rect 2973 14297 3007 14331
rect 3007 14297 3016 14331
rect 2964 14288 3016 14297
rect 3700 14288 3752 14340
rect 2872 14220 2924 14272
rect 4252 14263 4304 14272
rect 4252 14229 4261 14263
rect 4261 14229 4295 14263
rect 4295 14229 4304 14263
rect 4252 14220 4304 14229
rect 5448 14365 5457 14399
rect 5457 14365 5491 14399
rect 5491 14365 5500 14399
rect 5448 14356 5500 14365
rect 5356 14288 5408 14340
rect 5724 14433 5733 14467
rect 5733 14433 5767 14467
rect 5767 14433 5776 14467
rect 5724 14424 5776 14433
rect 6828 14424 6880 14476
rect 10416 14492 10468 14544
rect 11612 14560 11664 14612
rect 12808 14560 12860 14612
rect 13820 14560 13872 14612
rect 15844 14560 15896 14612
rect 15936 14560 15988 14612
rect 16580 14603 16632 14612
rect 11520 14492 11572 14544
rect 6460 14399 6512 14408
rect 6460 14365 6469 14399
rect 6469 14365 6503 14399
rect 6503 14365 6512 14399
rect 6460 14356 6512 14365
rect 5816 14220 5868 14272
rect 6828 14288 6880 14340
rect 7380 14356 7432 14408
rect 7748 14288 7800 14340
rect 9312 14356 9364 14408
rect 9864 14399 9916 14408
rect 9864 14365 9873 14399
rect 9873 14365 9907 14399
rect 9907 14365 9916 14399
rect 9864 14356 9916 14365
rect 11244 14399 11296 14408
rect 11244 14365 11253 14399
rect 11253 14365 11287 14399
rect 11287 14365 11296 14399
rect 11244 14356 11296 14365
rect 9128 14331 9180 14340
rect 9128 14297 9137 14331
rect 9137 14297 9171 14331
rect 9171 14297 9180 14331
rect 9128 14288 9180 14297
rect 11060 14288 11112 14340
rect 11704 14356 11756 14408
rect 12716 14356 12768 14408
rect 13084 14356 13136 14408
rect 14372 14399 14424 14408
rect 11796 14288 11848 14340
rect 12348 14331 12400 14340
rect 12348 14297 12357 14331
rect 12357 14297 12391 14331
rect 12391 14297 12400 14331
rect 12348 14288 12400 14297
rect 14372 14365 14381 14399
rect 14381 14365 14415 14399
rect 14415 14365 14424 14399
rect 14372 14356 14424 14365
rect 14464 14399 14516 14408
rect 14464 14365 14473 14399
rect 14473 14365 14507 14399
rect 14507 14365 14516 14399
rect 14740 14399 14792 14408
rect 14464 14356 14516 14365
rect 14740 14365 14749 14399
rect 14749 14365 14783 14399
rect 14783 14365 14792 14399
rect 14740 14356 14792 14365
rect 15568 14424 15620 14476
rect 16120 14492 16172 14544
rect 16580 14569 16589 14603
rect 16589 14569 16623 14603
rect 16623 14569 16632 14603
rect 16580 14560 16632 14569
rect 16672 14560 16724 14612
rect 18420 14560 18472 14612
rect 15384 14288 15436 14340
rect 15660 14399 15712 14408
rect 15660 14365 15669 14399
rect 15669 14365 15703 14399
rect 15703 14365 15712 14399
rect 15936 14399 15988 14408
rect 15660 14356 15712 14365
rect 15936 14365 15945 14399
rect 15945 14365 15979 14399
rect 15979 14365 15988 14399
rect 15936 14356 15988 14365
rect 16212 14356 16264 14408
rect 16672 14356 16724 14408
rect 15844 14288 15896 14340
rect 17040 14399 17092 14408
rect 17040 14365 17049 14399
rect 17049 14365 17083 14399
rect 17083 14365 17092 14399
rect 19984 14492 20036 14544
rect 19064 14424 19116 14476
rect 17040 14356 17092 14365
rect 18420 14356 18472 14408
rect 19708 14356 19760 14408
rect 20444 14356 20496 14408
rect 8116 14220 8168 14272
rect 9220 14220 9272 14272
rect 9956 14263 10008 14272
rect 9956 14229 9965 14263
rect 9965 14229 9999 14263
rect 9999 14229 10008 14263
rect 9956 14220 10008 14229
rect 13820 14220 13872 14272
rect 15292 14220 15344 14272
rect 15660 14220 15712 14272
rect 16212 14220 16264 14272
rect 16672 14220 16724 14272
rect 21640 14288 21692 14340
rect 18512 14263 18564 14272
rect 18512 14229 18521 14263
rect 18521 14229 18555 14263
rect 18555 14229 18564 14263
rect 18512 14220 18564 14229
rect 19156 14220 19208 14272
rect 19616 14220 19668 14272
rect 6630 14118 6682 14170
rect 6694 14118 6746 14170
rect 6758 14118 6810 14170
rect 6822 14118 6874 14170
rect 6886 14118 6938 14170
rect 12311 14118 12363 14170
rect 12375 14118 12427 14170
rect 12439 14118 12491 14170
rect 12503 14118 12555 14170
rect 12567 14118 12619 14170
rect 17992 14118 18044 14170
rect 18056 14118 18108 14170
rect 18120 14118 18172 14170
rect 18184 14118 18236 14170
rect 18248 14118 18300 14170
rect 23673 14118 23725 14170
rect 23737 14118 23789 14170
rect 23801 14118 23853 14170
rect 23865 14118 23917 14170
rect 23929 14118 23981 14170
rect 1860 14016 1912 14068
rect 2688 14016 2740 14068
rect 4896 14059 4948 14068
rect 4896 14025 4905 14059
rect 4905 14025 4939 14059
rect 4939 14025 4948 14059
rect 4896 14016 4948 14025
rect 2412 13991 2464 14000
rect 2412 13957 2421 13991
rect 2421 13957 2455 13991
rect 2455 13957 2464 13991
rect 2412 13948 2464 13957
rect 1768 13880 1820 13932
rect 2136 13880 2188 13932
rect 2872 13880 2924 13932
rect 3608 13948 3660 14000
rect 4528 13948 4580 14000
rect 5172 13991 5224 14000
rect 4160 13923 4212 13932
rect 4160 13889 4169 13923
rect 4169 13889 4203 13923
rect 4203 13889 4212 13923
rect 4160 13880 4212 13889
rect 4436 13880 4488 13932
rect 5172 13957 5181 13991
rect 5181 13957 5215 13991
rect 5215 13957 5224 13991
rect 5172 13948 5224 13957
rect 5724 13948 5776 14000
rect 6828 13991 6880 14000
rect 6828 13957 6837 13991
rect 6837 13957 6871 13991
rect 6871 13957 6880 13991
rect 6828 13948 6880 13957
rect 5908 13880 5960 13932
rect 6368 13880 6420 13932
rect 6920 13923 6972 13932
rect 6920 13889 6929 13923
rect 6929 13889 6963 13923
rect 6963 13889 6972 13923
rect 6920 13880 6972 13889
rect 7288 14016 7340 14068
rect 8300 14059 8352 14068
rect 8300 14025 8309 14059
rect 8309 14025 8343 14059
rect 8343 14025 8352 14059
rect 8300 14016 8352 14025
rect 9036 14059 9088 14068
rect 9036 14025 9045 14059
rect 9045 14025 9079 14059
rect 9079 14025 9088 14059
rect 9036 14016 9088 14025
rect 11336 14016 11388 14068
rect 13820 14016 13872 14068
rect 14464 14016 14516 14068
rect 15292 14016 15344 14068
rect 16672 14016 16724 14068
rect 17040 14016 17092 14068
rect 18788 14016 18840 14068
rect 19156 14059 19208 14068
rect 19156 14025 19165 14059
rect 19165 14025 19199 14059
rect 19199 14025 19208 14059
rect 19156 14016 19208 14025
rect 7104 13948 7156 14000
rect 7380 13948 7432 14000
rect 8024 13948 8076 14000
rect 12164 13948 12216 14000
rect 14740 13991 14792 14000
rect 7288 13880 7340 13932
rect 7748 13880 7800 13932
rect 9220 13923 9272 13932
rect 9220 13889 9229 13923
rect 9229 13889 9263 13923
rect 9263 13889 9272 13923
rect 9220 13880 9272 13889
rect 9312 13880 9364 13932
rect 10784 13880 10836 13932
rect 9036 13812 9088 13864
rect 10692 13812 10744 13864
rect 2688 13744 2740 13796
rect 5356 13744 5408 13796
rect 5448 13744 5500 13796
rect 3148 13719 3200 13728
rect 3148 13685 3157 13719
rect 3157 13685 3191 13719
rect 3191 13685 3200 13719
rect 3148 13676 3200 13685
rect 4804 13676 4856 13728
rect 7012 13744 7064 13796
rect 8116 13787 8168 13796
rect 8116 13753 8125 13787
rect 8125 13753 8159 13787
rect 8159 13753 8168 13787
rect 8116 13744 8168 13753
rect 10784 13744 10836 13796
rect 11520 13812 11572 13864
rect 13360 13880 13412 13932
rect 14740 13957 14749 13991
rect 14749 13957 14783 13991
rect 14783 13957 14792 13991
rect 14740 13948 14792 13957
rect 16764 13948 16816 14000
rect 16948 13948 17000 14000
rect 14556 13923 14608 13932
rect 14556 13889 14565 13923
rect 14565 13889 14599 13923
rect 14599 13889 14608 13923
rect 14556 13880 14608 13889
rect 15752 13880 15804 13932
rect 18328 13948 18380 14000
rect 18604 13948 18656 14000
rect 19524 13991 19576 14000
rect 19524 13957 19533 13991
rect 19533 13957 19567 13991
rect 19567 13957 19576 13991
rect 19524 13948 19576 13957
rect 12164 13855 12216 13864
rect 12164 13821 12173 13855
rect 12173 13821 12207 13855
rect 12207 13821 12216 13855
rect 12164 13812 12216 13821
rect 14004 13812 14056 13864
rect 15384 13855 15436 13864
rect 15384 13821 15393 13855
rect 15393 13821 15427 13855
rect 15427 13821 15436 13855
rect 15384 13812 15436 13821
rect 12992 13744 13044 13796
rect 16304 13812 16356 13864
rect 18420 13923 18472 13932
rect 17776 13812 17828 13864
rect 17868 13812 17920 13864
rect 18420 13889 18429 13923
rect 18429 13889 18463 13923
rect 18463 13889 18472 13923
rect 18420 13880 18472 13889
rect 19340 13923 19392 13932
rect 19340 13889 19349 13923
rect 19349 13889 19383 13923
rect 19383 13889 19392 13923
rect 19340 13880 19392 13889
rect 19432 13923 19484 13932
rect 19432 13889 19441 13923
rect 19441 13889 19475 13923
rect 19475 13889 19484 13923
rect 19708 13923 19760 13932
rect 19432 13880 19484 13889
rect 19708 13889 19717 13923
rect 19717 13889 19751 13923
rect 19751 13889 19760 13923
rect 19708 13880 19760 13889
rect 19984 13880 20036 13932
rect 20352 13923 20404 13932
rect 20352 13889 20361 13923
rect 20361 13889 20395 13923
rect 20395 13889 20404 13923
rect 20352 13880 20404 13889
rect 18328 13855 18380 13864
rect 18328 13821 18337 13855
rect 18337 13821 18371 13855
rect 18371 13821 18380 13855
rect 18328 13812 18380 13821
rect 6276 13676 6328 13728
rect 6736 13676 6788 13728
rect 10416 13676 10468 13728
rect 12440 13676 12492 13728
rect 13636 13676 13688 13728
rect 18420 13744 18472 13796
rect 15660 13676 15712 13728
rect 16212 13676 16264 13728
rect 17224 13676 17276 13728
rect 18696 13676 18748 13728
rect 3790 13574 3842 13626
rect 3854 13574 3906 13626
rect 3918 13574 3970 13626
rect 3982 13574 4034 13626
rect 4046 13574 4098 13626
rect 9471 13574 9523 13626
rect 9535 13574 9587 13626
rect 9599 13574 9651 13626
rect 9663 13574 9715 13626
rect 9727 13574 9779 13626
rect 15152 13574 15204 13626
rect 15216 13574 15268 13626
rect 15280 13574 15332 13626
rect 15344 13574 15396 13626
rect 15408 13574 15460 13626
rect 20833 13574 20885 13626
rect 20897 13574 20949 13626
rect 20961 13574 21013 13626
rect 21025 13574 21077 13626
rect 21089 13574 21141 13626
rect 3516 13472 3568 13524
rect 4436 13472 4488 13524
rect 4620 13472 4672 13524
rect 4712 13472 4764 13524
rect 4252 13404 4304 13456
rect 6276 13472 6328 13524
rect 6828 13472 6880 13524
rect 8852 13472 8904 13524
rect 10784 13472 10836 13524
rect 11244 13472 11296 13524
rect 11704 13472 11756 13524
rect 12164 13472 12216 13524
rect 5724 13404 5776 13456
rect 1860 13311 1912 13320
rect 1860 13277 1869 13311
rect 1869 13277 1903 13311
rect 1903 13277 1912 13311
rect 1860 13268 1912 13277
rect 2044 13311 2096 13320
rect 2044 13277 2053 13311
rect 2053 13277 2087 13311
rect 2087 13277 2096 13311
rect 2504 13311 2556 13320
rect 2044 13268 2096 13277
rect 2504 13277 2513 13311
rect 2513 13277 2547 13311
rect 2547 13277 2556 13311
rect 4896 13336 4948 13388
rect 6368 13379 6420 13388
rect 6368 13345 6377 13379
rect 6377 13345 6411 13379
rect 6411 13345 6420 13379
rect 6368 13336 6420 13345
rect 6460 13379 6512 13388
rect 6460 13345 6469 13379
rect 6469 13345 6503 13379
rect 6503 13345 6512 13379
rect 6460 13336 6512 13345
rect 9220 13336 9272 13388
rect 9588 13336 9640 13388
rect 2504 13268 2556 13277
rect 3792 13268 3844 13320
rect 2688 13200 2740 13252
rect 4344 13200 4396 13252
rect 5080 13311 5132 13320
rect 5080 13277 5089 13311
rect 5089 13277 5123 13311
rect 5123 13277 5132 13311
rect 5080 13268 5132 13277
rect 5356 13268 5408 13320
rect 6276 13268 6328 13320
rect 6644 13311 6696 13320
rect 6644 13277 6653 13311
rect 6653 13277 6687 13311
rect 6687 13277 6696 13311
rect 7472 13311 7524 13320
rect 6644 13268 6696 13277
rect 7472 13277 7481 13311
rect 7481 13277 7515 13311
rect 7515 13277 7524 13311
rect 7472 13268 7524 13277
rect 7564 13268 7616 13320
rect 8116 13311 8168 13320
rect 8116 13277 8125 13311
rect 8125 13277 8159 13311
rect 8159 13277 8168 13311
rect 8116 13268 8168 13277
rect 9312 13311 9364 13320
rect 9312 13277 9321 13311
rect 9321 13277 9355 13311
rect 9355 13277 9364 13311
rect 9312 13268 9364 13277
rect 11060 13336 11112 13388
rect 11336 13379 11388 13388
rect 11336 13345 11345 13379
rect 11345 13345 11379 13379
rect 11379 13345 11388 13379
rect 11336 13336 11388 13345
rect 12164 13336 12216 13388
rect 14372 13472 14424 13524
rect 15476 13472 15528 13524
rect 16764 13472 16816 13524
rect 18972 13472 19024 13524
rect 19432 13515 19484 13524
rect 19432 13481 19441 13515
rect 19441 13481 19475 13515
rect 19475 13481 19484 13515
rect 19432 13472 19484 13481
rect 19800 13472 19852 13524
rect 12992 13404 13044 13456
rect 14004 13404 14056 13456
rect 14924 13404 14976 13456
rect 15752 13404 15804 13456
rect 17316 13404 17368 13456
rect 11612 13311 11664 13320
rect 11612 13277 11621 13311
rect 11621 13277 11655 13311
rect 11655 13277 11664 13311
rect 11612 13268 11664 13277
rect 12440 13311 12492 13320
rect 12440 13277 12449 13311
rect 12449 13277 12483 13311
rect 12483 13277 12492 13311
rect 12440 13268 12492 13277
rect 13360 13268 13412 13320
rect 15844 13268 15896 13320
rect 16764 13311 16816 13320
rect 16764 13277 16773 13311
rect 16773 13277 16807 13311
rect 16807 13277 16816 13311
rect 16764 13268 16816 13277
rect 17500 13268 17552 13320
rect 19892 13404 19944 13456
rect 18236 13311 18288 13320
rect 18236 13277 18245 13311
rect 18245 13277 18279 13311
rect 18279 13277 18288 13311
rect 18236 13268 18288 13277
rect 18604 13268 18656 13320
rect 18880 13311 18932 13320
rect 18880 13277 18889 13311
rect 18889 13277 18923 13311
rect 18923 13277 18932 13311
rect 18880 13268 18932 13277
rect 18972 13268 19024 13320
rect 19708 13311 19760 13320
rect 19708 13277 19717 13311
rect 19717 13277 19751 13311
rect 19751 13277 19760 13311
rect 19708 13268 19760 13277
rect 5172 13200 5224 13252
rect 6736 13200 6788 13252
rect 2596 13175 2648 13184
rect 2596 13141 2605 13175
rect 2605 13141 2639 13175
rect 2639 13141 2648 13175
rect 2596 13132 2648 13141
rect 2780 13175 2832 13184
rect 2780 13141 2789 13175
rect 2789 13141 2823 13175
rect 2823 13141 2832 13175
rect 5264 13175 5316 13184
rect 2780 13132 2832 13141
rect 5264 13141 5273 13175
rect 5273 13141 5307 13175
rect 5307 13141 5316 13175
rect 5264 13132 5316 13141
rect 5448 13132 5500 13184
rect 7104 13132 7156 13184
rect 7748 13200 7800 13252
rect 9128 13132 9180 13184
rect 17316 13200 17368 13252
rect 20260 13268 20312 13320
rect 21272 13268 21324 13320
rect 21640 13311 21692 13320
rect 21640 13277 21649 13311
rect 21649 13277 21683 13311
rect 21683 13277 21692 13311
rect 21640 13268 21692 13277
rect 16212 13175 16264 13184
rect 16212 13141 16221 13175
rect 16221 13141 16255 13175
rect 16255 13141 16264 13175
rect 16212 13132 16264 13141
rect 17040 13132 17092 13184
rect 18604 13132 18656 13184
rect 18972 13132 19024 13184
rect 20536 13243 20588 13252
rect 20536 13209 20545 13243
rect 20545 13209 20579 13243
rect 20579 13209 20588 13243
rect 20536 13200 20588 13209
rect 20260 13132 20312 13184
rect 6630 13030 6682 13082
rect 6694 13030 6746 13082
rect 6758 13030 6810 13082
rect 6822 13030 6874 13082
rect 6886 13030 6938 13082
rect 12311 13030 12363 13082
rect 12375 13030 12427 13082
rect 12439 13030 12491 13082
rect 12503 13030 12555 13082
rect 12567 13030 12619 13082
rect 17992 13030 18044 13082
rect 18056 13030 18108 13082
rect 18120 13030 18172 13082
rect 18184 13030 18236 13082
rect 18248 13030 18300 13082
rect 23673 13030 23725 13082
rect 23737 13030 23789 13082
rect 23801 13030 23853 13082
rect 23865 13030 23917 13082
rect 23929 13030 23981 13082
rect 1860 12928 1912 12980
rect 2596 12928 2648 12980
rect 2504 12860 2556 12912
rect 1584 12835 1636 12844
rect 1584 12801 1593 12835
rect 1593 12801 1627 12835
rect 1627 12801 1636 12835
rect 1584 12792 1636 12801
rect 3240 12928 3292 12980
rect 4528 12971 4580 12980
rect 4528 12937 4537 12971
rect 4537 12937 4571 12971
rect 4571 12937 4580 12971
rect 4528 12928 4580 12937
rect 7840 12971 7892 12980
rect 2964 12860 3016 12912
rect 6460 12860 6512 12912
rect 6736 12860 6788 12912
rect 3148 12792 3200 12844
rect 3608 12792 3660 12844
rect 3792 12835 3844 12844
rect 3792 12801 3801 12835
rect 3801 12801 3835 12835
rect 3835 12801 3844 12835
rect 4068 12835 4120 12844
rect 3792 12792 3844 12801
rect 4068 12801 4077 12835
rect 4077 12801 4111 12835
rect 4111 12801 4120 12835
rect 4068 12792 4120 12801
rect 4712 12792 4764 12844
rect 6276 12792 6328 12844
rect 7840 12937 7849 12971
rect 7849 12937 7883 12971
rect 7883 12937 7892 12971
rect 7840 12928 7892 12937
rect 8024 12928 8076 12980
rect 15660 12928 15712 12980
rect 16488 12928 16540 12980
rect 7104 12860 7156 12912
rect 8576 12860 8628 12912
rect 9128 12860 9180 12912
rect 10048 12860 10100 12912
rect 11336 12860 11388 12912
rect 7564 12792 7616 12844
rect 9588 12835 9640 12844
rect 9588 12801 9597 12835
rect 9597 12801 9631 12835
rect 9631 12801 9640 12835
rect 9588 12792 9640 12801
rect 11704 12792 11756 12844
rect 14556 12860 14608 12912
rect 15752 12860 15804 12912
rect 18420 12928 18472 12980
rect 19340 12928 19392 12980
rect 15292 12835 15344 12844
rect 15292 12801 15301 12835
rect 15301 12801 15335 12835
rect 15335 12801 15344 12835
rect 15292 12792 15344 12801
rect 15568 12792 15620 12844
rect 17040 12835 17092 12844
rect 3148 12656 3200 12708
rect 3516 12724 3568 12776
rect 5724 12724 5776 12776
rect 6368 12724 6420 12776
rect 6736 12767 6788 12776
rect 6736 12733 6745 12767
rect 6745 12733 6779 12767
rect 6779 12733 6788 12767
rect 6736 12724 6788 12733
rect 7104 12724 7156 12776
rect 7748 12724 7800 12776
rect 8392 12724 8444 12776
rect 8668 12724 8720 12776
rect 9312 12724 9364 12776
rect 13820 12724 13872 12776
rect 4160 12656 4212 12708
rect 4528 12656 4580 12708
rect 7840 12656 7892 12708
rect 8760 12656 8812 12708
rect 13360 12656 13412 12708
rect 15660 12724 15712 12776
rect 2136 12588 2188 12640
rect 2504 12588 2556 12640
rect 4344 12588 4396 12640
rect 5356 12631 5408 12640
rect 5356 12597 5365 12631
rect 5365 12597 5399 12631
rect 5399 12597 5408 12631
rect 5356 12588 5408 12597
rect 7472 12588 7524 12640
rect 9312 12588 9364 12640
rect 14832 12631 14884 12640
rect 14832 12597 14841 12631
rect 14841 12597 14875 12631
rect 14875 12597 14884 12631
rect 14832 12588 14884 12597
rect 15752 12588 15804 12640
rect 16396 12588 16448 12640
rect 17040 12801 17049 12835
rect 17049 12801 17083 12835
rect 17083 12801 17092 12835
rect 17040 12792 17092 12801
rect 17224 12835 17276 12844
rect 17224 12801 17233 12835
rect 17233 12801 17267 12835
rect 17267 12801 17276 12835
rect 17224 12792 17276 12801
rect 18236 12792 18288 12844
rect 18604 12835 18656 12844
rect 17132 12724 17184 12776
rect 17684 12724 17736 12776
rect 18604 12801 18613 12835
rect 18613 12801 18647 12835
rect 18647 12801 18656 12835
rect 18604 12792 18656 12801
rect 18972 12792 19024 12844
rect 19340 12835 19392 12844
rect 19340 12801 19349 12835
rect 19349 12801 19383 12835
rect 19383 12801 19392 12835
rect 19340 12792 19392 12801
rect 19616 12792 19668 12844
rect 20168 12792 20220 12844
rect 20812 12835 20864 12844
rect 20812 12801 20821 12835
rect 20821 12801 20855 12835
rect 20855 12801 20864 12835
rect 20812 12792 20864 12801
rect 17224 12656 17276 12708
rect 18972 12656 19024 12708
rect 20536 12656 20588 12708
rect 18880 12588 18932 12640
rect 19432 12588 19484 12640
rect 20812 12588 20864 12640
rect 21732 12588 21784 12640
rect 22100 12631 22152 12640
rect 22100 12597 22109 12631
rect 22109 12597 22143 12631
rect 22143 12597 22152 12631
rect 22100 12588 22152 12597
rect 3790 12486 3842 12538
rect 3854 12486 3906 12538
rect 3918 12486 3970 12538
rect 3982 12486 4034 12538
rect 4046 12486 4098 12538
rect 9471 12486 9523 12538
rect 9535 12486 9587 12538
rect 9599 12486 9651 12538
rect 9663 12486 9715 12538
rect 9727 12486 9779 12538
rect 15152 12486 15204 12538
rect 15216 12486 15268 12538
rect 15280 12486 15332 12538
rect 15344 12486 15396 12538
rect 15408 12486 15460 12538
rect 20833 12486 20885 12538
rect 20897 12486 20949 12538
rect 20961 12486 21013 12538
rect 21025 12486 21077 12538
rect 21089 12486 21141 12538
rect 1952 12384 2004 12436
rect 5724 12427 5776 12436
rect 5724 12393 5733 12427
rect 5733 12393 5767 12427
rect 5767 12393 5776 12427
rect 5724 12384 5776 12393
rect 6184 12427 6236 12436
rect 6184 12393 6193 12427
rect 6193 12393 6227 12427
rect 6227 12393 6236 12427
rect 6184 12384 6236 12393
rect 7840 12384 7892 12436
rect 8208 12384 8260 12436
rect 11244 12384 11296 12436
rect 5172 12316 5224 12368
rect 6092 12316 6144 12368
rect 4712 12248 4764 12300
rect 5356 12291 5408 12300
rect 5356 12257 5365 12291
rect 5365 12257 5399 12291
rect 5399 12257 5408 12291
rect 5356 12248 5408 12257
rect 2228 12223 2280 12232
rect 2228 12189 2237 12223
rect 2237 12189 2271 12223
rect 2271 12189 2280 12223
rect 2228 12180 2280 12189
rect 4344 12180 4396 12232
rect 5172 12180 5224 12232
rect 5448 12223 5500 12232
rect 5448 12189 5457 12223
rect 5457 12189 5491 12223
rect 5491 12189 5500 12223
rect 5448 12180 5500 12189
rect 1768 12112 1820 12164
rect 2044 12087 2096 12096
rect 2044 12053 2053 12087
rect 2053 12053 2087 12087
rect 2087 12053 2096 12087
rect 2044 12044 2096 12053
rect 2596 12044 2648 12096
rect 3056 12044 3108 12096
rect 5448 12044 5500 12096
rect 7196 12248 7248 12300
rect 6828 12223 6880 12232
rect 6828 12189 6837 12223
rect 6837 12189 6871 12223
rect 6871 12189 6880 12223
rect 6828 12180 6880 12189
rect 6000 12112 6052 12164
rect 6552 12155 6604 12164
rect 6552 12121 6561 12155
rect 6561 12121 6595 12155
rect 6595 12121 6604 12155
rect 6552 12112 6604 12121
rect 8484 12291 8536 12300
rect 7472 12223 7524 12232
rect 7472 12189 7481 12223
rect 7481 12189 7515 12223
rect 7515 12189 7524 12223
rect 7472 12180 7524 12189
rect 8484 12257 8493 12291
rect 8493 12257 8527 12291
rect 8527 12257 8536 12291
rect 8484 12248 8536 12257
rect 8576 12248 8628 12300
rect 7564 12155 7616 12164
rect 7564 12121 7573 12155
rect 7573 12121 7607 12155
rect 7607 12121 7616 12155
rect 7564 12112 7616 12121
rect 9772 12223 9824 12232
rect 9772 12189 9781 12223
rect 9781 12189 9815 12223
rect 9815 12189 9824 12223
rect 9772 12180 9824 12189
rect 12072 12384 12124 12436
rect 12716 12384 12768 12436
rect 13636 12316 13688 12368
rect 15936 12384 15988 12436
rect 16580 12384 16632 12436
rect 17408 12384 17460 12436
rect 18328 12384 18380 12436
rect 12072 12180 12124 12232
rect 13820 12248 13872 12300
rect 12716 12223 12768 12232
rect 12716 12189 12725 12223
rect 12725 12189 12759 12223
rect 12759 12189 12768 12223
rect 12900 12223 12952 12232
rect 12716 12180 12768 12189
rect 12900 12189 12909 12223
rect 12909 12189 12943 12223
rect 12943 12189 12952 12223
rect 12900 12180 12952 12189
rect 13084 12180 13136 12232
rect 14280 12180 14332 12232
rect 7012 12044 7064 12096
rect 7196 12044 7248 12096
rect 8208 12112 8260 12164
rect 8576 12112 8628 12164
rect 9680 12112 9732 12164
rect 9864 12044 9916 12096
rect 10048 12044 10100 12096
rect 10600 12044 10652 12096
rect 11796 12044 11848 12096
rect 12072 12044 12124 12096
rect 12808 12044 12860 12096
rect 14556 12223 14608 12232
rect 14556 12189 14565 12223
rect 14565 12189 14599 12223
rect 14599 12189 14608 12223
rect 14832 12248 14884 12300
rect 14556 12180 14608 12189
rect 15568 12180 15620 12232
rect 15660 12223 15712 12232
rect 15660 12189 15669 12223
rect 15669 12189 15703 12223
rect 15703 12189 15712 12223
rect 16672 12316 16724 12368
rect 17316 12316 17368 12368
rect 15660 12180 15712 12189
rect 17868 12248 17920 12300
rect 18972 12384 19024 12436
rect 20168 12427 20220 12436
rect 20168 12393 20177 12427
rect 20177 12393 20211 12427
rect 20211 12393 20220 12427
rect 20168 12384 20220 12393
rect 17224 12180 17276 12232
rect 17592 12180 17644 12232
rect 18420 12223 18472 12232
rect 18420 12189 18429 12223
rect 18429 12189 18463 12223
rect 18463 12189 18472 12223
rect 18420 12180 18472 12189
rect 18880 12316 18932 12368
rect 19432 12180 19484 12232
rect 19892 12223 19944 12232
rect 19892 12189 19901 12223
rect 19901 12189 19935 12223
rect 19935 12189 19944 12223
rect 19892 12180 19944 12189
rect 20076 12180 20128 12232
rect 21088 12180 21140 12232
rect 21640 12180 21692 12232
rect 16948 12112 17000 12164
rect 15384 12044 15436 12096
rect 16396 12044 16448 12096
rect 16856 12044 16908 12096
rect 17408 12087 17460 12096
rect 17408 12053 17417 12087
rect 17417 12053 17451 12087
rect 17451 12053 17460 12087
rect 17408 12044 17460 12053
rect 17500 12044 17552 12096
rect 17868 12112 17920 12164
rect 20720 12112 20772 12164
rect 21180 12155 21232 12164
rect 21180 12121 21189 12155
rect 21189 12121 21223 12155
rect 21223 12121 21232 12155
rect 21180 12112 21232 12121
rect 22100 12112 22152 12164
rect 23112 12112 23164 12164
rect 21364 12044 21416 12096
rect 22560 12044 22612 12096
rect 6630 11942 6682 11994
rect 6694 11942 6746 11994
rect 6758 11942 6810 11994
rect 6822 11942 6874 11994
rect 6886 11942 6938 11994
rect 12311 11942 12363 11994
rect 12375 11942 12427 11994
rect 12439 11942 12491 11994
rect 12503 11942 12555 11994
rect 12567 11942 12619 11994
rect 17992 11942 18044 11994
rect 18056 11942 18108 11994
rect 18120 11942 18172 11994
rect 18184 11942 18236 11994
rect 18248 11942 18300 11994
rect 23673 11942 23725 11994
rect 23737 11942 23789 11994
rect 23801 11942 23853 11994
rect 23865 11942 23917 11994
rect 23929 11942 23981 11994
rect 2964 11883 3016 11892
rect 2964 11849 2973 11883
rect 2973 11849 3007 11883
rect 3007 11849 3016 11883
rect 2964 11840 3016 11849
rect 4252 11840 4304 11892
rect 4712 11883 4764 11892
rect 4712 11849 4721 11883
rect 4721 11849 4755 11883
rect 4755 11849 4764 11883
rect 4712 11840 4764 11849
rect 5356 11840 5408 11892
rect 6000 11883 6052 11892
rect 6000 11849 6009 11883
rect 6009 11849 6043 11883
rect 6043 11849 6052 11883
rect 6000 11840 6052 11849
rect 3240 11772 3292 11824
rect 2044 11747 2096 11756
rect 2044 11713 2053 11747
rect 2053 11713 2087 11747
rect 2087 11713 2096 11747
rect 2044 11704 2096 11713
rect 2596 11704 2648 11756
rect 2872 11636 2924 11688
rect 2964 11679 3016 11688
rect 2964 11645 2973 11679
rect 2973 11645 3007 11679
rect 3007 11645 3016 11679
rect 4160 11704 4212 11756
rect 4804 11747 4856 11756
rect 4804 11713 4813 11747
rect 4813 11713 4847 11747
rect 4847 11713 4856 11747
rect 4804 11704 4856 11713
rect 5632 11747 5684 11756
rect 5632 11713 5641 11747
rect 5641 11713 5675 11747
rect 5675 11713 5684 11747
rect 7196 11840 7248 11892
rect 7932 11883 7984 11892
rect 7932 11849 7941 11883
rect 7941 11849 7975 11883
rect 7975 11849 7984 11883
rect 7932 11840 7984 11849
rect 8116 11840 8168 11892
rect 8300 11840 8352 11892
rect 9036 11772 9088 11824
rect 5632 11704 5684 11713
rect 5448 11679 5500 11688
rect 2964 11636 3016 11645
rect 5448 11645 5457 11679
rect 5457 11645 5491 11679
rect 5491 11645 5500 11679
rect 5448 11636 5500 11645
rect 6184 11636 6236 11688
rect 7104 11704 7156 11756
rect 7748 11704 7800 11756
rect 8116 11747 8168 11756
rect 8116 11713 8125 11747
rect 8125 11713 8159 11747
rect 8159 11713 8168 11747
rect 8116 11704 8168 11713
rect 8300 11747 8352 11756
rect 8300 11713 8309 11747
rect 8309 11713 8343 11747
rect 8343 11713 8352 11747
rect 8300 11704 8352 11713
rect 9312 11704 9364 11756
rect 10968 11840 11020 11892
rect 13912 11840 13964 11892
rect 15476 11883 15528 11892
rect 15476 11849 15485 11883
rect 15485 11849 15519 11883
rect 15519 11849 15528 11883
rect 15476 11840 15528 11849
rect 16212 11840 16264 11892
rect 16304 11840 16356 11892
rect 10968 11704 11020 11756
rect 11428 11772 11480 11824
rect 13268 11772 13320 11824
rect 14096 11772 14148 11824
rect 11888 11747 11940 11756
rect 11888 11713 11897 11747
rect 11897 11713 11931 11747
rect 11931 11713 11940 11747
rect 11888 11704 11940 11713
rect 12164 11704 12216 11756
rect 12900 11747 12952 11756
rect 12900 11713 12909 11747
rect 12909 11713 12943 11747
rect 12943 11713 12952 11747
rect 12900 11704 12952 11713
rect 13636 11704 13688 11756
rect 14372 11704 14424 11756
rect 14556 11704 14608 11756
rect 15384 11747 15436 11756
rect 2780 11611 2832 11620
rect 2780 11577 2789 11611
rect 2789 11577 2823 11611
rect 2823 11577 2832 11611
rect 2780 11568 2832 11577
rect 5172 11568 5224 11620
rect 7288 11568 7340 11620
rect 8116 11568 8168 11620
rect 9680 11568 9732 11620
rect 10232 11611 10284 11620
rect 10232 11577 10241 11611
rect 10241 11577 10275 11611
rect 10275 11577 10284 11611
rect 10232 11568 10284 11577
rect 10600 11636 10652 11688
rect 10784 11568 10836 11620
rect 14280 11636 14332 11688
rect 14832 11679 14884 11688
rect 14832 11645 14841 11679
rect 14841 11645 14875 11679
rect 14875 11645 14884 11679
rect 14832 11636 14884 11645
rect 15384 11713 15393 11747
rect 15393 11713 15427 11747
rect 15427 11713 15436 11747
rect 15384 11704 15436 11713
rect 15568 11704 15620 11756
rect 16948 11772 17000 11824
rect 17316 11840 17368 11892
rect 17960 11883 18012 11892
rect 17960 11849 17969 11883
rect 17969 11849 18003 11883
rect 18003 11849 18012 11883
rect 17960 11840 18012 11849
rect 18328 11840 18380 11892
rect 18512 11840 18564 11892
rect 17500 11772 17552 11824
rect 19064 11772 19116 11824
rect 20076 11772 20128 11824
rect 20168 11772 20220 11824
rect 21824 11772 21876 11824
rect 17408 11704 17460 11756
rect 20260 11747 20312 11756
rect 20260 11713 20269 11747
rect 20269 11713 20303 11747
rect 20303 11713 20312 11747
rect 20260 11704 20312 11713
rect 20444 11704 20496 11756
rect 21180 11747 21232 11756
rect 16948 11636 17000 11688
rect 17132 11679 17184 11688
rect 17132 11645 17141 11679
rect 17141 11645 17175 11679
rect 17175 11645 17184 11679
rect 17132 11636 17184 11645
rect 18604 11679 18656 11688
rect 13452 11568 13504 11620
rect 15016 11568 15068 11620
rect 16028 11568 16080 11620
rect 18604 11645 18613 11679
rect 18613 11645 18647 11679
rect 18647 11645 18656 11679
rect 18604 11636 18656 11645
rect 17684 11568 17736 11620
rect 18328 11568 18380 11620
rect 20168 11636 20220 11688
rect 21180 11713 21189 11747
rect 21189 11713 21223 11747
rect 21223 11713 21232 11747
rect 21180 11704 21232 11713
rect 21640 11704 21692 11756
rect 21916 11636 21968 11688
rect 19248 11568 19300 11620
rect 19616 11568 19668 11620
rect 20444 11611 20496 11620
rect 20444 11577 20453 11611
rect 20453 11577 20487 11611
rect 20487 11577 20496 11611
rect 20444 11568 20496 11577
rect 3608 11500 3660 11552
rect 7564 11500 7616 11552
rect 7840 11500 7892 11552
rect 8392 11500 8444 11552
rect 10324 11543 10376 11552
rect 10324 11509 10333 11543
rect 10333 11509 10367 11543
rect 10367 11509 10376 11543
rect 10324 11500 10376 11509
rect 13084 11543 13136 11552
rect 13084 11509 13093 11543
rect 13093 11509 13127 11543
rect 13127 11509 13136 11543
rect 13084 11500 13136 11509
rect 14004 11543 14056 11552
rect 14004 11509 14013 11543
rect 14013 11509 14047 11543
rect 14047 11509 14056 11543
rect 14004 11500 14056 11509
rect 16672 11500 16724 11552
rect 17408 11500 17460 11552
rect 22008 11500 22060 11552
rect 22192 11704 22244 11756
rect 22560 11704 22612 11756
rect 22192 11500 22244 11552
rect 23112 11500 23164 11552
rect 3790 11398 3842 11450
rect 3854 11398 3906 11450
rect 3918 11398 3970 11450
rect 3982 11398 4034 11450
rect 4046 11398 4098 11450
rect 9471 11398 9523 11450
rect 9535 11398 9587 11450
rect 9599 11398 9651 11450
rect 9663 11398 9715 11450
rect 9727 11398 9779 11450
rect 15152 11398 15204 11450
rect 15216 11398 15268 11450
rect 15280 11398 15332 11450
rect 15344 11398 15396 11450
rect 15408 11398 15460 11450
rect 20833 11398 20885 11450
rect 20897 11398 20949 11450
rect 20961 11398 21013 11450
rect 21025 11398 21077 11450
rect 21089 11398 21141 11450
rect 1584 11296 1636 11348
rect 1768 11228 1820 11280
rect 2412 11228 2464 11280
rect 3148 11228 3200 11280
rect 3424 11228 3476 11280
rect 2872 11160 2924 11212
rect 3056 11160 3108 11212
rect 3240 11160 3292 11212
rect 2504 11092 2556 11144
rect 2780 11092 2832 11144
rect 3424 11135 3476 11144
rect 3424 11101 3433 11135
rect 3433 11101 3467 11135
rect 3467 11101 3476 11135
rect 3424 11092 3476 11101
rect 4068 11092 4120 11144
rect 4344 11092 4396 11144
rect 1492 11024 1544 11076
rect 2228 11024 2280 11076
rect 4988 11067 5040 11076
rect 4988 11033 4997 11067
rect 4997 11033 5031 11067
rect 5031 11033 5040 11067
rect 4988 11024 5040 11033
rect 5080 11024 5132 11076
rect 5448 11296 5500 11348
rect 6276 11339 6328 11348
rect 6276 11305 6285 11339
rect 6285 11305 6319 11339
rect 6319 11305 6328 11339
rect 6276 11296 6328 11305
rect 7656 11296 7708 11348
rect 8392 11339 8444 11348
rect 8392 11305 8401 11339
rect 8401 11305 8435 11339
rect 8435 11305 8444 11339
rect 8392 11296 8444 11305
rect 8576 11339 8628 11348
rect 8576 11305 8585 11339
rect 8585 11305 8619 11339
rect 8619 11305 8628 11339
rect 8576 11296 8628 11305
rect 9864 11296 9916 11348
rect 13084 11296 13136 11348
rect 14372 11296 14424 11348
rect 14832 11296 14884 11348
rect 16488 11339 16540 11348
rect 16488 11305 16497 11339
rect 16497 11305 16531 11339
rect 16531 11305 16540 11339
rect 16488 11296 16540 11305
rect 17224 11339 17276 11348
rect 17224 11305 17233 11339
rect 17233 11305 17267 11339
rect 17267 11305 17276 11339
rect 17224 11296 17276 11305
rect 17592 11296 17644 11348
rect 20352 11339 20404 11348
rect 20352 11305 20361 11339
rect 20361 11305 20395 11339
rect 20395 11305 20404 11339
rect 20352 11296 20404 11305
rect 20720 11296 20772 11348
rect 21732 11339 21784 11348
rect 21732 11305 21741 11339
rect 21741 11305 21775 11339
rect 21775 11305 21784 11339
rect 21732 11296 21784 11305
rect 9036 11228 9088 11280
rect 9220 11228 9272 11280
rect 9404 11228 9456 11280
rect 11336 11228 11388 11280
rect 11612 11228 11664 11280
rect 5632 11160 5684 11212
rect 6276 11160 6328 11212
rect 7104 11135 7156 11144
rect 5724 11024 5776 11076
rect 7104 11101 7113 11135
rect 7113 11101 7147 11135
rect 7147 11101 7156 11135
rect 7104 11092 7156 11101
rect 7196 11135 7248 11144
rect 7196 11101 7205 11135
rect 7205 11101 7239 11135
rect 7239 11101 7248 11135
rect 7564 11135 7616 11144
rect 7196 11092 7248 11101
rect 7564 11101 7573 11135
rect 7573 11101 7607 11135
rect 7607 11101 7616 11135
rect 7564 11092 7616 11101
rect 6184 11024 6236 11076
rect 7012 11024 7064 11076
rect 7288 11067 7340 11076
rect 7288 11033 7297 11067
rect 7297 11033 7331 11067
rect 7331 11033 7340 11067
rect 7288 11024 7340 11033
rect 8116 11024 8168 11076
rect 9128 11092 9180 11144
rect 9404 11135 9456 11144
rect 9404 11101 9413 11135
rect 9413 11101 9447 11135
rect 9447 11101 9456 11135
rect 10232 11160 10284 11212
rect 9404 11092 9456 11101
rect 10324 11135 10376 11144
rect 8484 11024 8536 11076
rect 9036 11024 9088 11076
rect 10324 11101 10333 11135
rect 10333 11101 10367 11135
rect 10367 11101 10376 11135
rect 10324 11092 10376 11101
rect 10600 11024 10652 11076
rect 11612 11092 11664 11144
rect 13176 11135 13228 11144
rect 13176 11101 13185 11135
rect 13185 11101 13219 11135
rect 13219 11101 13228 11135
rect 17868 11228 17920 11280
rect 18328 11228 18380 11280
rect 13820 11160 13872 11212
rect 14556 11203 14608 11212
rect 14556 11169 14565 11203
rect 14565 11169 14599 11203
rect 14599 11169 14608 11203
rect 14556 11160 14608 11169
rect 13176 11092 13228 11101
rect 11704 11024 11756 11076
rect 12716 11024 12768 11076
rect 12992 11024 13044 11076
rect 13084 11024 13136 11076
rect 14464 11135 14516 11144
rect 14464 11101 14473 11135
rect 14473 11101 14507 11135
rect 14507 11101 14516 11135
rect 14464 11092 14516 11101
rect 2780 10956 2832 11008
rect 4252 10956 4304 11008
rect 7840 10956 7892 11008
rect 13176 10999 13228 11008
rect 13176 10965 13185 10999
rect 13185 10965 13219 10999
rect 13219 10965 13228 10999
rect 13176 10956 13228 10965
rect 13636 11024 13688 11076
rect 14832 11092 14884 11144
rect 16120 11160 16172 11212
rect 15476 11092 15528 11144
rect 15752 11092 15804 11144
rect 16028 11135 16080 11144
rect 16028 11101 16037 11135
rect 16037 11101 16071 11135
rect 16071 11101 16080 11135
rect 16028 11092 16080 11101
rect 16396 11092 16448 11144
rect 16948 11135 17000 11144
rect 16948 11101 16957 11135
rect 16957 11101 16991 11135
rect 16991 11101 17000 11135
rect 16948 11092 17000 11101
rect 17684 11092 17736 11144
rect 19616 11228 19668 11280
rect 19892 11228 19944 11280
rect 19524 11160 19576 11212
rect 18512 11092 18564 11144
rect 18788 11092 18840 11144
rect 18972 11092 19024 11144
rect 19432 11135 19484 11144
rect 19432 11101 19441 11135
rect 19441 11101 19475 11135
rect 19475 11101 19484 11135
rect 19432 11092 19484 11101
rect 21180 11160 21232 11212
rect 19892 11135 19944 11144
rect 19892 11101 19901 11135
rect 19901 11101 19935 11135
rect 19935 11101 19944 11135
rect 19892 11092 19944 11101
rect 16672 11024 16724 11076
rect 17776 11024 17828 11076
rect 18328 11024 18380 11076
rect 19248 11024 19300 11076
rect 19708 11024 19760 11076
rect 20352 11024 20404 11076
rect 20720 11098 20726 11122
rect 20726 11098 20760 11122
rect 20760 11098 20772 11122
rect 20720 11070 20772 11098
rect 20812 11129 20864 11138
rect 20812 11095 20821 11129
rect 20821 11095 20855 11129
rect 20855 11095 20864 11129
rect 20812 11086 20864 11095
rect 20996 11135 21048 11144
rect 20996 11101 21005 11135
rect 21005 11101 21039 11135
rect 21039 11101 21048 11135
rect 20996 11092 21048 11101
rect 21640 11024 21692 11076
rect 21824 11135 21876 11144
rect 21824 11101 21833 11135
rect 21833 11101 21867 11135
rect 21867 11101 21876 11135
rect 21824 11092 21876 11101
rect 15568 10956 15620 11008
rect 15752 10956 15804 11008
rect 16488 10956 16540 11008
rect 19156 10956 19208 11008
rect 20536 10956 20588 11008
rect 6630 10854 6682 10906
rect 6694 10854 6746 10906
rect 6758 10854 6810 10906
rect 6822 10854 6874 10906
rect 6886 10854 6938 10906
rect 12311 10854 12363 10906
rect 12375 10854 12427 10906
rect 12439 10854 12491 10906
rect 12503 10854 12555 10906
rect 12567 10854 12619 10906
rect 17992 10854 18044 10906
rect 18056 10854 18108 10906
rect 18120 10854 18172 10906
rect 18184 10854 18236 10906
rect 18248 10854 18300 10906
rect 23673 10854 23725 10906
rect 23737 10854 23789 10906
rect 23801 10854 23853 10906
rect 23865 10854 23917 10906
rect 23929 10854 23981 10906
rect 2872 10752 2924 10804
rect 3700 10752 3752 10804
rect 1584 10616 1636 10668
rect 2228 10616 2280 10668
rect 2780 10616 2832 10668
rect 3608 10684 3660 10736
rect 5632 10752 5684 10804
rect 6552 10795 6604 10804
rect 6552 10761 6561 10795
rect 6561 10761 6595 10795
rect 6595 10761 6604 10795
rect 6552 10752 6604 10761
rect 8484 10795 8536 10804
rect 8484 10761 8493 10795
rect 8493 10761 8527 10795
rect 8527 10761 8536 10795
rect 8484 10752 8536 10761
rect 8944 10752 8996 10804
rect 9312 10752 9364 10804
rect 3056 10659 3108 10668
rect 3056 10625 3070 10659
rect 3070 10625 3104 10659
rect 3104 10625 3108 10659
rect 3056 10616 3108 10625
rect 3700 10616 3752 10668
rect 4620 10684 4672 10736
rect 8576 10684 8628 10736
rect 4528 10616 4580 10668
rect 4804 10616 4856 10668
rect 2964 10480 3016 10532
rect 6092 10616 6144 10668
rect 6276 10616 6328 10668
rect 8024 10659 8076 10668
rect 3240 10523 3292 10532
rect 3240 10489 3249 10523
rect 3249 10489 3283 10523
rect 3283 10489 3292 10523
rect 3240 10480 3292 10489
rect 3516 10480 3568 10532
rect 7196 10548 7248 10600
rect 8024 10625 8033 10659
rect 8033 10625 8067 10659
rect 8067 10625 8076 10659
rect 8024 10616 8076 10625
rect 8760 10659 8812 10668
rect 8760 10625 8769 10659
rect 8769 10625 8803 10659
rect 8803 10625 8812 10659
rect 8760 10616 8812 10625
rect 8392 10548 8444 10600
rect 8944 10659 8996 10668
rect 8944 10625 8953 10659
rect 8953 10625 8987 10659
rect 8987 10625 8996 10659
rect 8944 10616 8996 10625
rect 9404 10616 9456 10668
rect 1952 10455 2004 10464
rect 1952 10421 1961 10455
rect 1961 10421 1995 10455
rect 1995 10421 2004 10455
rect 1952 10412 2004 10421
rect 2504 10412 2556 10464
rect 3148 10412 3200 10464
rect 4252 10412 4304 10464
rect 4988 10412 5040 10464
rect 9312 10480 9364 10532
rect 9864 10591 9916 10600
rect 9864 10557 9873 10591
rect 9873 10557 9907 10591
rect 9907 10557 9916 10591
rect 9864 10548 9916 10557
rect 11152 10752 11204 10804
rect 11888 10752 11940 10804
rect 13084 10795 13136 10804
rect 13084 10761 13093 10795
rect 13093 10761 13127 10795
rect 13127 10761 13136 10795
rect 13084 10752 13136 10761
rect 13544 10752 13596 10804
rect 14372 10752 14424 10804
rect 16120 10752 16172 10804
rect 17592 10752 17644 10804
rect 18420 10752 18472 10804
rect 19340 10752 19392 10804
rect 20444 10752 20496 10804
rect 20536 10795 20588 10804
rect 20536 10761 20545 10795
rect 20545 10761 20579 10795
rect 20579 10761 20588 10795
rect 20536 10752 20588 10761
rect 20996 10752 21048 10804
rect 10968 10684 11020 10736
rect 11428 10616 11480 10668
rect 12808 10616 12860 10668
rect 13728 10684 13780 10736
rect 15292 10727 15344 10736
rect 15292 10693 15301 10727
rect 15301 10693 15335 10727
rect 15335 10693 15344 10727
rect 15292 10684 15344 10693
rect 15568 10684 15620 10736
rect 16948 10684 17000 10736
rect 14648 10659 14700 10668
rect 11060 10523 11112 10532
rect 11060 10489 11069 10523
rect 11069 10489 11103 10523
rect 11103 10489 11112 10523
rect 11060 10480 11112 10489
rect 11704 10480 11756 10532
rect 14648 10625 14657 10659
rect 14657 10625 14691 10659
rect 14691 10625 14700 10659
rect 14648 10616 14700 10625
rect 15844 10616 15896 10668
rect 16120 10659 16172 10668
rect 16120 10625 16129 10659
rect 16129 10625 16163 10659
rect 16163 10625 16172 10659
rect 16120 10616 16172 10625
rect 13912 10548 13964 10600
rect 17500 10616 17552 10668
rect 5724 10412 5776 10464
rect 6000 10412 6052 10464
rect 8208 10412 8260 10464
rect 10048 10412 10100 10464
rect 12348 10412 12400 10464
rect 13820 10412 13872 10464
rect 16672 10548 16724 10600
rect 17224 10548 17276 10600
rect 15844 10480 15896 10532
rect 14096 10412 14148 10464
rect 14556 10455 14608 10464
rect 14556 10421 14565 10455
rect 14565 10421 14599 10455
rect 14599 10421 14608 10455
rect 14556 10412 14608 10421
rect 15016 10412 15068 10464
rect 18420 10659 18472 10668
rect 18420 10625 18429 10659
rect 18429 10625 18463 10659
rect 18463 10625 18472 10659
rect 19432 10684 19484 10736
rect 18420 10616 18472 10625
rect 18788 10616 18840 10668
rect 19340 10616 19392 10668
rect 19892 10684 19944 10736
rect 20628 10659 20680 10668
rect 18880 10548 18932 10600
rect 19708 10591 19760 10600
rect 19708 10557 19717 10591
rect 19717 10557 19751 10591
rect 19751 10557 19760 10591
rect 19708 10548 19760 10557
rect 20628 10625 20637 10659
rect 20637 10625 20671 10659
rect 20671 10625 20680 10659
rect 20628 10616 20680 10625
rect 21364 10548 21416 10600
rect 18696 10412 18748 10464
rect 19432 10412 19484 10464
rect 21548 10480 21600 10532
rect 21456 10455 21508 10464
rect 21456 10421 21465 10455
rect 21465 10421 21499 10455
rect 21499 10421 21508 10455
rect 21456 10412 21508 10421
rect 3790 10310 3842 10362
rect 3854 10310 3906 10362
rect 3918 10310 3970 10362
rect 3982 10310 4034 10362
rect 4046 10310 4098 10362
rect 9471 10310 9523 10362
rect 9535 10310 9587 10362
rect 9599 10310 9651 10362
rect 9663 10310 9715 10362
rect 9727 10310 9779 10362
rect 15152 10310 15204 10362
rect 15216 10310 15268 10362
rect 15280 10310 15332 10362
rect 15344 10310 15396 10362
rect 15408 10310 15460 10362
rect 20833 10310 20885 10362
rect 20897 10310 20949 10362
rect 20961 10310 21013 10362
rect 21025 10310 21077 10362
rect 21089 10310 21141 10362
rect 2228 10251 2280 10260
rect 2228 10217 2237 10251
rect 2237 10217 2271 10251
rect 2271 10217 2280 10251
rect 2228 10208 2280 10217
rect 2412 10251 2464 10260
rect 2412 10217 2421 10251
rect 2421 10217 2455 10251
rect 2455 10217 2464 10251
rect 2412 10208 2464 10217
rect 3700 10208 3752 10260
rect 5080 10251 5132 10260
rect 5080 10217 5089 10251
rect 5089 10217 5123 10251
rect 5123 10217 5132 10251
rect 5080 10208 5132 10217
rect 5908 10251 5960 10260
rect 5908 10217 5917 10251
rect 5917 10217 5951 10251
rect 5951 10217 5960 10251
rect 5908 10208 5960 10217
rect 6184 10251 6236 10260
rect 6184 10217 6193 10251
rect 6193 10217 6227 10251
rect 6227 10217 6236 10251
rect 6184 10208 6236 10217
rect 8944 10208 8996 10260
rect 9128 10251 9180 10260
rect 9128 10217 9137 10251
rect 9137 10217 9171 10251
rect 9171 10217 9180 10251
rect 9128 10208 9180 10217
rect 4528 10140 4580 10192
rect 4620 10140 4672 10192
rect 3516 10072 3568 10124
rect 3332 10004 3384 10056
rect 4896 10072 4948 10124
rect 4988 10072 5040 10124
rect 7840 10140 7892 10192
rect 8024 10140 8076 10192
rect 5540 10072 5592 10124
rect 4252 10004 4304 10056
rect 5080 10047 5132 10056
rect 5080 10013 5089 10047
rect 5089 10013 5123 10047
rect 5123 10013 5132 10047
rect 5080 10004 5132 10013
rect 5816 10047 5868 10056
rect 5816 10013 5825 10047
rect 5825 10013 5859 10047
rect 5859 10013 5868 10047
rect 5816 10004 5868 10013
rect 4344 9979 4396 9988
rect 4344 9945 4353 9979
rect 4353 9945 4387 9979
rect 4387 9945 4396 9979
rect 4344 9936 4396 9945
rect 4988 9936 5040 9988
rect 4160 9868 4212 9920
rect 4804 9868 4856 9920
rect 6736 10047 6788 10056
rect 6736 10013 6745 10047
rect 6745 10013 6779 10047
rect 6779 10013 6788 10047
rect 6736 10004 6788 10013
rect 7748 10047 7800 10056
rect 7748 10013 7757 10047
rect 7757 10013 7791 10047
rect 7791 10013 7800 10047
rect 7748 10004 7800 10013
rect 6092 9868 6144 9920
rect 7472 9936 7524 9988
rect 7288 9868 7340 9920
rect 8484 10004 8536 10056
rect 8116 9979 8168 9988
rect 8116 9945 8125 9979
rect 8125 9945 8159 9979
rect 8159 9945 8168 9979
rect 8116 9936 8168 9945
rect 8484 9868 8536 9920
rect 9956 10208 10008 10260
rect 11704 10208 11756 10260
rect 12348 10208 12400 10260
rect 12716 10208 12768 10260
rect 9312 10140 9364 10192
rect 12532 10140 12584 10192
rect 11612 10115 11664 10124
rect 11612 10081 11621 10115
rect 11621 10081 11655 10115
rect 11655 10081 11664 10115
rect 11612 10072 11664 10081
rect 11704 10115 11756 10124
rect 11704 10081 11713 10115
rect 11713 10081 11747 10115
rect 11747 10081 11756 10115
rect 12624 10115 12676 10124
rect 11704 10072 11756 10081
rect 12624 10081 12633 10115
rect 12633 10081 12667 10115
rect 12667 10081 12676 10115
rect 12624 10072 12676 10081
rect 13176 10208 13228 10260
rect 13636 10251 13688 10260
rect 13636 10217 13645 10251
rect 13645 10217 13679 10251
rect 13679 10217 13688 10251
rect 13636 10208 13688 10217
rect 14648 10251 14700 10260
rect 14648 10217 14657 10251
rect 14657 10217 14691 10251
rect 14691 10217 14700 10251
rect 14648 10208 14700 10217
rect 18420 10208 18472 10260
rect 18604 10208 18656 10260
rect 19616 10251 19668 10260
rect 19616 10217 19625 10251
rect 19625 10217 19659 10251
rect 19659 10217 19668 10251
rect 19616 10208 19668 10217
rect 16672 10140 16724 10192
rect 20904 10251 20956 10260
rect 20904 10217 20913 10251
rect 20913 10217 20947 10251
rect 20947 10217 20956 10251
rect 20904 10208 20956 10217
rect 21180 10208 21232 10260
rect 12900 10115 12952 10124
rect 12900 10081 12909 10115
rect 12909 10081 12943 10115
rect 12943 10081 12952 10115
rect 12900 10072 12952 10081
rect 9312 10047 9364 10056
rect 9312 10013 9321 10047
rect 9321 10013 9355 10047
rect 9355 10013 9364 10047
rect 9312 10004 9364 10013
rect 9496 10047 9548 10056
rect 9496 10013 9505 10047
rect 9505 10013 9539 10047
rect 9539 10013 9548 10047
rect 9496 10004 9548 10013
rect 10968 10047 11020 10056
rect 9864 9936 9916 9988
rect 10968 10013 10977 10047
rect 10977 10013 11011 10047
rect 11011 10013 11020 10047
rect 10968 10004 11020 10013
rect 11520 10047 11572 10056
rect 11520 10013 11529 10047
rect 11529 10013 11563 10047
rect 11563 10013 11572 10047
rect 11520 10004 11572 10013
rect 11796 10047 11848 10056
rect 11796 10013 11805 10047
rect 11805 10013 11839 10047
rect 11839 10013 11848 10047
rect 11796 10004 11848 10013
rect 12532 10004 12584 10056
rect 13544 10072 13596 10124
rect 13636 10072 13688 10124
rect 14004 10004 14056 10056
rect 14280 10047 14332 10056
rect 14280 10013 14289 10047
rect 14289 10013 14323 10047
rect 14323 10013 14332 10047
rect 14280 10004 14332 10013
rect 15568 10047 15620 10056
rect 15568 10013 15575 10047
rect 15575 10013 15620 10047
rect 15568 10004 15620 10013
rect 16120 10072 16172 10124
rect 16396 10072 16448 10124
rect 17224 10072 17276 10124
rect 21272 10140 21324 10192
rect 19340 10072 19392 10124
rect 16764 10004 16816 10056
rect 18512 10004 18564 10056
rect 18696 10004 18748 10056
rect 20076 10072 20128 10124
rect 10048 9868 10100 9920
rect 10876 9868 10928 9920
rect 13820 9936 13872 9988
rect 15292 9936 15344 9988
rect 15660 9979 15712 9988
rect 15660 9945 15669 9979
rect 15669 9945 15703 9979
rect 15703 9945 15712 9979
rect 15660 9936 15712 9945
rect 16488 9979 16540 9988
rect 16488 9945 16497 9979
rect 16497 9945 16531 9979
rect 16531 9945 16540 9979
rect 16488 9936 16540 9945
rect 17132 9979 17184 9988
rect 17132 9945 17141 9979
rect 17141 9945 17175 9979
rect 17175 9945 17184 9979
rect 17132 9936 17184 9945
rect 17408 9979 17460 9988
rect 17408 9945 17417 9979
rect 17417 9945 17451 9979
rect 17451 9945 17460 9979
rect 17408 9936 17460 9945
rect 18880 9936 18932 9988
rect 19708 9936 19760 9988
rect 12532 9868 12584 9920
rect 12808 9868 12860 9920
rect 13636 9868 13688 9920
rect 16764 9868 16816 9920
rect 17224 9868 17276 9920
rect 17684 9868 17736 9920
rect 19432 9868 19484 9920
rect 20260 9936 20312 9988
rect 20444 9868 20496 9920
rect 21456 9868 21508 9920
rect 23112 9911 23164 9920
rect 23112 9877 23121 9911
rect 23121 9877 23155 9911
rect 23155 9877 23164 9911
rect 23112 9868 23164 9877
rect 6630 9766 6682 9818
rect 6694 9766 6746 9818
rect 6758 9766 6810 9818
rect 6822 9766 6874 9818
rect 6886 9766 6938 9818
rect 12311 9766 12363 9818
rect 12375 9766 12427 9818
rect 12439 9766 12491 9818
rect 12503 9766 12555 9818
rect 12567 9766 12619 9818
rect 17992 9766 18044 9818
rect 18056 9766 18108 9818
rect 18120 9766 18172 9818
rect 18184 9766 18236 9818
rect 18248 9766 18300 9818
rect 23673 9766 23725 9818
rect 23737 9766 23789 9818
rect 23801 9766 23853 9818
rect 23865 9766 23917 9818
rect 23929 9766 23981 9818
rect 1952 9707 2004 9716
rect 1952 9673 1961 9707
rect 1961 9673 1995 9707
rect 1995 9673 2004 9707
rect 1952 9664 2004 9673
rect 4252 9664 4304 9716
rect 5816 9664 5868 9716
rect 7288 9664 7340 9716
rect 11428 9664 11480 9716
rect 11612 9664 11664 9716
rect 12624 9664 12676 9716
rect 12992 9664 13044 9716
rect 13176 9664 13228 9716
rect 13360 9664 13412 9716
rect 13912 9664 13964 9716
rect 15568 9664 15620 9716
rect 15752 9664 15804 9716
rect 16120 9664 16172 9716
rect 17408 9664 17460 9716
rect 2780 9596 2832 9648
rect 3516 9596 3568 9648
rect 6460 9596 6512 9648
rect 2596 9571 2648 9580
rect 2596 9537 2605 9571
rect 2605 9537 2639 9571
rect 2639 9537 2648 9571
rect 4344 9571 4396 9580
rect 2596 9528 2648 9537
rect 1952 9460 2004 9512
rect 4344 9537 4353 9571
rect 4353 9537 4387 9571
rect 4387 9537 4396 9571
rect 4344 9528 4396 9537
rect 4988 9528 5040 9580
rect 5724 9528 5776 9580
rect 6828 9528 6880 9580
rect 7748 9596 7800 9648
rect 10232 9596 10284 9648
rect 11060 9596 11112 9648
rect 7288 9571 7340 9580
rect 7288 9537 7297 9571
rect 7297 9537 7331 9571
rect 7331 9537 7340 9571
rect 7288 9528 7340 9537
rect 7380 9528 7432 9580
rect 10048 9528 10100 9580
rect 10324 9571 10376 9580
rect 10324 9537 10333 9571
rect 10333 9537 10367 9571
rect 10367 9537 10376 9571
rect 10324 9528 10376 9537
rect 11612 9528 11664 9580
rect 12440 9528 12492 9580
rect 14556 9596 14608 9648
rect 18236 9664 18288 9716
rect 18604 9664 18656 9716
rect 19432 9664 19484 9716
rect 12992 9571 13044 9580
rect 12992 9537 13001 9571
rect 13001 9537 13035 9571
rect 13035 9537 13044 9571
rect 12992 9528 13044 9537
rect 5080 9460 5132 9512
rect 6368 9460 6420 9512
rect 3240 9392 3292 9444
rect 5264 9392 5316 9444
rect 8116 9460 8168 9512
rect 10508 9503 10560 9512
rect 10508 9469 10517 9503
rect 10517 9469 10551 9503
rect 10551 9469 10560 9503
rect 10508 9460 10560 9469
rect 10968 9460 11020 9512
rect 11980 9460 12032 9512
rect 3056 9324 3108 9376
rect 3700 9324 3752 9376
rect 4252 9324 4304 9376
rect 7012 9392 7064 9444
rect 13544 9528 13596 9580
rect 14648 9571 14700 9580
rect 14648 9537 14657 9571
rect 14657 9537 14691 9571
rect 14691 9537 14700 9571
rect 14648 9528 14700 9537
rect 17592 9596 17644 9648
rect 15384 9528 15436 9580
rect 6552 9367 6604 9376
rect 6552 9333 6561 9367
rect 6561 9333 6595 9367
rect 6595 9333 6604 9367
rect 6552 9324 6604 9333
rect 7564 9324 7616 9376
rect 7840 9367 7892 9376
rect 7840 9333 7849 9367
rect 7849 9333 7883 9367
rect 7883 9333 7892 9367
rect 7840 9324 7892 9333
rect 8852 9324 8904 9376
rect 9404 9324 9456 9376
rect 9864 9324 9916 9376
rect 10600 9324 10652 9376
rect 11888 9367 11940 9376
rect 11888 9333 11897 9367
rect 11897 9333 11931 9367
rect 11931 9333 11940 9367
rect 11888 9324 11940 9333
rect 11980 9367 12032 9376
rect 11980 9333 11989 9367
rect 11989 9333 12023 9367
rect 12023 9333 12032 9367
rect 14648 9392 14700 9444
rect 11980 9324 12032 9333
rect 13360 9324 13412 9376
rect 13912 9367 13964 9376
rect 13912 9333 13921 9367
rect 13921 9333 13955 9367
rect 13955 9333 13964 9367
rect 13912 9324 13964 9333
rect 14740 9324 14792 9376
rect 15752 9435 15804 9444
rect 15752 9401 15761 9435
rect 15761 9401 15795 9435
rect 15795 9401 15804 9435
rect 15752 9392 15804 9401
rect 15936 9503 15988 9512
rect 15936 9469 15945 9503
rect 15945 9469 15979 9503
rect 15979 9469 15988 9503
rect 16120 9537 16129 9542
rect 16129 9537 16163 9542
rect 16163 9537 16172 9542
rect 16120 9490 16172 9537
rect 17868 9571 17920 9580
rect 15936 9460 15988 9469
rect 16488 9460 16540 9512
rect 17224 9460 17276 9512
rect 17868 9537 17877 9571
rect 17877 9537 17911 9571
rect 17911 9537 17920 9571
rect 17868 9528 17920 9537
rect 17960 9528 18012 9580
rect 18420 9596 18472 9648
rect 18328 9528 18380 9580
rect 18604 9528 18656 9580
rect 19156 9528 19208 9580
rect 20444 9639 20496 9648
rect 19248 9460 19300 9512
rect 16396 9392 16448 9444
rect 16580 9392 16632 9444
rect 17592 9392 17644 9444
rect 19340 9392 19392 9444
rect 20444 9605 20453 9639
rect 20453 9605 20487 9639
rect 20487 9605 20496 9639
rect 20444 9596 20496 9605
rect 19892 9528 19944 9580
rect 20352 9571 20404 9580
rect 20352 9537 20359 9571
rect 20359 9537 20404 9571
rect 20076 9460 20128 9512
rect 20352 9528 20404 9537
rect 20536 9571 20588 9580
rect 20536 9537 20545 9571
rect 20545 9537 20579 9571
rect 20579 9537 20588 9571
rect 20536 9528 20588 9537
rect 21180 9528 21232 9580
rect 22192 9528 22244 9580
rect 23020 9571 23072 9580
rect 23020 9537 23029 9571
rect 23029 9537 23063 9571
rect 23063 9537 23072 9571
rect 23020 9528 23072 9537
rect 20444 9392 20496 9444
rect 20720 9392 20772 9444
rect 21732 9460 21784 9512
rect 22468 9460 22520 9512
rect 22376 9392 22428 9444
rect 18604 9367 18656 9376
rect 18604 9333 18613 9367
rect 18613 9333 18647 9367
rect 18647 9333 18656 9367
rect 18604 9324 18656 9333
rect 19248 9324 19300 9376
rect 19616 9324 19668 9376
rect 21180 9324 21232 9376
rect 21456 9324 21508 9376
rect 22192 9367 22244 9376
rect 22192 9333 22201 9367
rect 22201 9333 22235 9367
rect 22235 9333 22244 9367
rect 22192 9324 22244 9333
rect 3790 9222 3842 9274
rect 3854 9222 3906 9274
rect 3918 9222 3970 9274
rect 3982 9222 4034 9274
rect 4046 9222 4098 9274
rect 9471 9222 9523 9274
rect 9535 9222 9587 9274
rect 9599 9222 9651 9274
rect 9663 9222 9715 9274
rect 9727 9222 9779 9274
rect 15152 9222 15204 9274
rect 15216 9222 15268 9274
rect 15280 9222 15332 9274
rect 15344 9222 15396 9274
rect 15408 9222 15460 9274
rect 20833 9222 20885 9274
rect 20897 9222 20949 9274
rect 20961 9222 21013 9274
rect 21025 9222 21077 9274
rect 21089 9222 21141 9274
rect 3424 9120 3476 9172
rect 3976 9120 4028 9172
rect 5632 9120 5684 9172
rect 5908 9120 5960 9172
rect 6368 9163 6420 9172
rect 6368 9129 6377 9163
rect 6377 9129 6411 9163
rect 6411 9129 6420 9163
rect 6368 9120 6420 9129
rect 1584 9052 1636 9104
rect 2688 9052 2740 9104
rect 2872 9052 2924 9104
rect 2964 9027 3016 9036
rect 2964 8993 2973 9027
rect 2973 8993 3007 9027
rect 3007 8993 3016 9027
rect 2964 8984 3016 8993
rect 4988 9052 5040 9104
rect 6828 9120 6880 9172
rect 7196 9120 7248 9172
rect 8668 9120 8720 9172
rect 11244 9163 11296 9172
rect 11244 9129 11253 9163
rect 11253 9129 11287 9163
rect 11287 9129 11296 9163
rect 11244 9120 11296 9129
rect 11980 9120 12032 9172
rect 6644 9052 6696 9104
rect 6920 9052 6972 9104
rect 3516 8984 3568 9036
rect 2044 8916 2096 8968
rect 2872 8959 2924 8968
rect 2872 8925 2881 8959
rect 2881 8925 2915 8959
rect 2915 8925 2924 8959
rect 2872 8916 2924 8925
rect 3056 8959 3108 8968
rect 3056 8925 3065 8959
rect 3065 8925 3099 8959
rect 3099 8925 3108 8959
rect 3056 8916 3108 8925
rect 3240 8959 3292 8968
rect 3240 8925 3249 8959
rect 3249 8925 3283 8959
rect 3283 8925 3292 8959
rect 3240 8916 3292 8925
rect 4344 8916 4396 8968
rect 5264 8959 5316 8968
rect 3792 8848 3844 8900
rect 5264 8925 5273 8959
rect 5273 8925 5307 8959
rect 5307 8925 5316 8959
rect 5264 8916 5316 8925
rect 5724 8916 5776 8968
rect 6368 8916 6420 8968
rect 8392 8959 8444 8968
rect 8392 8925 8401 8959
rect 8401 8925 8435 8959
rect 8435 8925 8444 8959
rect 8392 8916 8444 8925
rect 11888 9052 11940 9104
rect 9496 8959 9548 8968
rect 9496 8925 9505 8959
rect 9505 8925 9539 8959
rect 9539 8925 9548 8959
rect 9496 8916 9548 8925
rect 10324 8916 10376 8968
rect 11428 8959 11480 8968
rect 11428 8925 11437 8959
rect 11437 8925 11471 8959
rect 11471 8925 11480 8959
rect 11428 8916 11480 8925
rect 12624 8984 12676 9036
rect 7012 8848 7064 8900
rect 10048 8848 10100 8900
rect 12164 8916 12216 8968
rect 13268 9052 13320 9104
rect 13912 9052 13964 9104
rect 1952 8780 2004 8832
rect 2596 8780 2648 8832
rect 4620 8780 4672 8832
rect 4896 8780 4948 8832
rect 6920 8780 6972 8832
rect 9956 8780 10008 8832
rect 10600 8823 10652 8832
rect 10600 8789 10609 8823
rect 10609 8789 10643 8823
rect 10643 8789 10652 8823
rect 10600 8780 10652 8789
rect 12256 8780 12308 8832
rect 12808 8780 12860 8832
rect 14188 9120 14240 9172
rect 14924 9120 14976 9172
rect 15752 9120 15804 9172
rect 16212 9120 16264 9172
rect 16304 9120 16356 9172
rect 17868 9120 17920 9172
rect 20352 9120 20404 9172
rect 20536 9120 20588 9172
rect 22008 9120 22060 9172
rect 16488 9052 16540 9104
rect 14464 9027 14516 9036
rect 13544 8959 13596 8968
rect 13544 8925 13568 8959
rect 13568 8925 13596 8959
rect 13544 8916 13596 8925
rect 14464 8993 14473 9027
rect 14473 8993 14507 9027
rect 14507 8993 14516 9027
rect 14464 8984 14516 8993
rect 14740 9027 14792 9036
rect 14740 8993 14749 9027
rect 14749 8993 14783 9027
rect 14783 8993 14792 9027
rect 14740 8984 14792 8993
rect 13912 8916 13964 8968
rect 14556 8959 14608 8968
rect 14556 8925 14566 8959
rect 14566 8925 14600 8959
rect 14600 8925 14608 8959
rect 14556 8916 14608 8925
rect 16672 9027 16724 9036
rect 16672 8993 16681 9027
rect 16681 8993 16715 9027
rect 16715 8993 16724 9027
rect 16672 8984 16724 8993
rect 16580 8959 16632 8968
rect 14832 8848 14884 8900
rect 14648 8780 14700 8832
rect 16580 8925 16589 8959
rect 16589 8925 16623 8959
rect 16623 8925 16632 8959
rect 16580 8916 16632 8925
rect 20996 9052 21048 9104
rect 17500 8916 17552 8968
rect 18512 8984 18564 9036
rect 18696 8984 18748 9036
rect 16488 8848 16540 8900
rect 17868 8925 17877 8946
rect 17877 8925 17911 8946
rect 17911 8925 17920 8946
rect 17868 8894 17920 8925
rect 19616 8916 19668 8968
rect 20444 8984 20496 9036
rect 21640 8984 21692 9036
rect 20536 8916 20588 8968
rect 20720 8959 20772 8968
rect 20720 8925 20729 8959
rect 20729 8925 20763 8959
rect 20763 8925 20772 8959
rect 20720 8916 20772 8925
rect 17776 8780 17828 8832
rect 18512 8823 18564 8832
rect 18512 8789 18521 8823
rect 18521 8789 18555 8823
rect 18555 8789 18564 8823
rect 18512 8780 18564 8789
rect 18696 8823 18748 8832
rect 18696 8789 18723 8823
rect 18723 8789 18748 8823
rect 18696 8780 18748 8789
rect 19892 8848 19944 8900
rect 20168 8848 20220 8900
rect 22284 8916 22336 8968
rect 23020 8916 23072 8968
rect 18972 8780 19024 8832
rect 19340 8780 19392 8832
rect 20536 8780 20588 8832
rect 20720 8780 20772 8832
rect 21180 8780 21232 8832
rect 21640 8823 21692 8832
rect 21640 8789 21649 8823
rect 21649 8789 21683 8823
rect 21683 8789 21692 8823
rect 21640 8780 21692 8789
rect 22100 8780 22152 8832
rect 22560 8780 22612 8832
rect 22836 8823 22888 8832
rect 22836 8789 22845 8823
rect 22845 8789 22879 8823
rect 22879 8789 22888 8823
rect 22836 8780 22888 8789
rect 6630 8678 6682 8730
rect 6694 8678 6746 8730
rect 6758 8678 6810 8730
rect 6822 8678 6874 8730
rect 6886 8678 6938 8730
rect 12311 8678 12363 8730
rect 12375 8678 12427 8730
rect 12439 8678 12491 8730
rect 12503 8678 12555 8730
rect 12567 8678 12619 8730
rect 17992 8678 18044 8730
rect 18056 8678 18108 8730
rect 18120 8678 18172 8730
rect 18184 8678 18236 8730
rect 18248 8678 18300 8730
rect 23673 8678 23725 8730
rect 23737 8678 23789 8730
rect 23801 8678 23853 8730
rect 23865 8678 23917 8730
rect 23929 8678 23981 8730
rect 2044 8619 2096 8628
rect 2044 8585 2053 8619
rect 2053 8585 2087 8619
rect 2087 8585 2096 8619
rect 2044 8576 2096 8585
rect 2688 8576 2740 8628
rect 3792 8576 3844 8628
rect 4712 8576 4764 8628
rect 5264 8576 5316 8628
rect 5356 8576 5408 8628
rect 7012 8576 7064 8628
rect 7104 8576 7156 8628
rect 8760 8576 8812 8628
rect 10232 8576 10284 8628
rect 2780 8508 2832 8560
rect 2320 8440 2372 8492
rect 2596 8440 2648 8492
rect 3240 8440 3292 8492
rect 3608 8440 3660 8492
rect 3976 8483 4028 8492
rect 3976 8449 3985 8483
rect 3985 8449 4019 8483
rect 4019 8449 4028 8483
rect 3976 8440 4028 8449
rect 4344 8440 4396 8492
rect 4896 8440 4948 8492
rect 7288 8508 7340 8560
rect 9864 8508 9916 8560
rect 2504 8415 2556 8424
rect 2504 8381 2513 8415
rect 2513 8381 2547 8415
rect 2547 8381 2556 8415
rect 2504 8372 2556 8381
rect 5540 8440 5592 8492
rect 7380 8440 7432 8492
rect 7564 8483 7616 8492
rect 7564 8449 7573 8483
rect 7573 8449 7607 8483
rect 7607 8449 7616 8483
rect 7564 8440 7616 8449
rect 7656 8483 7708 8492
rect 7656 8449 7665 8483
rect 7665 8449 7699 8483
rect 7699 8449 7708 8483
rect 7656 8440 7708 8449
rect 7840 8483 7892 8492
rect 7840 8449 7875 8483
rect 7875 8449 7892 8483
rect 8024 8483 8076 8492
rect 7840 8440 7892 8449
rect 8024 8449 8033 8483
rect 8033 8449 8067 8483
rect 8067 8449 8076 8483
rect 8024 8440 8076 8449
rect 8484 8483 8536 8492
rect 3700 8304 3752 8356
rect 5080 8304 5132 8356
rect 7012 8372 7064 8424
rect 8484 8449 8485 8483
rect 8485 8449 8519 8483
rect 8519 8449 8536 8483
rect 8484 8440 8536 8449
rect 8668 8440 8720 8492
rect 8944 8440 8996 8492
rect 10048 8508 10100 8560
rect 10416 8508 10468 8560
rect 12164 8576 12216 8628
rect 11612 8508 11664 8560
rect 11888 8508 11940 8560
rect 12072 8508 12124 8560
rect 12532 8551 12584 8560
rect 12532 8517 12541 8551
rect 12541 8517 12575 8551
rect 12575 8517 12584 8551
rect 12532 8508 12584 8517
rect 12992 8576 13044 8628
rect 14464 8576 14516 8628
rect 16028 8576 16080 8628
rect 16488 8576 16540 8628
rect 16580 8576 16632 8628
rect 12900 8440 12952 8492
rect 13636 8483 13688 8492
rect 13636 8449 13645 8483
rect 13645 8449 13679 8483
rect 13679 8449 13688 8483
rect 13636 8440 13688 8449
rect 13084 8372 13136 8424
rect 13176 8304 13228 8356
rect 1860 8236 1912 8288
rect 6368 8236 6420 8288
rect 7196 8236 7248 8288
rect 7656 8236 7708 8288
rect 9128 8279 9180 8288
rect 9128 8245 9137 8279
rect 9137 8245 9171 8279
rect 9171 8245 9180 8279
rect 9128 8236 9180 8245
rect 9312 8236 9364 8288
rect 9496 8236 9548 8288
rect 10416 8236 10468 8288
rect 12716 8236 12768 8288
rect 13544 8279 13596 8288
rect 13544 8245 13553 8279
rect 13553 8245 13587 8279
rect 13587 8245 13596 8279
rect 13544 8236 13596 8245
rect 14464 8440 14516 8492
rect 15752 8440 15804 8492
rect 14556 8372 14608 8424
rect 14832 8372 14884 8424
rect 14924 8304 14976 8356
rect 15476 8372 15528 8424
rect 16120 8440 16172 8492
rect 17316 8508 17368 8560
rect 17224 8483 17276 8492
rect 17224 8449 17233 8483
rect 17233 8449 17267 8483
rect 17267 8449 17276 8483
rect 17224 8440 17276 8449
rect 17684 8440 17736 8492
rect 18328 8576 18380 8628
rect 18696 8576 18748 8628
rect 20352 8576 20404 8628
rect 20628 8576 20680 8628
rect 22008 8576 22060 8628
rect 22284 8576 22336 8628
rect 22468 8619 22520 8628
rect 22468 8585 22477 8619
rect 22477 8585 22511 8619
rect 22511 8585 22520 8619
rect 22468 8576 22520 8585
rect 23020 8576 23072 8628
rect 18420 8508 18472 8560
rect 18236 8483 18288 8492
rect 18236 8449 18245 8483
rect 18245 8449 18279 8483
rect 18279 8449 18288 8483
rect 18236 8440 18288 8449
rect 18788 8440 18840 8492
rect 19524 8440 19576 8492
rect 22836 8508 22888 8560
rect 19892 8483 19944 8492
rect 19892 8449 19901 8483
rect 19901 8449 19935 8483
rect 19935 8449 19944 8483
rect 19892 8440 19944 8449
rect 20076 8483 20128 8492
rect 20076 8449 20085 8483
rect 20085 8449 20119 8483
rect 20119 8449 20128 8483
rect 20720 8483 20772 8492
rect 20076 8440 20128 8449
rect 20720 8449 20729 8483
rect 20729 8449 20763 8483
rect 20763 8449 20772 8483
rect 20720 8440 20772 8449
rect 20996 8483 21048 8492
rect 18420 8372 18472 8424
rect 17224 8304 17276 8356
rect 18236 8304 18288 8356
rect 14740 8236 14792 8288
rect 16304 8236 16356 8288
rect 18052 8236 18104 8288
rect 18972 8372 19024 8424
rect 20628 8372 20680 8424
rect 20996 8449 21005 8483
rect 21005 8449 21039 8483
rect 21039 8449 21048 8483
rect 20996 8440 21048 8449
rect 21640 8440 21692 8492
rect 21732 8440 21784 8492
rect 22376 8440 22428 8492
rect 21364 8372 21416 8424
rect 20812 8304 20864 8356
rect 19340 8236 19392 8288
rect 21088 8236 21140 8288
rect 22008 8304 22060 8356
rect 22192 8304 22244 8356
rect 22560 8236 22612 8288
rect 23020 8236 23072 8288
rect 3790 8134 3842 8186
rect 3854 8134 3906 8186
rect 3918 8134 3970 8186
rect 3982 8134 4034 8186
rect 4046 8134 4098 8186
rect 9471 8134 9523 8186
rect 9535 8134 9587 8186
rect 9599 8134 9651 8186
rect 9663 8134 9715 8186
rect 9727 8134 9779 8186
rect 15152 8134 15204 8186
rect 15216 8134 15268 8186
rect 15280 8134 15332 8186
rect 15344 8134 15396 8186
rect 15408 8134 15460 8186
rect 20833 8134 20885 8186
rect 20897 8134 20949 8186
rect 20961 8134 21013 8186
rect 21025 8134 21077 8186
rect 21089 8134 21141 8186
rect 1952 8032 2004 8084
rect 2872 8032 2924 8084
rect 3516 8032 3568 8084
rect 4344 8032 4396 8084
rect 5172 8032 5224 8084
rect 6460 8032 6512 8084
rect 2320 7871 2372 7880
rect 2320 7837 2345 7871
rect 2345 7837 2372 7871
rect 2320 7828 2372 7837
rect 2780 7964 2832 8016
rect 4712 8007 4764 8016
rect 4712 7973 4721 8007
rect 4721 7973 4755 8007
rect 4755 7973 4764 8007
rect 4712 7964 4764 7973
rect 6276 7964 6328 8016
rect 7564 8032 7616 8084
rect 9864 8032 9916 8084
rect 10784 8032 10836 8084
rect 13360 8032 13412 8084
rect 14648 8075 14700 8084
rect 14648 8041 14657 8075
rect 14657 8041 14691 8075
rect 14691 8041 14700 8075
rect 14648 8032 14700 8041
rect 15752 8075 15804 8084
rect 15752 8041 15761 8075
rect 15761 8041 15795 8075
rect 15795 8041 15804 8075
rect 15752 8032 15804 8041
rect 16488 8032 16540 8084
rect 17776 8075 17828 8084
rect 17776 8041 17785 8075
rect 17785 8041 17819 8075
rect 17819 8041 17828 8075
rect 17776 8032 17828 8041
rect 18788 8032 18840 8084
rect 19892 8032 19944 8084
rect 20260 8075 20312 8084
rect 20260 8041 20269 8075
rect 20269 8041 20303 8075
rect 20303 8041 20312 8075
rect 20260 8032 20312 8041
rect 4252 7896 4304 7948
rect 5632 7896 5684 7948
rect 2504 7871 2556 7880
rect 2504 7837 2513 7871
rect 2513 7837 2547 7871
rect 2547 7837 2556 7871
rect 2504 7828 2556 7837
rect 2688 7828 2740 7880
rect 3516 7828 3568 7880
rect 6000 7828 6052 7880
rect 6368 7896 6420 7948
rect 6552 7939 6604 7948
rect 6552 7905 6561 7939
rect 6561 7905 6595 7939
rect 6595 7905 6604 7939
rect 6552 7896 6604 7905
rect 6460 7871 6512 7880
rect 6460 7837 6469 7871
rect 6469 7837 6503 7871
rect 6503 7837 6512 7871
rect 6460 7828 6512 7837
rect 7196 7871 7248 7880
rect 7196 7837 7205 7871
rect 7205 7837 7239 7871
rect 7239 7837 7248 7871
rect 7196 7828 7248 7837
rect 5632 7760 5684 7812
rect 7656 7828 7708 7880
rect 11152 7964 11204 8016
rect 11520 7964 11572 8016
rect 16028 7964 16080 8016
rect 7932 7828 7984 7880
rect 8208 7871 8260 7880
rect 8208 7837 8217 7871
rect 8217 7837 8251 7871
rect 8251 7837 8260 7871
rect 8208 7828 8260 7837
rect 8392 7871 8444 7880
rect 8392 7837 8401 7871
rect 8401 7837 8435 7871
rect 8435 7837 8444 7871
rect 10416 7896 10468 7948
rect 12164 7896 12216 7948
rect 12900 7896 12952 7948
rect 14556 7896 14608 7948
rect 8392 7828 8444 7837
rect 8760 7760 8812 7812
rect 10048 7828 10100 7880
rect 10600 7828 10652 7880
rect 11796 7828 11848 7880
rect 11888 7871 11940 7880
rect 11888 7837 11897 7871
rect 11897 7837 11931 7871
rect 11931 7837 11940 7871
rect 11888 7828 11940 7837
rect 13360 7871 13412 7880
rect 11704 7803 11756 7812
rect 7288 7692 7340 7744
rect 7656 7692 7708 7744
rect 11704 7769 11713 7803
rect 11713 7769 11747 7803
rect 11747 7769 11756 7803
rect 11704 7760 11756 7769
rect 9588 7692 9640 7744
rect 13360 7837 13369 7871
rect 13369 7837 13403 7871
rect 13403 7837 13412 7871
rect 13360 7828 13412 7837
rect 13452 7871 13504 7880
rect 13452 7837 13461 7871
rect 13461 7837 13495 7871
rect 13495 7837 13504 7871
rect 15108 7896 15160 7948
rect 13452 7828 13504 7837
rect 14924 7871 14976 7880
rect 14924 7837 14933 7871
rect 14933 7837 14967 7871
rect 14967 7837 14976 7871
rect 14924 7828 14976 7837
rect 14372 7760 14424 7812
rect 14740 7760 14792 7812
rect 15384 7760 15436 7812
rect 15660 7760 15712 7812
rect 15936 7871 15988 7880
rect 15936 7837 15945 7871
rect 15945 7837 15979 7871
rect 15979 7837 15988 7871
rect 16856 8007 16908 8016
rect 16856 7973 16865 8007
rect 16865 7973 16899 8007
rect 16899 7973 16908 8007
rect 16856 7964 16908 7973
rect 15936 7828 15988 7837
rect 16212 7866 16264 7918
rect 16948 7896 17000 7948
rect 16304 7871 16356 7880
rect 16304 7837 16313 7871
rect 16313 7837 16347 7871
rect 16347 7837 16356 7871
rect 16304 7828 16356 7837
rect 16856 7828 16908 7880
rect 16212 7760 16264 7812
rect 22284 7964 22336 8016
rect 14004 7692 14056 7744
rect 14096 7692 14148 7744
rect 14924 7692 14976 7744
rect 16672 7692 16724 7744
rect 17684 7692 17736 7744
rect 18052 7871 18104 7880
rect 18052 7837 18061 7871
rect 18061 7837 18095 7871
rect 18095 7837 18104 7871
rect 19340 7896 19392 7948
rect 18052 7828 18104 7837
rect 18420 7828 18472 7880
rect 20168 7828 20220 7880
rect 18604 7760 18656 7812
rect 20536 7871 20588 7880
rect 20536 7837 20545 7871
rect 20545 7837 20579 7871
rect 20579 7837 20588 7871
rect 20536 7828 20588 7837
rect 20720 7760 20772 7812
rect 18328 7692 18380 7744
rect 19340 7692 19392 7744
rect 20352 7692 20404 7744
rect 21364 7828 21416 7880
rect 21732 7871 21784 7880
rect 21732 7837 21741 7871
rect 21741 7837 21775 7871
rect 21775 7837 21784 7871
rect 21732 7828 21784 7837
rect 22100 7760 22152 7812
rect 21640 7735 21692 7744
rect 21640 7701 21649 7735
rect 21649 7701 21683 7735
rect 21683 7701 21692 7735
rect 21640 7692 21692 7701
rect 22192 7692 22244 7744
rect 23020 7692 23072 7744
rect 6630 7590 6682 7642
rect 6694 7590 6746 7642
rect 6758 7590 6810 7642
rect 6822 7590 6874 7642
rect 6886 7590 6938 7642
rect 12311 7590 12363 7642
rect 12375 7590 12427 7642
rect 12439 7590 12491 7642
rect 12503 7590 12555 7642
rect 12567 7590 12619 7642
rect 17992 7590 18044 7642
rect 18056 7590 18108 7642
rect 18120 7590 18172 7642
rect 18184 7590 18236 7642
rect 18248 7590 18300 7642
rect 23673 7590 23725 7642
rect 23737 7590 23789 7642
rect 23801 7590 23853 7642
rect 23865 7590 23917 7642
rect 23929 7590 23981 7642
rect 3148 7488 3200 7540
rect 3240 7488 3292 7540
rect 2136 7420 2188 7472
rect 2688 7420 2740 7472
rect 5540 7488 5592 7540
rect 8116 7488 8168 7540
rect 8300 7488 8352 7540
rect 9312 7488 9364 7540
rect 6368 7420 6420 7472
rect 2412 7352 2464 7404
rect 2780 7395 2832 7404
rect 2780 7361 2789 7395
rect 2789 7361 2823 7395
rect 2823 7361 2832 7395
rect 2780 7352 2832 7361
rect 3516 7352 3568 7404
rect 4804 7395 4856 7404
rect 4804 7361 4813 7395
rect 4813 7361 4847 7395
rect 4847 7361 4856 7395
rect 4804 7352 4856 7361
rect 5356 7352 5408 7404
rect 5540 7352 5592 7404
rect 5724 7395 5776 7404
rect 5724 7361 5733 7395
rect 5733 7361 5767 7395
rect 5767 7361 5776 7395
rect 5724 7352 5776 7361
rect 5816 7395 5868 7404
rect 5816 7361 5825 7395
rect 5825 7361 5859 7395
rect 5859 7361 5868 7395
rect 5816 7352 5868 7361
rect 1860 7284 1912 7336
rect 2872 7284 2924 7336
rect 3056 7284 3108 7336
rect 6092 7284 6144 7336
rect 6368 7284 6420 7336
rect 7472 7352 7524 7404
rect 7932 7420 7984 7472
rect 8668 7420 8720 7472
rect 11704 7488 11756 7540
rect 12992 7531 13044 7540
rect 12992 7497 13001 7531
rect 13001 7497 13035 7531
rect 13035 7497 13044 7531
rect 12992 7488 13044 7497
rect 14004 7488 14056 7540
rect 15476 7488 15528 7540
rect 9312 7395 9364 7404
rect 7012 7327 7064 7336
rect 7012 7293 7043 7327
rect 7043 7293 7064 7327
rect 7012 7284 7064 7293
rect 7380 7284 7432 7336
rect 9312 7361 9321 7395
rect 9321 7361 9355 7395
rect 9355 7361 9364 7395
rect 9312 7352 9364 7361
rect 9588 7352 9640 7404
rect 11244 7420 11296 7472
rect 11980 7463 12032 7472
rect 11980 7429 11989 7463
rect 11989 7429 12023 7463
rect 12023 7429 12032 7463
rect 11980 7420 12032 7429
rect 13360 7420 13412 7472
rect 13544 7420 13596 7472
rect 15384 7420 15436 7472
rect 11152 7395 11204 7404
rect 7932 7284 7984 7336
rect 11152 7361 11161 7395
rect 11161 7361 11195 7395
rect 11195 7361 11204 7395
rect 11152 7352 11204 7361
rect 10416 7284 10468 7336
rect 12164 7352 12216 7404
rect 12900 7352 12952 7404
rect 13728 7352 13780 7404
rect 14188 7395 14240 7404
rect 14188 7361 14197 7395
rect 14197 7361 14231 7395
rect 14231 7361 14240 7395
rect 14188 7352 14240 7361
rect 14372 7395 14424 7404
rect 14372 7361 14381 7395
rect 14381 7361 14415 7395
rect 14415 7361 14424 7395
rect 14372 7352 14424 7361
rect 12716 7284 12768 7336
rect 14556 7395 14608 7404
rect 14556 7361 14565 7395
rect 14565 7361 14599 7395
rect 14599 7361 14608 7395
rect 14556 7352 14608 7361
rect 14740 7352 14792 7404
rect 15016 7284 15068 7336
rect 15108 7284 15160 7336
rect 2044 7148 2096 7200
rect 2504 7191 2556 7200
rect 2504 7157 2513 7191
rect 2513 7157 2547 7191
rect 2547 7157 2556 7191
rect 2504 7148 2556 7157
rect 3700 7191 3752 7200
rect 3700 7157 3709 7191
rect 3709 7157 3743 7191
rect 3743 7157 3752 7191
rect 3700 7148 3752 7157
rect 4528 7148 4580 7200
rect 5080 7148 5132 7200
rect 5908 7191 5960 7200
rect 5908 7157 5917 7191
rect 5917 7157 5951 7191
rect 5951 7157 5960 7191
rect 12072 7216 12124 7268
rect 13636 7216 13688 7268
rect 15660 7327 15712 7336
rect 15660 7293 15669 7327
rect 15669 7293 15703 7327
rect 15703 7293 15712 7327
rect 16488 7420 16540 7472
rect 17868 7488 17920 7540
rect 16672 7352 16724 7404
rect 18144 7420 18196 7472
rect 18604 7420 18656 7472
rect 18788 7420 18840 7472
rect 19616 7488 19668 7540
rect 21640 7488 21692 7540
rect 21916 7488 21968 7540
rect 23020 7531 23072 7540
rect 23020 7497 23029 7531
rect 23029 7497 23063 7531
rect 23063 7497 23072 7531
rect 23020 7488 23072 7497
rect 15660 7284 15712 7293
rect 16396 7284 16448 7336
rect 17224 7395 17276 7404
rect 17224 7361 17233 7395
rect 17233 7361 17267 7395
rect 17267 7361 17276 7395
rect 17224 7352 17276 7361
rect 17776 7284 17828 7336
rect 17960 7352 18012 7404
rect 18972 7395 19024 7404
rect 18972 7361 18981 7395
rect 18981 7361 19015 7395
rect 19015 7361 19024 7395
rect 18972 7352 19024 7361
rect 19340 7352 19392 7404
rect 19616 7352 19668 7404
rect 19800 7463 19852 7472
rect 19800 7429 19809 7463
rect 19809 7429 19843 7463
rect 19843 7429 19852 7463
rect 19800 7420 19852 7429
rect 21272 7420 21324 7472
rect 19984 7395 20036 7404
rect 18144 7284 18196 7336
rect 18236 7284 18288 7336
rect 18788 7284 18840 7336
rect 15844 7216 15896 7268
rect 16304 7216 16356 7268
rect 19432 7216 19484 7268
rect 19984 7361 19993 7395
rect 19993 7361 20027 7395
rect 20027 7361 20036 7395
rect 19984 7352 20036 7361
rect 20812 7395 20864 7404
rect 20812 7361 20821 7395
rect 20821 7361 20855 7395
rect 20855 7361 20864 7395
rect 20812 7352 20864 7361
rect 21732 7352 21784 7404
rect 22284 7395 22336 7404
rect 22284 7361 22293 7395
rect 22293 7361 22327 7395
rect 22327 7361 22336 7395
rect 22284 7352 22336 7361
rect 21272 7216 21324 7268
rect 21548 7216 21600 7268
rect 5908 7148 5960 7157
rect 8300 7148 8352 7200
rect 9128 7191 9180 7200
rect 9128 7157 9137 7191
rect 9137 7157 9171 7191
rect 9171 7157 9180 7191
rect 9128 7148 9180 7157
rect 9864 7148 9916 7200
rect 14188 7148 14240 7200
rect 15936 7148 15988 7200
rect 17500 7148 17552 7200
rect 18696 7148 18748 7200
rect 18972 7148 19024 7200
rect 22560 7395 22612 7404
rect 22560 7361 22569 7395
rect 22569 7361 22603 7395
rect 22603 7361 22612 7395
rect 22560 7352 22612 7361
rect 3790 7046 3842 7098
rect 3854 7046 3906 7098
rect 3918 7046 3970 7098
rect 3982 7046 4034 7098
rect 4046 7046 4098 7098
rect 9471 7046 9523 7098
rect 9535 7046 9587 7098
rect 9599 7046 9651 7098
rect 9663 7046 9715 7098
rect 9727 7046 9779 7098
rect 15152 7046 15204 7098
rect 15216 7046 15268 7098
rect 15280 7046 15332 7098
rect 15344 7046 15396 7098
rect 15408 7046 15460 7098
rect 20833 7046 20885 7098
rect 20897 7046 20949 7098
rect 20961 7046 21013 7098
rect 21025 7046 21077 7098
rect 21089 7046 21141 7098
rect 1768 6944 1820 6996
rect 3516 6944 3568 6996
rect 3700 6944 3752 6996
rect 2872 6876 2924 6928
rect 3332 6740 3384 6792
rect 5080 6944 5132 6996
rect 5264 6944 5316 6996
rect 6460 6944 6512 6996
rect 10600 6987 10652 6996
rect 4896 6876 4948 6928
rect 6000 6876 6052 6928
rect 4528 6783 4580 6792
rect 2136 6672 2188 6724
rect 3424 6672 3476 6724
rect 4528 6749 4537 6783
rect 4537 6749 4571 6783
rect 4571 6749 4580 6783
rect 4528 6740 4580 6749
rect 5356 6851 5408 6860
rect 5356 6817 5365 6851
rect 5365 6817 5399 6851
rect 5399 6817 5408 6851
rect 5356 6808 5408 6817
rect 5908 6808 5960 6860
rect 7748 6876 7800 6928
rect 10600 6953 10609 6987
rect 10609 6953 10643 6987
rect 10643 6953 10652 6987
rect 10600 6944 10652 6953
rect 11152 6987 11204 6996
rect 11152 6953 11161 6987
rect 11161 6953 11195 6987
rect 11195 6953 11204 6987
rect 11152 6944 11204 6953
rect 12992 6944 13044 6996
rect 14924 6987 14976 6996
rect 14924 6953 14933 6987
rect 14933 6953 14967 6987
rect 14967 6953 14976 6987
rect 14924 6944 14976 6953
rect 15476 6944 15528 6996
rect 16304 6944 16356 6996
rect 8484 6876 8536 6928
rect 8944 6876 8996 6928
rect 9496 6876 9548 6928
rect 11980 6876 12032 6928
rect 15936 6876 15988 6928
rect 16396 6876 16448 6928
rect 8208 6808 8260 6860
rect 8392 6808 8444 6860
rect 11244 6808 11296 6860
rect 4344 6672 4396 6724
rect 4804 6672 4856 6724
rect 7104 6740 7156 6792
rect 7472 6740 7524 6792
rect 8116 6740 8168 6792
rect 6000 6715 6052 6724
rect 6000 6681 6009 6715
rect 6009 6681 6043 6715
rect 6043 6681 6052 6715
rect 6000 6672 6052 6681
rect 7196 6672 7248 6724
rect 9496 6783 9548 6792
rect 9496 6749 9505 6783
rect 9505 6749 9539 6783
rect 9539 6749 9548 6783
rect 9496 6740 9548 6749
rect 2228 6647 2280 6656
rect 2228 6613 2237 6647
rect 2237 6613 2271 6647
rect 2271 6613 2280 6647
rect 2228 6604 2280 6613
rect 2688 6604 2740 6656
rect 5080 6604 5132 6656
rect 7012 6604 7064 6656
rect 7380 6604 7432 6656
rect 7472 6604 7524 6656
rect 8024 6604 8076 6656
rect 8208 6647 8260 6656
rect 8208 6613 8217 6647
rect 8217 6613 8251 6647
rect 8251 6613 8260 6647
rect 8208 6604 8260 6613
rect 8576 6604 8628 6656
rect 9404 6604 9456 6656
rect 11704 6783 11756 6792
rect 11704 6749 11713 6783
rect 11713 6749 11747 6783
rect 11747 6749 11756 6783
rect 11704 6740 11756 6749
rect 13544 6808 13596 6860
rect 13820 6808 13872 6860
rect 13912 6808 13964 6860
rect 17592 6944 17644 6996
rect 17776 6944 17828 6996
rect 20444 6944 20496 6996
rect 17500 6876 17552 6928
rect 18236 6876 18288 6928
rect 18972 6876 19024 6928
rect 13084 6783 13136 6792
rect 13084 6749 13093 6783
rect 13093 6749 13127 6783
rect 13127 6749 13136 6783
rect 13084 6740 13136 6749
rect 13176 6740 13228 6792
rect 14188 6740 14240 6792
rect 16580 6783 16632 6792
rect 11060 6672 11112 6724
rect 15936 6672 15988 6724
rect 10232 6604 10284 6656
rect 11428 6604 11480 6656
rect 14372 6604 14424 6656
rect 16580 6749 16589 6783
rect 16589 6749 16623 6783
rect 16623 6749 16632 6783
rect 16580 6740 16632 6749
rect 16856 6740 16908 6792
rect 17316 6783 17368 6792
rect 17316 6749 17325 6783
rect 17325 6749 17359 6783
rect 17359 6749 17368 6783
rect 17316 6740 17368 6749
rect 17408 6740 17460 6792
rect 18880 6808 18932 6860
rect 17684 6783 17736 6792
rect 17684 6749 17693 6783
rect 17693 6749 17727 6783
rect 17727 6749 17736 6783
rect 17684 6740 17736 6749
rect 18236 6740 18288 6792
rect 18420 6783 18472 6792
rect 18420 6749 18429 6783
rect 18429 6749 18463 6783
rect 18463 6749 18472 6783
rect 18420 6740 18472 6749
rect 18696 6740 18748 6792
rect 19800 6808 19852 6860
rect 20352 6851 20404 6860
rect 17040 6672 17092 6724
rect 19340 6740 19392 6792
rect 19892 6783 19944 6792
rect 19892 6749 19901 6783
rect 19901 6749 19935 6783
rect 19935 6749 19944 6783
rect 19892 6740 19944 6749
rect 20352 6817 20361 6851
rect 20361 6817 20395 6851
rect 20395 6817 20404 6851
rect 20352 6808 20404 6817
rect 21272 6876 21324 6928
rect 20536 6808 20588 6860
rect 20720 6808 20772 6860
rect 20076 6783 20128 6792
rect 20076 6749 20085 6783
rect 20085 6749 20119 6783
rect 20119 6749 20128 6783
rect 20076 6740 20128 6749
rect 20628 6740 20680 6792
rect 21456 6783 21508 6792
rect 18880 6715 18932 6724
rect 18880 6681 18889 6715
rect 18889 6681 18923 6715
rect 18923 6681 18932 6715
rect 18880 6672 18932 6681
rect 19800 6672 19852 6724
rect 21456 6749 21465 6783
rect 21465 6749 21499 6783
rect 21499 6749 21508 6783
rect 21456 6740 21508 6749
rect 18420 6604 18472 6656
rect 18788 6647 18840 6656
rect 18788 6613 18797 6647
rect 18797 6613 18831 6647
rect 18831 6613 18840 6647
rect 18788 6604 18840 6613
rect 19340 6604 19392 6656
rect 19708 6604 19760 6656
rect 6630 6502 6682 6554
rect 6694 6502 6746 6554
rect 6758 6502 6810 6554
rect 6822 6502 6874 6554
rect 6886 6502 6938 6554
rect 12311 6502 12363 6554
rect 12375 6502 12427 6554
rect 12439 6502 12491 6554
rect 12503 6502 12555 6554
rect 12567 6502 12619 6554
rect 17992 6502 18044 6554
rect 18056 6502 18108 6554
rect 18120 6502 18172 6554
rect 18184 6502 18236 6554
rect 18248 6502 18300 6554
rect 23673 6502 23725 6554
rect 23737 6502 23789 6554
rect 23801 6502 23853 6554
rect 23865 6502 23917 6554
rect 23929 6502 23981 6554
rect 3424 6400 3476 6452
rect 4344 6443 4396 6452
rect 4344 6409 4353 6443
rect 4353 6409 4387 6443
rect 4387 6409 4396 6443
rect 4344 6400 4396 6409
rect 4896 6400 4948 6452
rect 5172 6443 5224 6452
rect 5172 6409 5181 6443
rect 5181 6409 5215 6443
rect 5215 6409 5224 6443
rect 5172 6400 5224 6409
rect 5632 6400 5684 6452
rect 1860 6332 1912 6384
rect 2136 6332 2188 6384
rect 1768 6307 1820 6316
rect 1768 6273 1777 6307
rect 1777 6273 1811 6307
rect 1811 6273 1820 6307
rect 1768 6264 1820 6273
rect 1952 6307 2004 6316
rect 1952 6273 1961 6307
rect 1961 6273 1995 6307
rect 1995 6273 2004 6307
rect 1952 6264 2004 6273
rect 3608 6332 3660 6384
rect 4528 6332 4580 6384
rect 6552 6400 6604 6452
rect 7196 6443 7248 6452
rect 6460 6332 6512 6384
rect 7196 6409 7205 6443
rect 7205 6409 7239 6443
rect 7239 6409 7248 6443
rect 7196 6400 7248 6409
rect 9036 6443 9088 6452
rect 1584 6196 1636 6248
rect 2044 6196 2096 6248
rect 5816 6264 5868 6316
rect 4252 6196 4304 6248
rect 3700 6128 3752 6180
rect 3792 6171 3844 6180
rect 3792 6137 3801 6171
rect 3801 6137 3835 6171
rect 3835 6137 3844 6171
rect 3792 6128 3844 6137
rect 4896 6128 4948 6180
rect 6644 6307 6696 6316
rect 6644 6273 6654 6307
rect 6654 6273 6688 6307
rect 6688 6273 6696 6307
rect 6644 6264 6696 6273
rect 7104 6264 7156 6316
rect 7564 6264 7616 6316
rect 8024 6264 8076 6316
rect 6736 6196 6788 6248
rect 8484 6332 8536 6384
rect 9036 6409 9045 6443
rect 9045 6409 9079 6443
rect 9079 6409 9088 6443
rect 9036 6400 9088 6409
rect 9312 6400 9364 6452
rect 11796 6400 11848 6452
rect 16212 6443 16264 6452
rect 16212 6409 16221 6443
rect 16221 6409 16255 6443
rect 16255 6409 16264 6443
rect 16212 6400 16264 6409
rect 11704 6332 11756 6384
rect 12900 6332 12952 6384
rect 13912 6375 13964 6384
rect 13912 6341 13921 6375
rect 13921 6341 13955 6375
rect 13955 6341 13964 6375
rect 13912 6332 13964 6341
rect 8576 6307 8628 6316
rect 8576 6273 8585 6307
rect 8585 6273 8619 6307
rect 8619 6273 8628 6307
rect 8576 6264 8628 6273
rect 8668 6273 8677 6282
rect 8677 6273 8711 6282
rect 8711 6273 8720 6282
rect 8668 6230 8720 6273
rect 8760 6307 8812 6316
rect 8760 6273 8769 6307
rect 8769 6273 8803 6307
rect 8803 6273 8812 6307
rect 8760 6264 8812 6273
rect 10140 6264 10192 6316
rect 10232 6196 10284 6248
rect 10048 6128 10100 6180
rect 10876 6307 10928 6316
rect 10876 6273 10885 6307
rect 10885 6273 10919 6307
rect 10919 6273 10928 6307
rect 10876 6264 10928 6273
rect 12440 6264 12492 6316
rect 15752 6332 15804 6384
rect 15844 6332 15896 6384
rect 18144 6400 18196 6452
rect 19524 6400 19576 6452
rect 20536 6400 20588 6452
rect 21824 6400 21876 6452
rect 17684 6332 17736 6384
rect 19340 6375 19392 6384
rect 10508 6196 10560 6248
rect 11060 6196 11112 6248
rect 13084 6196 13136 6248
rect 13544 6239 13596 6248
rect 13544 6205 13553 6239
rect 13553 6205 13587 6239
rect 13587 6205 13596 6239
rect 13544 6196 13596 6205
rect 13636 6196 13688 6248
rect 15476 6264 15528 6316
rect 16120 6307 16172 6316
rect 16120 6273 16129 6307
rect 16129 6273 16163 6307
rect 16163 6273 16172 6307
rect 16120 6264 16172 6273
rect 16304 6307 16356 6316
rect 16304 6273 16313 6307
rect 16313 6273 16347 6307
rect 16347 6273 16356 6307
rect 16304 6264 16356 6273
rect 16396 6264 16448 6316
rect 17316 6264 17368 6316
rect 17776 6264 17828 6316
rect 19340 6341 19349 6375
rect 19349 6341 19383 6375
rect 19383 6341 19392 6375
rect 19340 6332 19392 6341
rect 18788 6264 18840 6316
rect 18972 6307 19024 6316
rect 18972 6273 18981 6307
rect 18981 6273 19015 6307
rect 19015 6273 19024 6307
rect 18972 6264 19024 6273
rect 19156 6264 19208 6316
rect 18052 6239 18104 6248
rect 11888 6128 11940 6180
rect 12900 6128 12952 6180
rect 18052 6205 18061 6239
rect 18061 6205 18095 6239
rect 18095 6205 18104 6239
rect 18052 6196 18104 6205
rect 14924 6128 14976 6180
rect 17960 6128 18012 6180
rect 18144 6128 18196 6180
rect 19984 6196 20036 6248
rect 20260 6307 20312 6316
rect 20260 6273 20269 6307
rect 20269 6273 20303 6307
rect 20303 6273 20312 6307
rect 20260 6264 20312 6273
rect 20720 6264 20772 6316
rect 21180 6196 21232 6248
rect 2044 6060 2096 6112
rect 5448 6060 5500 6112
rect 8024 6060 8076 6112
rect 10692 6060 10744 6112
rect 12808 6060 12860 6112
rect 13452 6103 13504 6112
rect 13452 6069 13461 6103
rect 13461 6069 13495 6103
rect 13495 6069 13504 6103
rect 14648 6103 14700 6112
rect 13452 6060 13504 6069
rect 14648 6069 14657 6103
rect 14657 6069 14691 6103
rect 14691 6069 14700 6103
rect 14648 6060 14700 6069
rect 16120 6060 16172 6112
rect 19892 6128 19944 6180
rect 20260 6128 20312 6180
rect 20444 6128 20496 6180
rect 18696 6060 18748 6112
rect 19340 6060 19392 6112
rect 19616 6060 19668 6112
rect 22100 6103 22152 6112
rect 22100 6069 22109 6103
rect 22109 6069 22143 6103
rect 22143 6069 22152 6103
rect 22100 6060 22152 6069
rect 3790 5958 3842 6010
rect 3854 5958 3906 6010
rect 3918 5958 3970 6010
rect 3982 5958 4034 6010
rect 4046 5958 4098 6010
rect 9471 5958 9523 6010
rect 9535 5958 9587 6010
rect 9599 5958 9651 6010
rect 9663 5958 9715 6010
rect 9727 5958 9779 6010
rect 15152 5958 15204 6010
rect 15216 5958 15268 6010
rect 15280 5958 15332 6010
rect 15344 5958 15396 6010
rect 15408 5958 15460 6010
rect 20833 5958 20885 6010
rect 20897 5958 20949 6010
rect 20961 5958 21013 6010
rect 21025 5958 21077 6010
rect 21089 5958 21141 6010
rect 5172 5856 5224 5908
rect 8116 5856 8168 5908
rect 8576 5856 8628 5908
rect 1492 5788 1544 5840
rect 1584 5720 1636 5772
rect 1952 5695 2004 5704
rect 1952 5661 1961 5695
rect 1961 5661 1995 5695
rect 1995 5661 2004 5695
rect 1952 5652 2004 5661
rect 2228 5695 2280 5704
rect 2228 5661 2237 5695
rect 2237 5661 2271 5695
rect 2271 5661 2280 5695
rect 2228 5652 2280 5661
rect 2320 5584 2372 5636
rect 2688 5720 2740 5772
rect 2228 5516 2280 5568
rect 2504 5516 2556 5568
rect 3608 5652 3660 5704
rect 4620 5720 4672 5772
rect 7472 5788 7524 5840
rect 9772 5788 9824 5840
rect 10048 5788 10100 5840
rect 10416 5831 10468 5840
rect 10416 5797 10425 5831
rect 10425 5797 10459 5831
rect 10459 5797 10468 5831
rect 10416 5788 10468 5797
rect 11244 5856 11296 5908
rect 11520 5856 11572 5908
rect 12808 5856 12860 5908
rect 12900 5856 12952 5908
rect 13360 5856 13412 5908
rect 13912 5856 13964 5908
rect 14832 5856 14884 5908
rect 16764 5856 16816 5908
rect 18328 5856 18380 5908
rect 18420 5856 18472 5908
rect 12992 5788 13044 5840
rect 17224 5788 17276 5840
rect 19616 5856 19668 5908
rect 20444 5899 20496 5908
rect 20444 5865 20453 5899
rect 20453 5865 20487 5899
rect 20487 5865 20496 5899
rect 20444 5856 20496 5865
rect 20628 5856 20680 5908
rect 4896 5695 4948 5704
rect 4896 5661 4905 5695
rect 4905 5661 4939 5695
rect 4939 5661 4948 5695
rect 4896 5652 4948 5661
rect 5080 5695 5132 5704
rect 5080 5661 5089 5695
rect 5089 5661 5123 5695
rect 5123 5661 5132 5695
rect 5080 5652 5132 5661
rect 5448 5695 5500 5704
rect 5448 5661 5457 5695
rect 5457 5661 5491 5695
rect 5491 5661 5500 5695
rect 5448 5652 5500 5661
rect 6092 5695 6144 5704
rect 6092 5661 6101 5695
rect 6101 5661 6135 5695
rect 6135 5661 6144 5695
rect 6092 5652 6144 5661
rect 6276 5695 6328 5704
rect 6276 5661 6285 5695
rect 6285 5661 6319 5695
rect 6319 5661 6328 5695
rect 6276 5652 6328 5661
rect 6644 5652 6696 5704
rect 7288 5695 7340 5704
rect 7288 5661 7297 5695
rect 7297 5661 7331 5695
rect 7331 5661 7340 5695
rect 7288 5652 7340 5661
rect 8208 5720 8260 5772
rect 7564 5695 7616 5704
rect 7564 5661 7573 5695
rect 7573 5661 7607 5695
rect 7607 5661 7616 5695
rect 7564 5652 7616 5661
rect 7656 5695 7708 5704
rect 7656 5661 7665 5695
rect 7665 5661 7699 5695
rect 7699 5661 7708 5695
rect 7656 5652 7708 5661
rect 8300 5652 8352 5704
rect 8576 5652 8628 5704
rect 13084 5720 13136 5772
rect 15016 5720 15068 5772
rect 15844 5720 15896 5772
rect 18972 5788 19024 5840
rect 19340 5788 19392 5840
rect 9496 5695 9548 5704
rect 9496 5661 9505 5695
rect 9505 5661 9539 5695
rect 9539 5661 9548 5695
rect 9496 5652 9548 5661
rect 9864 5652 9916 5704
rect 10048 5695 10100 5704
rect 10048 5661 10057 5695
rect 10057 5661 10091 5695
rect 10091 5661 10100 5695
rect 10048 5652 10100 5661
rect 10784 5652 10836 5704
rect 10968 5652 11020 5704
rect 8208 5584 8260 5636
rect 11428 5652 11480 5704
rect 13636 5652 13688 5704
rect 11888 5584 11940 5636
rect 12440 5584 12492 5636
rect 13820 5652 13872 5704
rect 16488 5695 16540 5704
rect 14648 5584 14700 5636
rect 4252 5516 4304 5568
rect 4436 5516 4488 5568
rect 6736 5516 6788 5568
rect 8300 5516 8352 5568
rect 9312 5516 9364 5568
rect 13176 5516 13228 5568
rect 16488 5661 16497 5695
rect 16497 5661 16531 5695
rect 16531 5661 16540 5695
rect 16488 5652 16540 5661
rect 16672 5695 16724 5704
rect 16672 5661 16681 5695
rect 16681 5661 16715 5695
rect 16715 5661 16724 5695
rect 16672 5652 16724 5661
rect 16948 5652 17000 5704
rect 18328 5652 18380 5704
rect 18696 5763 18748 5772
rect 18696 5729 18705 5763
rect 18705 5729 18739 5763
rect 18739 5729 18748 5763
rect 18696 5720 18748 5729
rect 19156 5720 19208 5772
rect 18696 5584 18748 5636
rect 19432 5584 19484 5636
rect 19340 5516 19392 5568
rect 20536 5584 20588 5636
rect 6630 5414 6682 5466
rect 6694 5414 6746 5466
rect 6758 5414 6810 5466
rect 6822 5414 6874 5466
rect 6886 5414 6938 5466
rect 12311 5414 12363 5466
rect 12375 5414 12427 5466
rect 12439 5414 12491 5466
rect 12503 5414 12555 5466
rect 12567 5414 12619 5466
rect 17992 5414 18044 5466
rect 18056 5414 18108 5466
rect 18120 5414 18172 5466
rect 18184 5414 18236 5466
rect 18248 5414 18300 5466
rect 23673 5414 23725 5466
rect 23737 5414 23789 5466
rect 23801 5414 23853 5466
rect 23865 5414 23917 5466
rect 23929 5414 23981 5466
rect 2780 5312 2832 5364
rect 3424 5355 3476 5364
rect 3424 5321 3433 5355
rect 3433 5321 3467 5355
rect 3467 5321 3476 5355
rect 3424 5312 3476 5321
rect 3516 5312 3568 5364
rect 2136 5244 2188 5296
rect 2228 5219 2280 5228
rect 2228 5185 2237 5219
rect 2237 5185 2271 5219
rect 2271 5185 2280 5219
rect 2228 5176 2280 5185
rect 3332 5176 3384 5228
rect 4712 5219 4764 5228
rect 4712 5185 4721 5219
rect 4721 5185 4755 5219
rect 4755 5185 4764 5219
rect 4712 5176 4764 5185
rect 6276 5312 6328 5364
rect 8668 5312 8720 5364
rect 8852 5355 8904 5364
rect 8852 5321 8861 5355
rect 8861 5321 8895 5355
rect 8895 5321 8904 5355
rect 8852 5312 8904 5321
rect 11888 5312 11940 5364
rect 13636 5312 13688 5364
rect 5632 5244 5684 5296
rect 4988 5219 5040 5228
rect 4988 5185 4997 5219
rect 4997 5185 5031 5219
rect 5031 5185 5040 5219
rect 4988 5176 5040 5185
rect 6552 5244 6604 5296
rect 7840 5244 7892 5296
rect 8116 5244 8168 5296
rect 10140 5244 10192 5296
rect 10508 5244 10560 5296
rect 11336 5244 11388 5296
rect 7380 5219 7432 5228
rect 2780 5108 2832 5160
rect 3700 5108 3752 5160
rect 5540 5108 5592 5160
rect 2320 5040 2372 5092
rect 7380 5185 7389 5219
rect 7389 5185 7423 5219
rect 7423 5185 7432 5219
rect 7380 5176 7432 5185
rect 6000 5040 6052 5092
rect 8024 5040 8076 5092
rect 8852 5176 8904 5228
rect 10784 5176 10836 5228
rect 11796 5219 11848 5228
rect 11796 5185 11805 5219
rect 11805 5185 11839 5219
rect 11839 5185 11848 5219
rect 11796 5176 11848 5185
rect 11980 5176 12032 5228
rect 12256 5287 12308 5296
rect 12256 5253 12265 5287
rect 12265 5253 12299 5287
rect 12299 5253 12308 5287
rect 12256 5244 12308 5253
rect 12716 5176 12768 5228
rect 13360 5244 13412 5296
rect 13820 5219 13872 5228
rect 8484 5108 8536 5160
rect 8760 5151 8812 5160
rect 8760 5117 8769 5151
rect 8769 5117 8803 5151
rect 8803 5117 8812 5151
rect 8760 5108 8812 5117
rect 9220 5108 9272 5160
rect 11520 5108 11572 5160
rect 13360 5108 13412 5160
rect 13820 5185 13829 5219
rect 13829 5185 13863 5219
rect 13863 5185 13872 5219
rect 13820 5176 13872 5185
rect 13912 5219 13964 5228
rect 13912 5185 13921 5219
rect 13921 5185 13955 5219
rect 13955 5185 13964 5219
rect 15476 5312 15528 5364
rect 15844 5312 15896 5364
rect 16396 5312 16448 5364
rect 17132 5312 17184 5364
rect 18420 5312 18472 5364
rect 18972 5312 19024 5364
rect 14740 5244 14792 5296
rect 15568 5287 15620 5296
rect 15568 5253 15577 5287
rect 15577 5253 15611 5287
rect 15611 5253 15620 5287
rect 15568 5244 15620 5253
rect 16580 5244 16632 5296
rect 13912 5176 13964 5185
rect 16488 5176 16540 5228
rect 16856 5219 16908 5228
rect 16856 5185 16865 5219
rect 16865 5185 16899 5219
rect 16899 5185 16908 5219
rect 16856 5176 16908 5185
rect 20628 5312 20680 5364
rect 18604 5219 18656 5228
rect 18604 5185 18613 5219
rect 18613 5185 18647 5219
rect 18647 5185 18656 5219
rect 18604 5176 18656 5185
rect 19616 5219 19668 5228
rect 19616 5185 19625 5219
rect 19625 5185 19659 5219
rect 19659 5185 19668 5219
rect 19616 5176 19668 5185
rect 20352 5219 20404 5228
rect 20352 5185 20361 5219
rect 20361 5185 20395 5219
rect 20395 5185 20404 5219
rect 20352 5176 20404 5185
rect 9036 5040 9088 5092
rect 9496 5040 9548 5092
rect 11244 5040 11296 5092
rect 12348 5040 12400 5092
rect 13176 5040 13228 5092
rect 19432 5108 19484 5160
rect 20720 5176 20772 5228
rect 17132 5040 17184 5092
rect 18696 5040 18748 5092
rect 20352 5040 20404 5092
rect 21180 5040 21232 5092
rect 6276 4972 6328 5024
rect 7288 4972 7340 5024
rect 9220 5015 9272 5024
rect 9220 4981 9229 5015
rect 9229 4981 9263 5015
rect 9263 4981 9272 5015
rect 9220 4972 9272 4981
rect 10876 5015 10928 5024
rect 10876 4981 10885 5015
rect 10885 4981 10919 5015
rect 10919 4981 10928 5015
rect 10876 4972 10928 4981
rect 13636 5015 13688 5024
rect 13636 4981 13645 5015
rect 13645 4981 13679 5015
rect 13679 4981 13688 5015
rect 13636 4972 13688 4981
rect 14648 5015 14700 5024
rect 14648 4981 14657 5015
rect 14657 4981 14691 5015
rect 14691 4981 14700 5015
rect 14648 4972 14700 4981
rect 15568 4972 15620 5024
rect 20536 4972 20588 5024
rect 3790 4870 3842 4922
rect 3854 4870 3906 4922
rect 3918 4870 3970 4922
rect 3982 4870 4034 4922
rect 4046 4870 4098 4922
rect 9471 4870 9523 4922
rect 9535 4870 9587 4922
rect 9599 4870 9651 4922
rect 9663 4870 9715 4922
rect 9727 4870 9779 4922
rect 15152 4870 15204 4922
rect 15216 4870 15268 4922
rect 15280 4870 15332 4922
rect 15344 4870 15396 4922
rect 15408 4870 15460 4922
rect 20833 4870 20885 4922
rect 20897 4870 20949 4922
rect 20961 4870 21013 4922
rect 21025 4870 21077 4922
rect 21089 4870 21141 4922
rect 1676 4811 1728 4820
rect 1676 4777 1685 4811
rect 1685 4777 1719 4811
rect 1719 4777 1728 4811
rect 1676 4768 1728 4777
rect 2320 4768 2372 4820
rect 2504 4811 2556 4820
rect 2504 4777 2513 4811
rect 2513 4777 2547 4811
rect 2547 4777 2556 4811
rect 2504 4768 2556 4777
rect 4068 4811 4120 4820
rect 4068 4777 4077 4811
rect 4077 4777 4111 4811
rect 4111 4777 4120 4811
rect 4068 4768 4120 4777
rect 7932 4768 7984 4820
rect 8024 4811 8076 4820
rect 8024 4777 8033 4811
rect 8033 4777 8067 4811
rect 8067 4777 8076 4811
rect 8392 4811 8444 4820
rect 8024 4768 8076 4777
rect 8392 4777 8401 4811
rect 8401 4777 8435 4811
rect 8435 4777 8444 4811
rect 8392 4768 8444 4777
rect 11520 4811 11572 4820
rect 11520 4777 11529 4811
rect 11529 4777 11563 4811
rect 11563 4777 11572 4811
rect 11520 4768 11572 4777
rect 12256 4811 12308 4820
rect 12256 4777 12265 4811
rect 12265 4777 12299 4811
rect 12299 4777 12308 4811
rect 12256 4768 12308 4777
rect 12348 4768 12400 4820
rect 15568 4768 15620 4820
rect 3240 4700 3292 4752
rect 3424 4700 3476 4752
rect 4252 4675 4304 4684
rect 2044 4564 2096 4616
rect 2780 4564 2832 4616
rect 4252 4641 4261 4675
rect 4261 4641 4295 4675
rect 4295 4641 4304 4675
rect 4252 4632 4304 4641
rect 3608 4564 3660 4616
rect 4068 4564 4120 4616
rect 4712 4700 4764 4752
rect 5356 4700 5408 4752
rect 5540 4700 5592 4752
rect 6092 4700 6144 4752
rect 5172 4607 5224 4616
rect 4528 4496 4580 4548
rect 4620 4496 4672 4548
rect 5172 4573 5181 4607
rect 5181 4573 5215 4607
rect 5215 4573 5224 4607
rect 5172 4564 5224 4573
rect 6552 4564 6604 4616
rect 6920 4700 6972 4752
rect 9864 4700 9916 4752
rect 10048 4700 10100 4752
rect 10600 4700 10652 4752
rect 11060 4700 11112 4752
rect 7196 4632 7248 4684
rect 7472 4564 7524 4616
rect 8116 4564 8168 4616
rect 9312 4564 9364 4616
rect 3240 4428 3292 4480
rect 5264 4471 5316 4480
rect 5264 4437 5273 4471
rect 5273 4437 5307 4471
rect 5307 4437 5316 4471
rect 5264 4428 5316 4437
rect 5356 4471 5408 4480
rect 5356 4437 5365 4471
rect 5365 4437 5399 4471
rect 5399 4437 5408 4471
rect 7196 4496 7248 4548
rect 7288 4496 7340 4548
rect 10232 4564 10284 4616
rect 10876 4607 10928 4616
rect 10876 4573 10885 4607
rect 10885 4573 10919 4607
rect 10919 4573 10928 4607
rect 10876 4564 10928 4573
rect 11888 4700 11940 4752
rect 12072 4632 12124 4684
rect 12716 4632 12768 4684
rect 11888 4564 11940 4616
rect 5356 4428 5408 4437
rect 7840 4428 7892 4480
rect 9496 4496 9548 4548
rect 10324 4539 10376 4548
rect 10324 4505 10333 4539
rect 10333 4505 10367 4539
rect 10367 4505 10376 4539
rect 10324 4496 10376 4505
rect 10508 4496 10560 4548
rect 11336 4496 11388 4548
rect 12256 4564 12308 4616
rect 13820 4632 13872 4684
rect 14924 4675 14976 4684
rect 14924 4641 14933 4675
rect 14933 4641 14967 4675
rect 14967 4641 14976 4675
rect 16856 4768 16908 4820
rect 18328 4768 18380 4820
rect 22100 4768 22152 4820
rect 16396 4743 16448 4752
rect 16396 4709 16405 4743
rect 16405 4709 16439 4743
rect 16439 4709 16448 4743
rect 16396 4700 16448 4709
rect 17132 4700 17184 4752
rect 18512 4700 18564 4752
rect 14924 4632 14976 4641
rect 17592 4632 17644 4684
rect 13912 4564 13964 4616
rect 20352 4564 20404 4616
rect 15016 4539 15068 4548
rect 15016 4505 15025 4539
rect 15025 4505 15059 4539
rect 15059 4505 15068 4539
rect 15016 4496 15068 4505
rect 15200 4496 15252 4548
rect 16488 4496 16540 4548
rect 11888 4428 11940 4480
rect 14556 4428 14608 4480
rect 6630 4326 6682 4378
rect 6694 4326 6746 4378
rect 6758 4326 6810 4378
rect 6822 4326 6874 4378
rect 6886 4326 6938 4378
rect 12311 4326 12363 4378
rect 12375 4326 12427 4378
rect 12439 4326 12491 4378
rect 12503 4326 12555 4378
rect 12567 4326 12619 4378
rect 17992 4326 18044 4378
rect 18056 4326 18108 4378
rect 18120 4326 18172 4378
rect 18184 4326 18236 4378
rect 18248 4326 18300 4378
rect 23673 4326 23725 4378
rect 23737 4326 23789 4378
rect 23801 4326 23853 4378
rect 23865 4326 23917 4378
rect 23929 4326 23981 4378
rect 1676 4267 1728 4276
rect 1676 4233 1685 4267
rect 1685 4233 1719 4267
rect 1719 4233 1728 4267
rect 1676 4224 1728 4233
rect 4068 4224 4120 4276
rect 4712 4224 4764 4276
rect 5264 4224 5316 4276
rect 7196 4267 7248 4276
rect 2044 4088 2096 4140
rect 2872 4131 2924 4140
rect 2872 4097 2881 4131
rect 2881 4097 2915 4131
rect 2915 4097 2924 4131
rect 2872 4088 2924 4097
rect 3424 4088 3476 4140
rect 5172 4156 5224 4208
rect 4344 4088 4396 4140
rect 4896 4131 4948 4140
rect 4896 4097 4905 4131
rect 4905 4097 4939 4131
rect 4939 4097 4948 4131
rect 4896 4088 4948 4097
rect 5080 4131 5132 4140
rect 5080 4097 5089 4131
rect 5089 4097 5123 4131
rect 5123 4097 5132 4131
rect 5080 4088 5132 4097
rect 7196 4233 7205 4267
rect 7205 4233 7239 4267
rect 7239 4233 7248 4267
rect 7196 4224 7248 4233
rect 10416 4224 10468 4276
rect 8484 4156 8536 4208
rect 6000 4063 6052 4072
rect 6000 4029 6009 4063
rect 6009 4029 6043 4063
rect 6043 4029 6052 4063
rect 6000 4020 6052 4029
rect 6552 4063 6604 4072
rect 6552 4029 6561 4063
rect 6561 4029 6595 4063
rect 6595 4029 6604 4063
rect 6552 4020 6604 4029
rect 6828 4131 6880 4140
rect 6828 4097 6837 4131
rect 6837 4097 6871 4131
rect 6871 4097 6880 4131
rect 6828 4088 6880 4097
rect 7840 4131 7892 4140
rect 7840 4097 7849 4131
rect 7849 4097 7883 4131
rect 7883 4097 7892 4131
rect 7840 4088 7892 4097
rect 6920 4020 6972 4072
rect 7104 4020 7156 4072
rect 8208 4088 8260 4140
rect 9128 4131 9180 4140
rect 9128 4097 9137 4131
rect 9137 4097 9171 4131
rect 9171 4097 9180 4131
rect 9128 4088 9180 4097
rect 11336 4156 11388 4208
rect 9956 4131 10008 4140
rect 9956 4097 9965 4131
rect 9965 4097 9999 4131
rect 9999 4097 10008 4131
rect 9956 4088 10008 4097
rect 8300 4020 8352 4072
rect 8576 4020 8628 4072
rect 9220 4020 9272 4072
rect 10876 4088 10928 4140
rect 11520 4088 11572 4140
rect 11888 4131 11940 4140
rect 11888 4097 11897 4131
rect 11897 4097 11931 4131
rect 11931 4097 11940 4131
rect 11888 4088 11940 4097
rect 15200 4267 15252 4276
rect 15200 4233 15209 4267
rect 15209 4233 15243 4267
rect 15243 4233 15252 4267
rect 15200 4224 15252 4233
rect 17132 4267 17184 4276
rect 17132 4233 17141 4267
rect 17141 4233 17175 4267
rect 17175 4233 17184 4267
rect 17132 4224 17184 4233
rect 12440 4156 12492 4208
rect 10232 4020 10284 4072
rect 11244 4020 11296 4072
rect 11428 4020 11480 4072
rect 11796 4020 11848 4072
rect 13544 4088 13596 4140
rect 16672 4156 16724 4208
rect 15752 4088 15804 4140
rect 13636 4020 13688 4072
rect 4160 3952 4212 4004
rect 4712 3952 4764 4004
rect 6092 3952 6144 4004
rect 10140 3952 10192 4004
rect 10324 3952 10376 4004
rect 12164 3952 12216 4004
rect 13452 3952 13504 4004
rect 5632 3884 5684 3936
rect 7472 3884 7524 3936
rect 11336 3884 11388 3936
rect 11520 3884 11572 3936
rect 12256 3884 12308 3936
rect 3790 3782 3842 3834
rect 3854 3782 3906 3834
rect 3918 3782 3970 3834
rect 3982 3782 4034 3834
rect 4046 3782 4098 3834
rect 9471 3782 9523 3834
rect 9535 3782 9587 3834
rect 9599 3782 9651 3834
rect 9663 3782 9715 3834
rect 9727 3782 9779 3834
rect 15152 3782 15204 3834
rect 15216 3782 15268 3834
rect 15280 3782 15332 3834
rect 15344 3782 15396 3834
rect 15408 3782 15460 3834
rect 20833 3782 20885 3834
rect 20897 3782 20949 3834
rect 20961 3782 21013 3834
rect 21025 3782 21077 3834
rect 21089 3782 21141 3834
rect 4160 3680 4212 3732
rect 4252 3680 4304 3732
rect 4528 3723 4580 3732
rect 4528 3689 4537 3723
rect 4537 3689 4571 3723
rect 4571 3689 4580 3723
rect 4528 3680 4580 3689
rect 4712 3680 4764 3732
rect 6368 3680 6420 3732
rect 6460 3680 6512 3732
rect 8760 3680 8812 3732
rect 10876 3680 10928 3732
rect 11060 3680 11112 3732
rect 11796 3680 11848 3732
rect 11888 3680 11940 3732
rect 12348 3680 12400 3732
rect 12716 3680 12768 3732
rect 13544 3680 13596 3732
rect 16672 3680 16724 3732
rect 4896 3655 4948 3664
rect 4896 3621 4905 3655
rect 4905 3621 4939 3655
rect 4939 3621 4948 3655
rect 4896 3612 4948 3621
rect 5356 3612 5408 3664
rect 3148 3544 3200 3596
rect 3424 3519 3476 3528
rect 2872 3408 2924 3460
rect 3424 3485 3433 3519
rect 3433 3485 3467 3519
rect 3467 3485 3476 3519
rect 3424 3476 3476 3485
rect 4436 3476 4488 3528
rect 4620 3519 4672 3528
rect 4620 3485 4629 3519
rect 4629 3485 4663 3519
rect 4663 3485 4672 3519
rect 4620 3476 4672 3485
rect 7748 3612 7800 3664
rect 10324 3612 10376 3664
rect 15016 3612 15068 3664
rect 6092 3587 6144 3596
rect 6092 3553 6101 3587
rect 6101 3553 6135 3587
rect 6135 3553 6144 3587
rect 6092 3544 6144 3553
rect 6828 3544 6880 3596
rect 8852 3544 8904 3596
rect 9220 3544 9272 3596
rect 10140 3544 10192 3596
rect 6460 3519 6512 3528
rect 6460 3485 6469 3519
rect 6469 3485 6503 3519
rect 6503 3485 6512 3519
rect 6460 3476 6512 3485
rect 7104 3476 7156 3528
rect 7288 3519 7340 3528
rect 7288 3485 7297 3519
rect 7297 3485 7331 3519
rect 7331 3485 7340 3519
rect 7288 3476 7340 3485
rect 7472 3519 7524 3528
rect 7472 3485 7481 3519
rect 7481 3485 7515 3519
rect 7515 3485 7524 3519
rect 7472 3476 7524 3485
rect 7840 3476 7892 3528
rect 8208 3476 8260 3528
rect 9128 3519 9180 3528
rect 2688 3383 2740 3392
rect 2688 3349 2697 3383
rect 2697 3349 2731 3383
rect 2731 3349 2740 3383
rect 2688 3340 2740 3349
rect 3240 3383 3292 3392
rect 3240 3349 3249 3383
rect 3249 3349 3283 3383
rect 3283 3349 3292 3383
rect 3240 3340 3292 3349
rect 5540 3340 5592 3392
rect 7748 3408 7800 3460
rect 8300 3451 8352 3460
rect 8300 3417 8309 3451
rect 8309 3417 8343 3451
rect 8343 3417 8352 3451
rect 8300 3408 8352 3417
rect 9128 3485 9137 3519
rect 9137 3485 9171 3519
rect 9171 3485 9180 3519
rect 9128 3476 9180 3485
rect 10232 3519 10284 3528
rect 10232 3485 10241 3519
rect 10241 3485 10275 3519
rect 10275 3485 10284 3519
rect 10232 3476 10284 3485
rect 10692 3544 10744 3596
rect 11612 3544 11664 3596
rect 12256 3587 12308 3596
rect 8576 3340 8628 3392
rect 9956 3408 10008 3460
rect 10600 3519 10652 3528
rect 10600 3485 10609 3519
rect 10609 3485 10643 3519
rect 10643 3485 10652 3519
rect 10600 3476 10652 3485
rect 11428 3519 11480 3528
rect 11428 3485 11437 3519
rect 11437 3485 11471 3519
rect 11471 3485 11480 3519
rect 11428 3476 11480 3485
rect 11520 3476 11572 3528
rect 11888 3476 11940 3528
rect 12256 3553 12265 3587
rect 12265 3553 12299 3587
rect 12299 3553 12308 3587
rect 12256 3544 12308 3553
rect 12348 3476 12400 3528
rect 13912 3476 13964 3528
rect 15752 3476 15804 3528
rect 23388 3476 23440 3528
rect 14372 3408 14424 3460
rect 17960 3451 18012 3460
rect 17960 3417 17969 3451
rect 17969 3417 18003 3451
rect 18003 3417 18012 3451
rect 17960 3408 18012 3417
rect 11980 3340 12032 3392
rect 17316 3383 17368 3392
rect 17316 3349 17325 3383
rect 17325 3349 17359 3383
rect 17359 3349 17368 3383
rect 17316 3340 17368 3349
rect 6630 3238 6682 3290
rect 6694 3238 6746 3290
rect 6758 3238 6810 3290
rect 6822 3238 6874 3290
rect 6886 3238 6938 3290
rect 12311 3238 12363 3290
rect 12375 3238 12427 3290
rect 12439 3238 12491 3290
rect 12503 3238 12555 3290
rect 12567 3238 12619 3290
rect 17992 3238 18044 3290
rect 18056 3238 18108 3290
rect 18120 3238 18172 3290
rect 18184 3238 18236 3290
rect 18248 3238 18300 3290
rect 23673 3238 23725 3290
rect 23737 3238 23789 3290
rect 23801 3238 23853 3290
rect 23865 3238 23917 3290
rect 23929 3238 23981 3290
rect 1676 3179 1728 3188
rect 1676 3145 1685 3179
rect 1685 3145 1719 3179
rect 1719 3145 1728 3179
rect 1676 3136 1728 3145
rect 4896 3136 4948 3188
rect 7380 3136 7432 3188
rect 9128 3136 9180 3188
rect 11520 3136 11572 3188
rect 11796 3136 11848 3188
rect 12072 3179 12124 3188
rect 12072 3145 12081 3179
rect 12081 3145 12115 3179
rect 12115 3145 12124 3179
rect 12072 3136 12124 3145
rect 13912 3179 13964 3188
rect 13912 3145 13921 3179
rect 13921 3145 13955 3179
rect 13955 3145 13964 3179
rect 13912 3136 13964 3145
rect 14372 3179 14424 3188
rect 14372 3145 14381 3179
rect 14381 3145 14415 3179
rect 14415 3145 14424 3179
rect 14372 3136 14424 3145
rect 17408 3179 17460 3188
rect 17408 3145 17417 3179
rect 17417 3145 17451 3179
rect 17451 3145 17460 3179
rect 17408 3136 17460 3145
rect 2504 3043 2556 3052
rect 2504 3009 2513 3043
rect 2513 3009 2547 3043
rect 2547 3009 2556 3043
rect 2504 3000 2556 3009
rect 7932 3068 7984 3120
rect 8484 3068 8536 3120
rect 8944 3068 8996 3120
rect 9220 3068 9272 3120
rect 10416 3111 10468 3120
rect 5632 3000 5684 3052
rect 5908 3000 5960 3052
rect 7288 3000 7340 3052
rect 8300 3000 8352 3052
rect 6460 2864 6512 2916
rect 2136 2796 2188 2848
rect 4528 2796 4580 2848
rect 7380 2932 7432 2984
rect 8484 2932 8536 2984
rect 8852 3000 8904 3052
rect 9312 3043 9364 3052
rect 9312 3009 9321 3043
rect 9321 3009 9355 3043
rect 9355 3009 9364 3043
rect 9312 3000 9364 3009
rect 10416 3077 10425 3111
rect 10425 3077 10459 3111
rect 10459 3077 10468 3111
rect 10416 3068 10468 3077
rect 11704 3111 11756 3120
rect 11704 3077 11713 3111
rect 11713 3077 11747 3111
rect 11747 3077 11756 3111
rect 11704 3068 11756 3077
rect 12164 3068 12216 3120
rect 10324 3043 10376 3052
rect 10324 3009 10333 3043
rect 10333 3009 10367 3043
rect 10367 3009 10376 3043
rect 10324 3000 10376 3009
rect 10968 3049 11020 3052
rect 10968 3015 10969 3049
rect 10969 3015 11003 3049
rect 11003 3015 11020 3049
rect 10968 3000 11020 3015
rect 6644 2907 6696 2916
rect 6644 2873 6653 2907
rect 6653 2873 6687 2907
rect 6687 2873 6696 2907
rect 6644 2864 6696 2873
rect 9864 2864 9916 2916
rect 11336 2796 11388 2848
rect 15660 2796 15712 2848
rect 16856 2839 16908 2848
rect 16856 2805 16865 2839
rect 16865 2805 16899 2839
rect 16899 2805 16908 2839
rect 16856 2796 16908 2805
rect 18328 2839 18380 2848
rect 18328 2805 18337 2839
rect 18337 2805 18371 2839
rect 18371 2805 18380 2839
rect 18328 2796 18380 2805
rect 20720 2796 20772 2848
rect 22744 2796 22796 2848
rect 3790 2694 3842 2746
rect 3854 2694 3906 2746
rect 3918 2694 3970 2746
rect 3982 2694 4034 2746
rect 4046 2694 4098 2746
rect 9471 2694 9523 2746
rect 9535 2694 9587 2746
rect 9599 2694 9651 2746
rect 9663 2694 9715 2746
rect 9727 2694 9779 2746
rect 15152 2694 15204 2746
rect 15216 2694 15268 2746
rect 15280 2694 15332 2746
rect 15344 2694 15396 2746
rect 15408 2694 15460 2746
rect 20833 2694 20885 2746
rect 20897 2694 20949 2746
rect 20961 2694 21013 2746
rect 21025 2694 21077 2746
rect 21089 2694 21141 2746
rect 7840 2635 7892 2644
rect 7840 2601 7849 2635
rect 7849 2601 7883 2635
rect 7883 2601 7892 2635
rect 7840 2592 7892 2601
rect 8484 2592 8536 2644
rect 1860 2431 1912 2440
rect 1860 2397 1869 2431
rect 1869 2397 1903 2431
rect 1903 2397 1912 2431
rect 1860 2388 1912 2397
rect 3240 2388 3292 2440
rect 3424 2431 3476 2440
rect 3424 2397 3433 2431
rect 3433 2397 3467 2431
rect 3467 2397 3476 2431
rect 3424 2388 3476 2397
rect 4252 2431 4304 2440
rect 4252 2397 4261 2431
rect 4261 2397 4295 2431
rect 4295 2397 4304 2431
rect 4252 2388 4304 2397
rect 5080 2524 5132 2576
rect 11152 2524 11204 2576
rect 11980 2592 12032 2644
rect 16856 2592 16908 2644
rect 8300 2456 8352 2508
rect 8944 2456 8996 2508
rect 5816 2388 5868 2440
rect 7380 2431 7432 2440
rect 1492 2252 1544 2304
rect 2780 2252 2832 2304
rect 3424 2252 3476 2304
rect 4068 2295 4120 2304
rect 4068 2261 4077 2295
rect 4077 2261 4111 2295
rect 4111 2261 4120 2295
rect 4068 2252 4120 2261
rect 4712 2252 4764 2304
rect 5356 2252 5408 2304
rect 6000 2252 6052 2304
rect 7380 2397 7389 2431
rect 7389 2397 7423 2431
rect 7423 2397 7432 2431
rect 7380 2388 7432 2397
rect 7472 2431 7524 2440
rect 7472 2397 7481 2431
rect 7481 2397 7515 2431
rect 7515 2397 7524 2431
rect 7656 2431 7708 2440
rect 7472 2388 7524 2397
rect 7656 2397 7665 2431
rect 7665 2397 7699 2431
rect 7699 2397 7708 2431
rect 7656 2388 7708 2397
rect 9036 2388 9088 2440
rect 10508 2320 10560 2372
rect 11612 2388 11664 2440
rect 11888 2431 11940 2440
rect 11888 2397 11897 2431
rect 11897 2397 11931 2431
rect 11931 2397 11940 2431
rect 11888 2388 11940 2397
rect 12716 2388 12768 2440
rect 13084 2388 13136 2440
rect 13728 2388 13780 2440
rect 14372 2388 14424 2440
rect 15016 2388 15068 2440
rect 11796 2320 11848 2372
rect 17316 2524 17368 2576
rect 16304 2388 16356 2440
rect 16948 2388 17000 2440
rect 17592 2388 17644 2440
rect 18880 2388 18932 2440
rect 19524 2388 19576 2440
rect 20168 2388 20220 2440
rect 21456 2388 21508 2440
rect 22100 2388 22152 2440
rect 16396 2320 16448 2372
rect 6630 2150 6682 2202
rect 6694 2150 6746 2202
rect 6758 2150 6810 2202
rect 6822 2150 6874 2202
rect 6886 2150 6938 2202
rect 12311 2150 12363 2202
rect 12375 2150 12427 2202
rect 12439 2150 12491 2202
rect 12503 2150 12555 2202
rect 12567 2150 12619 2202
rect 17992 2150 18044 2202
rect 18056 2150 18108 2202
rect 18120 2150 18172 2202
rect 18184 2150 18236 2202
rect 18248 2150 18300 2202
rect 23673 2150 23725 2202
rect 23737 2150 23789 2202
rect 23801 2150 23853 2202
rect 23865 2150 23917 2202
rect 23929 2150 23981 2202
rect 8208 2048 8260 2100
rect 16396 2048 16448 2100
<< metal2 >>
rect 2502 24200 2558 25000
rect 7470 24200 7526 25000
rect 12438 24200 12494 25000
rect 17406 24200 17462 25000
rect 22374 24200 22430 25000
rect 2516 21146 2544 24200
rect 3790 22332 4098 22341
rect 3790 22330 3796 22332
rect 3852 22330 3876 22332
rect 3932 22330 3956 22332
rect 4012 22330 4036 22332
rect 4092 22330 4098 22332
rect 3852 22278 3854 22330
rect 4034 22278 4036 22330
rect 3790 22276 3796 22278
rect 3852 22276 3876 22278
rect 3932 22276 3956 22278
rect 4012 22276 4036 22278
rect 4092 22276 4098 22278
rect 3790 22267 4098 22276
rect 7484 21962 7512 24200
rect 9471 22332 9779 22341
rect 9471 22330 9477 22332
rect 9533 22330 9557 22332
rect 9613 22330 9637 22332
rect 9693 22330 9717 22332
rect 9773 22330 9779 22332
rect 9533 22278 9535 22330
rect 9715 22278 9717 22330
rect 9471 22276 9477 22278
rect 9533 22276 9557 22278
rect 9613 22276 9637 22278
rect 9693 22276 9717 22278
rect 9773 22276 9779 22278
rect 9471 22267 9779 22276
rect 12452 22030 12480 24200
rect 15152 22332 15460 22341
rect 15152 22330 15158 22332
rect 15214 22330 15238 22332
rect 15294 22330 15318 22332
rect 15374 22330 15398 22332
rect 15454 22330 15460 22332
rect 15214 22278 15216 22330
rect 15396 22278 15398 22330
rect 15152 22276 15158 22278
rect 15214 22276 15238 22278
rect 15294 22276 15318 22278
rect 15374 22276 15398 22278
rect 15454 22276 15460 22278
rect 15152 22267 15460 22276
rect 17420 22030 17448 24200
rect 20833 22332 21141 22341
rect 20833 22330 20839 22332
rect 20895 22330 20919 22332
rect 20975 22330 20999 22332
rect 21055 22330 21079 22332
rect 21135 22330 21141 22332
rect 20895 22278 20897 22330
rect 21077 22278 21079 22330
rect 20833 22276 20839 22278
rect 20895 22276 20919 22278
rect 20975 22276 20999 22278
rect 21055 22276 21079 22278
rect 21135 22276 21141 22278
rect 20833 22267 21141 22276
rect 22388 22030 22416 24200
rect 9772 22024 9824 22030
rect 9772 21966 9824 21972
rect 12440 22024 12492 22030
rect 12440 21966 12492 21972
rect 13084 22024 13136 22030
rect 17408 22024 17460 22030
rect 13084 21966 13136 21972
rect 7472 21956 7524 21962
rect 7472 21898 7524 21904
rect 7564 21888 7616 21894
rect 7564 21830 7616 21836
rect 6630 21788 6938 21797
rect 6630 21786 6636 21788
rect 6692 21786 6716 21788
rect 6772 21786 6796 21788
rect 6852 21786 6876 21788
rect 6932 21786 6938 21788
rect 6692 21734 6694 21786
rect 6874 21734 6876 21786
rect 6630 21732 6636 21734
rect 6692 21732 6716 21734
rect 6772 21732 6796 21734
rect 6852 21732 6876 21734
rect 6932 21732 6938 21734
rect 6630 21723 6938 21732
rect 7104 21344 7156 21350
rect 7156 21292 7236 21298
rect 7104 21286 7236 21292
rect 7116 21270 7236 21286
rect 3790 21244 4098 21253
rect 3790 21242 3796 21244
rect 3852 21242 3876 21244
rect 3932 21242 3956 21244
rect 4012 21242 4036 21244
rect 4092 21242 4098 21244
rect 3852 21190 3854 21242
rect 4034 21190 4036 21242
rect 3790 21188 3796 21190
rect 3852 21188 3876 21190
rect 3932 21188 3956 21190
rect 4012 21188 4036 21190
rect 4092 21188 4098 21190
rect 3790 21179 4098 21188
rect 2504 21140 2556 21146
rect 2504 21082 2556 21088
rect 7104 21140 7156 21146
rect 7104 21082 7156 21088
rect 5540 20936 5592 20942
rect 5540 20878 5592 20884
rect 4896 20800 4948 20806
rect 4894 20768 4896 20777
rect 4948 20768 4950 20777
rect 4894 20703 4950 20712
rect 5552 20466 5580 20878
rect 6184 20868 6236 20874
rect 6184 20810 6236 20816
rect 4896 20460 4948 20466
rect 4896 20402 4948 20408
rect 5540 20460 5592 20466
rect 5540 20402 5592 20408
rect 4436 20256 4488 20262
rect 4436 20198 4488 20204
rect 3790 20156 4098 20165
rect 3790 20154 3796 20156
rect 3852 20154 3876 20156
rect 3932 20154 3956 20156
rect 4012 20154 4036 20156
rect 4092 20154 4098 20156
rect 3852 20102 3854 20154
rect 4034 20102 4036 20154
rect 3790 20100 3796 20102
rect 3852 20100 3876 20102
rect 3932 20100 3956 20102
rect 4012 20100 4036 20102
rect 4092 20100 4098 20102
rect 3790 20091 4098 20100
rect 4252 19780 4304 19786
rect 4252 19722 4304 19728
rect 2136 19712 2188 19718
rect 2136 19654 2188 19660
rect 1584 16108 1636 16114
rect 1584 16050 1636 16056
rect 1596 15706 1624 16050
rect 1584 15700 1636 15706
rect 1584 15642 1636 15648
rect 1952 15564 2004 15570
rect 1952 15506 2004 15512
rect 1860 15496 1912 15502
rect 1860 15438 1912 15444
rect 1872 15026 1900 15438
rect 1860 15020 1912 15026
rect 1860 14962 1912 14968
rect 1964 14822 1992 15506
rect 2044 14952 2096 14958
rect 2044 14894 2096 14900
rect 1860 14816 1912 14822
rect 1860 14758 1912 14764
rect 1952 14816 2004 14822
rect 1952 14758 2004 14764
rect 1768 14612 1820 14618
rect 1768 14554 1820 14560
rect 1584 14476 1636 14482
rect 1584 14418 1636 14424
rect 1596 12850 1624 14418
rect 1780 13938 1808 14554
rect 1872 14074 1900 14758
rect 1860 14068 1912 14074
rect 1860 14010 1912 14016
rect 1768 13932 1820 13938
rect 1768 13874 1820 13880
rect 1584 12844 1636 12850
rect 1584 12786 1636 12792
rect 1596 11354 1624 12786
rect 1780 12170 1808 13874
rect 1860 13320 1912 13326
rect 1860 13262 1912 13268
rect 1872 12986 1900 13262
rect 1860 12980 1912 12986
rect 1860 12922 1912 12928
rect 1964 12442 1992 14758
rect 2056 13326 2084 14894
rect 2148 14618 2176 19654
rect 3700 19508 3752 19514
rect 3700 19450 3752 19456
rect 3712 19417 3740 19450
rect 3698 19408 3754 19417
rect 3698 19343 3754 19352
rect 3790 19068 4098 19077
rect 3790 19066 3796 19068
rect 3852 19066 3876 19068
rect 3932 19066 3956 19068
rect 4012 19066 4036 19068
rect 4092 19066 4098 19068
rect 3852 19014 3854 19066
rect 4034 19014 4036 19066
rect 3790 19012 3796 19014
rect 3852 19012 3876 19014
rect 3932 19012 3956 19014
rect 4012 19012 4036 19014
rect 4092 19012 4098 19014
rect 3790 19003 4098 19012
rect 4264 18970 4292 19722
rect 4252 18964 4304 18970
rect 4252 18906 4304 18912
rect 2320 18760 2372 18766
rect 2320 18702 2372 18708
rect 2228 16992 2280 16998
rect 2228 16934 2280 16940
rect 2240 16726 2268 16934
rect 2228 16720 2280 16726
rect 2228 16662 2280 16668
rect 2136 14612 2188 14618
rect 2136 14554 2188 14560
rect 2136 13932 2188 13938
rect 2136 13874 2188 13880
rect 2044 13320 2096 13326
rect 2044 13262 2096 13268
rect 2148 12646 2176 13874
rect 2136 12640 2188 12646
rect 2136 12582 2188 12588
rect 1952 12436 2004 12442
rect 1952 12378 2004 12384
rect 1768 12164 1820 12170
rect 1768 12106 1820 12112
rect 1584 11348 1636 11354
rect 1584 11290 1636 11296
rect 1492 11076 1544 11082
rect 1492 11018 1544 11024
rect 1504 5846 1532 11018
rect 1596 10674 1624 11290
rect 1780 11286 1808 12106
rect 1768 11280 1820 11286
rect 1768 11222 1820 11228
rect 1584 10668 1636 10674
rect 1584 10610 1636 10616
rect 1596 9110 1624 10610
rect 1964 10554 1992 12378
rect 2044 12096 2096 12102
rect 2044 12038 2096 12044
rect 2056 11762 2084 12038
rect 2044 11756 2096 11762
rect 2044 11698 2096 11704
rect 1872 10526 1992 10554
rect 1584 9104 1636 9110
rect 1584 9046 1636 9052
rect 1596 6254 1624 9046
rect 1872 8294 1900 10526
rect 1952 10464 2004 10470
rect 1952 10406 2004 10412
rect 1964 9722 1992 10406
rect 1952 9716 2004 9722
rect 1952 9658 2004 9664
rect 1964 9518 1992 9658
rect 1952 9512 2004 9518
rect 1952 9454 2004 9460
rect 1964 8838 1992 9454
rect 2044 8968 2096 8974
rect 2044 8910 2096 8916
rect 1952 8832 2004 8838
rect 1952 8774 2004 8780
rect 1860 8288 1912 8294
rect 1860 8230 1912 8236
rect 1872 7342 1900 8230
rect 1964 8090 1992 8774
rect 2056 8634 2084 8910
rect 2044 8628 2096 8634
rect 2044 8570 2096 8576
rect 1952 8084 2004 8090
rect 1952 8026 2004 8032
rect 2148 7478 2176 12582
rect 2240 12238 2268 16662
rect 2332 16250 2360 18702
rect 4344 18284 4396 18290
rect 4344 18226 4396 18232
rect 3516 18080 3568 18086
rect 3516 18022 3568 18028
rect 2504 17604 2556 17610
rect 2504 17546 2556 17552
rect 2516 16794 2544 17546
rect 3424 17536 3476 17542
rect 3424 17478 3476 17484
rect 3240 17196 3292 17202
rect 3240 17138 3292 17144
rect 2504 16788 2556 16794
rect 2504 16730 2556 16736
rect 2504 16584 2556 16590
rect 2504 16526 2556 16532
rect 3056 16584 3108 16590
rect 3056 16526 3108 16532
rect 2320 16244 2372 16250
rect 2320 16186 2372 16192
rect 2516 15706 2544 16526
rect 2964 15972 3016 15978
rect 2964 15914 3016 15920
rect 2504 15700 2556 15706
rect 2504 15642 2556 15648
rect 2504 15360 2556 15366
rect 2504 15302 2556 15308
rect 2872 15360 2924 15366
rect 2872 15302 2924 15308
rect 2516 15094 2544 15302
rect 2504 15088 2556 15094
rect 2504 15030 2556 15036
rect 2516 14890 2544 15030
rect 2596 15020 2648 15026
rect 2596 14962 2648 14968
rect 2504 14884 2556 14890
rect 2504 14826 2556 14832
rect 2608 14618 2636 14962
rect 2688 14952 2740 14958
rect 2688 14894 2740 14900
rect 2700 14618 2728 14894
rect 2884 14822 2912 15302
rect 2872 14816 2924 14822
rect 2872 14758 2924 14764
rect 2596 14612 2648 14618
rect 2596 14554 2648 14560
rect 2688 14612 2740 14618
rect 2688 14554 2740 14560
rect 2412 14340 2464 14346
rect 2412 14282 2464 14288
rect 2424 14006 2452 14282
rect 2700 14074 2728 14554
rect 2884 14414 2912 14758
rect 2872 14408 2924 14414
rect 2872 14350 2924 14356
rect 2976 14346 3004 15914
rect 3068 15502 3096 16526
rect 3056 15496 3108 15502
rect 3056 15438 3108 15444
rect 2964 14340 3016 14346
rect 2964 14282 3016 14288
rect 2872 14272 2924 14278
rect 2872 14214 2924 14220
rect 2688 14068 2740 14074
rect 2688 14010 2740 14016
rect 2412 14000 2464 14006
rect 2412 13942 2464 13948
rect 2884 13938 2912 14214
rect 2872 13932 2924 13938
rect 2872 13874 2924 13880
rect 2688 13796 2740 13802
rect 2688 13738 2740 13744
rect 2504 13320 2556 13326
rect 2504 13262 2556 13268
rect 2516 12918 2544 13262
rect 2700 13258 2728 13738
rect 2688 13252 2740 13258
rect 2688 13194 2740 13200
rect 2596 13184 2648 13190
rect 2596 13126 2648 13132
rect 2608 12986 2636 13126
rect 2596 12980 2648 12986
rect 2596 12922 2648 12928
rect 2504 12912 2556 12918
rect 2504 12854 2556 12860
rect 2504 12640 2556 12646
rect 2504 12582 2556 12588
rect 2228 12232 2280 12238
rect 2228 12174 2280 12180
rect 2240 11082 2268 12174
rect 2412 11280 2464 11286
rect 2412 11222 2464 11228
rect 2228 11076 2280 11082
rect 2228 11018 2280 11024
rect 2228 10668 2280 10674
rect 2228 10610 2280 10616
rect 2240 10266 2268 10610
rect 2424 10266 2452 11222
rect 2516 11150 2544 12582
rect 2596 12096 2648 12102
rect 2596 12038 2648 12044
rect 2608 11762 2636 12038
rect 2596 11756 2648 11762
rect 2596 11698 2648 11704
rect 2608 11370 2636 11698
rect 2700 11506 2728 13194
rect 2780 13184 2832 13190
rect 2780 13126 2832 13132
rect 2792 11626 2820 13126
rect 2884 11694 2912 13874
rect 2964 12912 3016 12918
rect 2964 12854 3016 12860
rect 2976 11898 3004 12854
rect 3068 12102 3096 15438
rect 3148 15020 3200 15026
rect 3148 14962 3200 14968
rect 3160 14890 3188 14962
rect 3148 14884 3200 14890
rect 3148 14826 3200 14832
rect 3160 14618 3188 14826
rect 3148 14612 3200 14618
rect 3148 14554 3200 14560
rect 3148 13728 3200 13734
rect 3148 13670 3200 13676
rect 3160 12850 3188 13670
rect 3252 12986 3280 17138
rect 3436 16697 3464 17478
rect 3422 16688 3478 16697
rect 3422 16623 3478 16632
rect 3528 16590 3556 18022
rect 3790 17980 4098 17989
rect 3790 17978 3796 17980
rect 3852 17978 3876 17980
rect 3932 17978 3956 17980
rect 4012 17978 4036 17980
rect 4092 17978 4098 17980
rect 3852 17926 3854 17978
rect 4034 17926 4036 17978
rect 3790 17924 3796 17926
rect 3852 17924 3876 17926
rect 3932 17924 3956 17926
rect 4012 17924 4036 17926
rect 4092 17924 4098 17926
rect 3790 17915 4098 17924
rect 4252 17196 4304 17202
rect 4252 17138 4304 17144
rect 3790 16892 4098 16901
rect 3790 16890 3796 16892
rect 3852 16890 3876 16892
rect 3932 16890 3956 16892
rect 4012 16890 4036 16892
rect 4092 16890 4098 16892
rect 3852 16838 3854 16890
rect 4034 16838 4036 16890
rect 3790 16836 3796 16838
rect 3852 16836 3876 16838
rect 3932 16836 3956 16838
rect 4012 16836 4036 16838
rect 4092 16836 4098 16838
rect 3790 16827 4098 16836
rect 3516 16584 3568 16590
rect 3516 16526 3568 16532
rect 3700 16516 3752 16522
rect 3700 16458 3752 16464
rect 3712 16114 3740 16458
rect 3700 16108 3752 16114
rect 3700 16050 3752 16056
rect 3424 15564 3476 15570
rect 3424 15506 3476 15512
rect 3332 14884 3384 14890
rect 3332 14826 3384 14832
rect 3240 12980 3292 12986
rect 3240 12922 3292 12928
rect 3148 12844 3200 12850
rect 3148 12786 3200 12792
rect 3148 12708 3200 12714
rect 3148 12650 3200 12656
rect 3056 12096 3108 12102
rect 3056 12038 3108 12044
rect 2964 11892 3016 11898
rect 2964 11834 3016 11840
rect 2872 11688 2924 11694
rect 2872 11630 2924 11636
rect 2964 11688 3016 11694
rect 2964 11630 3016 11636
rect 2780 11620 2832 11626
rect 2780 11562 2832 11568
rect 2976 11506 3004 11630
rect 2700 11478 3004 11506
rect 3160 11370 3188 12650
rect 3240 11824 3292 11830
rect 3240 11766 3292 11772
rect 2608 11342 2820 11370
rect 2792 11150 2820 11342
rect 2976 11342 3188 11370
rect 2872 11212 2924 11218
rect 2872 11154 2924 11160
rect 2504 11144 2556 11150
rect 2504 11086 2556 11092
rect 2780 11144 2832 11150
rect 2780 11086 2832 11092
rect 2516 10470 2544 11086
rect 2780 11008 2832 11014
rect 2780 10950 2832 10956
rect 2792 10674 2820 10950
rect 2884 10810 2912 11154
rect 2872 10804 2924 10810
rect 2872 10746 2924 10752
rect 2780 10668 2832 10674
rect 2976 10656 3004 11342
rect 3148 11280 3200 11286
rect 3148 11222 3200 11228
rect 3056 11212 3108 11218
rect 3056 11154 3108 11160
rect 3068 10674 3096 11154
rect 2780 10610 2832 10616
rect 2884 10628 3004 10656
rect 3056 10668 3108 10674
rect 2504 10464 2556 10470
rect 2504 10406 2556 10412
rect 2228 10260 2280 10266
rect 2228 10202 2280 10208
rect 2412 10260 2464 10266
rect 2412 10202 2464 10208
rect 2424 9674 2452 10202
rect 2424 9646 2636 9674
rect 2608 9586 2636 9646
rect 2780 9648 2832 9654
rect 2780 9590 2832 9596
rect 2596 9580 2648 9586
rect 2596 9522 2648 9528
rect 2608 8838 2636 9522
rect 2688 9104 2740 9110
rect 2688 9046 2740 9052
rect 2596 8832 2648 8838
rect 2596 8774 2648 8780
rect 2608 8498 2636 8774
rect 2700 8634 2728 9046
rect 2688 8628 2740 8634
rect 2688 8570 2740 8576
rect 2792 8566 2820 9590
rect 2884 9110 2912 10628
rect 3056 10610 3108 10616
rect 3160 10554 3188 11222
rect 3252 11218 3280 11766
rect 3240 11212 3292 11218
rect 3240 11154 3292 11160
rect 2964 10532 3016 10538
rect 2964 10474 3016 10480
rect 3068 10526 3188 10554
rect 3238 10568 3294 10577
rect 2872 9104 2924 9110
rect 2872 9046 2924 9052
rect 2976 9042 3004 10474
rect 3068 9382 3096 10526
rect 3238 10503 3240 10512
rect 3292 10503 3294 10512
rect 3240 10474 3292 10480
rect 3148 10464 3200 10470
rect 3148 10406 3200 10412
rect 3056 9376 3108 9382
rect 3056 9318 3108 9324
rect 2964 9036 3016 9042
rect 2964 8978 3016 8984
rect 2872 8968 2924 8974
rect 2872 8910 2924 8916
rect 3056 8968 3108 8974
rect 3056 8910 3108 8916
rect 2780 8560 2832 8566
rect 2780 8502 2832 8508
rect 2320 8492 2372 8498
rect 2320 8434 2372 8440
rect 2596 8492 2648 8498
rect 2596 8434 2648 8440
rect 2332 7886 2360 8434
rect 2504 8424 2556 8430
rect 2504 8366 2556 8372
rect 2516 7886 2544 8366
rect 2792 8022 2820 8502
rect 2884 8090 2912 8910
rect 2872 8084 2924 8090
rect 2872 8026 2924 8032
rect 2780 8016 2832 8022
rect 2780 7958 2832 7964
rect 2320 7880 2372 7886
rect 2320 7822 2372 7828
rect 2504 7880 2556 7886
rect 2504 7822 2556 7828
rect 2688 7880 2740 7886
rect 2688 7822 2740 7828
rect 2136 7472 2188 7478
rect 2136 7414 2188 7420
rect 1860 7336 1912 7342
rect 1860 7278 1912 7284
rect 1768 6996 1820 7002
rect 1768 6938 1820 6944
rect 1780 6322 1808 6938
rect 1872 6390 1900 7278
rect 2044 7200 2096 7206
rect 2044 7142 2096 7148
rect 1860 6384 1912 6390
rect 1860 6326 1912 6332
rect 1768 6316 1820 6322
rect 1768 6258 1820 6264
rect 1952 6316 2004 6322
rect 1952 6258 2004 6264
rect 1584 6248 1636 6254
rect 1584 6190 1636 6196
rect 1492 5840 1544 5846
rect 1492 5782 1544 5788
rect 1596 5778 1624 6190
rect 1584 5772 1636 5778
rect 1584 5714 1636 5720
rect 1964 5710 1992 6258
rect 2056 6254 2084 7142
rect 2148 6730 2176 7414
rect 2136 6724 2188 6730
rect 2136 6666 2188 6672
rect 2148 6390 2176 6666
rect 2228 6656 2280 6662
rect 2228 6598 2280 6604
rect 2136 6384 2188 6390
rect 2136 6326 2188 6332
rect 2044 6248 2096 6254
rect 2044 6190 2096 6196
rect 2044 6112 2096 6118
rect 2044 6054 2096 6060
rect 1952 5704 2004 5710
rect 1952 5646 2004 5652
rect 1676 4820 1728 4826
rect 1676 4762 1728 4768
rect 1688 4282 1716 4762
rect 2056 4622 2084 6054
rect 2148 5302 2176 6326
rect 2240 5710 2268 6598
rect 2228 5704 2280 5710
rect 2228 5646 2280 5652
rect 2332 5642 2360 7822
rect 2412 7404 2464 7410
rect 2516 7392 2544 7822
rect 2700 7478 2728 7822
rect 2688 7472 2740 7478
rect 2688 7414 2740 7420
rect 2792 7410 2820 7958
rect 2464 7364 2544 7392
rect 2412 7346 2464 7352
rect 2516 7206 2544 7364
rect 2780 7404 2832 7410
rect 2780 7346 2832 7352
rect 2504 7200 2556 7206
rect 2504 7142 2556 7148
rect 2516 6914 2544 7142
rect 2516 6886 2728 6914
rect 2700 6662 2728 6886
rect 2688 6656 2740 6662
rect 2688 6598 2740 6604
rect 2700 5778 2728 6598
rect 2688 5772 2740 5778
rect 2688 5714 2740 5720
rect 2320 5636 2372 5642
rect 2320 5578 2372 5584
rect 2228 5568 2280 5574
rect 2228 5510 2280 5516
rect 2136 5296 2188 5302
rect 2136 5238 2188 5244
rect 2240 5234 2268 5510
rect 2228 5228 2280 5234
rect 2228 5170 2280 5176
rect 2332 5098 2360 5578
rect 2504 5568 2556 5574
rect 2504 5510 2556 5516
rect 2320 5092 2372 5098
rect 2320 5034 2372 5040
rect 2332 4826 2360 5034
rect 2516 4826 2544 5510
rect 2792 5370 2820 7346
rect 3068 7342 3096 8910
rect 3160 7546 3188 10406
rect 3344 10062 3372 14826
rect 3436 11286 3464 15506
rect 3712 15026 3740 16050
rect 4160 16040 4212 16046
rect 4160 15982 4212 15988
rect 3790 15804 4098 15813
rect 3790 15802 3796 15804
rect 3852 15802 3876 15804
rect 3932 15802 3956 15804
rect 4012 15802 4036 15804
rect 4092 15802 4098 15804
rect 3852 15750 3854 15802
rect 4034 15750 4036 15802
rect 3790 15748 3796 15750
rect 3852 15748 3876 15750
rect 3932 15748 3956 15750
rect 4012 15748 4036 15750
rect 4092 15748 4098 15750
rect 3790 15739 4098 15748
rect 4172 15434 4200 15982
rect 4160 15428 4212 15434
rect 4160 15370 4212 15376
rect 3976 15360 4028 15366
rect 3976 15302 4028 15308
rect 3516 15020 3568 15026
rect 3516 14962 3568 14968
rect 3700 15020 3752 15026
rect 3700 14962 3752 14968
rect 3528 13530 3556 14962
rect 3988 14958 4016 15302
rect 3976 14952 4028 14958
rect 3976 14894 4028 14900
rect 3700 14816 3752 14822
rect 3700 14758 3752 14764
rect 3712 14482 3740 14758
rect 3790 14716 4098 14725
rect 3790 14714 3796 14716
rect 3852 14714 3876 14716
rect 3932 14714 3956 14716
rect 4012 14714 4036 14716
rect 4092 14714 4098 14716
rect 3852 14662 3854 14714
rect 4034 14662 4036 14714
rect 3790 14660 3796 14662
rect 3852 14660 3876 14662
rect 3932 14660 3956 14662
rect 4012 14660 4036 14662
rect 4092 14660 4098 14662
rect 3790 14651 4098 14660
rect 4172 14618 4200 15370
rect 4264 15162 4292 17138
rect 4356 15162 4384 18226
rect 4252 15156 4304 15162
rect 4252 15098 4304 15104
rect 4344 15156 4396 15162
rect 4344 15098 4396 15104
rect 4448 15065 4476 20198
rect 4620 18080 4672 18086
rect 4620 18022 4672 18028
rect 4632 17678 4660 18022
rect 4620 17672 4672 17678
rect 4620 17614 4672 17620
rect 4632 17270 4660 17614
rect 4620 17264 4672 17270
rect 4620 17206 4672 17212
rect 4632 16658 4660 17206
rect 4620 16652 4672 16658
rect 4620 16594 4672 16600
rect 4632 16250 4660 16594
rect 4712 16448 4764 16454
rect 4712 16390 4764 16396
rect 4620 16244 4672 16250
rect 4620 16186 4672 16192
rect 4632 15502 4660 16186
rect 4724 15706 4752 16390
rect 4804 15904 4856 15910
rect 4804 15846 4856 15852
rect 4712 15700 4764 15706
rect 4712 15642 4764 15648
rect 4528 15496 4580 15502
rect 4528 15438 4580 15444
rect 4620 15496 4672 15502
rect 4620 15438 4672 15444
rect 4540 15162 4568 15438
rect 4724 15178 4752 15642
rect 4816 15434 4844 15846
rect 4804 15428 4856 15434
rect 4804 15370 4856 15376
rect 4528 15156 4580 15162
rect 4528 15098 4580 15104
rect 4632 15150 4752 15178
rect 4434 15056 4490 15065
rect 4632 15026 4660 15150
rect 4434 14991 4490 15000
rect 4528 15020 4580 15026
rect 4160 14612 4212 14618
rect 4160 14554 4212 14560
rect 3976 14544 4028 14550
rect 4344 14544 4396 14550
rect 4028 14492 4108 14498
rect 3976 14486 4108 14492
rect 3700 14476 3752 14482
rect 3988 14470 4108 14486
rect 3700 14418 3752 14424
rect 3700 14340 3752 14346
rect 3700 14282 3752 14288
rect 3608 14000 3660 14006
rect 3608 13942 3660 13948
rect 3516 13524 3568 13530
rect 3516 13466 3568 13472
rect 3620 12850 3648 13942
rect 3608 12844 3660 12850
rect 3608 12786 3660 12792
rect 3516 12776 3568 12782
rect 3516 12718 3568 12724
rect 3528 12434 3556 12718
rect 3528 12406 3648 12434
rect 3620 11558 3648 12406
rect 3608 11552 3660 11558
rect 3608 11494 3660 11500
rect 3424 11280 3476 11286
rect 3424 11222 3476 11228
rect 3424 11144 3476 11150
rect 3424 11086 3476 11092
rect 3332 10056 3384 10062
rect 3332 9998 3384 10004
rect 3240 9444 3292 9450
rect 3240 9386 3292 9392
rect 3252 8974 3280 9386
rect 3240 8968 3292 8974
rect 3240 8910 3292 8916
rect 3240 8492 3292 8498
rect 3240 8434 3292 8440
rect 3252 7546 3280 8434
rect 3148 7540 3200 7546
rect 3148 7482 3200 7488
rect 3240 7540 3292 7546
rect 3240 7482 3292 7488
rect 2872 7336 2924 7342
rect 2872 7278 2924 7284
rect 3056 7336 3108 7342
rect 3056 7278 3108 7284
rect 2884 6934 2912 7278
rect 2872 6928 2924 6934
rect 2872 6870 2924 6876
rect 2780 5364 2832 5370
rect 2780 5306 2832 5312
rect 2792 5166 2820 5306
rect 2780 5160 2832 5166
rect 2780 5102 2832 5108
rect 2320 4820 2372 4826
rect 2320 4762 2372 4768
rect 2504 4820 2556 4826
rect 2504 4762 2556 4768
rect 2792 4622 2820 5102
rect 2044 4616 2096 4622
rect 2044 4558 2096 4564
rect 2780 4616 2832 4622
rect 2780 4558 2832 4564
rect 1676 4276 1728 4282
rect 1676 4218 1728 4224
rect 1688 3194 1716 4218
rect 2056 4146 2084 4558
rect 2870 4176 2926 4185
rect 2044 4140 2096 4146
rect 2870 4111 2872 4120
rect 2044 4082 2096 4088
rect 2924 4111 2926 4120
rect 2872 4082 2924 4088
rect 2502 4040 2558 4049
rect 2502 3975 2558 3984
rect 1676 3188 1728 3194
rect 1676 3130 1728 3136
rect 2516 3058 2544 3975
rect 2884 3466 2912 4082
rect 3160 3602 3188 7482
rect 3344 6798 3372 9998
rect 3436 9178 3464 11086
rect 3620 10742 3648 11494
rect 3712 10810 3740 14282
rect 4080 13784 4108 14470
rect 4172 14492 4344 14498
rect 4172 14486 4396 14492
rect 4172 14470 4384 14486
rect 4172 13938 4200 14470
rect 4252 14272 4304 14278
rect 4252 14214 4304 14220
rect 4160 13932 4212 13938
rect 4160 13874 4212 13880
rect 4080 13756 4200 13784
rect 3790 13628 4098 13637
rect 3790 13626 3796 13628
rect 3852 13626 3876 13628
rect 3932 13626 3956 13628
rect 4012 13626 4036 13628
rect 4092 13626 4098 13628
rect 3852 13574 3854 13626
rect 4034 13574 4036 13626
rect 3790 13572 3796 13574
rect 3852 13572 3876 13574
rect 3932 13572 3956 13574
rect 4012 13572 4036 13574
rect 4092 13572 4098 13574
rect 3790 13563 4098 13572
rect 4172 13410 4200 13756
rect 4264 13462 4292 14214
rect 4080 13382 4200 13410
rect 4252 13456 4304 13462
rect 4252 13398 4304 13404
rect 3792 13320 3844 13326
rect 3792 13262 3844 13268
rect 3804 12850 3832 13262
rect 4080 12850 4108 13382
rect 4356 13258 4384 14470
rect 4448 13938 4476 14991
rect 4528 14962 4580 14968
rect 4620 15020 4672 15026
rect 4804 15020 4856 15026
rect 4620 14962 4672 14968
rect 4724 14980 4804 15008
rect 4540 14006 4568 14962
rect 4528 14000 4580 14006
rect 4528 13942 4580 13948
rect 4436 13932 4488 13938
rect 4436 13874 4488 13880
rect 4526 13832 4582 13841
rect 4526 13767 4582 13776
rect 4436 13524 4488 13530
rect 4436 13466 4488 13472
rect 4344 13252 4396 13258
rect 4344 13194 4396 13200
rect 3792 12844 3844 12850
rect 3792 12786 3844 12792
rect 4068 12844 4120 12850
rect 4068 12786 4120 12792
rect 4160 12708 4212 12714
rect 4160 12650 4212 12656
rect 3790 12540 4098 12549
rect 3790 12538 3796 12540
rect 3852 12538 3876 12540
rect 3932 12538 3956 12540
rect 4012 12538 4036 12540
rect 4092 12538 4098 12540
rect 3852 12486 3854 12538
rect 4034 12486 4036 12538
rect 3790 12484 3796 12486
rect 3852 12484 3876 12486
rect 3932 12484 3956 12486
rect 4012 12484 4036 12486
rect 4092 12484 4098 12486
rect 3790 12475 4098 12484
rect 4172 11762 4200 12650
rect 4356 12646 4384 13194
rect 4344 12640 4396 12646
rect 4344 12582 4396 12588
rect 4448 12434 4476 13466
rect 4540 12986 4568 13767
rect 4632 13530 4660 14962
rect 4724 13530 4752 14980
rect 4804 14962 4856 14968
rect 4908 14074 4936 20402
rect 5552 19854 5580 20402
rect 5540 19848 5592 19854
rect 5540 19790 5592 19796
rect 5552 19378 5580 19790
rect 5908 19440 5960 19446
rect 5908 19382 5960 19388
rect 5540 19372 5592 19378
rect 5540 19314 5592 19320
rect 5552 18766 5580 19314
rect 5540 18760 5592 18766
rect 5540 18702 5592 18708
rect 5080 18624 5132 18630
rect 5080 18566 5132 18572
rect 4988 15360 5040 15366
rect 4988 15302 5040 15308
rect 5000 14550 5028 15302
rect 4988 14544 5040 14550
rect 4988 14486 5040 14492
rect 5092 14113 5120 18566
rect 5552 17882 5580 18702
rect 5540 17876 5592 17882
rect 5540 17818 5592 17824
rect 5356 16992 5408 16998
rect 5356 16934 5408 16940
rect 5172 16108 5224 16114
rect 5172 16050 5224 16056
rect 5184 15094 5212 16050
rect 5264 15428 5316 15434
rect 5264 15370 5316 15376
rect 5172 15088 5224 15094
rect 5172 15030 5224 15036
rect 5276 14634 5304 15370
rect 5368 14822 5396 16934
rect 5540 16788 5592 16794
rect 5540 16730 5592 16736
rect 5448 15632 5500 15638
rect 5448 15574 5500 15580
rect 5460 15366 5488 15574
rect 5448 15360 5500 15366
rect 5448 15302 5500 15308
rect 5552 15162 5580 16730
rect 5920 16250 5948 19382
rect 6092 18692 6144 18698
rect 6092 18634 6144 18640
rect 6000 17536 6052 17542
rect 6000 17478 6052 17484
rect 5908 16244 5960 16250
rect 5908 16186 5960 16192
rect 6012 16114 6040 17478
rect 5724 16108 5776 16114
rect 5644 16068 5724 16096
rect 5540 15156 5592 15162
rect 5540 15098 5592 15104
rect 5448 15020 5500 15026
rect 5644 15008 5672 16068
rect 6000 16108 6052 16114
rect 5776 16068 6000 16096
rect 5724 16050 5776 16056
rect 6000 16050 6052 16056
rect 5816 15972 5868 15978
rect 5816 15914 5868 15920
rect 5500 14980 5672 15008
rect 5448 14962 5500 14968
rect 5356 14816 5408 14822
rect 5356 14758 5408 14764
rect 5184 14606 5304 14634
rect 5644 14618 5672 14980
rect 5632 14612 5684 14618
rect 5078 14104 5134 14113
rect 4896 14068 4948 14074
rect 5078 14039 5134 14048
rect 4896 14010 4948 14016
rect 5184 14006 5212 14606
rect 5632 14554 5684 14560
rect 5264 14544 5316 14550
rect 5264 14486 5316 14492
rect 5172 14000 5224 14006
rect 5000 13960 5172 13988
rect 4804 13728 4856 13734
rect 4804 13670 4856 13676
rect 4620 13524 4672 13530
rect 4620 13466 4672 13472
rect 4712 13524 4764 13530
rect 4712 13466 4764 13472
rect 4528 12980 4580 12986
rect 4528 12922 4580 12928
rect 4540 12714 4568 12922
rect 4712 12844 4764 12850
rect 4712 12786 4764 12792
rect 4528 12708 4580 12714
rect 4528 12650 4580 12656
rect 4540 12617 4568 12650
rect 4526 12608 4582 12617
rect 4526 12543 4582 12552
rect 4356 12406 4476 12434
rect 4356 12238 4384 12406
rect 4724 12306 4752 12786
rect 4712 12300 4764 12306
rect 4712 12242 4764 12248
rect 4344 12232 4396 12238
rect 4344 12174 4396 12180
rect 4250 11928 4306 11937
rect 4250 11863 4252 11872
rect 4304 11863 4306 11872
rect 4252 11834 4304 11840
rect 4160 11756 4212 11762
rect 4160 11698 4212 11704
rect 3790 11452 4098 11461
rect 3790 11450 3796 11452
rect 3852 11450 3876 11452
rect 3932 11450 3956 11452
rect 4012 11450 4036 11452
rect 4092 11450 4098 11452
rect 3852 11398 3854 11450
rect 4034 11398 4036 11450
rect 3790 11396 3796 11398
rect 3852 11396 3876 11398
rect 3932 11396 3956 11398
rect 4012 11396 4036 11398
rect 4092 11396 4098 11398
rect 3790 11387 4098 11396
rect 4068 11144 4120 11150
rect 4172 11132 4200 11698
rect 4356 11150 4384 12174
rect 4724 11898 4752 12242
rect 4712 11892 4764 11898
rect 4712 11834 4764 11840
rect 4816 11762 4844 13670
rect 4896 13388 4948 13394
rect 5000 13376 5028 13960
rect 5172 13942 5224 13948
rect 4948 13348 5028 13376
rect 4896 13330 4948 13336
rect 4804 11756 4856 11762
rect 4804 11698 4856 11704
rect 4120 11104 4200 11132
rect 4068 11086 4120 11092
rect 3700 10804 3752 10810
rect 3700 10746 3752 10752
rect 3608 10736 3660 10742
rect 3608 10678 3660 10684
rect 3516 10532 3568 10538
rect 3516 10474 3568 10480
rect 3528 10130 3556 10474
rect 3516 10124 3568 10130
rect 3516 10066 3568 10072
rect 3528 9654 3556 10066
rect 3516 9648 3568 9654
rect 3516 9590 3568 9596
rect 3424 9172 3476 9178
rect 3424 9114 3476 9120
rect 3332 6792 3384 6798
rect 3332 6734 3384 6740
rect 3344 5234 3372 6734
rect 3436 6730 3464 9114
rect 3516 9036 3568 9042
rect 3516 8978 3568 8984
rect 3528 8090 3556 8978
rect 3620 8498 3648 10678
rect 3700 10668 3752 10674
rect 3700 10610 3752 10616
rect 3712 10266 3740 10610
rect 3790 10364 4098 10373
rect 3790 10362 3796 10364
rect 3852 10362 3876 10364
rect 3932 10362 3956 10364
rect 4012 10362 4036 10364
rect 4092 10362 4098 10364
rect 3852 10310 3854 10362
rect 4034 10310 4036 10362
rect 3790 10308 3796 10310
rect 3852 10308 3876 10310
rect 3932 10308 3956 10310
rect 4012 10308 4036 10310
rect 4092 10308 4098 10310
rect 3790 10299 4098 10308
rect 3700 10260 3752 10266
rect 3700 10202 3752 10208
rect 4172 10044 4200 11104
rect 4344 11144 4396 11150
rect 4344 11086 4396 11092
rect 4252 11008 4304 11014
rect 4252 10950 4304 10956
rect 4264 10470 4292 10950
rect 4252 10464 4304 10470
rect 4252 10406 4304 10412
rect 4252 10056 4304 10062
rect 4172 10016 4252 10044
rect 4252 9998 4304 10004
rect 4160 9920 4212 9926
rect 4160 9862 4212 9868
rect 3700 9376 3752 9382
rect 3700 9318 3752 9324
rect 3608 8492 3660 8498
rect 3608 8434 3660 8440
rect 3516 8084 3568 8090
rect 3516 8026 3568 8032
rect 3516 7880 3568 7886
rect 3620 7868 3648 8434
rect 3712 8362 3740 9318
rect 3790 9276 4098 9285
rect 3790 9274 3796 9276
rect 3852 9274 3876 9276
rect 3932 9274 3956 9276
rect 4012 9274 4036 9276
rect 4092 9274 4098 9276
rect 3852 9222 3854 9274
rect 4034 9222 4036 9274
rect 3790 9220 3796 9222
rect 3852 9220 3876 9222
rect 3932 9220 3956 9222
rect 4012 9220 4036 9222
rect 4092 9220 4098 9222
rect 3790 9211 4098 9220
rect 3976 9172 4028 9178
rect 3976 9114 4028 9120
rect 3792 8900 3844 8906
rect 3792 8842 3844 8848
rect 3804 8634 3832 8842
rect 3792 8628 3844 8634
rect 3792 8570 3844 8576
rect 3988 8498 4016 9114
rect 3976 8492 4028 8498
rect 3976 8434 4028 8440
rect 3700 8356 3752 8362
rect 3700 8298 3752 8304
rect 3790 8188 4098 8197
rect 3790 8186 3796 8188
rect 3852 8186 3876 8188
rect 3932 8186 3956 8188
rect 4012 8186 4036 8188
rect 4092 8186 4098 8188
rect 3852 8134 3854 8186
rect 4034 8134 4036 8186
rect 3790 8132 3796 8134
rect 3852 8132 3876 8134
rect 3932 8132 3956 8134
rect 4012 8132 4036 8134
rect 4092 8132 4098 8134
rect 3790 8123 4098 8132
rect 3568 7840 3648 7868
rect 3516 7822 3568 7828
rect 3528 7410 3556 7822
rect 3516 7404 3568 7410
rect 3516 7346 3568 7352
rect 3528 7002 3556 7346
rect 3700 7200 3752 7206
rect 3700 7142 3752 7148
rect 3712 7002 3740 7142
rect 3790 7100 4098 7109
rect 3790 7098 3796 7100
rect 3852 7098 3876 7100
rect 3932 7098 3956 7100
rect 4012 7098 4036 7100
rect 4092 7098 4098 7100
rect 3852 7046 3854 7098
rect 4034 7046 4036 7098
rect 3790 7044 3796 7046
rect 3852 7044 3876 7046
rect 3932 7044 3956 7046
rect 4012 7044 4036 7046
rect 4092 7044 4098 7046
rect 3790 7035 4098 7044
rect 3516 6996 3568 7002
rect 3516 6938 3568 6944
rect 3700 6996 3752 7002
rect 3700 6938 3752 6944
rect 3424 6724 3476 6730
rect 3424 6666 3476 6672
rect 3436 6458 3464 6666
rect 3424 6452 3476 6458
rect 3424 6394 3476 6400
rect 3528 5370 3556 6938
rect 3608 6384 3660 6390
rect 3608 6326 3660 6332
rect 3620 5710 3648 6326
rect 3712 6270 3740 6938
rect 3712 6242 3832 6270
rect 3804 6186 3832 6242
rect 3700 6180 3752 6186
rect 3700 6122 3752 6128
rect 3792 6180 3844 6186
rect 3792 6122 3844 6128
rect 3608 5704 3660 5710
rect 3608 5646 3660 5652
rect 3424 5364 3476 5370
rect 3424 5306 3476 5312
rect 3516 5364 3568 5370
rect 3516 5306 3568 5312
rect 3332 5228 3384 5234
rect 3332 5170 3384 5176
rect 3436 4758 3464 5306
rect 3240 4752 3292 4758
rect 3240 4694 3292 4700
rect 3424 4752 3476 4758
rect 3424 4694 3476 4700
rect 3252 4486 3280 4694
rect 3240 4480 3292 4486
rect 3240 4422 3292 4428
rect 3436 4146 3464 4694
rect 3620 4622 3648 5646
rect 3712 5166 3740 6122
rect 3790 6012 4098 6021
rect 3790 6010 3796 6012
rect 3852 6010 3876 6012
rect 3932 6010 3956 6012
rect 4012 6010 4036 6012
rect 4092 6010 4098 6012
rect 3852 5958 3854 6010
rect 4034 5958 4036 6010
rect 3790 5956 3796 5958
rect 3852 5956 3876 5958
rect 3932 5956 3956 5958
rect 4012 5956 4036 5958
rect 4092 5956 4098 5958
rect 3790 5947 4098 5956
rect 3700 5160 3752 5166
rect 3700 5102 3752 5108
rect 3790 4924 4098 4933
rect 3790 4922 3796 4924
rect 3852 4922 3876 4924
rect 3932 4922 3956 4924
rect 4012 4922 4036 4924
rect 4092 4922 4098 4924
rect 3852 4870 3854 4922
rect 4034 4870 4036 4922
rect 3790 4868 3796 4870
rect 3852 4868 3876 4870
rect 3932 4868 3956 4870
rect 4012 4868 4036 4870
rect 4092 4868 4098 4870
rect 3790 4859 4098 4868
rect 4068 4820 4120 4826
rect 4068 4762 4120 4768
rect 4080 4729 4108 4762
rect 4066 4720 4122 4729
rect 4066 4655 4122 4664
rect 3608 4616 3660 4622
rect 3608 4558 3660 4564
rect 4068 4616 4120 4622
rect 4068 4558 4120 4564
rect 4080 4282 4108 4558
rect 4068 4276 4120 4282
rect 4068 4218 4120 4224
rect 3424 4140 3476 4146
rect 3424 4082 3476 4088
rect 4172 4010 4200 9862
rect 4264 9722 4292 9998
rect 4356 9994 4384 11086
rect 4620 10736 4672 10742
rect 4620 10678 4672 10684
rect 4528 10668 4580 10674
rect 4528 10610 4580 10616
rect 4540 10198 4568 10610
rect 4632 10198 4660 10678
rect 4816 10674 4844 11698
rect 5000 11082 5028 13348
rect 5080 13320 5132 13326
rect 5080 13262 5132 13268
rect 5170 13288 5226 13297
rect 5092 11082 5120 13262
rect 5170 13223 5172 13232
rect 5224 13223 5226 13232
rect 5172 13194 5224 13200
rect 5184 12374 5212 13194
rect 5276 13190 5304 14486
rect 5724 14476 5776 14482
rect 5724 14418 5776 14424
rect 5448 14408 5500 14414
rect 5448 14350 5500 14356
rect 5356 14340 5408 14346
rect 5356 14282 5408 14288
rect 5368 13802 5396 14282
rect 5460 13802 5488 14350
rect 5736 14006 5764 14418
rect 5828 14278 5856 15914
rect 5908 15360 5960 15366
rect 5908 15302 5960 15308
rect 5816 14272 5868 14278
rect 5816 14214 5868 14220
rect 5724 14000 5776 14006
rect 5724 13942 5776 13948
rect 5356 13796 5408 13802
rect 5356 13738 5408 13744
rect 5448 13796 5500 13802
rect 5448 13738 5500 13744
rect 5368 13326 5396 13738
rect 5356 13320 5408 13326
rect 5356 13262 5408 13268
rect 5264 13184 5316 13190
rect 5264 13126 5316 13132
rect 5172 12368 5224 12374
rect 5172 12310 5224 12316
rect 5172 12232 5224 12238
rect 5172 12174 5224 12180
rect 5184 11626 5212 12174
rect 5172 11620 5224 11626
rect 5172 11562 5224 11568
rect 4988 11076 5040 11082
rect 4988 11018 5040 11024
rect 5080 11076 5132 11082
rect 5080 11018 5132 11024
rect 4804 10668 4856 10674
rect 4804 10610 4856 10616
rect 5000 10470 5028 11018
rect 4988 10464 5040 10470
rect 4908 10424 4988 10452
rect 4528 10192 4580 10198
rect 4528 10134 4580 10140
rect 4620 10192 4672 10198
rect 4620 10134 4672 10140
rect 4344 9988 4396 9994
rect 4344 9930 4396 9936
rect 4252 9716 4304 9722
rect 4252 9658 4304 9664
rect 4264 9382 4292 9658
rect 4344 9580 4396 9586
rect 4344 9522 4396 9528
rect 4356 9489 4384 9522
rect 4342 9480 4398 9489
rect 4342 9415 4398 9424
rect 4252 9376 4304 9382
rect 4252 9318 4304 9324
rect 4356 8974 4384 9415
rect 4344 8968 4396 8974
rect 4344 8910 4396 8916
rect 4356 8498 4384 8910
rect 4344 8492 4396 8498
rect 4344 8434 4396 8440
rect 4356 8090 4384 8434
rect 4344 8084 4396 8090
rect 4344 8026 4396 8032
rect 4540 7970 4568 10134
rect 4908 10130 4936 10424
rect 4988 10406 5040 10412
rect 5092 10266 5120 11018
rect 5080 10260 5132 10266
rect 5080 10202 5132 10208
rect 4896 10124 4948 10130
rect 4896 10066 4948 10072
rect 4988 10124 5040 10130
rect 4988 10066 5040 10072
rect 5000 9994 5028 10066
rect 5080 10056 5132 10062
rect 5080 9998 5132 10004
rect 4988 9988 5040 9994
rect 4988 9930 5040 9936
rect 4804 9920 4856 9926
rect 4804 9862 4856 9868
rect 4620 8832 4672 8838
rect 4620 8774 4672 8780
rect 4252 7948 4304 7954
rect 4252 7890 4304 7896
rect 4448 7942 4568 7970
rect 4264 6254 4292 7890
rect 4344 6724 4396 6730
rect 4344 6666 4396 6672
rect 4356 6458 4384 6666
rect 4344 6452 4396 6458
rect 4344 6394 4396 6400
rect 4252 6248 4304 6254
rect 4252 6190 4304 6196
rect 4448 5574 4476 7942
rect 4528 7200 4580 7206
rect 4528 7142 4580 7148
rect 4540 6798 4568 7142
rect 4528 6792 4580 6798
rect 4528 6734 4580 6740
rect 4540 6390 4568 6734
rect 4528 6384 4580 6390
rect 4528 6326 4580 6332
rect 4632 5778 4660 8774
rect 4712 8628 4764 8634
rect 4712 8570 4764 8576
rect 4724 8022 4752 8570
rect 4712 8016 4764 8022
rect 4712 7958 4764 7964
rect 4816 7868 4844 9862
rect 5000 9586 5028 9930
rect 4988 9580 5040 9586
rect 4988 9522 5040 9528
rect 5000 9110 5028 9522
rect 5092 9518 5120 9998
rect 5080 9512 5132 9518
rect 5132 9472 5212 9500
rect 5080 9454 5132 9460
rect 4988 9104 5040 9110
rect 4988 9046 5040 9052
rect 4894 8936 4950 8945
rect 4894 8871 4950 8880
rect 4908 8838 4936 8871
rect 4896 8832 4948 8838
rect 4896 8774 4948 8780
rect 4896 8492 4948 8498
rect 4896 8434 4948 8440
rect 4724 7840 4844 7868
rect 4620 5772 4672 5778
rect 4620 5714 4672 5720
rect 4724 5658 4752 7840
rect 4802 7440 4858 7449
rect 4802 7375 4804 7384
rect 4856 7375 4858 7384
rect 4804 7346 4856 7352
rect 4908 6934 4936 8434
rect 4896 6928 4948 6934
rect 4896 6870 4948 6876
rect 4802 6760 4858 6769
rect 4802 6695 4804 6704
rect 4856 6695 4858 6704
rect 4804 6666 4856 6672
rect 4908 6458 4936 6870
rect 4896 6452 4948 6458
rect 4896 6394 4948 6400
rect 4896 6180 4948 6186
rect 4896 6122 4948 6128
rect 4908 5710 4936 6122
rect 4632 5630 4752 5658
rect 4896 5704 4948 5710
rect 4896 5646 4948 5652
rect 4252 5568 4304 5574
rect 4252 5510 4304 5516
rect 4436 5568 4488 5574
rect 4436 5510 4488 5516
rect 4264 4690 4292 5510
rect 4252 4684 4304 4690
rect 4252 4626 4304 4632
rect 4160 4004 4212 4010
rect 4160 3946 4212 3952
rect 3790 3836 4098 3845
rect 3790 3834 3796 3836
rect 3852 3834 3876 3836
rect 3932 3834 3956 3836
rect 4012 3834 4036 3836
rect 4092 3834 4098 3836
rect 3852 3782 3854 3834
rect 4034 3782 4036 3834
rect 3790 3780 3796 3782
rect 3852 3780 3876 3782
rect 3932 3780 3956 3782
rect 4012 3780 4036 3782
rect 4092 3780 4098 3782
rect 3790 3771 4098 3780
rect 4264 3738 4292 4626
rect 4344 4140 4396 4146
rect 4344 4082 4396 4088
rect 4160 3732 4212 3738
rect 4160 3674 4212 3680
rect 4252 3732 4304 3738
rect 4252 3674 4304 3680
rect 4172 3618 4200 3674
rect 4356 3618 4384 4082
rect 3148 3596 3200 3602
rect 4172 3590 4384 3618
rect 3148 3538 3200 3544
rect 4448 3534 4476 5510
rect 4632 4554 4660 5630
rect 4712 5228 4764 5234
rect 4712 5170 4764 5176
rect 4724 4758 4752 5170
rect 4712 4752 4764 4758
rect 4712 4694 4764 4700
rect 4528 4548 4580 4554
rect 4528 4490 4580 4496
rect 4620 4548 4672 4554
rect 4620 4490 4672 4496
rect 4540 3738 4568 4490
rect 4724 4434 4752 4694
rect 4632 4406 4752 4434
rect 4528 3732 4580 3738
rect 4528 3674 4580 3680
rect 3424 3528 3476 3534
rect 3422 3496 3424 3505
rect 4436 3528 4488 3534
rect 3476 3496 3478 3505
rect 2872 3460 2924 3466
rect 4436 3470 4488 3476
rect 3422 3431 3478 3440
rect 2872 3402 2924 3408
rect 2688 3392 2740 3398
rect 2688 3334 2740 3340
rect 3240 3392 3292 3398
rect 3240 3334 3292 3340
rect 2504 3052 2556 3058
rect 2504 2994 2556 3000
rect 2700 2961 2728 3334
rect 2686 2952 2742 2961
rect 2686 2887 2742 2896
rect 2136 2848 2188 2854
rect 2136 2790 2188 2796
rect 1860 2440 1912 2446
rect 1860 2382 1912 2388
rect 1492 2304 1544 2310
rect 1492 2246 1544 2252
rect 1504 800 1532 2246
rect 1872 2009 1900 2382
rect 1858 2000 1914 2009
rect 1858 1935 1914 1944
rect 2148 800 2176 2790
rect 3252 2446 3280 3334
rect 4540 2854 4568 3674
rect 4632 3534 4660 4406
rect 4712 4276 4764 4282
rect 4712 4218 4764 4224
rect 4724 4010 4752 4218
rect 4908 4146 4936 5646
rect 5000 5234 5028 9046
rect 5080 8356 5132 8362
rect 5080 8298 5132 8304
rect 5092 7206 5120 8298
rect 5184 8242 5212 9472
rect 5276 9450 5304 13126
rect 5368 12646 5396 13262
rect 5460 13190 5488 13738
rect 5736 13462 5764 13942
rect 5920 13938 5948 15302
rect 5908 13932 5960 13938
rect 5908 13874 5960 13880
rect 5724 13456 5776 13462
rect 5724 13398 5776 13404
rect 5448 13184 5500 13190
rect 5448 13126 5500 13132
rect 5724 12776 5776 12782
rect 5724 12718 5776 12724
rect 5356 12640 5408 12646
rect 5356 12582 5408 12588
rect 5736 12442 5764 12718
rect 5724 12436 5776 12442
rect 5724 12378 5776 12384
rect 6104 12374 6132 18634
rect 6196 12442 6224 20810
rect 6630 20700 6938 20709
rect 6630 20698 6636 20700
rect 6692 20698 6716 20700
rect 6772 20698 6796 20700
rect 6852 20698 6876 20700
rect 6932 20698 6938 20700
rect 6692 20646 6694 20698
rect 6874 20646 6876 20698
rect 6630 20644 6636 20646
rect 6692 20644 6716 20646
rect 6772 20644 6796 20646
rect 6852 20644 6876 20646
rect 6932 20644 6938 20646
rect 6630 20635 6938 20644
rect 6368 19712 6420 19718
rect 6368 19654 6420 19660
rect 6380 19417 6408 19654
rect 6630 19612 6938 19621
rect 6630 19610 6636 19612
rect 6692 19610 6716 19612
rect 6772 19610 6796 19612
rect 6852 19610 6876 19612
rect 6932 19610 6938 19612
rect 6692 19558 6694 19610
rect 6874 19558 6876 19610
rect 6630 19556 6636 19558
rect 6692 19556 6716 19558
rect 6772 19556 6796 19558
rect 6852 19556 6876 19558
rect 6932 19556 6938 19558
rect 6630 19547 6938 19556
rect 7116 19514 7144 21082
rect 7104 19508 7156 19514
rect 7104 19450 7156 19456
rect 6366 19408 6422 19417
rect 6366 19343 6422 19352
rect 6630 18524 6938 18533
rect 6630 18522 6636 18524
rect 6692 18522 6716 18524
rect 6772 18522 6796 18524
rect 6852 18522 6876 18524
rect 6932 18522 6938 18524
rect 6692 18470 6694 18522
rect 6874 18470 6876 18522
rect 6630 18468 6636 18470
rect 6692 18468 6716 18470
rect 6772 18468 6796 18470
rect 6852 18468 6876 18470
rect 6932 18468 6938 18470
rect 6630 18459 6938 18468
rect 7104 18216 7156 18222
rect 7104 18158 7156 18164
rect 7012 17604 7064 17610
rect 7012 17546 7064 17552
rect 6630 17436 6938 17445
rect 6630 17434 6636 17436
rect 6692 17434 6716 17436
rect 6772 17434 6796 17436
rect 6852 17434 6876 17436
rect 6932 17434 6938 17436
rect 6692 17382 6694 17434
rect 6874 17382 6876 17434
rect 6630 17380 6636 17382
rect 6692 17380 6716 17382
rect 6772 17380 6796 17382
rect 6852 17380 6876 17382
rect 6932 17380 6938 17382
rect 6630 17371 6938 17380
rect 6630 16348 6938 16357
rect 6630 16346 6636 16348
rect 6692 16346 6716 16348
rect 6772 16346 6796 16348
rect 6852 16346 6876 16348
rect 6932 16346 6938 16348
rect 6692 16294 6694 16346
rect 6874 16294 6876 16346
rect 6630 16292 6636 16294
rect 6692 16292 6716 16294
rect 6772 16292 6796 16294
rect 6852 16292 6876 16294
rect 6932 16292 6938 16294
rect 6630 16283 6938 16292
rect 7024 16250 7052 17546
rect 7116 17202 7144 18158
rect 7104 17196 7156 17202
rect 7104 17138 7156 17144
rect 7012 16244 7064 16250
rect 7012 16186 7064 16192
rect 7104 16108 7156 16114
rect 7104 16050 7156 16056
rect 6552 15904 6604 15910
rect 6552 15846 6604 15852
rect 6276 15496 6328 15502
rect 6276 15438 6328 15444
rect 6288 13734 6316 15438
rect 6460 14816 6512 14822
rect 6460 14758 6512 14764
rect 6368 14612 6420 14618
rect 6368 14554 6420 14560
rect 6380 13938 6408 14554
rect 6472 14414 6500 14758
rect 6460 14408 6512 14414
rect 6460 14350 6512 14356
rect 6368 13932 6420 13938
rect 6368 13874 6420 13880
rect 6276 13728 6328 13734
rect 6276 13670 6328 13676
rect 6288 13530 6316 13670
rect 6276 13524 6328 13530
rect 6276 13466 6328 13472
rect 6368 13388 6420 13394
rect 6368 13330 6420 13336
rect 6460 13388 6512 13394
rect 6460 13330 6512 13336
rect 6276 13320 6328 13326
rect 6276 13262 6328 13268
rect 6288 12850 6316 13262
rect 6276 12844 6328 12850
rect 6276 12786 6328 12792
rect 6184 12436 6236 12442
rect 6184 12378 6236 12384
rect 6092 12368 6144 12374
rect 6092 12310 6144 12316
rect 5356 12300 5408 12306
rect 5356 12242 5408 12248
rect 5368 11898 5396 12242
rect 5448 12232 5500 12238
rect 5500 12192 5580 12220
rect 5448 12174 5500 12180
rect 5448 12096 5500 12102
rect 5448 12038 5500 12044
rect 5356 11892 5408 11898
rect 5356 11834 5408 11840
rect 5460 11694 5488 12038
rect 5448 11688 5500 11694
rect 5448 11630 5500 11636
rect 5460 11354 5488 11630
rect 5448 11348 5500 11354
rect 5448 11290 5500 11296
rect 5552 10713 5580 12192
rect 6000 12164 6052 12170
rect 6000 12106 6052 12112
rect 6012 11898 6040 12106
rect 6000 11892 6052 11898
rect 6000 11834 6052 11840
rect 5632 11756 5684 11762
rect 5632 11698 5684 11704
rect 5644 11218 5672 11698
rect 6184 11688 6236 11694
rect 6184 11630 6236 11636
rect 5632 11212 5684 11218
rect 5632 11154 5684 11160
rect 5644 10810 5672 11154
rect 6196 11082 6224 11630
rect 6288 11354 6316 12786
rect 6380 12782 6408 13330
rect 6472 12918 6500 13330
rect 6460 12912 6512 12918
rect 6460 12854 6512 12860
rect 6368 12776 6420 12782
rect 6368 12718 6420 12724
rect 6564 12434 6592 15846
rect 7116 15706 7144 16050
rect 7208 16046 7236 21270
rect 7288 20460 7340 20466
rect 7288 20402 7340 20408
rect 7196 16040 7248 16046
rect 7196 15982 7248 15988
rect 7104 15700 7156 15706
rect 7104 15642 7156 15648
rect 7196 15564 7248 15570
rect 7196 15506 7248 15512
rect 6630 15260 6938 15269
rect 6630 15258 6636 15260
rect 6692 15258 6716 15260
rect 6772 15258 6796 15260
rect 6852 15258 6876 15260
rect 6932 15258 6938 15260
rect 6692 15206 6694 15258
rect 6874 15206 6876 15258
rect 6630 15204 6636 15206
rect 6692 15204 6716 15206
rect 6772 15204 6796 15206
rect 6852 15204 6876 15206
rect 6932 15204 6938 15206
rect 6630 15195 6938 15204
rect 6644 15088 6696 15094
rect 6642 15056 6644 15065
rect 6696 15056 6698 15065
rect 6642 14991 6698 15000
rect 7012 14816 7064 14822
rect 7012 14758 7064 14764
rect 6828 14612 6880 14618
rect 6828 14554 6880 14560
rect 6840 14482 6868 14554
rect 6828 14476 6880 14482
rect 6828 14418 6880 14424
rect 6840 14346 6868 14418
rect 6828 14340 6880 14346
rect 6828 14282 6880 14288
rect 6630 14172 6938 14181
rect 6630 14170 6636 14172
rect 6692 14170 6716 14172
rect 6772 14170 6796 14172
rect 6852 14170 6876 14172
rect 6932 14170 6938 14172
rect 6692 14118 6694 14170
rect 6874 14118 6876 14170
rect 6630 14116 6636 14118
rect 6692 14116 6716 14118
rect 6772 14116 6796 14118
rect 6852 14116 6876 14118
rect 6932 14116 6938 14118
rect 6630 14107 6938 14116
rect 6828 14000 6880 14006
rect 6828 13942 6880 13948
rect 6736 13728 6788 13734
rect 6736 13670 6788 13676
rect 6644 13320 6696 13326
rect 6642 13288 6644 13297
rect 6696 13288 6698 13297
rect 6748 13258 6776 13670
rect 6840 13530 6868 13942
rect 6920 13932 6972 13938
rect 6920 13874 6972 13880
rect 6828 13524 6880 13530
rect 6828 13466 6880 13472
rect 6642 13223 6698 13232
rect 6736 13252 6788 13258
rect 6736 13194 6788 13200
rect 6932 13172 6960 13874
rect 7024 13802 7052 14758
rect 7104 14000 7156 14006
rect 7104 13942 7156 13948
rect 7208 13954 7236 15506
rect 7300 14074 7328 20402
rect 7380 18284 7432 18290
rect 7380 18226 7432 18232
rect 7392 18057 7420 18226
rect 7378 18048 7434 18057
rect 7378 17983 7434 17992
rect 7472 17672 7524 17678
rect 7472 17614 7524 17620
rect 7484 16522 7512 17614
rect 7472 16516 7524 16522
rect 7472 16458 7524 16464
rect 7380 16108 7432 16114
rect 7380 16050 7432 16056
rect 7392 15638 7420 16050
rect 7380 15632 7432 15638
rect 7380 15574 7432 15580
rect 7484 15434 7512 16458
rect 7576 15978 7604 21830
rect 9312 21548 9364 21554
rect 9312 21490 9364 21496
rect 9324 21078 9352 21490
rect 9784 21486 9812 21966
rect 10140 21956 10192 21962
rect 10140 21898 10192 21904
rect 11336 21956 11388 21962
rect 11336 21898 11388 21904
rect 9772 21480 9824 21486
rect 9824 21428 9904 21434
rect 9772 21422 9904 21428
rect 9784 21406 9904 21422
rect 9471 21244 9779 21253
rect 9471 21242 9477 21244
rect 9533 21242 9557 21244
rect 9613 21242 9637 21244
rect 9693 21242 9717 21244
rect 9773 21242 9779 21244
rect 9533 21190 9535 21242
rect 9715 21190 9717 21242
rect 9471 21188 9477 21190
rect 9533 21188 9557 21190
rect 9613 21188 9637 21190
rect 9693 21188 9717 21190
rect 9773 21188 9779 21190
rect 9471 21179 9779 21188
rect 9876 21146 9904 21406
rect 9864 21140 9916 21146
rect 9864 21082 9916 21088
rect 9312 21072 9364 21078
rect 9312 21014 9364 21020
rect 7656 20868 7708 20874
rect 7656 20810 7708 20816
rect 8944 20868 8996 20874
rect 8944 20810 8996 20816
rect 7564 15972 7616 15978
rect 7564 15914 7616 15920
rect 7576 15502 7604 15914
rect 7564 15496 7616 15502
rect 7564 15438 7616 15444
rect 7472 15428 7524 15434
rect 7472 15370 7524 15376
rect 7380 14408 7432 14414
rect 7380 14350 7432 14356
rect 7288 14068 7340 14074
rect 7288 14010 7340 14016
rect 7392 14006 7420 14350
rect 7380 14000 7432 14006
rect 7012 13796 7064 13802
rect 7012 13738 7064 13744
rect 7116 13308 7144 13942
rect 7208 13938 7328 13954
rect 7380 13942 7432 13948
rect 7208 13932 7340 13938
rect 7208 13926 7288 13932
rect 7288 13874 7340 13880
rect 7300 13818 7328 13874
rect 7300 13790 7420 13818
rect 7116 13280 7236 13308
rect 7208 13274 7236 13280
rect 7208 13246 7328 13274
rect 7104 13184 7156 13190
rect 6932 13144 7052 13172
rect 6630 13084 6938 13093
rect 6630 13082 6636 13084
rect 6692 13082 6716 13084
rect 6772 13082 6796 13084
rect 6852 13082 6876 13084
rect 6932 13082 6938 13084
rect 6692 13030 6694 13082
rect 6874 13030 6876 13082
rect 6630 13028 6636 13030
rect 6692 13028 6716 13030
rect 6772 13028 6796 13030
rect 6852 13028 6876 13030
rect 6932 13028 6938 13030
rect 6630 13019 6938 13028
rect 6736 12912 6788 12918
rect 6736 12854 6788 12860
rect 6748 12782 6776 12854
rect 6736 12776 6788 12782
rect 6736 12718 6788 12724
rect 6472 12406 6592 12434
rect 6276 11348 6328 11354
rect 6276 11290 6328 11296
rect 6276 11212 6328 11218
rect 6276 11154 6328 11160
rect 5724 11076 5776 11082
rect 5724 11018 5776 11024
rect 6184 11076 6236 11082
rect 6184 11018 6236 11024
rect 5632 10804 5684 10810
rect 5632 10746 5684 10752
rect 5538 10704 5594 10713
rect 5538 10639 5594 10648
rect 5736 10470 5764 11018
rect 6092 10668 6144 10674
rect 6092 10610 6144 10616
rect 5724 10464 5776 10470
rect 5724 10406 5776 10412
rect 6000 10464 6052 10470
rect 6000 10406 6052 10412
rect 5908 10260 5960 10266
rect 5908 10202 5960 10208
rect 5540 10124 5592 10130
rect 5540 10066 5592 10072
rect 5552 9674 5580 10066
rect 5816 10056 5868 10062
rect 5816 9998 5868 10004
rect 5828 9722 5856 9998
rect 5816 9716 5868 9722
rect 5552 9646 5764 9674
rect 5816 9658 5868 9664
rect 5736 9586 5764 9646
rect 5724 9580 5776 9586
rect 5724 9522 5776 9528
rect 5264 9444 5316 9450
rect 5264 9386 5316 9392
rect 5632 9172 5684 9178
rect 5632 9114 5684 9120
rect 5264 8968 5316 8974
rect 5264 8910 5316 8916
rect 5446 8936 5502 8945
rect 5276 8634 5304 8910
rect 5446 8871 5502 8880
rect 5264 8628 5316 8634
rect 5264 8570 5316 8576
rect 5356 8628 5408 8634
rect 5356 8570 5408 8576
rect 5184 8214 5304 8242
rect 5172 8084 5224 8090
rect 5172 8026 5224 8032
rect 5080 7200 5132 7206
rect 5080 7142 5132 7148
rect 5080 6996 5132 7002
rect 5080 6938 5132 6944
rect 5092 6662 5120 6938
rect 5080 6656 5132 6662
rect 5080 6598 5132 6604
rect 5184 6458 5212 8026
rect 5276 7002 5304 8214
rect 5368 7410 5396 8570
rect 5356 7404 5408 7410
rect 5356 7346 5408 7352
rect 5264 6996 5316 7002
rect 5264 6938 5316 6944
rect 5356 6860 5408 6866
rect 5460 6848 5488 8871
rect 5540 8492 5592 8498
rect 5540 8434 5592 8440
rect 5552 7546 5580 8434
rect 5644 7954 5672 9114
rect 5736 8974 5764 9522
rect 5920 9178 5948 10202
rect 5908 9172 5960 9178
rect 5908 9114 5960 9120
rect 5724 8968 5776 8974
rect 5724 8910 5776 8916
rect 5632 7948 5684 7954
rect 5632 7890 5684 7896
rect 5632 7812 5684 7818
rect 5632 7754 5684 7760
rect 5540 7540 5592 7546
rect 5540 7482 5592 7488
rect 5540 7404 5592 7410
rect 5540 7346 5592 7352
rect 5408 6820 5488 6848
rect 5356 6802 5408 6808
rect 5172 6452 5224 6458
rect 5172 6394 5224 6400
rect 5184 5914 5212 6394
rect 5448 6112 5500 6118
rect 5448 6054 5500 6060
rect 5172 5908 5224 5914
rect 5172 5850 5224 5856
rect 5460 5710 5488 6054
rect 5080 5704 5132 5710
rect 5080 5646 5132 5652
rect 5448 5704 5500 5710
rect 5448 5646 5500 5652
rect 4988 5228 5040 5234
rect 4988 5170 5040 5176
rect 5092 4146 5120 5646
rect 5552 5166 5580 7346
rect 5644 6458 5672 7754
rect 5736 7410 5764 8910
rect 6012 7886 6040 10406
rect 6104 9926 6132 10610
rect 6196 10266 6224 11018
rect 6288 10674 6316 11154
rect 6276 10668 6328 10674
rect 6276 10610 6328 10616
rect 6184 10260 6236 10266
rect 6184 10202 6236 10208
rect 6092 9920 6144 9926
rect 6092 9862 6144 9868
rect 6000 7880 6052 7886
rect 6000 7822 6052 7828
rect 5724 7404 5776 7410
rect 5724 7346 5776 7352
rect 5816 7404 5868 7410
rect 5816 7346 5868 7352
rect 5632 6452 5684 6458
rect 5632 6394 5684 6400
rect 5644 5302 5672 6394
rect 5828 6322 5856 7346
rect 5908 7200 5960 7206
rect 5908 7142 5960 7148
rect 5920 6866 5948 7142
rect 6012 6934 6040 7822
rect 6104 7342 6132 9862
rect 6288 8022 6316 10610
rect 6472 9654 6500 12406
rect 6826 12336 6882 12345
rect 6826 12271 6882 12280
rect 6840 12238 6868 12271
rect 6828 12232 6880 12238
rect 6828 12174 6880 12180
rect 6552 12164 6604 12170
rect 6552 12106 6604 12112
rect 6564 10810 6592 12106
rect 7024 12102 7052 13144
rect 7104 13126 7156 13132
rect 7116 12918 7144 13126
rect 7104 12912 7156 12918
rect 7104 12854 7156 12860
rect 7104 12776 7156 12782
rect 7104 12718 7156 12724
rect 7012 12096 7064 12102
rect 7012 12038 7064 12044
rect 6630 11996 6938 12005
rect 6630 11994 6636 11996
rect 6692 11994 6716 11996
rect 6772 11994 6796 11996
rect 6852 11994 6876 11996
rect 6932 11994 6938 11996
rect 6692 11942 6694 11994
rect 6874 11942 6876 11994
rect 6630 11940 6636 11942
rect 6692 11940 6716 11942
rect 6772 11940 6796 11942
rect 6852 11940 6876 11942
rect 6932 11940 6938 11942
rect 6630 11931 6938 11940
rect 7116 11762 7144 12718
rect 7196 12300 7248 12306
rect 7196 12242 7248 12248
rect 7208 12102 7236 12242
rect 7196 12096 7248 12102
rect 7196 12038 7248 12044
rect 7208 11898 7236 12038
rect 7196 11892 7248 11898
rect 7196 11834 7248 11840
rect 7104 11756 7156 11762
rect 7104 11698 7156 11704
rect 7208 11150 7236 11834
rect 7300 11626 7328 13246
rect 7288 11620 7340 11626
rect 7288 11562 7340 11568
rect 7104 11144 7156 11150
rect 7104 11086 7156 11092
rect 7196 11144 7248 11150
rect 7196 11086 7248 11092
rect 7012 11076 7064 11082
rect 7012 11018 7064 11024
rect 6630 10908 6938 10917
rect 6630 10906 6636 10908
rect 6692 10906 6716 10908
rect 6772 10906 6796 10908
rect 6852 10906 6876 10908
rect 6932 10906 6938 10908
rect 6692 10854 6694 10906
rect 6874 10854 6876 10906
rect 6630 10852 6636 10854
rect 6692 10852 6716 10854
rect 6772 10852 6796 10854
rect 6852 10852 6876 10854
rect 6932 10852 6938 10854
rect 6630 10843 6938 10852
rect 6552 10804 6604 10810
rect 6552 10746 6604 10752
rect 6736 10056 6788 10062
rect 6734 10024 6736 10033
rect 6788 10024 6790 10033
rect 6564 9982 6734 10010
rect 6564 9674 6592 9982
rect 6734 9959 6790 9968
rect 6630 9820 6938 9829
rect 6630 9818 6636 9820
rect 6692 9818 6716 9820
rect 6772 9818 6796 9820
rect 6852 9818 6876 9820
rect 6932 9818 6938 9820
rect 6692 9766 6694 9818
rect 6874 9766 6876 9818
rect 6630 9764 6636 9766
rect 6692 9764 6716 9766
rect 6772 9764 6796 9766
rect 6852 9764 6876 9766
rect 6932 9764 6938 9766
rect 6630 9755 6938 9764
rect 7024 9704 7052 11018
rect 6932 9676 7052 9704
rect 6460 9648 6512 9654
rect 6460 9590 6512 9596
rect 6564 9646 6684 9674
rect 6368 9512 6420 9518
rect 6564 9466 6592 9646
rect 6368 9454 6420 9460
rect 6380 9178 6408 9454
rect 6472 9438 6592 9466
rect 6368 9172 6420 9178
rect 6368 9114 6420 9120
rect 6368 8968 6420 8974
rect 6366 8936 6368 8945
rect 6420 8936 6422 8945
rect 6366 8871 6422 8880
rect 6368 8288 6420 8294
rect 6368 8230 6420 8236
rect 6276 8016 6328 8022
rect 6276 7958 6328 7964
rect 6380 7954 6408 8230
rect 6472 8090 6500 9438
rect 6552 9376 6604 9382
rect 6552 9318 6604 9324
rect 6460 8084 6512 8090
rect 6460 8026 6512 8032
rect 6564 7954 6592 9318
rect 6656 9110 6684 9646
rect 6828 9580 6880 9586
rect 6828 9522 6880 9528
rect 6840 9178 6868 9522
rect 6828 9172 6880 9178
rect 6828 9114 6880 9120
rect 6932 9110 6960 9676
rect 7010 9480 7066 9489
rect 7010 9415 7012 9424
rect 7064 9415 7066 9424
rect 7012 9386 7064 9392
rect 6644 9104 6696 9110
rect 6644 9046 6696 9052
rect 6920 9104 6972 9110
rect 6920 9046 6972 9052
rect 6932 8838 6960 9046
rect 7012 8900 7064 8906
rect 7012 8842 7064 8848
rect 6920 8832 6972 8838
rect 6920 8774 6972 8780
rect 6630 8732 6938 8741
rect 6630 8730 6636 8732
rect 6692 8730 6716 8732
rect 6772 8730 6796 8732
rect 6852 8730 6876 8732
rect 6932 8730 6938 8732
rect 6692 8678 6694 8730
rect 6874 8678 6876 8730
rect 6630 8676 6636 8678
rect 6692 8676 6716 8678
rect 6772 8676 6796 8678
rect 6852 8676 6876 8678
rect 6932 8676 6938 8678
rect 6630 8667 6938 8676
rect 7024 8634 7052 8842
rect 7116 8634 7144 11086
rect 7300 11082 7328 11562
rect 7288 11076 7340 11082
rect 7288 11018 7340 11024
rect 7196 10600 7248 10606
rect 7196 10542 7248 10548
rect 7208 9178 7236 10542
rect 7288 9920 7340 9926
rect 7288 9862 7340 9868
rect 7300 9722 7328 9862
rect 7288 9716 7340 9722
rect 7288 9658 7340 9664
rect 7392 9586 7420 13790
rect 7484 13326 7512 15370
rect 7472 13320 7524 13326
rect 7472 13262 7524 13268
rect 7564 13320 7616 13326
rect 7564 13262 7616 13268
rect 7576 12850 7604 13262
rect 7564 12844 7616 12850
rect 7564 12786 7616 12792
rect 7472 12640 7524 12646
rect 7472 12582 7524 12588
rect 7484 12238 7512 12582
rect 7472 12232 7524 12238
rect 7472 12174 7524 12180
rect 7564 12164 7616 12170
rect 7564 12106 7616 12112
rect 7576 11558 7604 12106
rect 7564 11552 7616 11558
rect 7564 11494 7616 11500
rect 7668 11354 7696 20810
rect 8116 20800 8168 20806
rect 8114 20768 8116 20777
rect 8168 20768 8170 20777
rect 8114 20703 8170 20712
rect 8116 20256 8168 20262
rect 8116 20198 8168 20204
rect 8024 18624 8076 18630
rect 8024 18566 8076 18572
rect 7748 17196 7800 17202
rect 7748 17138 7800 17144
rect 7760 15162 7788 17138
rect 7932 16516 7984 16522
rect 7932 16458 7984 16464
rect 7840 16448 7892 16454
rect 7840 16390 7892 16396
rect 7748 15156 7800 15162
rect 7748 15098 7800 15104
rect 7748 14340 7800 14346
rect 7748 14282 7800 14288
rect 7760 13938 7788 14282
rect 7748 13932 7800 13938
rect 7748 13874 7800 13880
rect 7748 13252 7800 13258
rect 7748 13194 7800 13200
rect 7760 12782 7788 13194
rect 7852 12986 7880 16390
rect 7840 12980 7892 12986
rect 7840 12922 7892 12928
rect 7748 12776 7800 12782
rect 7748 12718 7800 12724
rect 7840 12708 7892 12714
rect 7840 12650 7892 12656
rect 7852 12442 7880 12650
rect 7840 12436 7892 12442
rect 7840 12378 7892 12384
rect 7944 11898 7972 16458
rect 8036 15570 8064 18566
rect 8128 17882 8156 20198
rect 8300 19848 8352 19854
rect 8300 19790 8352 19796
rect 8208 19712 8260 19718
rect 8208 19654 8260 19660
rect 8116 17876 8168 17882
rect 8116 17818 8168 17824
rect 8128 16114 8156 17818
rect 8116 16108 8168 16114
rect 8116 16050 8168 16056
rect 8024 15564 8076 15570
rect 8024 15506 8076 15512
rect 8024 15360 8076 15366
rect 8024 15302 8076 15308
rect 8036 15026 8064 15302
rect 8024 15020 8076 15026
rect 8024 14962 8076 14968
rect 8036 14618 8064 14962
rect 8024 14612 8076 14618
rect 8024 14554 8076 14560
rect 8036 14006 8064 14554
rect 8116 14272 8168 14278
rect 8116 14214 8168 14220
rect 8024 14000 8076 14006
rect 8024 13942 8076 13948
rect 8128 13802 8156 14214
rect 8116 13796 8168 13802
rect 8116 13738 8168 13744
rect 8116 13320 8168 13326
rect 8116 13262 8168 13268
rect 8024 12980 8076 12986
rect 8024 12922 8076 12928
rect 7932 11892 7984 11898
rect 8036 11880 8064 12922
rect 8128 12322 8156 13262
rect 8220 12442 8248 19654
rect 8312 18766 8340 19790
rect 8956 19174 8984 20810
rect 9471 20156 9779 20165
rect 9471 20154 9477 20156
rect 9533 20154 9557 20156
rect 9613 20154 9637 20156
rect 9693 20154 9717 20156
rect 9773 20154 9779 20156
rect 9533 20102 9535 20154
rect 9715 20102 9717 20154
rect 9471 20100 9477 20102
rect 9533 20100 9557 20102
rect 9613 20100 9637 20102
rect 9693 20100 9717 20102
rect 9773 20100 9779 20102
rect 9471 20091 9779 20100
rect 8944 19168 8996 19174
rect 8944 19110 8996 19116
rect 8300 18760 8352 18766
rect 8300 18702 8352 18708
rect 8392 18760 8444 18766
rect 8392 18702 8444 18708
rect 8312 18290 8340 18702
rect 8300 18284 8352 18290
rect 8300 18226 8352 18232
rect 8300 16652 8352 16658
rect 8300 16594 8352 16600
rect 8312 16250 8340 16594
rect 8300 16244 8352 16250
rect 8300 16186 8352 16192
rect 8404 15706 8432 18702
rect 8484 16992 8536 16998
rect 8484 16934 8536 16940
rect 8392 15700 8444 15706
rect 8392 15642 8444 15648
rect 8300 15428 8352 15434
rect 8300 15370 8352 15376
rect 8312 15094 8340 15370
rect 8300 15088 8352 15094
rect 8300 15030 8352 15036
rect 8312 14074 8340 15030
rect 8496 15026 8524 16934
rect 8956 16182 8984 19110
rect 9471 19068 9779 19077
rect 9471 19066 9477 19068
rect 9533 19066 9557 19068
rect 9613 19066 9637 19068
rect 9693 19066 9717 19068
rect 9773 19066 9779 19068
rect 9533 19014 9535 19066
rect 9715 19014 9717 19066
rect 9471 19012 9477 19014
rect 9533 19012 9557 19014
rect 9613 19012 9637 19014
rect 9693 19012 9717 19014
rect 9773 19012 9779 19014
rect 9471 19003 9779 19012
rect 9312 18284 9364 18290
rect 9312 18226 9364 18232
rect 9128 18080 9180 18086
rect 9128 18022 9180 18028
rect 8944 16176 8996 16182
rect 8944 16118 8996 16124
rect 9140 15502 9168 18022
rect 9324 17678 9352 18226
rect 9471 17980 9779 17989
rect 9471 17978 9477 17980
rect 9533 17978 9557 17980
rect 9613 17978 9637 17980
rect 9693 17978 9717 17980
rect 9773 17978 9779 17980
rect 9533 17926 9535 17978
rect 9715 17926 9717 17978
rect 9471 17924 9477 17926
rect 9533 17924 9557 17926
rect 9613 17924 9637 17926
rect 9693 17924 9717 17926
rect 9773 17924 9779 17926
rect 9471 17915 9779 17924
rect 9312 17672 9364 17678
rect 9312 17614 9364 17620
rect 9324 17202 9352 17614
rect 9312 17196 9364 17202
rect 9312 17138 9364 17144
rect 9324 16658 9352 17138
rect 9471 16892 9779 16901
rect 9471 16890 9477 16892
rect 9533 16890 9557 16892
rect 9613 16890 9637 16892
rect 9693 16890 9717 16892
rect 9773 16890 9779 16892
rect 9533 16838 9535 16890
rect 9715 16838 9717 16890
rect 9471 16836 9477 16838
rect 9533 16836 9557 16838
rect 9613 16836 9637 16838
rect 9693 16836 9717 16838
rect 9773 16836 9779 16838
rect 9471 16827 9779 16836
rect 9312 16652 9364 16658
rect 9312 16594 9364 16600
rect 9312 16448 9364 16454
rect 9312 16390 9364 16396
rect 9324 15910 9352 16390
rect 9312 15904 9364 15910
rect 9312 15846 9364 15852
rect 9220 15564 9272 15570
rect 9220 15506 9272 15512
rect 9128 15496 9180 15502
rect 9128 15438 9180 15444
rect 8392 15020 8444 15026
rect 8392 14962 8444 14968
rect 8484 15020 8536 15026
rect 8484 14962 8536 14968
rect 8300 14068 8352 14074
rect 8300 14010 8352 14016
rect 8404 12782 8432 14962
rect 8852 14884 8904 14890
rect 8852 14826 8904 14832
rect 8864 13530 8892 14826
rect 9232 14822 9260 15506
rect 9324 15484 9352 15846
rect 9471 15804 9779 15813
rect 9471 15802 9477 15804
rect 9533 15802 9557 15804
rect 9613 15802 9637 15804
rect 9693 15802 9717 15804
rect 9773 15802 9779 15804
rect 9533 15750 9535 15802
rect 9715 15750 9717 15802
rect 9471 15748 9477 15750
rect 9533 15748 9557 15750
rect 9613 15748 9637 15750
rect 9693 15748 9717 15750
rect 9773 15748 9779 15750
rect 9471 15739 9779 15748
rect 9404 15496 9456 15502
rect 9324 15456 9404 15484
rect 9404 15438 9456 15444
rect 9312 15020 9364 15026
rect 9312 14962 9364 14968
rect 8944 14816 8996 14822
rect 8944 14758 8996 14764
rect 9220 14816 9272 14822
rect 9220 14758 9272 14764
rect 8852 13524 8904 13530
rect 8852 13466 8904 13472
rect 8576 12912 8628 12918
rect 8576 12854 8628 12860
rect 8392 12776 8444 12782
rect 8392 12718 8444 12724
rect 8208 12436 8260 12442
rect 8208 12378 8260 12384
rect 8128 12294 8340 12322
rect 8588 12306 8616 12854
rect 8668 12776 8720 12782
rect 8668 12718 8720 12724
rect 8208 12164 8260 12170
rect 8208 12106 8260 12112
rect 8114 11928 8170 11937
rect 8036 11872 8114 11880
rect 8036 11852 8116 11872
rect 7932 11834 7984 11840
rect 8168 11863 8170 11872
rect 8116 11834 8168 11840
rect 7748 11756 7800 11762
rect 7748 11698 7800 11704
rect 8116 11756 8168 11762
rect 8220 11744 8248 12106
rect 8312 11898 8340 12294
rect 8484 12300 8536 12306
rect 8484 12242 8536 12248
rect 8576 12300 8628 12306
rect 8576 12242 8628 12248
rect 8496 12073 8524 12242
rect 8576 12164 8628 12170
rect 8576 12106 8628 12112
rect 8482 12064 8538 12073
rect 8482 11999 8538 12008
rect 8300 11892 8352 11898
rect 8300 11834 8352 11840
rect 8168 11716 8248 11744
rect 8300 11756 8352 11762
rect 8116 11698 8168 11704
rect 8300 11698 8352 11704
rect 7656 11348 7708 11354
rect 7656 11290 7708 11296
rect 7562 11248 7618 11257
rect 7562 11183 7618 11192
rect 7576 11150 7604 11183
rect 7564 11144 7616 11150
rect 7564 11086 7616 11092
rect 7472 9988 7524 9994
rect 7472 9930 7524 9936
rect 7288 9580 7340 9586
rect 7288 9522 7340 9528
rect 7380 9580 7432 9586
rect 7380 9522 7432 9528
rect 7196 9172 7248 9178
rect 7196 9114 7248 9120
rect 7012 8628 7064 8634
rect 7012 8570 7064 8576
rect 7104 8628 7156 8634
rect 7104 8570 7156 8576
rect 7300 8566 7328 9522
rect 7288 8560 7340 8566
rect 7288 8502 7340 8508
rect 7012 8424 7064 8430
rect 7012 8366 7064 8372
rect 6368 7948 6420 7954
rect 6368 7890 6420 7896
rect 6552 7948 6604 7954
rect 6552 7890 6604 7896
rect 6460 7880 6512 7886
rect 6460 7822 6512 7828
rect 6368 7472 6420 7478
rect 6368 7414 6420 7420
rect 6380 7342 6408 7414
rect 6092 7336 6144 7342
rect 6092 7278 6144 7284
rect 6368 7336 6420 7342
rect 6368 7278 6420 7284
rect 6472 7002 6500 7822
rect 6630 7644 6938 7653
rect 6630 7642 6636 7644
rect 6692 7642 6716 7644
rect 6772 7642 6796 7644
rect 6852 7642 6876 7644
rect 6932 7642 6938 7644
rect 6692 7590 6694 7642
rect 6874 7590 6876 7642
rect 6630 7588 6636 7590
rect 6692 7588 6716 7590
rect 6772 7588 6796 7590
rect 6852 7588 6876 7590
rect 6932 7588 6938 7590
rect 6630 7579 6938 7588
rect 7024 7342 7052 8366
rect 7196 8288 7248 8294
rect 7196 8230 7248 8236
rect 7208 7886 7236 8230
rect 7196 7880 7248 7886
rect 7194 7848 7196 7857
rect 7248 7848 7250 7857
rect 7300 7834 7328 8502
rect 7380 8492 7432 8498
rect 7484 8480 7512 9930
rect 7576 9382 7604 11086
rect 7760 10062 7788 11698
rect 8128 11626 8156 11698
rect 8116 11620 8168 11626
rect 8116 11562 8168 11568
rect 7840 11552 7892 11558
rect 7840 11494 7892 11500
rect 7852 11014 7880 11494
rect 8128 11082 8156 11562
rect 8116 11076 8168 11082
rect 8116 11018 8168 11024
rect 7840 11008 7892 11014
rect 7840 10950 7892 10956
rect 8024 10668 8076 10674
rect 8024 10610 8076 10616
rect 8036 10577 8064 10610
rect 8022 10568 8078 10577
rect 8022 10503 8078 10512
rect 8208 10464 8260 10470
rect 8208 10406 8260 10412
rect 7840 10192 7892 10198
rect 8024 10192 8076 10198
rect 7892 10152 8024 10180
rect 7840 10134 7892 10140
rect 8220 10146 8248 10406
rect 8024 10134 8076 10140
rect 7748 10056 7800 10062
rect 7800 10016 7972 10044
rect 7748 9998 7800 10004
rect 7748 9648 7800 9654
rect 7748 9590 7800 9596
rect 7564 9376 7616 9382
rect 7564 9318 7616 9324
rect 7432 8452 7512 8480
rect 7380 8434 7432 8440
rect 7300 7806 7420 7834
rect 7194 7783 7250 7792
rect 7288 7744 7340 7750
rect 7288 7686 7340 7692
rect 7012 7336 7064 7342
rect 7012 7278 7064 7284
rect 6460 6996 6512 7002
rect 6460 6938 6512 6944
rect 6000 6928 6052 6934
rect 6000 6870 6052 6876
rect 5908 6860 5960 6866
rect 5908 6802 5960 6808
rect 7104 6792 7156 6798
rect 5998 6760 6054 6769
rect 7104 6734 7156 6740
rect 5920 6704 5998 6712
rect 5920 6684 6000 6704
rect 5816 6316 5868 6322
rect 5816 6258 5868 6264
rect 5632 5296 5684 5302
rect 5632 5238 5684 5244
rect 5540 5160 5592 5166
rect 5540 5102 5592 5108
rect 5356 4752 5408 4758
rect 5356 4694 5408 4700
rect 5540 4752 5592 4758
rect 5540 4694 5592 4700
rect 5172 4616 5224 4622
rect 5172 4558 5224 4564
rect 5184 4214 5212 4558
rect 5368 4486 5396 4694
rect 5264 4480 5316 4486
rect 5264 4422 5316 4428
rect 5356 4480 5408 4486
rect 5356 4422 5408 4428
rect 5276 4282 5304 4422
rect 5264 4276 5316 4282
rect 5264 4218 5316 4224
rect 5172 4208 5224 4214
rect 5172 4150 5224 4156
rect 4896 4140 4948 4146
rect 4896 4082 4948 4088
rect 5080 4140 5132 4146
rect 5080 4082 5132 4088
rect 4712 4004 4764 4010
rect 4712 3946 4764 3952
rect 4724 3738 4752 3946
rect 4908 3777 4936 4082
rect 4894 3768 4950 3777
rect 4712 3732 4764 3738
rect 4894 3703 4950 3712
rect 4712 3674 4764 3680
rect 5368 3670 5396 4422
rect 4896 3664 4948 3670
rect 4896 3606 4948 3612
rect 5356 3664 5408 3670
rect 5356 3606 5408 3612
rect 4620 3528 4672 3534
rect 4620 3470 4672 3476
rect 4908 3194 4936 3606
rect 5552 3398 5580 4694
rect 5920 4185 5948 6684
rect 6052 6695 6054 6704
rect 6000 6666 6052 6672
rect 7012 6656 7064 6662
rect 7012 6598 7064 6604
rect 6630 6556 6938 6565
rect 6630 6554 6636 6556
rect 6692 6554 6716 6556
rect 6772 6554 6796 6556
rect 6852 6554 6876 6556
rect 6932 6554 6938 6556
rect 6692 6502 6694 6554
rect 6874 6502 6876 6554
rect 6630 6500 6636 6502
rect 6692 6500 6716 6502
rect 6772 6500 6796 6502
rect 6852 6500 6876 6502
rect 6932 6500 6938 6502
rect 6630 6491 6938 6500
rect 6552 6452 6604 6458
rect 6552 6394 6604 6400
rect 6460 6384 6512 6390
rect 6460 6326 6512 6332
rect 6092 5704 6144 5710
rect 6092 5646 6144 5652
rect 6276 5704 6328 5710
rect 6276 5646 6328 5652
rect 6000 5092 6052 5098
rect 6000 5034 6052 5040
rect 5906 4176 5962 4185
rect 5906 4111 5962 4120
rect 5632 3936 5684 3942
rect 5632 3878 5684 3884
rect 5540 3392 5592 3398
rect 5540 3334 5592 3340
rect 4896 3188 4948 3194
rect 4896 3130 4948 3136
rect 5644 3058 5672 3878
rect 5814 3496 5870 3505
rect 5814 3431 5870 3440
rect 5632 3052 5684 3058
rect 5632 2994 5684 3000
rect 4528 2848 4580 2854
rect 4528 2790 4580 2796
rect 3790 2748 4098 2757
rect 3790 2746 3796 2748
rect 3852 2746 3876 2748
rect 3932 2746 3956 2748
rect 4012 2746 4036 2748
rect 4092 2746 4098 2748
rect 3852 2694 3854 2746
rect 4034 2694 4036 2746
rect 3790 2692 3796 2694
rect 3852 2692 3876 2694
rect 3932 2692 3956 2694
rect 4012 2692 4036 2694
rect 4092 2692 4098 2694
rect 3790 2683 4098 2692
rect 5078 2680 5134 2689
rect 5078 2615 5134 2624
rect 5092 2582 5120 2615
rect 5080 2576 5132 2582
rect 4250 2544 4306 2553
rect 5080 2518 5132 2524
rect 4250 2479 4306 2488
rect 4264 2446 4292 2479
rect 5828 2446 5856 3431
rect 5920 3058 5948 4111
rect 6012 4078 6040 5034
rect 6104 4758 6132 5646
rect 6288 5370 6316 5646
rect 6276 5364 6328 5370
rect 6276 5306 6328 5312
rect 6276 5024 6328 5030
rect 6276 4966 6328 4972
rect 6092 4752 6144 4758
rect 6092 4694 6144 4700
rect 6000 4072 6052 4078
rect 6000 4014 6052 4020
rect 6092 4004 6144 4010
rect 6092 3946 6144 3952
rect 6104 3602 6132 3946
rect 6092 3596 6144 3602
rect 6092 3538 6144 3544
rect 6288 3074 6316 4966
rect 6472 3738 6500 6326
rect 6564 5302 6592 6394
rect 6644 6316 6696 6322
rect 6644 6258 6696 6264
rect 6656 5710 6684 6258
rect 6736 6248 6788 6254
rect 6736 6190 6788 6196
rect 6644 5704 6696 5710
rect 6644 5646 6696 5652
rect 6748 5574 6776 6190
rect 6736 5568 6788 5574
rect 6736 5510 6788 5516
rect 6630 5468 6938 5477
rect 6630 5466 6636 5468
rect 6692 5466 6716 5468
rect 6772 5466 6796 5468
rect 6852 5466 6876 5468
rect 6932 5466 6938 5468
rect 6692 5414 6694 5466
rect 6874 5414 6876 5466
rect 6630 5412 6636 5414
rect 6692 5412 6716 5414
rect 6772 5412 6796 5414
rect 6852 5412 6876 5414
rect 6932 5412 6938 5414
rect 6630 5403 6938 5412
rect 6552 5296 6604 5302
rect 6552 5238 6604 5244
rect 6564 4622 6592 5238
rect 6920 4752 6972 4758
rect 6920 4694 6972 4700
rect 7024 4706 7052 6598
rect 7116 6322 7144 6734
rect 7196 6724 7248 6730
rect 7196 6666 7248 6672
rect 7208 6458 7236 6666
rect 7196 6452 7248 6458
rect 7196 6394 7248 6400
rect 7104 6316 7156 6322
rect 7104 6258 7156 6264
rect 7300 5710 7328 7686
rect 7392 7342 7420 7806
rect 7484 7410 7512 8452
rect 7564 8492 7616 8498
rect 7564 8434 7616 8440
rect 7656 8492 7708 8498
rect 7656 8434 7708 8440
rect 7576 8090 7604 8434
rect 7668 8401 7696 8434
rect 7654 8392 7710 8401
rect 7654 8327 7710 8336
rect 7656 8288 7708 8294
rect 7656 8230 7708 8236
rect 7564 8084 7616 8090
rect 7564 8026 7616 8032
rect 7668 7886 7696 8230
rect 7656 7880 7708 7886
rect 7656 7822 7708 7828
rect 7656 7744 7708 7750
rect 7656 7686 7708 7692
rect 7472 7404 7524 7410
rect 7472 7346 7524 7352
rect 7380 7336 7432 7342
rect 7380 7278 7432 7284
rect 7472 6792 7524 6798
rect 7472 6734 7524 6740
rect 7484 6662 7512 6734
rect 7380 6656 7432 6662
rect 7380 6598 7432 6604
rect 7472 6656 7524 6662
rect 7472 6598 7524 6604
rect 7288 5704 7340 5710
rect 7288 5646 7340 5652
rect 7392 5556 7420 6598
rect 7484 5846 7512 6598
rect 7564 6316 7616 6322
rect 7564 6258 7616 6264
rect 7472 5840 7524 5846
rect 7472 5782 7524 5788
rect 7576 5710 7604 6258
rect 7668 5710 7696 7686
rect 7760 6934 7788 9590
rect 7840 9376 7892 9382
rect 7838 9344 7840 9353
rect 7892 9344 7894 9353
rect 7838 9279 7894 9288
rect 7840 8492 7892 8498
rect 7840 8434 7892 8440
rect 7748 6928 7800 6934
rect 7748 6870 7800 6876
rect 7564 5704 7616 5710
rect 7564 5646 7616 5652
rect 7656 5704 7708 5710
rect 7656 5646 7708 5652
rect 7300 5528 7420 5556
rect 7300 5030 7328 5528
rect 7380 5228 7432 5234
rect 7380 5170 7432 5176
rect 7288 5024 7340 5030
rect 7288 4966 7340 4972
rect 6552 4616 6604 4622
rect 6552 4558 6604 4564
rect 6564 4078 6592 4558
rect 6932 4468 6960 4694
rect 7024 4690 7236 4706
rect 7024 4684 7248 4690
rect 7024 4678 7196 4684
rect 7196 4626 7248 4632
rect 7300 4554 7328 4966
rect 7196 4548 7248 4554
rect 7196 4490 7248 4496
rect 7288 4548 7340 4554
rect 7288 4490 7340 4496
rect 6932 4440 7052 4468
rect 6630 4380 6938 4389
rect 6630 4378 6636 4380
rect 6692 4378 6716 4380
rect 6772 4378 6796 4380
rect 6852 4378 6876 4380
rect 6932 4378 6938 4380
rect 6692 4326 6694 4378
rect 6874 4326 6876 4378
rect 6630 4324 6636 4326
rect 6692 4324 6716 4326
rect 6772 4324 6796 4326
rect 6852 4324 6876 4326
rect 6932 4324 6938 4326
rect 6630 4315 6938 4324
rect 7024 4162 7052 4440
rect 7208 4282 7236 4490
rect 7196 4276 7248 4282
rect 7196 4218 7248 4224
rect 6828 4140 6880 4146
rect 6828 4082 6880 4088
rect 6932 4134 7052 4162
rect 6552 4072 6604 4078
rect 6552 4014 6604 4020
rect 6368 3732 6420 3738
rect 6368 3674 6420 3680
rect 6460 3732 6512 3738
rect 6460 3674 6512 3680
rect 6380 3618 6408 3674
rect 6380 3590 6500 3618
rect 6840 3602 6868 4082
rect 6932 4078 6960 4134
rect 6920 4072 6972 4078
rect 6920 4014 6972 4020
rect 7104 4072 7156 4078
rect 7104 4014 7156 4020
rect 6472 3534 6500 3590
rect 6828 3596 6880 3602
rect 6828 3538 6880 3544
rect 7116 3534 7144 4014
rect 7286 3768 7342 3777
rect 7286 3703 7342 3712
rect 7300 3534 7328 3703
rect 6460 3528 6512 3534
rect 6460 3470 6512 3476
rect 7104 3528 7156 3534
rect 7104 3470 7156 3476
rect 7288 3528 7340 3534
rect 7288 3470 7340 3476
rect 6630 3292 6938 3301
rect 6630 3290 6636 3292
rect 6692 3290 6716 3292
rect 6772 3290 6796 3292
rect 6852 3290 6876 3292
rect 6932 3290 6938 3292
rect 6692 3238 6694 3290
rect 6874 3238 6876 3290
rect 6630 3236 6636 3238
rect 6692 3236 6716 3238
rect 6772 3236 6796 3238
rect 6852 3236 6876 3238
rect 6932 3236 6938 3238
rect 6630 3227 6938 3236
rect 7392 3194 7420 5170
rect 7472 4616 7524 4622
rect 7472 4558 7524 4564
rect 7484 3942 7512 4558
rect 7472 3936 7524 3942
rect 7472 3878 7524 3884
rect 7760 3670 7788 6870
rect 7852 5302 7880 8434
rect 7944 8378 7972 10016
rect 8036 8498 8064 10134
rect 8128 10118 8248 10146
rect 8128 9994 8156 10118
rect 8116 9988 8168 9994
rect 8116 9930 8168 9936
rect 8116 9512 8168 9518
rect 8116 9454 8168 9460
rect 8024 8492 8076 8498
rect 8024 8434 8076 8440
rect 7944 8350 8064 8378
rect 7932 7880 7984 7886
rect 7932 7822 7984 7828
rect 7944 7478 7972 7822
rect 7932 7472 7984 7478
rect 7932 7414 7984 7420
rect 7932 7336 7984 7342
rect 7932 7278 7984 7284
rect 7840 5296 7892 5302
rect 7840 5238 7892 5244
rect 7944 4826 7972 7278
rect 8036 6662 8064 8350
rect 8128 7546 8156 9454
rect 8208 7880 8260 7886
rect 8208 7822 8260 7828
rect 8116 7540 8168 7546
rect 8116 7482 8168 7488
rect 8220 6866 8248 7822
rect 8312 7546 8340 11698
rect 8392 11552 8444 11558
rect 8392 11494 8444 11500
rect 8404 11354 8432 11494
rect 8588 11354 8616 12106
rect 8392 11348 8444 11354
rect 8392 11290 8444 11296
rect 8576 11348 8628 11354
rect 8576 11290 8628 11296
rect 8484 11076 8536 11082
rect 8484 11018 8536 11024
rect 8496 10810 8524 11018
rect 8484 10804 8536 10810
rect 8484 10746 8536 10752
rect 8576 10736 8628 10742
rect 8576 10678 8628 10684
rect 8392 10600 8444 10606
rect 8392 10542 8444 10548
rect 8404 9761 8432 10542
rect 8484 10056 8536 10062
rect 8482 10024 8484 10033
rect 8536 10024 8538 10033
rect 8482 9959 8538 9968
rect 8484 9920 8536 9926
rect 8484 9862 8536 9868
rect 8390 9752 8446 9761
rect 8390 9687 8446 9696
rect 8392 8968 8444 8974
rect 8392 8910 8444 8916
rect 8404 7886 8432 8910
rect 8496 8498 8524 9862
rect 8484 8492 8536 8498
rect 8484 8434 8536 8440
rect 8392 7880 8444 7886
rect 8390 7848 8392 7857
rect 8444 7848 8446 7857
rect 8390 7783 8446 7792
rect 8300 7540 8352 7546
rect 8300 7482 8352 7488
rect 8300 7200 8352 7206
rect 8300 7142 8352 7148
rect 8208 6860 8260 6866
rect 8208 6802 8260 6808
rect 8116 6792 8168 6798
rect 8116 6734 8168 6740
rect 8024 6656 8076 6662
rect 8024 6598 8076 6604
rect 8024 6316 8076 6322
rect 8024 6258 8076 6264
rect 8036 6118 8064 6258
rect 8024 6112 8076 6118
rect 8024 6054 8076 6060
rect 8036 5098 8064 6054
rect 8128 5914 8156 6734
rect 8208 6656 8260 6662
rect 8208 6598 8260 6604
rect 8116 5908 8168 5914
rect 8116 5850 8168 5856
rect 8220 5778 8248 6598
rect 8208 5772 8260 5778
rect 8208 5714 8260 5720
rect 8312 5710 8340 7142
rect 8484 6928 8536 6934
rect 8484 6870 8536 6876
rect 8392 6860 8444 6866
rect 8392 6802 8444 6808
rect 8300 5704 8352 5710
rect 8300 5646 8352 5652
rect 8208 5636 8260 5642
rect 8208 5578 8260 5584
rect 8116 5296 8168 5302
rect 8116 5238 8168 5244
rect 8024 5092 8076 5098
rect 8024 5034 8076 5040
rect 8036 4826 8064 5034
rect 7932 4820 7984 4826
rect 7932 4762 7984 4768
rect 8024 4820 8076 4826
rect 8024 4762 8076 4768
rect 8128 4622 8156 5238
rect 8116 4616 8168 4622
rect 8116 4558 8168 4564
rect 7840 4480 7892 4486
rect 7840 4422 7892 4428
rect 7852 4146 7880 4422
rect 8220 4146 8248 5578
rect 8300 5568 8352 5574
rect 8300 5510 8352 5516
rect 8312 4706 8340 5510
rect 8404 4826 8432 6802
rect 8496 6390 8524 6870
rect 8588 6662 8616 10678
rect 8680 9178 8708 12718
rect 8760 12708 8812 12714
rect 8760 12650 8812 12656
rect 8772 10713 8800 12650
rect 8956 10826 8984 14758
rect 9128 14340 9180 14346
rect 9128 14282 9180 14288
rect 9036 14068 9088 14074
rect 9036 14010 9088 14016
rect 9048 13870 9076 14010
rect 9036 13864 9088 13870
rect 9036 13806 9088 13812
rect 9048 11830 9076 13806
rect 9140 13190 9168 14282
rect 9232 14278 9260 14758
rect 9324 14414 9352 14962
rect 9416 14890 9444 15438
rect 9864 15428 9916 15434
rect 9864 15370 9916 15376
rect 9404 14884 9456 14890
rect 9404 14826 9456 14832
rect 9471 14716 9779 14725
rect 9471 14714 9477 14716
rect 9533 14714 9557 14716
rect 9613 14714 9637 14716
rect 9693 14714 9717 14716
rect 9773 14714 9779 14716
rect 9533 14662 9535 14714
rect 9715 14662 9717 14714
rect 9471 14660 9477 14662
rect 9533 14660 9557 14662
rect 9613 14660 9637 14662
rect 9693 14660 9717 14662
rect 9773 14660 9779 14662
rect 9471 14651 9779 14660
rect 9876 14414 9904 15370
rect 9312 14408 9364 14414
rect 9312 14350 9364 14356
rect 9864 14408 9916 14414
rect 9864 14350 9916 14356
rect 9220 14272 9272 14278
rect 9220 14214 9272 14220
rect 9232 13938 9260 14214
rect 9324 13938 9352 14350
rect 9956 14272 10008 14278
rect 9956 14214 10008 14220
rect 9220 13932 9272 13938
rect 9220 13874 9272 13880
rect 9312 13932 9364 13938
rect 9312 13874 9364 13880
rect 9232 13394 9260 13874
rect 9220 13388 9272 13394
rect 9220 13330 9272 13336
rect 9324 13326 9352 13874
rect 9471 13628 9779 13637
rect 9471 13626 9477 13628
rect 9533 13626 9557 13628
rect 9613 13626 9637 13628
rect 9693 13626 9717 13628
rect 9773 13626 9779 13628
rect 9533 13574 9535 13626
rect 9715 13574 9717 13626
rect 9471 13572 9477 13574
rect 9533 13572 9557 13574
rect 9613 13572 9637 13574
rect 9693 13572 9717 13574
rect 9773 13572 9779 13574
rect 9471 13563 9779 13572
rect 9588 13388 9640 13394
rect 9588 13330 9640 13336
rect 9312 13320 9364 13326
rect 9312 13262 9364 13268
rect 9128 13184 9180 13190
rect 9128 13126 9180 13132
rect 9140 12918 9168 13126
rect 9128 12912 9180 12918
rect 9128 12854 9180 12860
rect 9324 12782 9352 13262
rect 9600 12850 9628 13330
rect 9588 12844 9640 12850
rect 9588 12786 9640 12792
rect 9312 12776 9364 12782
rect 9312 12718 9364 12724
rect 9324 12646 9352 12718
rect 9312 12640 9364 12646
rect 9312 12582 9364 12588
rect 9471 12540 9779 12549
rect 9471 12538 9477 12540
rect 9533 12538 9557 12540
rect 9613 12538 9637 12540
rect 9693 12538 9717 12540
rect 9773 12538 9779 12540
rect 9533 12486 9535 12538
rect 9715 12486 9717 12538
rect 9471 12484 9477 12486
rect 9533 12484 9557 12486
rect 9613 12484 9637 12486
rect 9693 12484 9717 12486
rect 9773 12484 9779 12486
rect 9471 12475 9779 12484
rect 9772 12232 9824 12238
rect 9772 12174 9824 12180
rect 9680 12164 9732 12170
rect 9680 12106 9732 12112
rect 9036 11824 9088 11830
rect 9036 11766 9088 11772
rect 9048 11286 9076 11766
rect 9312 11756 9364 11762
rect 9312 11698 9364 11704
rect 9036 11280 9088 11286
rect 9036 11222 9088 11228
rect 9220 11280 9272 11286
rect 9220 11222 9272 11228
rect 9128 11144 9180 11150
rect 9128 11086 9180 11092
rect 9036 11076 9088 11082
rect 9036 11018 9088 11024
rect 8864 10810 8984 10826
rect 8864 10804 8996 10810
rect 8864 10798 8944 10804
rect 8758 10704 8814 10713
rect 8758 10639 8760 10648
rect 8812 10639 8814 10648
rect 8760 10610 8812 10616
rect 8668 9172 8720 9178
rect 8668 9114 8720 9120
rect 8772 8634 8800 10610
rect 8864 9466 8892 10798
rect 8944 10746 8996 10752
rect 8944 10668 8996 10674
rect 8944 10610 8996 10616
rect 8956 10266 8984 10610
rect 8944 10260 8996 10266
rect 8944 10202 8996 10208
rect 8864 9438 8984 9466
rect 8852 9376 8904 9382
rect 8852 9318 8904 9324
rect 8760 8628 8812 8634
rect 8760 8570 8812 8576
rect 8668 8492 8720 8498
rect 8668 8434 8720 8440
rect 8680 7478 8708 8434
rect 8772 7818 8800 8570
rect 8760 7812 8812 7818
rect 8760 7754 8812 7760
rect 8668 7472 8720 7478
rect 8668 7414 8720 7420
rect 8576 6656 8628 6662
rect 8576 6598 8628 6604
rect 8484 6384 8536 6390
rect 8484 6326 8536 6332
rect 8496 5166 8524 6326
rect 8772 6322 8800 7754
rect 8576 6316 8628 6322
rect 8760 6316 8812 6322
rect 8576 6258 8628 6264
rect 8668 6282 8720 6288
rect 8588 5914 8616 6258
rect 8760 6258 8812 6264
rect 8668 6224 8720 6230
rect 8576 5908 8628 5914
rect 8576 5850 8628 5856
rect 8576 5704 8628 5710
rect 8576 5646 8628 5652
rect 8484 5160 8536 5166
rect 8484 5102 8536 5108
rect 8392 4820 8444 4826
rect 8392 4762 8444 4768
rect 8312 4678 8432 4706
rect 7840 4140 7892 4146
rect 7840 4082 7892 4088
rect 8208 4140 8260 4146
rect 8208 4082 8260 4088
rect 7748 3664 7800 3670
rect 7748 3606 7800 3612
rect 7472 3528 7524 3534
rect 7472 3470 7524 3476
rect 7380 3188 7432 3194
rect 7380 3130 7432 3136
rect 5908 3052 5960 3058
rect 6288 3046 6684 3074
rect 5908 2994 5960 3000
rect 6656 2922 6684 3046
rect 7288 3052 7340 3058
rect 7288 2994 7340 3000
rect 6460 2916 6512 2922
rect 6460 2858 6512 2864
rect 6644 2916 6696 2922
rect 6644 2858 6696 2864
rect 3240 2440 3292 2446
rect 3424 2440 3476 2446
rect 3240 2382 3292 2388
rect 3422 2408 3424 2417
rect 4252 2440 4304 2446
rect 3476 2408 3478 2417
rect 4252 2382 4304 2388
rect 5816 2440 5868 2446
rect 5816 2382 5868 2388
rect 3422 2343 3478 2352
rect 2780 2304 2832 2310
rect 2780 2246 2832 2252
rect 3424 2304 3476 2310
rect 3424 2246 3476 2252
rect 4068 2304 4120 2310
rect 4068 2246 4120 2252
rect 4712 2304 4764 2310
rect 4712 2246 4764 2252
rect 5356 2304 5408 2310
rect 5356 2246 5408 2252
rect 6000 2304 6052 2310
rect 6000 2246 6052 2252
rect 2792 800 2820 2246
rect 3436 800 3464 2246
rect 4080 800 4108 2246
rect 4724 800 4752 2246
rect 5368 800 5396 2246
rect 6012 800 6040 2246
rect 6472 1442 6500 2858
rect 6630 2204 6938 2213
rect 6630 2202 6636 2204
rect 6692 2202 6716 2204
rect 6772 2202 6796 2204
rect 6852 2202 6876 2204
rect 6932 2202 6938 2204
rect 6692 2150 6694 2202
rect 6874 2150 6876 2202
rect 6630 2148 6636 2150
rect 6692 2148 6716 2150
rect 6772 2148 6796 2150
rect 6852 2148 6876 2150
rect 6932 2148 6938 2150
rect 6630 2139 6938 2148
rect 6472 1414 6684 1442
rect 6656 800 6684 1414
rect 7300 800 7328 2994
rect 7380 2984 7432 2990
rect 7380 2926 7432 2932
rect 7392 2446 7420 2926
rect 7484 2446 7512 3470
rect 7760 3466 7788 3606
rect 7852 3534 7880 4082
rect 8220 3534 8248 4082
rect 8300 4072 8352 4078
rect 8300 4014 8352 4020
rect 7840 3528 7892 3534
rect 7840 3470 7892 3476
rect 8208 3528 8260 3534
rect 8208 3470 8260 3476
rect 8312 3466 8340 4014
rect 7748 3460 7800 3466
rect 7748 3402 7800 3408
rect 8300 3460 8352 3466
rect 8300 3402 8352 3408
rect 7932 3120 7984 3126
rect 7932 3062 7984 3068
rect 7654 2952 7710 2961
rect 7654 2887 7710 2896
rect 7668 2446 7696 2887
rect 7838 2680 7894 2689
rect 7838 2615 7840 2624
rect 7892 2615 7894 2624
rect 7840 2586 7892 2592
rect 7380 2440 7432 2446
rect 7380 2382 7432 2388
rect 7472 2440 7524 2446
rect 7472 2382 7524 2388
rect 7656 2440 7708 2446
rect 7656 2382 7708 2388
rect 7944 800 7972 3062
rect 8300 3052 8352 3058
rect 8300 2994 8352 3000
rect 8312 2961 8340 2994
rect 8298 2952 8354 2961
rect 8298 2887 8354 2896
rect 8404 2774 8432 4678
rect 8484 4208 8536 4214
rect 8484 4150 8536 4156
rect 8496 3126 8524 4150
rect 8588 4078 8616 5646
rect 8680 5370 8708 6224
rect 8864 5370 8892 9318
rect 8956 8498 8984 9438
rect 8944 8492 8996 8498
rect 8944 8434 8996 8440
rect 8956 6934 8984 8434
rect 8944 6928 8996 6934
rect 8944 6870 8996 6876
rect 9048 6458 9076 11018
rect 9140 10266 9168 11086
rect 9128 10260 9180 10266
rect 9128 10202 9180 10208
rect 9128 8288 9180 8294
rect 9128 8230 9180 8236
rect 9140 7206 9168 8230
rect 9128 7200 9180 7206
rect 9128 7142 9180 7148
rect 9036 6452 9088 6458
rect 9036 6394 9088 6400
rect 8668 5364 8720 5370
rect 8668 5306 8720 5312
rect 8852 5364 8904 5370
rect 8852 5306 8904 5312
rect 8864 5234 8892 5306
rect 8852 5228 8904 5234
rect 8852 5170 8904 5176
rect 9232 5166 9260 11222
rect 9324 10810 9352 11698
rect 9692 11626 9720 12106
rect 9784 12073 9812 12174
rect 9864 12096 9916 12102
rect 9770 12064 9826 12073
rect 9864 12038 9916 12044
rect 9770 11999 9826 12008
rect 9680 11620 9732 11626
rect 9680 11562 9732 11568
rect 9471 11452 9779 11461
rect 9471 11450 9477 11452
rect 9533 11450 9557 11452
rect 9613 11450 9637 11452
rect 9693 11450 9717 11452
rect 9773 11450 9779 11452
rect 9533 11398 9535 11450
rect 9715 11398 9717 11450
rect 9471 11396 9477 11398
rect 9533 11396 9557 11398
rect 9613 11396 9637 11398
rect 9693 11396 9717 11398
rect 9773 11396 9779 11398
rect 9471 11387 9779 11396
rect 9876 11354 9904 12038
rect 9864 11348 9916 11354
rect 9864 11290 9916 11296
rect 9404 11280 9456 11286
rect 9404 11222 9456 11228
rect 9416 11150 9444 11222
rect 9404 11144 9456 11150
rect 9404 11086 9456 11092
rect 9312 10804 9364 10810
rect 9312 10746 9364 10752
rect 9402 10704 9458 10713
rect 9402 10639 9404 10648
rect 9456 10639 9458 10648
rect 9404 10610 9456 10616
rect 9864 10600 9916 10606
rect 9864 10542 9916 10548
rect 9312 10532 9364 10538
rect 9312 10474 9364 10480
rect 9324 10198 9352 10474
rect 9471 10364 9779 10373
rect 9471 10362 9477 10364
rect 9533 10362 9557 10364
rect 9613 10362 9637 10364
rect 9693 10362 9717 10364
rect 9773 10362 9779 10364
rect 9533 10310 9535 10362
rect 9715 10310 9717 10362
rect 9471 10308 9477 10310
rect 9533 10308 9557 10310
rect 9613 10308 9637 10310
rect 9693 10308 9717 10310
rect 9773 10308 9779 10310
rect 9471 10299 9779 10308
rect 9312 10192 9364 10198
rect 9312 10134 9364 10140
rect 9494 10160 9550 10169
rect 9494 10095 9550 10104
rect 9508 10062 9536 10095
rect 9312 10056 9364 10062
rect 9312 9998 9364 10004
rect 9496 10056 9548 10062
rect 9496 9998 9548 10004
rect 9324 9761 9352 9998
rect 9310 9752 9366 9761
rect 9310 9687 9366 9696
rect 9508 9674 9536 9998
rect 9876 9994 9904 10542
rect 9968 10266 9996 14214
rect 10048 12912 10100 12918
rect 10048 12854 10100 12860
rect 10060 12102 10088 12854
rect 10048 12096 10100 12102
rect 10048 12038 10100 12044
rect 10048 10464 10100 10470
rect 10048 10406 10100 10412
rect 9956 10260 10008 10266
rect 9956 10202 10008 10208
rect 9864 9988 9916 9994
rect 9864 9930 9916 9936
rect 10060 9926 10088 10406
rect 10048 9920 10100 9926
rect 10048 9862 10100 9868
rect 9416 9646 9536 9674
rect 9416 9382 9444 9646
rect 10048 9580 10100 9586
rect 10048 9522 10100 9528
rect 9404 9376 9456 9382
rect 9404 9318 9456 9324
rect 9864 9376 9916 9382
rect 9864 9318 9916 9324
rect 9471 9276 9779 9285
rect 9471 9274 9477 9276
rect 9533 9274 9557 9276
rect 9613 9274 9637 9276
rect 9693 9274 9717 9276
rect 9773 9274 9779 9276
rect 9533 9222 9535 9274
rect 9715 9222 9717 9274
rect 9471 9220 9477 9222
rect 9533 9220 9557 9222
rect 9613 9220 9637 9222
rect 9693 9220 9717 9222
rect 9773 9220 9779 9222
rect 9471 9211 9779 9220
rect 9496 8968 9548 8974
rect 9496 8910 9548 8916
rect 9508 8294 9536 8910
rect 9876 8809 9904 9318
rect 10060 8906 10088 9522
rect 10152 9217 10180 21898
rect 11244 21548 11296 21554
rect 11244 21490 11296 21496
rect 11060 21412 11112 21418
rect 11060 21354 11112 21360
rect 10416 20256 10468 20262
rect 10416 20198 10468 20204
rect 10428 14550 10456 20198
rect 10784 19712 10836 19718
rect 10784 19654 10836 19660
rect 10968 19712 11020 19718
rect 10968 19654 11020 19660
rect 10692 15360 10744 15366
rect 10692 15302 10744 15308
rect 10508 14816 10560 14822
rect 10508 14758 10560 14764
rect 10416 14544 10468 14550
rect 10416 14486 10468 14492
rect 10416 13728 10468 13734
rect 10416 13670 10468 13676
rect 10232 11620 10284 11626
rect 10232 11562 10284 11568
rect 10244 11218 10272 11562
rect 10324 11552 10376 11558
rect 10324 11494 10376 11500
rect 10232 11212 10284 11218
rect 10232 11154 10284 11160
rect 10336 11150 10364 11494
rect 10324 11144 10376 11150
rect 10324 11086 10376 11092
rect 10232 9648 10284 9654
rect 10232 9590 10284 9596
rect 10138 9208 10194 9217
rect 10138 9143 10194 9152
rect 10048 8900 10100 8906
rect 10048 8842 10100 8848
rect 9956 8832 10008 8838
rect 9862 8800 9918 8809
rect 9956 8774 10008 8780
rect 9862 8735 9918 8744
rect 9864 8560 9916 8566
rect 9864 8502 9916 8508
rect 9312 8288 9364 8294
rect 9312 8230 9364 8236
rect 9496 8288 9548 8294
rect 9496 8230 9548 8236
rect 9324 7546 9352 8230
rect 9471 8188 9779 8197
rect 9471 8186 9477 8188
rect 9533 8186 9557 8188
rect 9613 8186 9637 8188
rect 9693 8186 9717 8188
rect 9773 8186 9779 8188
rect 9533 8134 9535 8186
rect 9715 8134 9717 8186
rect 9471 8132 9477 8134
rect 9533 8132 9557 8134
rect 9613 8132 9637 8134
rect 9693 8132 9717 8134
rect 9773 8132 9779 8134
rect 9471 8123 9779 8132
rect 9876 8090 9904 8502
rect 9864 8084 9916 8090
rect 9864 8026 9916 8032
rect 9588 7744 9640 7750
rect 9588 7686 9640 7692
rect 9312 7540 9364 7546
rect 9312 7482 9364 7488
rect 9600 7410 9628 7686
rect 9312 7404 9364 7410
rect 9312 7346 9364 7352
rect 9588 7404 9640 7410
rect 9588 7346 9640 7352
rect 9324 6458 9352 7346
rect 9864 7200 9916 7206
rect 9864 7142 9916 7148
rect 9471 7100 9779 7109
rect 9471 7098 9477 7100
rect 9533 7098 9557 7100
rect 9613 7098 9637 7100
rect 9693 7098 9717 7100
rect 9773 7098 9779 7100
rect 9533 7046 9535 7098
rect 9715 7046 9717 7098
rect 9471 7044 9477 7046
rect 9533 7044 9557 7046
rect 9613 7044 9637 7046
rect 9693 7044 9717 7046
rect 9773 7044 9779 7046
rect 9471 7035 9779 7044
rect 9496 6928 9548 6934
rect 9496 6870 9548 6876
rect 9508 6798 9536 6870
rect 9496 6792 9548 6798
rect 9496 6734 9548 6740
rect 9404 6656 9456 6662
rect 9404 6598 9456 6604
rect 9312 6452 9364 6458
rect 9312 6394 9364 6400
rect 9416 6338 9444 6598
rect 9324 6310 9444 6338
rect 9324 5574 9352 6310
rect 9471 6012 9779 6021
rect 9471 6010 9477 6012
rect 9533 6010 9557 6012
rect 9613 6010 9637 6012
rect 9693 6010 9717 6012
rect 9773 6010 9779 6012
rect 9533 5958 9535 6010
rect 9715 5958 9717 6010
rect 9471 5956 9477 5958
rect 9533 5956 9557 5958
rect 9613 5956 9637 5958
rect 9693 5956 9717 5958
rect 9773 5956 9779 5958
rect 9471 5947 9779 5956
rect 9772 5840 9824 5846
rect 9494 5808 9550 5817
rect 9772 5782 9824 5788
rect 9494 5743 9550 5752
rect 9508 5710 9536 5743
rect 9496 5704 9548 5710
rect 9496 5646 9548 5652
rect 9312 5568 9364 5574
rect 9312 5510 9364 5516
rect 8760 5160 8812 5166
rect 8760 5102 8812 5108
rect 9220 5160 9272 5166
rect 9272 5108 9352 5114
rect 9220 5102 9352 5108
rect 8576 4072 8628 4078
rect 8576 4014 8628 4020
rect 8772 3738 8800 5102
rect 9036 5092 9088 5098
rect 9232 5086 9352 5102
rect 9508 5098 9536 5646
rect 9036 5034 9088 5040
rect 8760 3732 8812 3738
rect 8760 3674 8812 3680
rect 8852 3596 8904 3602
rect 8852 3538 8904 3544
rect 8576 3392 8628 3398
rect 8576 3334 8628 3340
rect 8484 3120 8536 3126
rect 8484 3062 8536 3068
rect 8484 2984 8536 2990
rect 8484 2926 8536 2932
rect 8312 2746 8432 2774
rect 8312 2514 8340 2746
rect 8496 2650 8524 2926
rect 8484 2644 8536 2650
rect 8484 2586 8536 2592
rect 8300 2508 8352 2514
rect 8300 2450 8352 2456
rect 8206 2408 8262 2417
rect 8206 2343 8262 2352
rect 8220 2106 8248 2343
rect 8208 2100 8260 2106
rect 8208 2042 8260 2048
rect 8588 800 8616 3334
rect 8864 3058 8892 3538
rect 8944 3120 8996 3126
rect 8944 3062 8996 3068
rect 8852 3052 8904 3058
rect 8852 2994 8904 3000
rect 8956 2514 8984 3062
rect 8944 2508 8996 2514
rect 8944 2450 8996 2456
rect 9048 2446 9076 5034
rect 9220 5024 9272 5030
rect 9220 4966 9272 4972
rect 9128 4140 9180 4146
rect 9128 4082 9180 4088
rect 9140 3534 9168 4082
rect 9232 4078 9260 4966
rect 9324 4622 9352 5086
rect 9496 5092 9548 5098
rect 9784 5080 9812 5782
rect 9876 5710 9904 7142
rect 9864 5704 9916 5710
rect 9864 5646 9916 5652
rect 9784 5052 9904 5080
rect 9496 5034 9548 5040
rect 9471 4924 9779 4933
rect 9471 4922 9477 4924
rect 9533 4922 9557 4924
rect 9613 4922 9637 4924
rect 9693 4922 9717 4924
rect 9773 4922 9779 4924
rect 9533 4870 9535 4922
rect 9715 4870 9717 4922
rect 9471 4868 9477 4870
rect 9533 4868 9557 4870
rect 9613 4868 9637 4870
rect 9693 4868 9717 4870
rect 9773 4868 9779 4870
rect 9471 4859 9779 4868
rect 9876 4758 9904 5052
rect 9864 4752 9916 4758
rect 9864 4694 9916 4700
rect 9312 4616 9364 4622
rect 9364 4564 9536 4570
rect 9312 4558 9536 4564
rect 9324 4554 9536 4558
rect 9324 4548 9548 4554
rect 9324 4542 9496 4548
rect 9220 4072 9272 4078
rect 9220 4014 9272 4020
rect 9232 3602 9260 4014
rect 9220 3596 9272 3602
rect 9220 3538 9272 3544
rect 9128 3528 9180 3534
rect 9128 3470 9180 3476
rect 9140 3194 9168 3470
rect 9128 3188 9180 3194
rect 9128 3130 9180 3136
rect 9220 3120 9272 3126
rect 9220 3062 9272 3068
rect 9036 2440 9088 2446
rect 9036 2382 9088 2388
rect 9232 800 9260 3062
rect 9324 3058 9352 4542
rect 9496 4490 9548 4496
rect 9968 4146 9996 8774
rect 10244 8634 10272 9590
rect 10336 9586 10364 11086
rect 10324 9580 10376 9586
rect 10324 9522 10376 9528
rect 10336 8974 10364 9522
rect 10324 8968 10376 8974
rect 10324 8910 10376 8916
rect 10322 8800 10378 8809
rect 10322 8735 10378 8744
rect 10232 8628 10284 8634
rect 10232 8570 10284 8576
rect 10048 8560 10100 8566
rect 10048 8502 10100 8508
rect 10060 7886 10088 8502
rect 10048 7880 10100 7886
rect 10048 7822 10100 7828
rect 10060 6186 10088 7822
rect 10244 6662 10272 8570
rect 10232 6656 10284 6662
rect 10232 6598 10284 6604
rect 10140 6316 10192 6322
rect 10140 6258 10192 6264
rect 10048 6180 10100 6186
rect 10048 6122 10100 6128
rect 10060 5846 10088 6122
rect 10048 5840 10100 5846
rect 10048 5782 10100 5788
rect 10048 5704 10100 5710
rect 10048 5646 10100 5652
rect 10060 4758 10088 5646
rect 10152 5302 10180 6258
rect 10232 6248 10284 6254
rect 10232 6190 10284 6196
rect 10140 5296 10192 5302
rect 10140 5238 10192 5244
rect 10048 4752 10100 4758
rect 10048 4694 10100 4700
rect 10244 4622 10272 6190
rect 10232 4616 10284 4622
rect 10232 4558 10284 4564
rect 10336 4554 10364 8735
rect 10428 8566 10456 13670
rect 10520 12434 10548 14758
rect 10704 13870 10732 15302
rect 10796 15094 10824 19654
rect 10876 17536 10928 17542
rect 10876 17478 10928 17484
rect 10784 15088 10836 15094
rect 10784 15030 10836 15036
rect 10784 14816 10836 14822
rect 10784 14758 10836 14764
rect 10796 14618 10824 14758
rect 10784 14612 10836 14618
rect 10784 14554 10836 14560
rect 10796 13938 10824 14554
rect 10784 13932 10836 13938
rect 10784 13874 10836 13880
rect 10692 13864 10744 13870
rect 10692 13806 10744 13812
rect 10784 13796 10836 13802
rect 10784 13738 10836 13744
rect 10796 13530 10824 13738
rect 10784 13524 10836 13530
rect 10784 13466 10836 13472
rect 10520 12406 10732 12434
rect 10600 12096 10652 12102
rect 10600 12038 10652 12044
rect 10612 11694 10640 12038
rect 10600 11688 10652 11694
rect 10600 11630 10652 11636
rect 10612 11082 10640 11630
rect 10600 11076 10652 11082
rect 10600 11018 10652 11024
rect 10508 9512 10560 9518
rect 10508 9454 10560 9460
rect 10416 8560 10468 8566
rect 10416 8502 10468 8508
rect 10416 8288 10468 8294
rect 10416 8230 10468 8236
rect 10428 7954 10456 8230
rect 10416 7948 10468 7954
rect 10416 7890 10468 7896
rect 10416 7336 10468 7342
rect 10416 7278 10468 7284
rect 10428 5846 10456 7278
rect 10520 6254 10548 9454
rect 10612 9382 10640 11018
rect 10600 9376 10652 9382
rect 10600 9318 10652 9324
rect 10600 8832 10652 8838
rect 10600 8774 10652 8780
rect 10612 7886 10640 8774
rect 10600 7880 10652 7886
rect 10600 7822 10652 7828
rect 10612 7002 10640 7822
rect 10600 6996 10652 7002
rect 10600 6938 10652 6944
rect 10508 6248 10560 6254
rect 10508 6190 10560 6196
rect 10416 5840 10468 5846
rect 10416 5782 10468 5788
rect 10520 5302 10548 6190
rect 10704 6118 10732 12406
rect 10784 11620 10836 11626
rect 10784 11562 10836 11568
rect 10796 8090 10824 11562
rect 10888 9926 10916 17478
rect 10980 11898 11008 19654
rect 11072 16046 11100 21354
rect 11152 21140 11204 21146
rect 11152 21082 11204 21088
rect 11164 20466 11192 21082
rect 11152 20460 11204 20466
rect 11152 20402 11204 20408
rect 11164 19922 11192 20402
rect 11256 20262 11284 21490
rect 11244 20256 11296 20262
rect 11244 20198 11296 20204
rect 11152 19916 11204 19922
rect 11152 19858 11204 19864
rect 11152 17672 11204 17678
rect 11152 17614 11204 17620
rect 11060 16040 11112 16046
rect 11060 15982 11112 15988
rect 11060 15904 11112 15910
rect 11060 15846 11112 15852
rect 11072 15502 11100 15846
rect 11164 15570 11192 17614
rect 11152 15564 11204 15570
rect 11152 15506 11204 15512
rect 11060 15496 11112 15502
rect 11060 15438 11112 15444
rect 11072 14958 11100 15438
rect 11152 15360 11204 15366
rect 11152 15302 11204 15308
rect 11060 14952 11112 14958
rect 11060 14894 11112 14900
rect 11060 14340 11112 14346
rect 11060 14282 11112 14288
rect 11072 13394 11100 14282
rect 11060 13388 11112 13394
rect 11060 13330 11112 13336
rect 10968 11892 11020 11898
rect 10968 11834 11020 11840
rect 10968 11756 11020 11762
rect 10968 11698 11020 11704
rect 10980 10742 11008 11698
rect 11164 10810 11192 15302
rect 11256 14890 11284 20198
rect 11244 14884 11296 14890
rect 11244 14826 11296 14832
rect 11244 14408 11296 14414
rect 11244 14350 11296 14356
rect 11256 13530 11284 14350
rect 11348 14074 11376 21898
rect 11428 21888 11480 21894
rect 11428 21830 11480 21836
rect 11440 15570 11468 21830
rect 12311 21788 12619 21797
rect 12311 21786 12317 21788
rect 12373 21786 12397 21788
rect 12453 21786 12477 21788
rect 12533 21786 12557 21788
rect 12613 21786 12619 21788
rect 12373 21734 12375 21786
rect 12555 21734 12557 21786
rect 12311 21732 12317 21734
rect 12373 21732 12397 21734
rect 12453 21732 12477 21734
rect 12533 21732 12557 21734
rect 12613 21732 12619 21734
rect 12311 21723 12619 21732
rect 13096 21486 13124 21966
rect 14384 21962 14596 21978
rect 17408 21966 17460 21972
rect 22376 22024 22428 22030
rect 22376 21966 22428 21972
rect 14372 21956 14608 21962
rect 14424 21950 14556 21956
rect 14372 21898 14424 21904
rect 14556 21898 14608 21904
rect 13544 21888 13596 21894
rect 13544 21830 13596 21836
rect 13728 21888 13780 21894
rect 13728 21830 13780 21836
rect 13084 21480 13136 21486
rect 13084 21422 13136 21428
rect 13360 21412 13412 21418
rect 13360 21354 13412 21360
rect 11520 21344 11572 21350
rect 11520 21286 11572 21292
rect 11796 21344 11848 21350
rect 11796 21286 11848 21292
rect 11428 15564 11480 15570
rect 11428 15506 11480 15512
rect 11532 15026 11560 21286
rect 11808 21146 11836 21286
rect 11796 21140 11848 21146
rect 11796 21082 11848 21088
rect 13372 20942 13400 21354
rect 13452 21344 13504 21350
rect 13452 21286 13504 21292
rect 13464 21010 13492 21286
rect 13452 21004 13504 21010
rect 13452 20946 13504 20952
rect 13360 20936 13412 20942
rect 13360 20878 13412 20884
rect 12311 20700 12619 20709
rect 12311 20698 12317 20700
rect 12373 20698 12397 20700
rect 12453 20698 12477 20700
rect 12533 20698 12557 20700
rect 12613 20698 12619 20700
rect 12373 20646 12375 20698
rect 12555 20646 12557 20698
rect 12311 20644 12317 20646
rect 12373 20644 12397 20646
rect 12453 20644 12477 20646
rect 12533 20644 12557 20646
rect 12613 20644 12619 20646
rect 12311 20635 12619 20644
rect 12716 20528 12768 20534
rect 12716 20470 12768 20476
rect 11704 19848 11756 19854
rect 11704 19790 11756 19796
rect 11612 19712 11664 19718
rect 11612 19654 11664 19660
rect 11624 15162 11652 19654
rect 11716 18834 11744 19790
rect 12311 19612 12619 19621
rect 12311 19610 12317 19612
rect 12373 19610 12397 19612
rect 12453 19610 12477 19612
rect 12533 19610 12557 19612
rect 12613 19610 12619 19612
rect 12373 19558 12375 19610
rect 12555 19558 12557 19610
rect 12311 19556 12317 19558
rect 12373 19556 12397 19558
rect 12453 19556 12477 19558
rect 12533 19556 12557 19558
rect 12613 19556 12619 19558
rect 12311 19547 12619 19556
rect 11704 18828 11756 18834
rect 11704 18770 11756 18776
rect 11704 18624 11756 18630
rect 11704 18566 11756 18572
rect 11612 15156 11664 15162
rect 11612 15098 11664 15104
rect 11520 15020 11572 15026
rect 11520 14962 11572 14968
rect 11428 14884 11480 14890
rect 11428 14826 11480 14832
rect 11336 14068 11388 14074
rect 11336 14010 11388 14016
rect 11244 13524 11296 13530
rect 11244 13466 11296 13472
rect 11336 13388 11388 13394
rect 11336 13330 11388 13336
rect 11348 12918 11376 13330
rect 11336 12912 11388 12918
rect 11336 12854 11388 12860
rect 11244 12436 11296 12442
rect 11244 12378 11296 12384
rect 11152 10804 11204 10810
rect 11256 10792 11284 12378
rect 11348 11286 11376 12854
rect 11440 11830 11468 14826
rect 11532 14550 11560 14962
rect 11612 14612 11664 14618
rect 11612 14554 11664 14560
rect 11520 14544 11572 14550
rect 11520 14486 11572 14492
rect 11520 13864 11572 13870
rect 11520 13806 11572 13812
rect 11428 11824 11480 11830
rect 11428 11766 11480 11772
rect 11336 11280 11388 11286
rect 11336 11222 11388 11228
rect 11256 10764 11376 10792
rect 11152 10746 11204 10752
rect 10968 10736 11020 10742
rect 10968 10678 11020 10684
rect 11060 10532 11112 10538
rect 11060 10474 11112 10480
rect 10968 10056 11020 10062
rect 10968 9998 11020 10004
rect 10876 9920 10928 9926
rect 10876 9862 10928 9868
rect 10980 9761 11008 9998
rect 10966 9752 11022 9761
rect 10966 9687 11022 9696
rect 11072 9654 11100 10474
rect 11348 9674 11376 10764
rect 11440 10674 11468 11766
rect 11428 10668 11480 10674
rect 11428 10610 11480 10616
rect 11440 9722 11468 10610
rect 11532 10062 11560 13806
rect 11624 13326 11652 14554
rect 11716 14414 11744 18566
rect 12311 18524 12619 18533
rect 12311 18522 12317 18524
rect 12373 18522 12397 18524
rect 12453 18522 12477 18524
rect 12533 18522 12557 18524
rect 12613 18522 12619 18524
rect 12373 18470 12375 18522
rect 12555 18470 12557 18522
rect 12311 18468 12317 18470
rect 12373 18468 12397 18470
rect 12453 18468 12477 18470
rect 12533 18468 12557 18470
rect 12613 18468 12619 18470
rect 12311 18459 12619 18468
rect 12072 18284 12124 18290
rect 12072 18226 12124 18232
rect 11888 18148 11940 18154
rect 11888 18090 11940 18096
rect 11796 18080 11848 18086
rect 11796 18022 11848 18028
rect 11808 17610 11836 18022
rect 11796 17604 11848 17610
rect 11796 17546 11848 17552
rect 11808 17338 11836 17546
rect 11796 17332 11848 17338
rect 11796 17274 11848 17280
rect 11796 17196 11848 17202
rect 11796 17138 11848 17144
rect 11808 16998 11836 17138
rect 11796 16992 11848 16998
rect 11796 16934 11848 16940
rect 11808 15910 11836 16934
rect 11796 15904 11848 15910
rect 11796 15846 11848 15852
rect 11704 14408 11756 14414
rect 11704 14350 11756 14356
rect 11796 14340 11848 14346
rect 11796 14282 11848 14288
rect 11704 13524 11756 13530
rect 11704 13466 11756 13472
rect 11612 13320 11664 13326
rect 11612 13262 11664 13268
rect 11716 12850 11744 13466
rect 11704 12844 11756 12850
rect 11704 12786 11756 12792
rect 11612 11280 11664 11286
rect 11612 11222 11664 11228
rect 11624 11150 11652 11222
rect 11612 11144 11664 11150
rect 11612 11086 11664 11092
rect 11624 10130 11652 11086
rect 11716 11082 11744 12786
rect 11808 12102 11836 14282
rect 11900 12434 11928 18090
rect 11980 16448 12032 16454
rect 11980 16390 12032 16396
rect 11992 15502 12020 16390
rect 11980 15496 12032 15502
rect 11980 15438 12032 15444
rect 12084 12442 12112 18226
rect 12311 17436 12619 17445
rect 12311 17434 12317 17436
rect 12373 17434 12397 17436
rect 12453 17434 12477 17436
rect 12533 17434 12557 17436
rect 12613 17434 12619 17436
rect 12373 17382 12375 17434
rect 12555 17382 12557 17434
rect 12311 17380 12317 17382
rect 12373 17380 12397 17382
rect 12453 17380 12477 17382
rect 12533 17380 12557 17382
rect 12613 17380 12619 17382
rect 12311 17371 12619 17380
rect 12311 16348 12619 16357
rect 12311 16346 12317 16348
rect 12373 16346 12397 16348
rect 12453 16346 12477 16348
rect 12533 16346 12557 16348
rect 12613 16346 12619 16348
rect 12373 16294 12375 16346
rect 12555 16294 12557 16346
rect 12311 16292 12317 16294
rect 12373 16292 12397 16294
rect 12453 16292 12477 16294
rect 12533 16292 12557 16294
rect 12613 16292 12619 16294
rect 12311 16283 12619 16292
rect 12176 15570 12296 15586
rect 12176 15564 12308 15570
rect 12176 15558 12256 15564
rect 12176 14006 12204 15558
rect 12256 15506 12308 15512
rect 12311 15260 12619 15269
rect 12311 15258 12317 15260
rect 12373 15258 12397 15260
rect 12453 15258 12477 15260
rect 12533 15258 12557 15260
rect 12613 15258 12619 15260
rect 12373 15206 12375 15258
rect 12555 15206 12557 15258
rect 12311 15204 12317 15206
rect 12373 15204 12397 15206
rect 12453 15204 12477 15206
rect 12533 15204 12557 15206
rect 12613 15204 12619 15206
rect 12311 15195 12619 15204
rect 12348 14816 12400 14822
rect 12348 14758 12400 14764
rect 12360 14346 12388 14758
rect 12728 14414 12756 20470
rect 13452 18624 13504 18630
rect 13452 18566 13504 18572
rect 12992 17604 13044 17610
rect 12992 17546 13044 17552
rect 12808 16108 12860 16114
rect 12808 16050 12860 16056
rect 12820 15706 12848 16050
rect 12808 15700 12860 15706
rect 12808 15642 12860 15648
rect 12808 15496 12860 15502
rect 12808 15438 12860 15444
rect 12820 15026 12848 15438
rect 12808 15020 12860 15026
rect 12808 14962 12860 14968
rect 12820 14618 12848 14962
rect 12808 14612 12860 14618
rect 12808 14554 12860 14560
rect 12716 14408 12768 14414
rect 12716 14350 12768 14356
rect 12348 14340 12400 14346
rect 12348 14282 12400 14288
rect 12311 14172 12619 14181
rect 12311 14170 12317 14172
rect 12373 14170 12397 14172
rect 12453 14170 12477 14172
rect 12533 14170 12557 14172
rect 12613 14170 12619 14172
rect 12373 14118 12375 14170
rect 12555 14118 12557 14170
rect 12311 14116 12317 14118
rect 12373 14116 12397 14118
rect 12453 14116 12477 14118
rect 12533 14116 12557 14118
rect 12613 14116 12619 14118
rect 12311 14107 12619 14116
rect 12164 14000 12216 14006
rect 12164 13942 12216 13948
rect 12164 13864 12216 13870
rect 12164 13806 12216 13812
rect 12176 13530 12204 13806
rect 13004 13802 13032 17546
rect 13084 17060 13136 17066
rect 13084 17002 13136 17008
rect 13096 15502 13124 17002
rect 13084 15496 13136 15502
rect 13084 15438 13136 15444
rect 13268 15496 13320 15502
rect 13268 15438 13320 15444
rect 13096 15094 13124 15438
rect 13280 15162 13308 15438
rect 13268 15156 13320 15162
rect 13268 15098 13320 15104
rect 13084 15088 13136 15094
rect 13084 15030 13136 15036
rect 13464 14634 13492 18566
rect 13556 14822 13584 21830
rect 13740 20466 13768 21830
rect 14188 21480 14240 21486
rect 14188 21422 14240 21428
rect 14200 20602 14228 21422
rect 14188 20596 14240 20602
rect 14188 20538 14240 20544
rect 14384 20534 14412 21898
rect 14648 21888 14700 21894
rect 14648 21830 14700 21836
rect 17500 21888 17552 21894
rect 17500 21830 17552 21836
rect 14660 21554 14688 21830
rect 14648 21548 14700 21554
rect 14648 21490 14700 21496
rect 17512 21418 17540 21830
rect 17992 21788 18300 21797
rect 17992 21786 17998 21788
rect 18054 21786 18078 21788
rect 18134 21786 18158 21788
rect 18214 21786 18238 21788
rect 18294 21786 18300 21788
rect 18054 21734 18056 21786
rect 18236 21734 18238 21786
rect 17992 21732 17998 21734
rect 18054 21732 18078 21734
rect 18134 21732 18158 21734
rect 18214 21732 18238 21734
rect 18294 21732 18300 21734
rect 17992 21723 18300 21732
rect 23673 21788 23981 21797
rect 23673 21786 23679 21788
rect 23735 21786 23759 21788
rect 23815 21786 23839 21788
rect 23895 21786 23919 21788
rect 23975 21786 23981 21788
rect 23735 21734 23737 21786
rect 23917 21734 23919 21786
rect 23673 21732 23679 21734
rect 23735 21732 23759 21734
rect 23815 21732 23839 21734
rect 23895 21732 23919 21734
rect 23975 21732 23981 21734
rect 23673 21723 23981 21732
rect 17500 21412 17552 21418
rect 17500 21354 17552 21360
rect 15152 21244 15460 21253
rect 15152 21242 15158 21244
rect 15214 21242 15238 21244
rect 15294 21242 15318 21244
rect 15374 21242 15398 21244
rect 15454 21242 15460 21244
rect 15214 21190 15216 21242
rect 15396 21190 15398 21242
rect 15152 21188 15158 21190
rect 15214 21188 15238 21190
rect 15294 21188 15318 21190
rect 15374 21188 15398 21190
rect 15454 21188 15460 21190
rect 15152 21179 15460 21188
rect 20833 21244 21141 21253
rect 20833 21242 20839 21244
rect 20895 21242 20919 21244
rect 20975 21242 20999 21244
rect 21055 21242 21079 21244
rect 21135 21242 21141 21244
rect 20895 21190 20897 21242
rect 21077 21190 21079 21242
rect 20833 21188 20839 21190
rect 20895 21188 20919 21190
rect 20975 21188 20999 21190
rect 21055 21188 21079 21190
rect 21135 21188 21141 21190
rect 20833 21179 21141 21188
rect 17992 20700 18300 20709
rect 17992 20698 17998 20700
rect 18054 20698 18078 20700
rect 18134 20698 18158 20700
rect 18214 20698 18238 20700
rect 18294 20698 18300 20700
rect 18054 20646 18056 20698
rect 18236 20646 18238 20698
rect 17992 20644 17998 20646
rect 18054 20644 18078 20646
rect 18134 20644 18158 20646
rect 18214 20644 18238 20646
rect 18294 20644 18300 20646
rect 17992 20635 18300 20644
rect 23673 20700 23981 20709
rect 23673 20698 23679 20700
rect 23735 20698 23759 20700
rect 23815 20698 23839 20700
rect 23895 20698 23919 20700
rect 23975 20698 23981 20700
rect 23735 20646 23737 20698
rect 23917 20646 23919 20698
rect 23673 20644 23679 20646
rect 23735 20644 23759 20646
rect 23815 20644 23839 20646
rect 23895 20644 23919 20646
rect 23975 20644 23981 20646
rect 23673 20635 23981 20644
rect 14372 20528 14424 20534
rect 14372 20470 14424 20476
rect 13728 20460 13780 20466
rect 13728 20402 13780 20408
rect 15152 20156 15460 20165
rect 15152 20154 15158 20156
rect 15214 20154 15238 20156
rect 15294 20154 15318 20156
rect 15374 20154 15398 20156
rect 15454 20154 15460 20156
rect 15214 20102 15216 20154
rect 15396 20102 15398 20154
rect 15152 20100 15158 20102
rect 15214 20100 15238 20102
rect 15294 20100 15318 20102
rect 15374 20100 15398 20102
rect 15454 20100 15460 20102
rect 15152 20091 15460 20100
rect 20833 20156 21141 20165
rect 20833 20154 20839 20156
rect 20895 20154 20919 20156
rect 20975 20154 20999 20156
rect 21055 20154 21079 20156
rect 21135 20154 21141 20156
rect 20895 20102 20897 20154
rect 21077 20102 21079 20154
rect 20833 20100 20839 20102
rect 20895 20100 20919 20102
rect 20975 20100 20999 20102
rect 21055 20100 21079 20102
rect 21135 20100 21141 20102
rect 20833 20091 21141 20100
rect 18328 19780 18380 19786
rect 18328 19722 18380 19728
rect 17992 19612 18300 19621
rect 17992 19610 17998 19612
rect 18054 19610 18078 19612
rect 18134 19610 18158 19612
rect 18214 19610 18238 19612
rect 18294 19610 18300 19612
rect 18054 19558 18056 19610
rect 18236 19558 18238 19610
rect 17992 19556 17998 19558
rect 18054 19556 18078 19558
rect 18134 19556 18158 19558
rect 18214 19556 18238 19558
rect 18294 19556 18300 19558
rect 17992 19547 18300 19556
rect 15152 19068 15460 19077
rect 15152 19066 15158 19068
rect 15214 19066 15238 19068
rect 15294 19066 15318 19068
rect 15374 19066 15398 19068
rect 15454 19066 15460 19068
rect 15214 19014 15216 19066
rect 15396 19014 15398 19066
rect 15152 19012 15158 19014
rect 15214 19012 15238 19014
rect 15294 19012 15318 19014
rect 15374 19012 15398 19014
rect 15454 19012 15460 19014
rect 15152 19003 15460 19012
rect 18340 18970 18368 19722
rect 23673 19612 23981 19621
rect 23673 19610 23679 19612
rect 23735 19610 23759 19612
rect 23815 19610 23839 19612
rect 23895 19610 23919 19612
rect 23975 19610 23981 19612
rect 23735 19558 23737 19610
rect 23917 19558 23919 19610
rect 23673 19556 23679 19558
rect 23735 19556 23759 19558
rect 23815 19556 23839 19558
rect 23895 19556 23919 19558
rect 23975 19556 23981 19558
rect 23673 19547 23981 19556
rect 20833 19068 21141 19077
rect 20833 19066 20839 19068
rect 20895 19066 20919 19068
rect 20975 19066 20999 19068
rect 21055 19066 21079 19068
rect 21135 19066 21141 19068
rect 20895 19014 20897 19066
rect 21077 19014 21079 19066
rect 20833 19012 20839 19014
rect 20895 19012 20919 19014
rect 20975 19012 20999 19014
rect 21055 19012 21079 19014
rect 21135 19012 21141 19014
rect 20833 19003 21141 19012
rect 18328 18964 18380 18970
rect 18328 18906 18380 18912
rect 18420 18760 18472 18766
rect 18420 18702 18472 18708
rect 17992 18524 18300 18533
rect 17992 18522 17998 18524
rect 18054 18522 18078 18524
rect 18134 18522 18158 18524
rect 18214 18522 18238 18524
rect 18294 18522 18300 18524
rect 18054 18470 18056 18522
rect 18236 18470 18238 18522
rect 17992 18468 17998 18470
rect 18054 18468 18078 18470
rect 18134 18468 18158 18470
rect 18214 18468 18238 18470
rect 18294 18468 18300 18470
rect 17992 18459 18300 18468
rect 15152 17980 15460 17989
rect 15152 17978 15158 17980
rect 15214 17978 15238 17980
rect 15294 17978 15318 17980
rect 15374 17978 15398 17980
rect 15454 17978 15460 17980
rect 15214 17926 15216 17978
rect 15396 17926 15398 17978
rect 15152 17924 15158 17926
rect 15214 17924 15238 17926
rect 15294 17924 15318 17926
rect 15374 17924 15398 17926
rect 15454 17924 15460 17926
rect 15152 17915 15460 17924
rect 16028 17536 16080 17542
rect 16028 17478 16080 17484
rect 14004 17332 14056 17338
rect 14004 17274 14056 17280
rect 13636 15564 13688 15570
rect 13636 15506 13688 15512
rect 13544 14816 13596 14822
rect 13544 14758 13596 14764
rect 13464 14606 13584 14634
rect 13084 14408 13136 14414
rect 13084 14350 13136 14356
rect 12992 13796 13044 13802
rect 12992 13738 13044 13744
rect 12440 13728 12492 13734
rect 12440 13670 12492 13676
rect 12164 13524 12216 13530
rect 12164 13466 12216 13472
rect 12164 13388 12216 13394
rect 12164 13330 12216 13336
rect 12072 12436 12124 12442
rect 11900 12406 12020 12434
rect 11796 12096 11848 12102
rect 11796 12038 11848 12044
rect 11888 11756 11940 11762
rect 11888 11698 11940 11704
rect 11704 11076 11756 11082
rect 11756 11036 11836 11064
rect 11704 11018 11756 11024
rect 11704 10532 11756 10538
rect 11704 10474 11756 10480
rect 11716 10266 11744 10474
rect 11704 10260 11756 10266
rect 11704 10202 11756 10208
rect 11808 10146 11836 11036
rect 11900 10810 11928 11698
rect 11888 10804 11940 10810
rect 11888 10746 11940 10752
rect 11716 10130 11836 10146
rect 11612 10124 11664 10130
rect 11612 10066 11664 10072
rect 11704 10124 11836 10130
rect 11756 10118 11836 10124
rect 11704 10066 11756 10072
rect 11520 10056 11572 10062
rect 11520 9998 11572 10004
rect 11060 9648 11112 9654
rect 11060 9590 11112 9596
rect 11256 9646 11376 9674
rect 11428 9716 11480 9722
rect 11428 9658 11480 9664
rect 11256 9568 11284 9646
rect 11164 9540 11284 9568
rect 10968 9512 11020 9518
rect 10968 9454 11020 9460
rect 10784 8084 10836 8090
rect 10784 8026 10836 8032
rect 10692 6112 10744 6118
rect 10692 6054 10744 6060
rect 10796 5710 10824 8026
rect 10876 6316 10928 6322
rect 10876 6258 10928 6264
rect 10784 5704 10836 5710
rect 10784 5646 10836 5652
rect 10508 5296 10560 5302
rect 10508 5238 10560 5244
rect 10520 4554 10548 5238
rect 10796 5234 10824 5646
rect 10784 5228 10836 5234
rect 10704 5188 10784 5216
rect 10600 4752 10652 4758
rect 10600 4694 10652 4700
rect 10324 4548 10376 4554
rect 10324 4490 10376 4496
rect 10508 4548 10560 4554
rect 10508 4490 10560 4496
rect 9956 4140 10008 4146
rect 9956 4082 10008 4088
rect 9471 3836 9779 3845
rect 9471 3834 9477 3836
rect 9533 3834 9557 3836
rect 9613 3834 9637 3836
rect 9693 3834 9717 3836
rect 9773 3834 9779 3836
rect 9533 3782 9535 3834
rect 9715 3782 9717 3834
rect 9471 3780 9477 3782
rect 9533 3780 9557 3782
rect 9613 3780 9637 3782
rect 9693 3780 9717 3782
rect 9773 3780 9779 3782
rect 9471 3771 9779 3780
rect 9968 3466 9996 4082
rect 10232 4072 10284 4078
rect 10232 4014 10284 4020
rect 10140 4004 10192 4010
rect 10140 3946 10192 3952
rect 10152 3602 10180 3946
rect 10140 3596 10192 3602
rect 10140 3538 10192 3544
rect 10244 3534 10272 4014
rect 10336 4010 10364 4490
rect 10416 4276 10468 4282
rect 10416 4218 10468 4224
rect 10324 4004 10376 4010
rect 10324 3946 10376 3952
rect 10324 3664 10376 3670
rect 10324 3606 10376 3612
rect 10232 3528 10284 3534
rect 10232 3470 10284 3476
rect 9956 3460 10008 3466
rect 9956 3402 10008 3408
rect 10336 3058 10364 3606
rect 10428 3126 10456 4218
rect 10612 3534 10640 4694
rect 10704 3602 10732 5188
rect 10784 5170 10836 5176
rect 10888 5030 10916 6258
rect 10980 5710 11008 9454
rect 11164 8022 11192 9540
rect 11242 9480 11298 9489
rect 11242 9415 11298 9424
rect 11256 9178 11284 9415
rect 11244 9172 11296 9178
rect 11244 9114 11296 9120
rect 11428 8968 11480 8974
rect 11426 8936 11428 8945
rect 11480 8936 11482 8945
rect 11426 8871 11482 8880
rect 11532 8022 11560 9998
rect 11612 9716 11664 9722
rect 11612 9658 11664 9664
rect 11624 9586 11652 9658
rect 11612 9580 11664 9586
rect 11612 9522 11664 9528
rect 11624 8566 11652 9522
rect 11612 8560 11664 8566
rect 11612 8502 11664 8508
rect 11152 8016 11204 8022
rect 11520 8016 11572 8022
rect 11204 7976 11284 8004
rect 11152 7958 11204 7964
rect 11256 7478 11284 7976
rect 11520 7958 11572 7964
rect 11244 7472 11296 7478
rect 11244 7414 11296 7420
rect 11152 7404 11204 7410
rect 11152 7346 11204 7352
rect 11164 7002 11192 7346
rect 11152 6996 11204 7002
rect 11152 6938 11204 6944
rect 11244 6860 11296 6866
rect 11244 6802 11296 6808
rect 11060 6724 11112 6730
rect 11060 6666 11112 6672
rect 11072 6254 11100 6666
rect 11060 6248 11112 6254
rect 11060 6190 11112 6196
rect 10968 5704 11020 5710
rect 10968 5646 11020 5652
rect 10876 5024 10928 5030
rect 10876 4966 10928 4972
rect 10888 4622 10916 4966
rect 10876 4616 10928 4622
rect 10876 4558 10928 4564
rect 10888 4146 10916 4558
rect 10876 4140 10928 4146
rect 10876 4082 10928 4088
rect 10888 3738 10916 4082
rect 10876 3732 10928 3738
rect 10876 3674 10928 3680
rect 10692 3596 10744 3602
rect 10692 3538 10744 3544
rect 10600 3528 10652 3534
rect 10600 3470 10652 3476
rect 10416 3120 10468 3126
rect 10416 3062 10468 3068
rect 10980 3058 11008 5646
rect 11072 4758 11100 6190
rect 11256 5914 11284 6802
rect 11428 6656 11480 6662
rect 11428 6598 11480 6604
rect 11244 5908 11296 5914
rect 11244 5850 11296 5856
rect 11256 5098 11284 5850
rect 11440 5710 11468 6598
rect 11532 5914 11560 7958
rect 11716 7818 11744 10066
rect 11796 10056 11848 10062
rect 11796 9998 11848 10004
rect 11808 7886 11836 9998
rect 11992 9518 12020 12406
rect 12072 12378 12124 12384
rect 12072 12232 12124 12238
rect 12070 12200 12072 12209
rect 12124 12200 12126 12209
rect 12070 12135 12126 12144
rect 12072 12096 12124 12102
rect 12072 12038 12124 12044
rect 11980 9512 12032 9518
rect 12084 9489 12112 12038
rect 12176 11762 12204 13330
rect 12452 13326 12480 13670
rect 13004 13462 13032 13738
rect 12992 13456 13044 13462
rect 12992 13398 13044 13404
rect 12440 13320 12492 13326
rect 12440 13262 12492 13268
rect 12311 13084 12619 13093
rect 12311 13082 12317 13084
rect 12373 13082 12397 13084
rect 12453 13082 12477 13084
rect 12533 13082 12557 13084
rect 12613 13082 12619 13084
rect 12373 13030 12375 13082
rect 12555 13030 12557 13082
rect 12311 13028 12317 13030
rect 12373 13028 12397 13030
rect 12453 13028 12477 13030
rect 12533 13028 12557 13030
rect 12613 13028 12619 13030
rect 12311 13019 12619 13028
rect 12898 12472 12954 12481
rect 12716 12436 12768 12442
rect 12898 12407 12954 12416
rect 12716 12378 12768 12384
rect 12728 12238 12756 12378
rect 12912 12238 12940 12407
rect 13096 12238 13124 14350
rect 13360 13932 13412 13938
rect 13360 13874 13412 13880
rect 13372 13326 13400 13874
rect 13360 13320 13412 13326
rect 13360 13262 13412 13268
rect 13372 12714 13400 13262
rect 13360 12708 13412 12714
rect 13360 12650 13412 12656
rect 12716 12232 12768 12238
rect 12716 12174 12768 12180
rect 12900 12232 12952 12238
rect 12900 12174 12952 12180
rect 13084 12232 13136 12238
rect 13136 12192 13216 12220
rect 13084 12174 13136 12180
rect 12311 11996 12619 12005
rect 12311 11994 12317 11996
rect 12373 11994 12397 11996
rect 12453 11994 12477 11996
rect 12533 11994 12557 11996
rect 12613 11994 12619 11996
rect 12373 11942 12375 11994
rect 12555 11942 12557 11994
rect 12311 11940 12317 11942
rect 12373 11940 12397 11942
rect 12453 11940 12477 11942
rect 12533 11940 12557 11942
rect 12613 11940 12619 11942
rect 12311 11931 12619 11940
rect 12164 11756 12216 11762
rect 12164 11698 12216 11704
rect 12176 9674 12204 11698
rect 12728 11082 12756 12174
rect 12808 12096 12860 12102
rect 12808 12038 12860 12044
rect 12716 11076 12768 11082
rect 12716 11018 12768 11024
rect 12311 10908 12619 10917
rect 12311 10906 12317 10908
rect 12373 10906 12397 10908
rect 12453 10906 12477 10908
rect 12533 10906 12557 10908
rect 12613 10906 12619 10908
rect 12373 10854 12375 10906
rect 12555 10854 12557 10906
rect 12311 10852 12317 10854
rect 12373 10852 12397 10854
rect 12453 10852 12477 10854
rect 12533 10852 12557 10854
rect 12613 10852 12619 10854
rect 12311 10843 12619 10852
rect 12820 10674 12848 12038
rect 12900 11756 12952 11762
rect 12900 11698 12952 11704
rect 12808 10668 12860 10674
rect 12808 10610 12860 10616
rect 12348 10464 12400 10470
rect 12912 10418 12940 11698
rect 13084 11552 13136 11558
rect 13084 11494 13136 11500
rect 13096 11354 13124 11494
rect 13084 11348 13136 11354
rect 13084 11290 13136 11296
rect 13188 11150 13216 12192
rect 13268 11824 13320 11830
rect 13268 11766 13320 11772
rect 13176 11144 13228 11150
rect 13176 11086 13228 11092
rect 12992 11076 13044 11082
rect 12992 11018 13044 11024
rect 13084 11076 13136 11082
rect 13084 11018 13136 11024
rect 12348 10406 12400 10412
rect 12360 10266 12388 10406
rect 12544 10390 12940 10418
rect 12348 10260 12400 10266
rect 12348 10202 12400 10208
rect 12544 10198 12572 10390
rect 12716 10260 12768 10266
rect 12716 10202 12768 10208
rect 12532 10192 12584 10198
rect 12532 10134 12584 10140
rect 12622 10160 12678 10169
rect 12622 10095 12624 10104
rect 12676 10095 12678 10104
rect 12624 10066 12676 10072
rect 12532 10056 12584 10062
rect 12532 9998 12584 10004
rect 12544 9926 12572 9998
rect 12532 9920 12584 9926
rect 12532 9862 12584 9868
rect 12311 9820 12619 9829
rect 12311 9818 12317 9820
rect 12373 9818 12397 9820
rect 12453 9818 12477 9820
rect 12533 9818 12557 9820
rect 12613 9818 12619 9820
rect 12373 9766 12375 9818
rect 12555 9766 12557 9818
rect 12311 9764 12317 9766
rect 12373 9764 12397 9766
rect 12453 9764 12477 9766
rect 12533 9764 12557 9766
rect 12613 9764 12619 9766
rect 12311 9755 12619 9764
rect 12624 9716 12676 9722
rect 12176 9646 12296 9674
rect 11980 9454 12032 9460
rect 12070 9480 12126 9489
rect 12070 9415 12126 9424
rect 11888 9376 11940 9382
rect 11888 9318 11940 9324
rect 11980 9376 12032 9382
rect 11980 9318 12032 9324
rect 11900 9110 11928 9318
rect 11992 9178 12020 9318
rect 11980 9172 12032 9178
rect 11980 9114 12032 9120
rect 11888 9104 11940 9110
rect 11888 9046 11940 9052
rect 12084 8566 12112 9415
rect 12164 8968 12216 8974
rect 12164 8910 12216 8916
rect 12176 8634 12204 8910
rect 12268 8838 12296 9646
rect 12544 9664 12624 9674
rect 12544 9658 12676 9664
rect 12544 9646 12664 9658
rect 12438 9616 12494 9625
rect 12438 9551 12440 9560
rect 12492 9551 12494 9560
rect 12440 9522 12492 9528
rect 12256 8832 12308 8838
rect 12544 8820 12572 9646
rect 12728 9568 12756 10202
rect 12912 10130 12940 10390
rect 12900 10124 12952 10130
rect 12900 10066 12952 10072
rect 12808 9920 12860 9926
rect 12808 9862 12860 9868
rect 12898 9888 12954 9897
rect 12636 9540 12756 9568
rect 12636 9042 12664 9540
rect 12624 9036 12676 9042
rect 12624 8978 12676 8984
rect 12820 8838 12848 9862
rect 12898 9823 12954 9832
rect 12808 8832 12860 8838
rect 12544 8792 12756 8820
rect 12256 8774 12308 8780
rect 12311 8732 12619 8741
rect 12311 8730 12317 8732
rect 12373 8730 12397 8732
rect 12453 8730 12477 8732
rect 12533 8730 12557 8732
rect 12613 8730 12619 8732
rect 12373 8678 12375 8730
rect 12555 8678 12557 8730
rect 12311 8676 12317 8678
rect 12373 8676 12397 8678
rect 12453 8676 12477 8678
rect 12533 8676 12557 8678
rect 12613 8676 12619 8678
rect 12311 8667 12619 8676
rect 12164 8628 12216 8634
rect 12164 8570 12216 8576
rect 11888 8560 11940 8566
rect 11886 8528 11888 8537
rect 12072 8560 12124 8566
rect 11940 8528 11942 8537
rect 12072 8502 12124 8508
rect 12532 8560 12584 8566
rect 12728 8548 12756 8792
rect 12808 8774 12860 8780
rect 12584 8520 12756 8548
rect 12532 8502 12584 8508
rect 11886 8463 11942 8472
rect 11796 7880 11848 7886
rect 11796 7822 11848 7828
rect 11888 7880 11940 7886
rect 11888 7822 11940 7828
rect 11704 7812 11756 7818
rect 11704 7754 11756 7760
rect 11716 7546 11744 7754
rect 11704 7540 11756 7546
rect 11704 7482 11756 7488
rect 11704 6792 11756 6798
rect 11704 6734 11756 6740
rect 11716 6390 11744 6734
rect 11808 6458 11836 7822
rect 11796 6452 11848 6458
rect 11796 6394 11848 6400
rect 11704 6384 11756 6390
rect 11624 6344 11704 6372
rect 11520 5908 11572 5914
rect 11520 5850 11572 5856
rect 11428 5704 11480 5710
rect 11428 5646 11480 5652
rect 11336 5296 11388 5302
rect 11336 5238 11388 5244
rect 11244 5092 11296 5098
rect 11244 5034 11296 5040
rect 11060 4752 11112 4758
rect 11060 4694 11112 4700
rect 11072 3738 11100 4694
rect 11256 4078 11284 5034
rect 11348 4554 11376 5238
rect 11520 5160 11572 5166
rect 11520 5102 11572 5108
rect 11532 4826 11560 5102
rect 11520 4820 11572 4826
rect 11520 4762 11572 4768
rect 11336 4548 11388 4554
rect 11336 4490 11388 4496
rect 11348 4214 11376 4490
rect 11336 4208 11388 4214
rect 11336 4150 11388 4156
rect 11520 4140 11572 4146
rect 11520 4082 11572 4088
rect 11244 4072 11296 4078
rect 11244 4014 11296 4020
rect 11428 4072 11480 4078
rect 11428 4014 11480 4020
rect 11336 3936 11388 3942
rect 11336 3878 11388 3884
rect 11060 3732 11112 3738
rect 11060 3674 11112 3680
rect 9312 3052 9364 3058
rect 9312 2994 9364 3000
rect 10324 3052 10376 3058
rect 10324 2994 10376 3000
rect 10968 3052 11020 3058
rect 10968 2994 11020 3000
rect 9864 2916 9916 2922
rect 9864 2858 9916 2864
rect 9471 2748 9779 2757
rect 9471 2746 9477 2748
rect 9533 2746 9557 2748
rect 9613 2746 9637 2748
rect 9693 2746 9717 2748
rect 9773 2746 9779 2748
rect 9533 2694 9535 2746
rect 9715 2694 9717 2746
rect 9471 2692 9477 2694
rect 9533 2692 9557 2694
rect 9613 2692 9637 2694
rect 9693 2692 9717 2694
rect 9773 2692 9779 2694
rect 9471 2683 9779 2692
rect 9876 800 9904 2858
rect 11348 2854 11376 3878
rect 11440 3534 11468 4014
rect 11532 3942 11560 4082
rect 11520 3936 11572 3942
rect 11520 3878 11572 3884
rect 11624 3602 11652 6344
rect 11704 6326 11756 6332
rect 11900 6186 11928 7822
rect 11980 7472 12032 7478
rect 11980 7414 12032 7420
rect 11992 6934 12020 7414
rect 12084 7274 12112 8502
rect 12728 8294 12756 8520
rect 12912 8498 12940 9823
rect 13004 9722 13032 11018
rect 13096 10810 13124 11018
rect 13176 11008 13228 11014
rect 13176 10950 13228 10956
rect 13084 10804 13136 10810
rect 13084 10746 13136 10752
rect 12992 9716 13044 9722
rect 12992 9658 13044 9664
rect 12992 9580 13044 9586
rect 12992 9522 13044 9528
rect 13004 8634 13032 9522
rect 12992 8628 13044 8634
rect 12992 8570 13044 8576
rect 13096 8514 13124 10746
rect 13188 10266 13216 10950
rect 13176 10260 13228 10266
rect 13176 10202 13228 10208
rect 13176 9716 13228 9722
rect 13176 9658 13228 9664
rect 12900 8492 12952 8498
rect 12900 8434 12952 8440
rect 13004 8486 13124 8514
rect 12716 8288 12768 8294
rect 12716 8230 12768 8236
rect 12164 7948 12216 7954
rect 12164 7890 12216 7896
rect 12176 7410 12204 7890
rect 12311 7644 12619 7653
rect 12311 7642 12317 7644
rect 12373 7642 12397 7644
rect 12453 7642 12477 7644
rect 12533 7642 12557 7644
rect 12613 7642 12619 7644
rect 12373 7590 12375 7642
rect 12555 7590 12557 7642
rect 12311 7588 12317 7590
rect 12373 7588 12397 7590
rect 12453 7588 12477 7590
rect 12533 7588 12557 7590
rect 12613 7588 12619 7590
rect 12311 7579 12619 7588
rect 12164 7404 12216 7410
rect 12164 7346 12216 7352
rect 12728 7342 12756 8230
rect 12912 7954 12940 8434
rect 12900 7948 12952 7954
rect 12900 7890 12952 7896
rect 13004 7546 13032 8486
rect 13084 8424 13136 8430
rect 13084 8366 13136 8372
rect 13096 7721 13124 8366
rect 13188 8362 13216 9658
rect 13280 9110 13308 11766
rect 13372 9722 13400 12650
rect 13452 11620 13504 11626
rect 13452 11562 13504 11568
rect 13464 10112 13492 11562
rect 13556 10810 13584 14606
rect 13648 13734 13676 15506
rect 13912 15496 13964 15502
rect 13912 15438 13964 15444
rect 13820 15020 13872 15026
rect 13820 14962 13872 14968
rect 13832 14618 13860 14962
rect 13820 14612 13872 14618
rect 13820 14554 13872 14560
rect 13820 14272 13872 14278
rect 13820 14214 13872 14220
rect 13832 14074 13860 14214
rect 13820 14068 13872 14074
rect 13820 14010 13872 14016
rect 13636 13728 13688 13734
rect 13636 13670 13688 13676
rect 13648 12374 13676 13670
rect 13820 12776 13872 12782
rect 13820 12718 13872 12724
rect 13636 12368 13688 12374
rect 13636 12310 13688 12316
rect 13648 11762 13676 12310
rect 13832 12306 13860 12718
rect 13820 12300 13872 12306
rect 13820 12242 13872 12248
rect 13924 11898 13952 15438
rect 14016 13870 14044 17274
rect 15152 16892 15460 16901
rect 15152 16890 15158 16892
rect 15214 16890 15238 16892
rect 15294 16890 15318 16892
rect 15374 16890 15398 16892
rect 15454 16890 15460 16892
rect 15214 16838 15216 16890
rect 15396 16838 15398 16890
rect 15152 16836 15158 16838
rect 15214 16836 15238 16838
rect 15294 16836 15318 16838
rect 15374 16836 15398 16838
rect 15454 16836 15460 16838
rect 15152 16827 15460 16836
rect 14188 15904 14240 15910
rect 14188 15846 14240 15852
rect 14200 15570 14228 15846
rect 15152 15804 15460 15813
rect 15152 15802 15158 15804
rect 15214 15802 15238 15804
rect 15294 15802 15318 15804
rect 15374 15802 15398 15804
rect 15454 15802 15460 15804
rect 15214 15750 15216 15802
rect 15396 15750 15398 15802
rect 15152 15748 15158 15750
rect 15214 15748 15238 15750
rect 15294 15748 15318 15750
rect 15374 15748 15398 15750
rect 15454 15748 15460 15750
rect 15152 15739 15460 15748
rect 14188 15564 14240 15570
rect 14188 15506 14240 15512
rect 14556 15496 14608 15502
rect 14556 15438 14608 15444
rect 15292 15496 15344 15502
rect 15292 15438 15344 15444
rect 14568 15162 14596 15438
rect 15304 15162 15332 15438
rect 14556 15156 14608 15162
rect 14556 15098 14608 15104
rect 15292 15156 15344 15162
rect 15292 15098 15344 15104
rect 14096 15088 14148 15094
rect 14096 15030 14148 15036
rect 15476 15088 15528 15094
rect 15476 15030 15528 15036
rect 14004 13864 14056 13870
rect 14004 13806 14056 13812
rect 14016 13462 14044 13806
rect 14004 13456 14056 13462
rect 14004 13398 14056 13404
rect 14108 12730 14136 15030
rect 14280 15020 14332 15026
rect 14280 14962 14332 14968
rect 14188 14884 14240 14890
rect 14188 14826 14240 14832
rect 14016 12702 14136 12730
rect 13912 11892 13964 11898
rect 13912 11834 13964 11840
rect 13636 11756 13688 11762
rect 13636 11698 13688 11704
rect 14016 11558 14044 12702
rect 14096 11824 14148 11830
rect 14096 11766 14148 11772
rect 14004 11552 14056 11558
rect 14004 11494 14056 11500
rect 13820 11212 13872 11218
rect 13820 11154 13872 11160
rect 13636 11076 13688 11082
rect 13636 11018 13688 11024
rect 13544 10804 13596 10810
rect 13544 10746 13596 10752
rect 13648 10266 13676 11018
rect 13728 10736 13780 10742
rect 13728 10678 13780 10684
rect 13636 10260 13688 10266
rect 13636 10202 13688 10208
rect 13648 10130 13676 10202
rect 13544 10124 13596 10130
rect 13464 10084 13544 10112
rect 13360 9716 13412 9722
rect 13360 9658 13412 9664
rect 13360 9376 13412 9382
rect 13360 9318 13412 9324
rect 13268 9104 13320 9110
rect 13268 9046 13320 9052
rect 13176 8356 13228 8362
rect 13176 8298 13228 8304
rect 13082 7712 13138 7721
rect 13082 7647 13138 7656
rect 12992 7540 13044 7546
rect 12992 7482 13044 7488
rect 12900 7404 12952 7410
rect 12900 7346 12952 7352
rect 12716 7336 12768 7342
rect 12716 7278 12768 7284
rect 12072 7268 12124 7274
rect 12072 7210 12124 7216
rect 11980 6928 12032 6934
rect 11980 6870 12032 6876
rect 12311 6556 12619 6565
rect 12311 6554 12317 6556
rect 12373 6554 12397 6556
rect 12453 6554 12477 6556
rect 12533 6554 12557 6556
rect 12613 6554 12619 6556
rect 12373 6502 12375 6554
rect 12555 6502 12557 6554
rect 12311 6500 12317 6502
rect 12373 6500 12397 6502
rect 12453 6500 12477 6502
rect 12533 6500 12557 6502
rect 12613 6500 12619 6502
rect 12311 6491 12619 6500
rect 12912 6390 12940 7346
rect 13004 7002 13032 7482
rect 12992 6996 13044 7002
rect 12992 6938 13044 6944
rect 13096 6882 13124 7647
rect 13004 6854 13124 6882
rect 12900 6384 12952 6390
rect 12900 6326 12952 6332
rect 12440 6316 12492 6322
rect 12440 6258 12492 6264
rect 11888 6180 11940 6186
rect 11888 6122 11940 6128
rect 11900 5642 11928 6122
rect 12452 5642 12480 6258
rect 12900 6180 12952 6186
rect 12900 6122 12952 6128
rect 12808 6112 12860 6118
rect 12808 6054 12860 6060
rect 12820 5914 12848 6054
rect 12912 5914 12940 6122
rect 12808 5908 12860 5914
rect 12808 5850 12860 5856
rect 12900 5908 12952 5914
rect 12900 5850 12952 5856
rect 13004 5846 13032 6854
rect 13188 6798 13216 8298
rect 13372 8090 13400 9318
rect 13360 8084 13412 8090
rect 13360 8026 13412 8032
rect 13464 7886 13492 10084
rect 13544 10066 13596 10072
rect 13636 10124 13688 10130
rect 13636 10066 13688 10072
rect 13648 9926 13676 10066
rect 13636 9920 13688 9926
rect 13636 9862 13688 9868
rect 13648 9674 13676 9862
rect 13556 9646 13676 9674
rect 13556 9586 13584 9646
rect 13544 9580 13596 9586
rect 13544 9522 13596 9528
rect 13556 8974 13584 9522
rect 13544 8968 13596 8974
rect 13544 8910 13596 8916
rect 13634 8664 13690 8673
rect 13634 8599 13690 8608
rect 13648 8498 13676 8599
rect 13636 8492 13688 8498
rect 13636 8434 13688 8440
rect 13544 8288 13596 8294
rect 13544 8230 13596 8236
rect 13360 7880 13412 7886
rect 13360 7822 13412 7828
rect 13452 7880 13504 7886
rect 13452 7822 13504 7828
rect 13372 7478 13400 7822
rect 13556 7478 13584 8230
rect 13360 7472 13412 7478
rect 13360 7414 13412 7420
rect 13544 7472 13596 7478
rect 13544 7414 13596 7420
rect 13648 7274 13676 8434
rect 13740 7410 13768 10678
rect 13832 10470 13860 11154
rect 14108 10826 14136 11766
rect 14016 10798 14136 10826
rect 13912 10600 13964 10606
rect 13912 10542 13964 10548
rect 13820 10464 13872 10470
rect 13820 10406 13872 10412
rect 13820 9988 13872 9994
rect 13820 9930 13872 9936
rect 13728 7404 13780 7410
rect 13728 7346 13780 7352
rect 13636 7268 13688 7274
rect 13636 7210 13688 7216
rect 13832 6866 13860 9930
rect 13924 9722 13952 10542
rect 14016 10062 14044 10798
rect 14096 10464 14148 10470
rect 14096 10406 14148 10412
rect 14004 10056 14056 10062
rect 14004 9998 14056 10004
rect 13912 9716 13964 9722
rect 13912 9658 13964 9664
rect 13912 9376 13964 9382
rect 13912 9318 13964 9324
rect 13924 9110 13952 9318
rect 13912 9104 13964 9110
rect 13912 9046 13964 9052
rect 13912 8968 13964 8974
rect 13912 8910 13964 8916
rect 13924 8537 13952 8910
rect 14016 8673 14044 9998
rect 14002 8664 14058 8673
rect 14002 8599 14058 8608
rect 13910 8528 13966 8537
rect 13910 8463 13966 8472
rect 13924 6866 13952 8463
rect 14108 7750 14136 10406
rect 14200 9178 14228 14826
rect 14292 12238 14320 14962
rect 14556 14884 14608 14890
rect 14556 14826 14608 14832
rect 14372 14816 14424 14822
rect 14372 14758 14424 14764
rect 14384 14414 14412 14758
rect 14372 14408 14424 14414
rect 14372 14350 14424 14356
rect 14464 14408 14516 14414
rect 14464 14350 14516 14356
rect 14384 13530 14412 14350
rect 14476 14074 14504 14350
rect 14464 14068 14516 14074
rect 14464 14010 14516 14016
rect 14568 13938 14596 14826
rect 15152 14716 15460 14725
rect 15152 14714 15158 14716
rect 15214 14714 15238 14716
rect 15294 14714 15318 14716
rect 15374 14714 15398 14716
rect 15454 14714 15460 14716
rect 15214 14662 15216 14714
rect 15396 14662 15398 14714
rect 15152 14660 15158 14662
rect 15214 14660 15238 14662
rect 15294 14660 15318 14662
rect 15374 14660 15398 14662
rect 15454 14660 15460 14662
rect 15152 14651 15460 14660
rect 14740 14408 14792 14414
rect 14740 14350 14792 14356
rect 14752 14006 14780 14350
rect 15384 14340 15436 14346
rect 15384 14282 15436 14288
rect 15292 14272 15344 14278
rect 15292 14214 15344 14220
rect 15304 14074 15332 14214
rect 15292 14068 15344 14074
rect 15292 14010 15344 14016
rect 14740 14000 14792 14006
rect 14740 13942 14792 13948
rect 14556 13932 14608 13938
rect 14556 13874 14608 13880
rect 14372 13524 14424 13530
rect 14372 13466 14424 13472
rect 14568 12918 14596 13874
rect 15396 13870 15424 14282
rect 15384 13864 15436 13870
rect 15382 13832 15384 13841
rect 15436 13832 15438 13841
rect 15382 13767 15438 13776
rect 15152 13628 15460 13637
rect 15152 13626 15158 13628
rect 15214 13626 15238 13628
rect 15294 13626 15318 13628
rect 15374 13626 15398 13628
rect 15454 13626 15460 13628
rect 15214 13574 15216 13626
rect 15396 13574 15398 13626
rect 15152 13572 15158 13574
rect 15214 13572 15238 13574
rect 15294 13572 15318 13574
rect 15374 13572 15398 13574
rect 15454 13572 15460 13574
rect 15152 13563 15460 13572
rect 15488 13530 15516 15030
rect 15844 14884 15896 14890
rect 15844 14826 15896 14832
rect 15856 14618 15884 14826
rect 15844 14612 15896 14618
rect 15844 14554 15896 14560
rect 15936 14612 15988 14618
rect 15936 14554 15988 14560
rect 15948 14498 15976 14554
rect 15568 14476 15620 14482
rect 15568 14418 15620 14424
rect 15856 14470 15976 14498
rect 15476 13524 15528 13530
rect 15476 13466 15528 13472
rect 14924 13456 14976 13462
rect 14924 13398 14976 13404
rect 14556 12912 14608 12918
rect 14608 12872 14688 12900
rect 14556 12854 14608 12860
rect 14554 12336 14610 12345
rect 14554 12271 14610 12280
rect 14568 12238 14596 12271
rect 14280 12232 14332 12238
rect 14280 12174 14332 12180
rect 14556 12232 14608 12238
rect 14556 12174 14608 12180
rect 14660 12073 14688 12872
rect 14832 12640 14884 12646
rect 14832 12582 14884 12588
rect 14844 12306 14872 12582
rect 14832 12300 14884 12306
rect 14832 12242 14884 12248
rect 14646 12064 14702 12073
rect 14646 11999 14702 12008
rect 14372 11756 14424 11762
rect 14372 11698 14424 11704
rect 14556 11756 14608 11762
rect 14556 11698 14608 11704
rect 14280 11688 14332 11694
rect 14280 11630 14332 11636
rect 14292 10062 14320 11630
rect 14384 11354 14412 11698
rect 14372 11348 14424 11354
rect 14372 11290 14424 11296
rect 14568 11218 14596 11698
rect 14832 11688 14884 11694
rect 14830 11656 14832 11665
rect 14884 11656 14886 11665
rect 14830 11591 14886 11600
rect 14832 11348 14884 11354
rect 14832 11290 14884 11296
rect 14738 11248 14794 11257
rect 14556 11212 14608 11218
rect 14738 11183 14794 11192
rect 14556 11154 14608 11160
rect 14464 11144 14516 11150
rect 14752 11098 14780 11183
rect 14844 11150 14872 11290
rect 14832 11144 14884 11150
rect 14516 11092 14780 11098
rect 14464 11086 14780 11092
rect 14476 11070 14780 11086
rect 14372 10804 14424 10810
rect 14372 10746 14424 10752
rect 14280 10056 14332 10062
rect 14280 9998 14332 10004
rect 14188 9172 14240 9178
rect 14188 9114 14240 9120
rect 14292 8537 14320 9998
rect 14384 9625 14412 10746
rect 14648 10668 14700 10674
rect 14648 10610 14700 10616
rect 14556 10464 14608 10470
rect 14556 10406 14608 10412
rect 14462 9888 14518 9897
rect 14462 9823 14518 9832
rect 14370 9616 14426 9625
rect 14370 9551 14426 9560
rect 14278 8528 14334 8537
rect 14278 8463 14334 8472
rect 14384 7818 14412 9551
rect 14476 9489 14504 9823
rect 14568 9654 14596 10406
rect 14660 10266 14688 10610
rect 14648 10260 14700 10266
rect 14648 10202 14700 10208
rect 14752 9674 14780 11070
rect 14830 11112 14832 11121
rect 14884 11112 14886 11121
rect 14830 11047 14886 11056
rect 14556 9648 14608 9654
rect 14556 9590 14608 9596
rect 14660 9646 14780 9674
rect 14462 9480 14518 9489
rect 14462 9415 14518 9424
rect 14568 9160 14596 9590
rect 14660 9586 14688 9646
rect 14648 9580 14700 9586
rect 14648 9522 14700 9528
rect 14660 9450 14688 9522
rect 14648 9444 14700 9450
rect 14648 9386 14700 9392
rect 14740 9376 14792 9382
rect 14740 9318 14792 9324
rect 14568 9132 14688 9160
rect 14554 9072 14610 9081
rect 14464 9036 14516 9042
rect 14554 9007 14610 9016
rect 14464 8978 14516 8984
rect 14476 8634 14504 8978
rect 14568 8974 14596 9007
rect 14556 8968 14608 8974
rect 14556 8910 14608 8916
rect 14660 8934 14688 9132
rect 14752 9042 14780 9318
rect 14830 9208 14886 9217
rect 14936 9178 14964 13398
rect 15580 12850 15608 14418
rect 15660 14408 15712 14414
rect 15660 14350 15712 14356
rect 15672 14278 15700 14350
rect 15856 14346 15884 14470
rect 15936 14408 15988 14414
rect 15936 14350 15988 14356
rect 15844 14340 15896 14346
rect 15844 14282 15896 14288
rect 15660 14272 15712 14278
rect 15660 14214 15712 14220
rect 15752 13932 15804 13938
rect 15752 13874 15804 13880
rect 15660 13728 15712 13734
rect 15660 13670 15712 13676
rect 15672 12986 15700 13670
rect 15764 13462 15792 13874
rect 15752 13456 15804 13462
rect 15752 13398 15804 13404
rect 15660 12980 15712 12986
rect 15660 12922 15712 12928
rect 15292 12844 15344 12850
rect 15028 12804 15292 12832
rect 15028 12481 15056 12804
rect 15292 12786 15344 12792
rect 15568 12844 15620 12850
rect 15568 12786 15620 12792
rect 15672 12782 15700 12922
rect 15764 12918 15792 13398
rect 15856 13326 15884 14282
rect 15844 13320 15896 13326
rect 15844 13262 15896 13268
rect 15752 12912 15804 12918
rect 15752 12854 15804 12860
rect 15660 12776 15712 12782
rect 15660 12718 15712 12724
rect 15752 12640 15804 12646
rect 15752 12582 15804 12588
rect 15152 12540 15460 12549
rect 15152 12538 15158 12540
rect 15214 12538 15238 12540
rect 15294 12538 15318 12540
rect 15374 12538 15398 12540
rect 15454 12538 15460 12540
rect 15214 12486 15216 12538
rect 15396 12486 15398 12538
rect 15152 12484 15158 12486
rect 15214 12484 15238 12486
rect 15294 12484 15318 12486
rect 15374 12484 15398 12486
rect 15454 12484 15460 12486
rect 15014 12472 15070 12481
rect 15152 12475 15460 12484
rect 15014 12407 15070 12416
rect 15028 11626 15056 12407
rect 15568 12232 15620 12238
rect 15660 12232 15712 12238
rect 15568 12174 15620 12180
rect 15658 12200 15660 12209
rect 15712 12200 15714 12209
rect 15384 12096 15436 12102
rect 15384 12038 15436 12044
rect 15396 11762 15424 12038
rect 15476 11892 15528 11898
rect 15476 11834 15528 11840
rect 15384 11756 15436 11762
rect 15384 11698 15436 11704
rect 15016 11620 15068 11626
rect 15016 11562 15068 11568
rect 15028 10470 15056 11562
rect 15152 11452 15460 11461
rect 15152 11450 15158 11452
rect 15214 11450 15238 11452
rect 15294 11450 15318 11452
rect 15374 11450 15398 11452
rect 15454 11450 15460 11452
rect 15214 11398 15216 11450
rect 15396 11398 15398 11450
rect 15152 11396 15158 11398
rect 15214 11396 15238 11398
rect 15294 11396 15318 11398
rect 15374 11396 15398 11398
rect 15454 11396 15460 11398
rect 15152 11387 15460 11396
rect 15488 11234 15516 11834
rect 15580 11762 15608 12174
rect 15658 12135 15714 12144
rect 15568 11756 15620 11762
rect 15620 11716 15700 11744
rect 15568 11698 15620 11704
rect 15488 11206 15608 11234
rect 15476 11144 15528 11150
rect 15476 11086 15528 11092
rect 15290 10840 15346 10849
rect 15290 10775 15346 10784
rect 15304 10742 15332 10775
rect 15292 10736 15344 10742
rect 15292 10678 15344 10684
rect 15016 10464 15068 10470
rect 15016 10406 15068 10412
rect 15152 10364 15460 10373
rect 15152 10362 15158 10364
rect 15214 10362 15238 10364
rect 15294 10362 15318 10364
rect 15374 10362 15398 10364
rect 15454 10362 15460 10364
rect 15214 10310 15216 10362
rect 15396 10310 15398 10362
rect 15152 10308 15158 10310
rect 15214 10308 15238 10310
rect 15294 10308 15318 10310
rect 15374 10308 15398 10310
rect 15454 10308 15460 10310
rect 15152 10299 15460 10308
rect 15290 10024 15346 10033
rect 15290 9959 15292 9968
rect 15344 9959 15346 9968
rect 15292 9930 15344 9936
rect 15384 9580 15436 9586
rect 15384 9522 15436 9528
rect 15396 9489 15424 9522
rect 15382 9480 15438 9489
rect 15382 9415 15438 9424
rect 15152 9276 15460 9285
rect 15152 9274 15158 9276
rect 15214 9274 15238 9276
rect 15294 9274 15318 9276
rect 15374 9274 15398 9276
rect 15454 9274 15460 9276
rect 15214 9222 15216 9274
rect 15396 9222 15398 9274
rect 15152 9220 15158 9222
rect 15214 9220 15238 9222
rect 15294 9220 15318 9222
rect 15374 9220 15398 9222
rect 15454 9220 15460 9222
rect 15152 9211 15460 9220
rect 14830 9143 14886 9152
rect 14924 9172 14976 9178
rect 14740 9036 14792 9042
rect 14740 8978 14792 8984
rect 14660 8906 14780 8934
rect 14844 8906 14872 9143
rect 14976 9132 15056 9160
rect 14924 9114 14976 9120
rect 14648 8832 14700 8838
rect 14648 8774 14700 8780
rect 14464 8628 14516 8634
rect 14464 8570 14516 8576
rect 14462 8528 14518 8537
rect 14462 8463 14464 8472
rect 14516 8463 14518 8472
rect 14464 8434 14516 8440
rect 14556 8424 14608 8430
rect 14556 8366 14608 8372
rect 14568 7970 14596 8366
rect 14660 8090 14688 8774
rect 14752 8294 14780 8906
rect 14832 8900 14884 8906
rect 14832 8842 14884 8848
rect 14832 8424 14884 8430
rect 14832 8366 14884 8372
rect 14740 8288 14792 8294
rect 14740 8230 14792 8236
rect 14648 8084 14700 8090
rect 14648 8026 14700 8032
rect 14568 7954 14688 7970
rect 14556 7948 14688 7954
rect 14608 7942 14688 7948
rect 14556 7890 14608 7896
rect 14568 7859 14596 7890
rect 14372 7812 14424 7818
rect 14372 7754 14424 7760
rect 14004 7744 14056 7750
rect 14004 7686 14056 7692
rect 14096 7744 14148 7750
rect 14096 7686 14148 7692
rect 14016 7546 14044 7686
rect 14004 7540 14056 7546
rect 14004 7482 14056 7488
rect 14660 7449 14688 7942
rect 14740 7812 14792 7818
rect 14740 7754 14792 7760
rect 14646 7440 14702 7449
rect 14188 7404 14240 7410
rect 14188 7346 14240 7352
rect 14372 7404 14424 7410
rect 14372 7346 14424 7352
rect 14556 7404 14608 7410
rect 14752 7410 14780 7754
rect 14646 7375 14702 7384
rect 14740 7404 14792 7410
rect 14556 7346 14608 7352
rect 14740 7346 14792 7352
rect 14200 7206 14228 7346
rect 14188 7200 14240 7206
rect 14188 7142 14240 7148
rect 13544 6860 13596 6866
rect 13544 6802 13596 6808
rect 13820 6860 13872 6866
rect 13820 6802 13872 6808
rect 13912 6860 13964 6866
rect 13912 6802 13964 6808
rect 13084 6792 13136 6798
rect 13084 6734 13136 6740
rect 13176 6792 13228 6798
rect 13176 6734 13228 6740
rect 13096 6254 13124 6734
rect 13084 6248 13136 6254
rect 13084 6190 13136 6196
rect 12992 5840 13044 5846
rect 12992 5782 13044 5788
rect 13096 5778 13124 6190
rect 13084 5772 13136 5778
rect 13084 5714 13136 5720
rect 11888 5636 11940 5642
rect 11888 5578 11940 5584
rect 12440 5636 12492 5642
rect 12440 5578 12492 5584
rect 11900 5370 11928 5578
rect 13188 5574 13216 6734
rect 13556 6254 13584 6802
rect 14200 6798 14228 7142
rect 14188 6792 14240 6798
rect 14188 6734 14240 6740
rect 14384 6662 14412 7346
rect 14372 6656 14424 6662
rect 14372 6598 14424 6604
rect 13910 6488 13966 6497
rect 13910 6423 13966 6432
rect 13924 6390 13952 6423
rect 13912 6384 13964 6390
rect 13912 6326 13964 6332
rect 13544 6248 13596 6254
rect 13544 6190 13596 6196
rect 13636 6248 13688 6254
rect 13636 6190 13688 6196
rect 13452 6112 13504 6118
rect 13452 6054 13504 6060
rect 13360 5908 13412 5914
rect 13464 5896 13492 6054
rect 13412 5868 13492 5896
rect 13360 5850 13412 5856
rect 13176 5568 13228 5574
rect 13176 5510 13228 5516
rect 12311 5468 12619 5477
rect 12311 5466 12317 5468
rect 12373 5466 12397 5468
rect 12453 5466 12477 5468
rect 12533 5466 12557 5468
rect 12613 5466 12619 5468
rect 12373 5414 12375 5466
rect 12555 5414 12557 5466
rect 12311 5412 12317 5414
rect 12373 5412 12397 5414
rect 12453 5412 12477 5414
rect 12533 5412 12557 5414
rect 12613 5412 12619 5414
rect 12311 5403 12619 5412
rect 11888 5364 11940 5370
rect 11888 5306 11940 5312
rect 11796 5228 11848 5234
rect 11796 5170 11848 5176
rect 11808 4078 11836 5170
rect 11900 4758 11928 5306
rect 12256 5296 12308 5302
rect 12256 5238 12308 5244
rect 11980 5228 12032 5234
rect 12032 5188 12204 5216
rect 11980 5170 12032 5176
rect 11888 4752 11940 4758
rect 11888 4694 11940 4700
rect 11888 4616 11940 4622
rect 11886 4584 11888 4593
rect 11940 4584 11942 4593
rect 11886 4519 11942 4528
rect 11888 4480 11940 4486
rect 11888 4422 11940 4428
rect 11900 4146 11928 4422
rect 11888 4140 11940 4146
rect 11888 4082 11940 4088
rect 11796 4072 11848 4078
rect 11796 4014 11848 4020
rect 11900 3890 11928 4082
rect 11716 3862 11928 3890
rect 11612 3596 11664 3602
rect 11612 3538 11664 3544
rect 11428 3528 11480 3534
rect 11428 3470 11480 3476
rect 11520 3528 11572 3534
rect 11520 3470 11572 3476
rect 11532 3194 11560 3470
rect 11520 3188 11572 3194
rect 11520 3130 11572 3136
rect 11336 2848 11388 2854
rect 11336 2790 11388 2796
rect 11152 2576 11204 2582
rect 11152 2518 11204 2524
rect 10508 2372 10560 2378
rect 10508 2314 10560 2320
rect 10520 800 10548 2314
rect 11164 800 11192 2518
rect 11624 2446 11652 3538
rect 11716 3126 11744 3862
rect 11900 3738 11928 3862
rect 11796 3732 11848 3738
rect 11796 3674 11848 3680
rect 11888 3732 11940 3738
rect 11888 3674 11940 3680
rect 11808 3194 11836 3674
rect 11888 3528 11940 3534
rect 11888 3470 11940 3476
rect 11796 3188 11848 3194
rect 11796 3130 11848 3136
rect 11704 3120 11756 3126
rect 11704 3062 11756 3068
rect 11900 2446 11928 3470
rect 11992 3398 12020 5170
rect 12072 4684 12124 4690
rect 12072 4626 12124 4632
rect 11980 3392 12032 3398
rect 11980 3334 12032 3340
rect 11992 2650 12020 3334
rect 12084 3194 12112 4626
rect 12176 4604 12204 5188
rect 12268 4826 12296 5238
rect 12716 5228 12768 5234
rect 12716 5170 12768 5176
rect 12348 5092 12400 5098
rect 12348 5034 12400 5040
rect 12360 4826 12388 5034
rect 12256 4820 12308 4826
rect 12256 4762 12308 4768
rect 12348 4820 12400 4826
rect 12348 4762 12400 4768
rect 12728 4690 12756 5170
rect 13188 5098 13216 5510
rect 13360 5296 13412 5302
rect 13360 5238 13412 5244
rect 13372 5166 13400 5238
rect 13360 5160 13412 5166
rect 13360 5102 13412 5108
rect 13176 5092 13228 5098
rect 13176 5034 13228 5040
rect 12716 4684 12768 4690
rect 12716 4626 12768 4632
rect 12256 4616 12308 4622
rect 12176 4576 12256 4604
rect 12256 4558 12308 4564
rect 12714 4584 12770 4593
rect 12714 4519 12770 4528
rect 12311 4380 12619 4389
rect 12311 4378 12317 4380
rect 12373 4378 12397 4380
rect 12453 4378 12477 4380
rect 12533 4378 12557 4380
rect 12613 4378 12619 4380
rect 12373 4326 12375 4378
rect 12555 4326 12557 4378
rect 12311 4324 12317 4326
rect 12373 4324 12397 4326
rect 12453 4324 12477 4326
rect 12533 4324 12557 4326
rect 12613 4324 12619 4326
rect 12311 4315 12619 4324
rect 12440 4208 12492 4214
rect 12440 4150 12492 4156
rect 12164 4004 12216 4010
rect 12164 3946 12216 3952
rect 12072 3188 12124 3194
rect 12072 3130 12124 3136
rect 12176 3126 12204 3946
rect 12256 3936 12308 3942
rect 12256 3878 12308 3884
rect 12268 3602 12296 3878
rect 12348 3732 12400 3738
rect 12452 3720 12480 4150
rect 12728 3738 12756 4519
rect 13464 4010 13492 5868
rect 13556 4146 13584 6190
rect 13648 5710 13676 6190
rect 13912 5908 13964 5914
rect 13912 5850 13964 5856
rect 13636 5704 13688 5710
rect 13636 5646 13688 5652
rect 13820 5704 13872 5710
rect 13820 5646 13872 5652
rect 13648 5370 13676 5646
rect 13636 5364 13688 5370
rect 13636 5306 13688 5312
rect 13648 5030 13676 5306
rect 13832 5234 13860 5646
rect 13924 5234 13952 5850
rect 13820 5228 13872 5234
rect 13820 5170 13872 5176
rect 13912 5228 13964 5234
rect 13912 5170 13964 5176
rect 13636 5024 13688 5030
rect 13636 4966 13688 4972
rect 13544 4140 13596 4146
rect 13544 4082 13596 4088
rect 13452 4004 13504 4010
rect 13452 3946 13504 3952
rect 13556 3738 13584 4082
rect 13648 4078 13676 4966
rect 13832 4690 13860 5170
rect 13820 4684 13872 4690
rect 13820 4626 13872 4632
rect 13924 4622 13952 5170
rect 13912 4616 13964 4622
rect 13912 4558 13964 4564
rect 14568 4486 14596 7346
rect 14648 6112 14700 6118
rect 14648 6054 14700 6060
rect 14660 5642 14688 6054
rect 14648 5636 14700 5642
rect 14648 5578 14700 5584
rect 14660 5030 14688 5578
rect 14752 5302 14780 7346
rect 14844 6202 14872 8366
rect 14924 8356 14976 8362
rect 14924 8298 14976 8304
rect 14936 7886 14964 8298
rect 14924 7880 14976 7886
rect 14924 7822 14976 7828
rect 14924 7744 14976 7750
rect 14924 7686 14976 7692
rect 14936 7002 14964 7686
rect 15028 7342 15056 9132
rect 15488 8430 15516 11086
rect 15580 11014 15608 11206
rect 15568 11008 15620 11014
rect 15568 10950 15620 10956
rect 15568 10736 15620 10742
rect 15568 10678 15620 10684
rect 15580 10062 15608 10678
rect 15568 10056 15620 10062
rect 15568 9998 15620 10004
rect 15672 9994 15700 11716
rect 15764 11150 15792 12582
rect 15948 12442 15976 14350
rect 15936 12436 15988 12442
rect 15936 12378 15988 12384
rect 16040 12186 16068 17478
rect 17992 17436 18300 17445
rect 17992 17434 17998 17436
rect 18054 17434 18078 17436
rect 18134 17434 18158 17436
rect 18214 17434 18238 17436
rect 18294 17434 18300 17436
rect 18054 17382 18056 17434
rect 18236 17382 18238 17434
rect 17992 17380 17998 17382
rect 18054 17380 18078 17382
rect 18134 17380 18158 17382
rect 18214 17380 18238 17382
rect 18294 17380 18300 17382
rect 17992 17371 18300 17380
rect 16580 16584 16632 16590
rect 16580 16526 16632 16532
rect 16592 15706 16620 16526
rect 17992 16348 18300 16357
rect 17992 16346 17998 16348
rect 18054 16346 18078 16348
rect 18134 16346 18158 16348
rect 18214 16346 18238 16348
rect 18294 16346 18300 16348
rect 18054 16294 18056 16346
rect 18236 16294 18238 16346
rect 17992 16292 17998 16294
rect 18054 16292 18078 16294
rect 18134 16292 18158 16294
rect 18214 16292 18238 16294
rect 18294 16292 18300 16294
rect 17992 16283 18300 16292
rect 16580 15700 16632 15706
rect 16580 15642 16632 15648
rect 16948 15360 17000 15366
rect 16948 15302 17000 15308
rect 17040 15360 17092 15366
rect 17040 15302 17092 15308
rect 16764 15088 16816 15094
rect 16762 15056 16764 15065
rect 16816 15056 16818 15065
rect 16212 15020 16264 15026
rect 16212 14962 16264 14968
rect 16580 15020 16632 15026
rect 16762 14991 16818 15000
rect 16580 14962 16632 14968
rect 16120 14544 16172 14550
rect 16120 14486 16172 14492
rect 15856 12158 16068 12186
rect 15752 11144 15804 11150
rect 15752 11086 15804 11092
rect 15752 11008 15804 11014
rect 15752 10950 15804 10956
rect 15660 9988 15712 9994
rect 15660 9930 15712 9936
rect 15568 9716 15620 9722
rect 15568 9658 15620 9664
rect 15476 8424 15528 8430
rect 15476 8366 15528 8372
rect 15152 8188 15460 8197
rect 15152 8186 15158 8188
rect 15214 8186 15238 8188
rect 15294 8186 15318 8188
rect 15374 8186 15398 8188
rect 15454 8186 15460 8188
rect 15214 8134 15216 8186
rect 15396 8134 15398 8186
rect 15152 8132 15158 8134
rect 15214 8132 15238 8134
rect 15294 8132 15318 8134
rect 15374 8132 15398 8134
rect 15454 8132 15460 8134
rect 15152 8123 15460 8132
rect 15108 7948 15160 7954
rect 15108 7890 15160 7896
rect 15120 7342 15148 7890
rect 15384 7812 15436 7818
rect 15384 7754 15436 7760
rect 15396 7478 15424 7754
rect 15488 7546 15516 8366
rect 15476 7540 15528 7546
rect 15476 7482 15528 7488
rect 15384 7472 15436 7478
rect 15384 7414 15436 7420
rect 15016 7336 15068 7342
rect 15016 7278 15068 7284
rect 15108 7336 15160 7342
rect 15108 7278 15160 7284
rect 14924 6996 14976 7002
rect 14924 6938 14976 6944
rect 14844 6186 14964 6202
rect 14844 6180 14976 6186
rect 14844 6174 14924 6180
rect 14844 5914 14872 6174
rect 14924 6122 14976 6128
rect 14832 5908 14884 5914
rect 14832 5850 14884 5856
rect 15028 5778 15056 7278
rect 15152 7100 15460 7109
rect 15152 7098 15158 7100
rect 15214 7098 15238 7100
rect 15294 7098 15318 7100
rect 15374 7098 15398 7100
rect 15454 7098 15460 7100
rect 15214 7046 15216 7098
rect 15396 7046 15398 7098
rect 15152 7044 15158 7046
rect 15214 7044 15238 7046
rect 15294 7044 15318 7046
rect 15374 7044 15398 7046
rect 15454 7044 15460 7046
rect 15152 7035 15460 7044
rect 15488 7002 15516 7482
rect 15580 7324 15608 9658
rect 15672 7818 15700 9930
rect 15764 9722 15792 10950
rect 15856 10674 15884 12158
rect 15934 12064 15990 12073
rect 15934 11999 15990 12008
rect 15844 10668 15896 10674
rect 15844 10610 15896 10616
rect 15856 10538 15884 10610
rect 15844 10532 15896 10538
rect 15844 10474 15896 10480
rect 15752 9716 15804 9722
rect 15752 9658 15804 9664
rect 15752 9444 15804 9450
rect 15752 9386 15804 9392
rect 15764 9178 15792 9386
rect 15752 9172 15804 9178
rect 15752 9114 15804 9120
rect 15752 8492 15804 8498
rect 15752 8434 15804 8440
rect 15764 8090 15792 8434
rect 15752 8084 15804 8090
rect 15752 8026 15804 8032
rect 15660 7812 15712 7818
rect 15660 7754 15712 7760
rect 15856 7392 15884 10474
rect 15948 9518 15976 11999
rect 16132 11778 16160 14486
rect 16224 14414 16252 14962
rect 16592 14618 16620 14962
rect 16580 14612 16632 14618
rect 16580 14554 16632 14560
rect 16672 14612 16724 14618
rect 16672 14554 16724 14560
rect 16684 14414 16712 14554
rect 16212 14408 16264 14414
rect 16212 14350 16264 14356
rect 16672 14408 16724 14414
rect 16672 14350 16724 14356
rect 16212 14272 16264 14278
rect 16212 14214 16264 14220
rect 16672 14272 16724 14278
rect 16672 14214 16724 14220
rect 16224 13734 16252 14214
rect 16684 14074 16712 14214
rect 16672 14068 16724 14074
rect 16672 14010 16724 14016
rect 16960 14006 16988 15302
rect 17052 14890 17080 15302
rect 17992 15260 18300 15269
rect 17992 15258 17998 15260
rect 18054 15258 18078 15260
rect 18134 15258 18158 15260
rect 18214 15258 18238 15260
rect 18294 15258 18300 15260
rect 18054 15206 18056 15258
rect 18236 15206 18238 15258
rect 17992 15204 17998 15206
rect 18054 15204 18078 15206
rect 18134 15204 18158 15206
rect 18214 15204 18238 15206
rect 18294 15204 18300 15206
rect 17992 15195 18300 15204
rect 17132 15020 17184 15026
rect 17132 14962 17184 14968
rect 17040 14884 17092 14890
rect 17040 14826 17092 14832
rect 17040 14408 17092 14414
rect 17040 14350 17092 14356
rect 17052 14074 17080 14350
rect 17040 14068 17092 14074
rect 17040 14010 17092 14016
rect 16764 14000 16816 14006
rect 16764 13942 16816 13948
rect 16948 14000 17000 14006
rect 16948 13942 17000 13948
rect 16304 13864 16356 13870
rect 16304 13806 16356 13812
rect 16212 13728 16264 13734
rect 16212 13670 16264 13676
rect 16212 13184 16264 13190
rect 16212 13126 16264 13132
rect 16224 11898 16252 13126
rect 16316 11898 16344 13806
rect 16776 13530 16804 13942
rect 16764 13524 16816 13530
rect 16764 13466 16816 13472
rect 16776 13326 16804 13466
rect 16764 13320 16816 13326
rect 16764 13262 16816 13268
rect 16488 12980 16540 12986
rect 16488 12922 16540 12928
rect 16396 12640 16448 12646
rect 16396 12582 16448 12588
rect 16408 12102 16436 12582
rect 16396 12096 16448 12102
rect 16396 12038 16448 12044
rect 16212 11892 16264 11898
rect 16212 11834 16264 11840
rect 16304 11892 16356 11898
rect 16304 11834 16356 11840
rect 16132 11750 16252 11778
rect 16028 11620 16080 11626
rect 16028 11562 16080 11568
rect 16040 11257 16068 11562
rect 16026 11248 16082 11257
rect 16026 11183 16082 11192
rect 16120 11212 16172 11218
rect 16224 11200 16252 11750
rect 16172 11172 16252 11200
rect 16120 11154 16172 11160
rect 16028 11144 16080 11150
rect 16028 11086 16080 11092
rect 15936 9512 15988 9518
rect 15936 9454 15988 9460
rect 15948 7886 15976 9454
rect 16040 8634 16068 11086
rect 16132 10810 16160 11154
rect 16408 11150 16436 12038
rect 16500 11354 16528 12922
rect 16580 12436 16632 12442
rect 16580 12378 16632 12384
rect 16488 11348 16540 11354
rect 16488 11290 16540 11296
rect 16396 11144 16448 11150
rect 16224 11104 16396 11132
rect 16120 10804 16172 10810
rect 16120 10746 16172 10752
rect 16120 10668 16172 10674
rect 16224 10656 16252 11104
rect 16396 11086 16448 11092
rect 16488 11008 16540 11014
rect 16488 10950 16540 10956
rect 16394 10840 16450 10849
rect 16394 10775 16450 10784
rect 16172 10628 16252 10656
rect 16120 10610 16172 10616
rect 16120 10124 16172 10130
rect 16120 10066 16172 10072
rect 16132 9722 16160 10066
rect 16120 9716 16172 9722
rect 16120 9658 16172 9664
rect 16132 9548 16160 9658
rect 16120 9542 16172 9548
rect 16120 9484 16172 9490
rect 16224 9330 16252 10628
rect 16408 10130 16436 10775
rect 16500 10169 16528 10950
rect 16486 10160 16542 10169
rect 16396 10124 16448 10130
rect 16486 10095 16542 10104
rect 16396 10066 16448 10072
rect 16486 10024 16542 10033
rect 16486 9959 16488 9968
rect 16540 9959 16542 9968
rect 16488 9930 16540 9936
rect 16486 9616 16542 9625
rect 16486 9551 16542 9560
rect 16500 9518 16528 9551
rect 16488 9512 16540 9518
rect 16488 9454 16540 9460
rect 16592 9450 16620 12378
rect 16672 12368 16724 12374
rect 16672 12310 16724 12316
rect 16684 11558 16712 12310
rect 16672 11552 16724 11558
rect 16672 11494 16724 11500
rect 16672 11076 16724 11082
rect 16672 11018 16724 11024
rect 16684 10606 16712 11018
rect 16672 10600 16724 10606
rect 16672 10542 16724 10548
rect 16672 10192 16724 10198
rect 16672 10134 16724 10140
rect 16396 9444 16448 9450
rect 16396 9386 16448 9392
rect 16580 9444 16632 9450
rect 16580 9386 16632 9392
rect 16224 9302 16344 9330
rect 16316 9178 16344 9302
rect 16212 9172 16264 9178
rect 16212 9114 16264 9120
rect 16304 9172 16356 9178
rect 16304 9114 16356 9120
rect 16028 8628 16080 8634
rect 16028 8570 16080 8576
rect 16120 8492 16172 8498
rect 16120 8434 16172 8440
rect 16028 8016 16080 8022
rect 16028 7958 16080 7964
rect 15936 7880 15988 7886
rect 15936 7822 15988 7828
rect 15764 7364 15884 7392
rect 15660 7336 15712 7342
rect 15580 7296 15660 7324
rect 15660 7278 15712 7284
rect 15476 6996 15528 7002
rect 15476 6938 15528 6944
rect 15476 6316 15528 6322
rect 15476 6258 15528 6264
rect 15152 6012 15460 6021
rect 15152 6010 15158 6012
rect 15214 6010 15238 6012
rect 15294 6010 15318 6012
rect 15374 6010 15398 6012
rect 15454 6010 15460 6012
rect 15214 5958 15216 6010
rect 15396 5958 15398 6010
rect 15152 5956 15158 5958
rect 15214 5956 15238 5958
rect 15294 5956 15318 5958
rect 15374 5956 15398 5958
rect 15454 5956 15460 5958
rect 15152 5947 15460 5956
rect 15016 5772 15068 5778
rect 15016 5714 15068 5720
rect 15488 5370 15516 6258
rect 15476 5364 15528 5370
rect 15476 5306 15528 5312
rect 14740 5296 14792 5302
rect 14740 5238 14792 5244
rect 15568 5296 15620 5302
rect 15568 5238 15620 5244
rect 15580 5030 15608 5238
rect 14648 5024 14700 5030
rect 14648 4966 14700 4972
rect 15568 5024 15620 5030
rect 15568 4966 15620 4972
rect 15152 4924 15460 4933
rect 15152 4922 15158 4924
rect 15214 4922 15238 4924
rect 15294 4922 15318 4924
rect 15374 4922 15398 4924
rect 15454 4922 15460 4924
rect 15214 4870 15216 4922
rect 15396 4870 15398 4922
rect 15152 4868 15158 4870
rect 15214 4868 15238 4870
rect 15294 4868 15318 4870
rect 15374 4868 15398 4870
rect 15454 4868 15460 4870
rect 15152 4859 15460 4868
rect 15568 4820 15620 4826
rect 15672 4808 15700 7278
rect 15764 6390 15792 7364
rect 15844 7268 15896 7274
rect 15844 7210 15896 7216
rect 15856 6390 15884 7210
rect 15948 7206 15976 7822
rect 15936 7200 15988 7206
rect 15936 7142 15988 7148
rect 15936 6928 15988 6934
rect 16040 6905 16068 7958
rect 15936 6870 15988 6876
rect 16026 6896 16082 6905
rect 15948 6730 15976 6870
rect 16026 6831 16082 6840
rect 15936 6724 15988 6730
rect 15936 6666 15988 6672
rect 15752 6384 15804 6390
rect 15752 6326 15804 6332
rect 15844 6384 15896 6390
rect 15844 6326 15896 6332
rect 15620 4780 15700 4808
rect 15568 4762 15620 4768
rect 14924 4684 14976 4690
rect 14924 4626 14976 4632
rect 14936 4593 14964 4626
rect 14922 4584 14978 4593
rect 14922 4519 14978 4528
rect 15016 4548 15068 4554
rect 15016 4490 15068 4496
rect 15200 4548 15252 4554
rect 15200 4490 15252 4496
rect 14556 4480 14608 4486
rect 14556 4422 14608 4428
rect 13636 4072 13688 4078
rect 13636 4014 13688 4020
rect 12400 3692 12480 3720
rect 12716 3732 12768 3738
rect 12348 3674 12400 3680
rect 12716 3674 12768 3680
rect 13544 3732 13596 3738
rect 13544 3674 13596 3680
rect 12256 3596 12308 3602
rect 12256 3538 12308 3544
rect 12360 3534 12388 3674
rect 15028 3670 15056 4490
rect 15212 4282 15240 4490
rect 15200 4276 15252 4282
rect 15200 4218 15252 4224
rect 15764 4146 15792 6326
rect 16132 6322 16160 8434
rect 16224 7924 16252 9114
rect 16316 8294 16344 9114
rect 16304 8288 16356 8294
rect 16304 8230 16356 8236
rect 16212 7918 16264 7924
rect 16212 7860 16264 7866
rect 16304 7880 16356 7886
rect 16304 7822 16356 7828
rect 16212 7812 16264 7818
rect 16212 7754 16264 7760
rect 16224 6458 16252 7754
rect 16316 7721 16344 7822
rect 16302 7712 16358 7721
rect 16302 7647 16358 7656
rect 16408 7342 16436 9386
rect 16486 9208 16542 9217
rect 16486 9143 16542 9152
rect 16500 9110 16528 9143
rect 16488 9104 16540 9110
rect 16488 9046 16540 9052
rect 16684 9042 16712 10134
rect 16776 10062 16804 13262
rect 17040 13184 17092 13190
rect 17040 13126 17092 13132
rect 17052 12850 17080 13126
rect 17040 12844 17092 12850
rect 17040 12786 17092 12792
rect 17144 12782 17172 14962
rect 18328 14816 18380 14822
rect 18328 14758 18380 14764
rect 17992 14172 18300 14181
rect 17992 14170 17998 14172
rect 18054 14170 18078 14172
rect 18134 14170 18158 14172
rect 18214 14170 18238 14172
rect 18294 14170 18300 14172
rect 18054 14118 18056 14170
rect 18236 14118 18238 14170
rect 17992 14116 17998 14118
rect 18054 14116 18078 14118
rect 18134 14116 18158 14118
rect 18214 14116 18238 14118
rect 18294 14116 18300 14118
rect 17992 14107 18300 14116
rect 18340 14006 18368 14758
rect 18432 14618 18460 18702
rect 23673 18524 23981 18533
rect 23673 18522 23679 18524
rect 23735 18522 23759 18524
rect 23815 18522 23839 18524
rect 23895 18522 23919 18524
rect 23975 18522 23981 18524
rect 23735 18470 23737 18522
rect 23917 18470 23919 18522
rect 23673 18468 23679 18470
rect 23735 18468 23759 18470
rect 23815 18468 23839 18470
rect 23895 18468 23919 18470
rect 23975 18468 23981 18470
rect 23673 18459 23981 18468
rect 20833 17980 21141 17989
rect 20833 17978 20839 17980
rect 20895 17978 20919 17980
rect 20975 17978 20999 17980
rect 21055 17978 21079 17980
rect 21135 17978 21141 17980
rect 20895 17926 20897 17978
rect 21077 17926 21079 17978
rect 20833 17924 20839 17926
rect 20895 17924 20919 17926
rect 20975 17924 20999 17926
rect 21055 17924 21079 17926
rect 21135 17924 21141 17926
rect 20833 17915 21141 17924
rect 23673 17436 23981 17445
rect 23673 17434 23679 17436
rect 23735 17434 23759 17436
rect 23815 17434 23839 17436
rect 23895 17434 23919 17436
rect 23975 17434 23981 17436
rect 23735 17382 23737 17434
rect 23917 17382 23919 17434
rect 23673 17380 23679 17382
rect 23735 17380 23759 17382
rect 23815 17380 23839 17382
rect 23895 17380 23919 17382
rect 23975 17380 23981 17382
rect 23673 17371 23981 17380
rect 20833 16892 21141 16901
rect 20833 16890 20839 16892
rect 20895 16890 20919 16892
rect 20975 16890 20999 16892
rect 21055 16890 21079 16892
rect 21135 16890 21141 16892
rect 20895 16838 20897 16890
rect 21077 16838 21079 16890
rect 20833 16836 20839 16838
rect 20895 16836 20919 16838
rect 20975 16836 20999 16838
rect 21055 16836 21079 16838
rect 21135 16836 21141 16838
rect 20833 16827 21141 16836
rect 23673 16348 23981 16357
rect 23673 16346 23679 16348
rect 23735 16346 23759 16348
rect 23815 16346 23839 16348
rect 23895 16346 23919 16348
rect 23975 16346 23981 16348
rect 23735 16294 23737 16346
rect 23917 16294 23919 16346
rect 23673 16292 23679 16294
rect 23735 16292 23759 16294
rect 23815 16292 23839 16294
rect 23895 16292 23919 16294
rect 23975 16292 23981 16294
rect 23673 16283 23981 16292
rect 20833 15804 21141 15813
rect 20833 15802 20839 15804
rect 20895 15802 20919 15804
rect 20975 15802 20999 15804
rect 21055 15802 21079 15804
rect 21135 15802 21141 15804
rect 20895 15750 20897 15802
rect 21077 15750 21079 15802
rect 20833 15748 20839 15750
rect 20895 15748 20919 15750
rect 20975 15748 20999 15750
rect 21055 15748 21079 15750
rect 21135 15748 21141 15750
rect 20833 15739 21141 15748
rect 19064 15428 19116 15434
rect 19064 15370 19116 15376
rect 18696 15360 18748 15366
rect 18696 15302 18748 15308
rect 18708 15026 18736 15302
rect 18696 15020 18748 15026
rect 18696 14962 18748 14968
rect 18604 14952 18656 14958
rect 18604 14894 18656 14900
rect 18420 14612 18472 14618
rect 18420 14554 18472 14560
rect 18420 14408 18472 14414
rect 18420 14350 18472 14356
rect 18328 14000 18380 14006
rect 18328 13942 18380 13948
rect 18432 13938 18460 14350
rect 18512 14272 18564 14278
rect 18512 14214 18564 14220
rect 18420 13932 18472 13938
rect 18420 13874 18472 13880
rect 17776 13864 17828 13870
rect 17776 13806 17828 13812
rect 17868 13864 17920 13870
rect 17868 13806 17920 13812
rect 18328 13864 18380 13870
rect 18328 13806 18380 13812
rect 17224 13728 17276 13734
rect 17224 13670 17276 13676
rect 17236 12850 17264 13670
rect 17316 13456 17368 13462
rect 17316 13398 17368 13404
rect 17328 13258 17356 13398
rect 17500 13320 17552 13326
rect 17788 13297 17816 13806
rect 17500 13262 17552 13268
rect 17774 13288 17830 13297
rect 17316 13252 17368 13258
rect 17316 13194 17368 13200
rect 17224 12844 17276 12850
rect 17224 12786 17276 12792
rect 17132 12776 17184 12782
rect 17132 12718 17184 12724
rect 17224 12708 17276 12714
rect 17224 12650 17276 12656
rect 17236 12238 17264 12650
rect 17328 12434 17356 13194
rect 17408 12436 17460 12442
rect 17328 12406 17408 12434
rect 17512 12434 17540 13262
rect 17774 13223 17830 13232
rect 17684 12776 17736 12782
rect 17684 12718 17736 12724
rect 17512 12406 17632 12434
rect 17408 12378 17460 12384
rect 17316 12368 17368 12374
rect 17316 12310 17368 12316
rect 17224 12232 17276 12238
rect 17224 12174 17276 12180
rect 16948 12164 17000 12170
rect 16948 12106 17000 12112
rect 16856 12096 16908 12102
rect 16856 12038 16908 12044
rect 16764 10056 16816 10062
rect 16764 9998 16816 10004
rect 16764 9920 16816 9926
rect 16764 9862 16816 9868
rect 16672 9036 16724 9042
rect 16672 8978 16724 8984
rect 16580 8968 16632 8974
rect 16580 8910 16632 8916
rect 16488 8900 16540 8906
rect 16488 8842 16540 8848
rect 16500 8634 16528 8842
rect 16592 8634 16620 8910
rect 16488 8628 16540 8634
rect 16488 8570 16540 8576
rect 16580 8628 16632 8634
rect 16580 8570 16632 8576
rect 16776 8242 16804 9862
rect 16592 8214 16804 8242
rect 16488 8084 16540 8090
rect 16488 8026 16540 8032
rect 16500 7478 16528 8026
rect 16488 7472 16540 7478
rect 16488 7414 16540 7420
rect 16396 7336 16448 7342
rect 16396 7278 16448 7284
rect 16304 7268 16356 7274
rect 16304 7210 16356 7216
rect 16316 7002 16344 7210
rect 16304 6996 16356 7002
rect 16304 6938 16356 6944
rect 16212 6452 16264 6458
rect 16212 6394 16264 6400
rect 16316 6322 16344 6938
rect 16396 6928 16448 6934
rect 16592 6916 16620 8214
rect 16868 8106 16896 12038
rect 16960 11830 16988 12106
rect 16948 11824 17000 11830
rect 16946 11792 16948 11801
rect 17000 11792 17002 11801
rect 16946 11727 17002 11736
rect 16948 11688 17000 11694
rect 17132 11688 17184 11694
rect 16948 11630 17000 11636
rect 17038 11656 17094 11665
rect 16960 11150 16988 11630
rect 17132 11630 17184 11636
rect 17038 11591 17094 11600
rect 16948 11144 17000 11150
rect 16948 11086 17000 11092
rect 16948 10736 17000 10742
rect 16948 10678 17000 10684
rect 16776 8078 16896 8106
rect 16672 7744 16724 7750
rect 16672 7686 16724 7692
rect 16684 7410 16712 7686
rect 16672 7404 16724 7410
rect 16672 7346 16724 7352
rect 16448 6888 16712 6916
rect 16396 6870 16448 6876
rect 16580 6792 16632 6798
rect 16580 6734 16632 6740
rect 16120 6316 16172 6322
rect 16120 6258 16172 6264
rect 16304 6316 16356 6322
rect 16304 6258 16356 6264
rect 16396 6316 16448 6322
rect 16396 6258 16448 6264
rect 16132 6118 16160 6258
rect 16120 6112 16172 6118
rect 16120 6054 16172 6060
rect 15844 5772 15896 5778
rect 15844 5714 15896 5720
rect 15856 5370 15884 5714
rect 16408 5370 16436 6258
rect 16488 5704 16540 5710
rect 16488 5646 16540 5652
rect 15844 5364 15896 5370
rect 15844 5306 15896 5312
rect 16396 5364 16448 5370
rect 16396 5306 16448 5312
rect 16408 4758 16436 5306
rect 16500 5234 16528 5646
rect 16592 5302 16620 6734
rect 16684 5710 16712 6888
rect 16776 5914 16804 8078
rect 16856 8016 16908 8022
rect 16854 7984 16856 7993
rect 16908 7984 16910 7993
rect 16960 7954 16988 10678
rect 16854 7919 16910 7928
rect 16948 7948 17000 7954
rect 16948 7890 17000 7896
rect 16856 7880 16908 7886
rect 16856 7822 16908 7828
rect 16868 6798 16896 7822
rect 16946 7712 17002 7721
rect 16946 7647 17002 7656
rect 16856 6792 16908 6798
rect 16856 6734 16908 6740
rect 16764 5908 16816 5914
rect 16764 5850 16816 5856
rect 16776 5817 16804 5850
rect 16762 5808 16818 5817
rect 16762 5743 16818 5752
rect 16672 5704 16724 5710
rect 16672 5646 16724 5652
rect 16580 5296 16632 5302
rect 16580 5238 16632 5244
rect 16488 5228 16540 5234
rect 16488 5170 16540 5176
rect 16396 4752 16448 4758
rect 16396 4694 16448 4700
rect 16500 4554 16528 5170
rect 16488 4548 16540 4554
rect 16488 4490 16540 4496
rect 16684 4214 16712 5646
rect 16868 5234 16896 6734
rect 16960 5710 16988 7647
rect 17052 6730 17080 11591
rect 17144 10849 17172 11630
rect 17236 11354 17264 12174
rect 17328 11898 17356 12310
rect 17604 12238 17632 12406
rect 17592 12232 17644 12238
rect 17592 12174 17644 12180
rect 17408 12096 17460 12102
rect 17408 12038 17460 12044
rect 17500 12096 17552 12102
rect 17500 12038 17552 12044
rect 17316 11892 17368 11898
rect 17316 11834 17368 11840
rect 17224 11348 17276 11354
rect 17224 11290 17276 11296
rect 17130 10840 17186 10849
rect 17130 10775 17186 10784
rect 17328 10713 17356 11834
rect 17420 11762 17448 12038
rect 17512 11830 17540 12038
rect 17500 11824 17552 11830
rect 17500 11766 17552 11772
rect 17408 11756 17460 11762
rect 17408 11698 17460 11704
rect 17408 11552 17460 11558
rect 17408 11494 17460 11500
rect 17314 10704 17370 10713
rect 17314 10639 17370 10648
rect 17224 10600 17276 10606
rect 17224 10542 17276 10548
rect 17236 10130 17264 10542
rect 17224 10124 17276 10130
rect 17224 10066 17276 10072
rect 17132 9988 17184 9994
rect 17132 9930 17184 9936
rect 17144 9897 17172 9930
rect 17236 9926 17264 10066
rect 17224 9920 17276 9926
rect 17130 9888 17186 9897
rect 17224 9862 17276 9868
rect 17130 9823 17186 9832
rect 17224 9512 17276 9518
rect 17130 9480 17186 9489
rect 17224 9454 17276 9460
rect 17130 9415 17186 9424
rect 17040 6724 17092 6730
rect 17040 6666 17092 6672
rect 16948 5704 17000 5710
rect 16948 5646 17000 5652
rect 17144 5370 17172 9415
rect 17236 9217 17264 9454
rect 17222 9208 17278 9217
rect 17222 9143 17278 9152
rect 17236 8498 17264 9143
rect 17328 8566 17356 10639
rect 17420 9994 17448 11494
rect 17604 11354 17632 12174
rect 17696 11626 17724 12718
rect 17684 11620 17736 11626
rect 17684 11562 17736 11568
rect 17592 11348 17644 11354
rect 17592 11290 17644 11296
rect 17604 10810 17632 11290
rect 17684 11144 17736 11150
rect 17684 11086 17736 11092
rect 17592 10804 17644 10810
rect 17592 10746 17644 10752
rect 17500 10668 17552 10674
rect 17500 10610 17552 10616
rect 17408 9988 17460 9994
rect 17408 9930 17460 9936
rect 17408 9716 17460 9722
rect 17408 9658 17460 9664
rect 17316 8560 17368 8566
rect 17316 8502 17368 8508
rect 17224 8492 17276 8498
rect 17224 8434 17276 8440
rect 17224 8356 17276 8362
rect 17224 8298 17276 8304
rect 17236 7721 17264 8298
rect 17222 7712 17278 7721
rect 17222 7647 17278 7656
rect 17224 7404 17276 7410
rect 17224 7346 17276 7352
rect 17236 5846 17264 7346
rect 17420 6798 17448 9658
rect 17512 9636 17540 10610
rect 17696 9926 17724 11086
rect 17788 11082 17816 13223
rect 17880 12306 17908 13806
rect 18236 13320 18288 13326
rect 18234 13288 18236 13297
rect 18288 13288 18290 13297
rect 18234 13223 18290 13232
rect 17992 13084 18300 13093
rect 17992 13082 17998 13084
rect 18054 13082 18078 13084
rect 18134 13082 18158 13084
rect 18214 13082 18238 13084
rect 18294 13082 18300 13084
rect 18054 13030 18056 13082
rect 18236 13030 18238 13082
rect 17992 13028 17998 13030
rect 18054 13028 18078 13030
rect 18134 13028 18158 13030
rect 18214 13028 18238 13030
rect 18294 13028 18300 13030
rect 17992 13019 18300 13028
rect 18236 12844 18288 12850
rect 18236 12786 18288 12792
rect 17868 12300 17920 12306
rect 17868 12242 17920 12248
rect 17868 12164 17920 12170
rect 17868 12106 17920 12112
rect 17880 11286 17908 12106
rect 18248 12084 18276 12786
rect 18340 12442 18368 13806
rect 18420 13796 18472 13802
rect 18420 13738 18472 13744
rect 18432 12986 18460 13738
rect 18420 12980 18472 12986
rect 18420 12922 18472 12928
rect 18328 12436 18380 12442
rect 18328 12378 18380 12384
rect 18420 12232 18472 12238
rect 18420 12174 18472 12180
rect 18248 12056 18368 12084
rect 17992 11996 18300 12005
rect 17992 11994 17998 11996
rect 18054 11994 18078 11996
rect 18134 11994 18158 11996
rect 18214 11994 18238 11996
rect 18294 11994 18300 11996
rect 18054 11942 18056 11994
rect 18236 11942 18238 11994
rect 17992 11940 17998 11942
rect 18054 11940 18078 11942
rect 18134 11940 18158 11942
rect 18214 11940 18238 11942
rect 18294 11940 18300 11942
rect 17992 11931 18300 11940
rect 18340 11898 18368 12056
rect 17960 11892 18012 11898
rect 17960 11834 18012 11840
rect 18328 11892 18380 11898
rect 18328 11834 18380 11840
rect 17868 11280 17920 11286
rect 17868 11222 17920 11228
rect 17776 11076 17828 11082
rect 17776 11018 17828 11024
rect 17972 10996 18000 11834
rect 18328 11620 18380 11626
rect 18328 11562 18380 11568
rect 18340 11286 18368 11562
rect 18328 11280 18380 11286
rect 18328 11222 18380 11228
rect 18328 11076 18380 11082
rect 18328 11018 18380 11024
rect 17880 10968 18000 10996
rect 17684 9920 17736 9926
rect 17684 9862 17736 9868
rect 17592 9648 17644 9654
rect 17512 9608 17592 9636
rect 17592 9590 17644 9596
rect 17604 9450 17632 9590
rect 17696 9489 17724 9862
rect 17880 9674 17908 10968
rect 17992 10908 18300 10917
rect 17992 10906 17998 10908
rect 18054 10906 18078 10908
rect 18134 10906 18158 10908
rect 18214 10906 18238 10908
rect 18294 10906 18300 10908
rect 18054 10854 18056 10906
rect 18236 10854 18238 10906
rect 17992 10852 17998 10854
rect 18054 10852 18078 10854
rect 18134 10852 18158 10854
rect 18214 10852 18238 10854
rect 18294 10852 18300 10854
rect 17992 10843 18300 10852
rect 17992 9820 18300 9829
rect 17992 9818 17998 9820
rect 18054 9818 18078 9820
rect 18134 9818 18158 9820
rect 18214 9818 18238 9820
rect 18294 9818 18300 9820
rect 18054 9766 18056 9818
rect 18236 9766 18238 9818
rect 17992 9764 17998 9766
rect 18054 9764 18078 9766
rect 18134 9764 18158 9766
rect 18214 9764 18238 9766
rect 18294 9764 18300 9766
rect 17992 9755 18300 9764
rect 17788 9646 17908 9674
rect 18236 9716 18288 9722
rect 18236 9658 18288 9664
rect 17682 9480 17738 9489
rect 17592 9444 17644 9450
rect 17682 9415 17738 9424
rect 17592 9386 17644 9392
rect 17500 8968 17552 8974
rect 17552 8928 17632 8956
rect 17500 8910 17552 8916
rect 17604 7857 17632 8928
rect 17788 8922 17816 9646
rect 17868 9580 17920 9586
rect 17868 9522 17920 9528
rect 17960 9580 18012 9586
rect 17960 9522 18012 9528
rect 17880 9178 17908 9522
rect 17972 9353 18000 9522
rect 17958 9344 18014 9353
rect 17958 9279 18014 9288
rect 17868 9172 17920 9178
rect 17868 9114 17920 9120
rect 17696 8894 17816 8922
rect 17868 8946 17920 8952
rect 17696 8498 17724 8894
rect 17868 8888 17920 8894
rect 17776 8832 17828 8838
rect 17776 8774 17828 8780
rect 17684 8492 17736 8498
rect 17684 8434 17736 8440
rect 17590 7848 17646 7857
rect 17590 7783 17646 7792
rect 17500 7200 17552 7206
rect 17500 7142 17552 7148
rect 17512 6934 17540 7142
rect 17604 7002 17632 7783
rect 17696 7750 17724 8434
rect 17788 8090 17816 8774
rect 17776 8084 17828 8090
rect 17776 8026 17828 8032
rect 17684 7744 17736 7750
rect 17684 7686 17736 7692
rect 17880 7546 17908 8888
rect 18248 8820 18276 9658
rect 18340 9586 18368 11018
rect 18432 10810 18460 12174
rect 18524 11898 18552 14214
rect 18616 14006 18644 14894
rect 18604 14000 18656 14006
rect 18604 13942 18656 13948
rect 18708 13734 18736 14962
rect 19076 14482 19104 15370
rect 23673 15260 23981 15269
rect 23673 15258 23679 15260
rect 23735 15258 23759 15260
rect 23815 15258 23839 15260
rect 23895 15258 23919 15260
rect 23975 15258 23981 15260
rect 23735 15206 23737 15258
rect 23917 15206 23919 15258
rect 23673 15204 23679 15206
rect 23735 15204 23759 15206
rect 23815 15204 23839 15206
rect 23895 15204 23919 15206
rect 23975 15204 23981 15206
rect 23673 15195 23981 15204
rect 19248 15156 19300 15162
rect 19248 15098 19300 15104
rect 19064 14476 19116 14482
rect 19064 14418 19116 14424
rect 18788 14068 18840 14074
rect 18788 14010 18840 14016
rect 18696 13728 18748 13734
rect 18696 13670 18748 13676
rect 18604 13320 18656 13326
rect 18800 13274 18828 14010
rect 19076 13920 19104 14418
rect 19156 14272 19208 14278
rect 19156 14214 19208 14220
rect 19168 14074 19196 14214
rect 19156 14068 19208 14074
rect 19156 14010 19208 14016
rect 19076 13892 19196 13920
rect 18972 13524 19024 13530
rect 18972 13466 19024 13472
rect 18984 13326 19012 13466
rect 18656 13268 18828 13274
rect 18604 13262 18828 13268
rect 18880 13320 18932 13326
rect 18880 13262 18932 13268
rect 18972 13320 19024 13326
rect 18972 13262 19024 13268
rect 18616 13246 18828 13262
rect 18604 13184 18656 13190
rect 18604 13126 18656 13132
rect 18616 12850 18644 13126
rect 18604 12844 18656 12850
rect 18604 12786 18656 12792
rect 18512 11892 18564 11898
rect 18512 11834 18564 11840
rect 18616 11778 18644 12786
rect 18616 11750 18736 11778
rect 18604 11688 18656 11694
rect 18604 11630 18656 11636
rect 18512 11144 18564 11150
rect 18512 11086 18564 11092
rect 18420 10804 18472 10810
rect 18420 10746 18472 10752
rect 18420 10668 18472 10674
rect 18420 10610 18472 10616
rect 18432 10266 18460 10610
rect 18420 10260 18472 10266
rect 18420 10202 18472 10208
rect 18432 9654 18460 10202
rect 18524 10146 18552 11086
rect 18616 10266 18644 11630
rect 18708 10656 18736 11750
rect 18800 11665 18828 13246
rect 18892 12646 18920 13262
rect 18972 13184 19024 13190
rect 18972 13126 19024 13132
rect 18984 12850 19012 13126
rect 18972 12844 19024 12850
rect 18972 12786 19024 12792
rect 18972 12708 19024 12714
rect 18972 12650 19024 12656
rect 18880 12640 18932 12646
rect 18880 12582 18932 12588
rect 18984 12442 19012 12650
rect 18972 12436 19024 12442
rect 18972 12378 19024 12384
rect 18880 12368 18932 12374
rect 18880 12310 18932 12316
rect 18892 11801 18920 12310
rect 18878 11792 18934 11801
rect 18878 11727 18934 11736
rect 18786 11656 18842 11665
rect 18786 11591 18842 11600
rect 18800 11150 18828 11591
rect 18788 11144 18840 11150
rect 18788 11086 18840 11092
rect 18892 10962 18920 11727
rect 18984 11150 19012 12378
rect 19064 11824 19116 11830
rect 19064 11766 19116 11772
rect 19076 11665 19104 11766
rect 19062 11656 19118 11665
rect 19062 11591 19118 11600
rect 18972 11144 19024 11150
rect 18972 11086 19024 11092
rect 19168 11014 19196 13892
rect 19260 11626 19288 15098
rect 19616 15020 19668 15026
rect 19616 14962 19668 14968
rect 19628 14278 19656 14962
rect 20833 14716 21141 14725
rect 20833 14714 20839 14716
rect 20895 14714 20919 14716
rect 20975 14714 20999 14716
rect 21055 14714 21079 14716
rect 21135 14714 21141 14716
rect 20895 14662 20897 14714
rect 21077 14662 21079 14714
rect 20833 14660 20839 14662
rect 20895 14660 20919 14662
rect 20975 14660 20999 14662
rect 21055 14660 21079 14662
rect 21135 14660 21141 14662
rect 20833 14651 21141 14660
rect 19984 14544 20036 14550
rect 19984 14486 20036 14492
rect 19708 14408 19760 14414
rect 19708 14350 19760 14356
rect 19616 14272 19668 14278
rect 19616 14214 19668 14220
rect 19524 14000 19576 14006
rect 19524 13942 19576 13948
rect 19340 13932 19392 13938
rect 19340 13874 19392 13880
rect 19432 13932 19484 13938
rect 19432 13874 19484 13880
rect 19352 12986 19380 13874
rect 19444 13530 19472 13874
rect 19536 13841 19564 13942
rect 19522 13832 19578 13841
rect 19522 13767 19578 13776
rect 19432 13524 19484 13530
rect 19432 13466 19484 13472
rect 19340 12980 19392 12986
rect 19340 12922 19392 12928
rect 19628 12850 19656 14214
rect 19720 13938 19748 14350
rect 19996 13938 20024 14486
rect 20444 14408 20496 14414
rect 20444 14350 20496 14356
rect 19708 13932 19760 13938
rect 19708 13874 19760 13880
rect 19984 13932 20036 13938
rect 19984 13874 20036 13880
rect 20352 13932 20404 13938
rect 20352 13874 20404 13880
rect 19800 13524 19852 13530
rect 19800 13466 19852 13472
rect 19708 13320 19760 13326
rect 19708 13262 19760 13268
rect 19720 12889 19748 13262
rect 19706 12880 19762 12889
rect 19340 12844 19392 12850
rect 19340 12786 19392 12792
rect 19616 12844 19668 12850
rect 19706 12815 19762 12824
rect 19616 12786 19668 12792
rect 19248 11620 19300 11626
rect 19248 11562 19300 11568
rect 19246 11112 19302 11121
rect 19246 11047 19248 11056
rect 19300 11047 19302 11056
rect 19248 11018 19300 11024
rect 19156 11008 19208 11014
rect 18892 10934 19012 10962
rect 19156 10950 19208 10956
rect 18788 10668 18840 10674
rect 18708 10628 18788 10656
rect 18788 10610 18840 10616
rect 18696 10464 18748 10470
rect 18696 10406 18748 10412
rect 18604 10260 18656 10266
rect 18604 10202 18656 10208
rect 18524 10118 18644 10146
rect 18512 10056 18564 10062
rect 18512 9998 18564 10004
rect 18420 9648 18472 9654
rect 18420 9590 18472 9596
rect 18328 9580 18380 9586
rect 18328 9522 18380 9528
rect 18248 8792 18368 8820
rect 17992 8732 18300 8741
rect 17992 8730 17998 8732
rect 18054 8730 18078 8732
rect 18134 8730 18158 8732
rect 18214 8730 18238 8732
rect 18294 8730 18300 8732
rect 18054 8678 18056 8730
rect 18236 8678 18238 8730
rect 17992 8676 17998 8678
rect 18054 8676 18078 8678
rect 18134 8676 18158 8678
rect 18214 8676 18238 8678
rect 18294 8676 18300 8678
rect 17992 8667 18300 8676
rect 18340 8634 18368 8792
rect 18328 8628 18380 8634
rect 18328 8570 18380 8576
rect 18432 8566 18460 9590
rect 18524 9042 18552 9998
rect 18616 9761 18644 10118
rect 18708 10062 18736 10406
rect 18696 10056 18748 10062
rect 18696 9998 18748 10004
rect 18602 9752 18658 9761
rect 18602 9687 18604 9696
rect 18656 9687 18658 9696
rect 18604 9658 18656 9664
rect 18604 9580 18656 9586
rect 18604 9522 18656 9528
rect 18616 9382 18644 9522
rect 18604 9376 18656 9382
rect 18604 9318 18656 9324
rect 18512 9036 18564 9042
rect 18512 8978 18564 8984
rect 18510 8936 18566 8945
rect 18510 8871 18566 8880
rect 18524 8838 18552 8871
rect 18512 8832 18564 8838
rect 18512 8774 18564 8780
rect 18420 8560 18472 8566
rect 18420 8502 18472 8508
rect 18236 8492 18288 8498
rect 18236 8434 18288 8440
rect 18248 8362 18276 8434
rect 18420 8424 18472 8430
rect 18420 8366 18472 8372
rect 18236 8356 18288 8362
rect 18236 8298 18288 8304
rect 18052 8288 18104 8294
rect 18052 8230 18104 8236
rect 18064 7886 18092 8230
rect 18432 7886 18460 8366
rect 18052 7880 18104 7886
rect 18050 7848 18052 7857
rect 18420 7880 18472 7886
rect 18104 7848 18106 7857
rect 18420 7822 18472 7828
rect 18050 7783 18106 7792
rect 18328 7744 18380 7750
rect 18328 7686 18380 7692
rect 17992 7644 18300 7653
rect 17992 7642 17998 7644
rect 18054 7642 18078 7644
rect 18134 7642 18158 7644
rect 18214 7642 18238 7644
rect 18294 7642 18300 7644
rect 18054 7590 18056 7642
rect 18236 7590 18238 7642
rect 17992 7588 17998 7590
rect 18054 7588 18078 7590
rect 18134 7588 18158 7590
rect 18214 7588 18238 7590
rect 18294 7588 18300 7590
rect 17992 7579 18300 7588
rect 17868 7540 17920 7546
rect 17868 7482 17920 7488
rect 18144 7472 18196 7478
rect 18144 7414 18196 7420
rect 17960 7404 18012 7410
rect 17960 7346 18012 7352
rect 17776 7336 17828 7342
rect 17776 7278 17828 7284
rect 17788 7002 17816 7278
rect 17592 6996 17644 7002
rect 17592 6938 17644 6944
rect 17776 6996 17828 7002
rect 17776 6938 17828 6944
rect 17500 6928 17552 6934
rect 17500 6870 17552 6876
rect 17316 6792 17368 6798
rect 17316 6734 17368 6740
rect 17408 6792 17460 6798
rect 17408 6734 17460 6740
rect 17328 6322 17356 6734
rect 17316 6316 17368 6322
rect 17316 6258 17368 6264
rect 17224 5840 17276 5846
rect 17224 5782 17276 5788
rect 17132 5364 17184 5370
rect 17132 5306 17184 5312
rect 16856 5228 16908 5234
rect 16856 5170 16908 5176
rect 16868 4826 16896 5170
rect 17132 5092 17184 5098
rect 17132 5034 17184 5040
rect 16856 4820 16908 4826
rect 16856 4762 16908 4768
rect 17144 4758 17172 5034
rect 17132 4752 17184 4758
rect 17132 4694 17184 4700
rect 17144 4282 17172 4694
rect 17604 4690 17632 6938
rect 17682 6896 17738 6905
rect 17682 6831 17738 6840
rect 17696 6798 17724 6831
rect 17684 6792 17736 6798
rect 17684 6734 17736 6740
rect 17682 6488 17738 6497
rect 17682 6423 17738 6432
rect 17696 6390 17724 6423
rect 17684 6384 17736 6390
rect 17684 6326 17736 6332
rect 17788 6322 17816 6938
rect 17972 6746 18000 7346
rect 18156 7342 18184 7414
rect 18144 7336 18196 7342
rect 18144 7278 18196 7284
rect 18236 7336 18288 7342
rect 18236 7278 18288 7284
rect 18248 6934 18276 7278
rect 18236 6928 18288 6934
rect 18236 6870 18288 6876
rect 18248 6798 18276 6870
rect 17880 6718 18000 6746
rect 18236 6792 18288 6798
rect 18236 6734 18288 6740
rect 17880 6440 17908 6718
rect 17992 6556 18300 6565
rect 17992 6554 17998 6556
rect 18054 6554 18078 6556
rect 18134 6554 18158 6556
rect 18214 6554 18238 6556
rect 18294 6554 18300 6556
rect 18054 6502 18056 6554
rect 18236 6502 18238 6554
rect 17992 6500 17998 6502
rect 18054 6500 18078 6502
rect 18134 6500 18158 6502
rect 18214 6500 18238 6502
rect 18294 6500 18300 6502
rect 17992 6491 18300 6500
rect 18144 6452 18196 6458
rect 17880 6412 18000 6440
rect 17776 6316 17828 6322
rect 17776 6258 17828 6264
rect 17972 6186 18000 6412
rect 18144 6394 18196 6400
rect 18050 6352 18106 6361
rect 18050 6287 18106 6296
rect 18064 6254 18092 6287
rect 18052 6248 18104 6254
rect 18052 6190 18104 6196
rect 18156 6186 18184 6394
rect 17960 6180 18012 6186
rect 17960 6122 18012 6128
rect 18144 6180 18196 6186
rect 18144 6122 18196 6128
rect 18340 5914 18368 7686
rect 18432 6798 18460 7822
rect 18616 7818 18644 9318
rect 18694 9208 18750 9217
rect 18694 9143 18750 9152
rect 18708 9042 18736 9143
rect 18696 9036 18748 9042
rect 18696 8978 18748 8984
rect 18696 8832 18748 8838
rect 18696 8774 18748 8780
rect 18708 8634 18736 8774
rect 18696 8628 18748 8634
rect 18696 8570 18748 8576
rect 18800 8498 18828 10610
rect 18880 10600 18932 10606
rect 18880 10542 18932 10548
rect 18892 9994 18920 10542
rect 18880 9988 18932 9994
rect 18880 9930 18932 9936
rect 18892 9625 18920 9930
rect 18878 9616 18934 9625
rect 18878 9551 18934 9560
rect 18788 8492 18840 8498
rect 18788 8434 18840 8440
rect 18800 8090 18828 8434
rect 18788 8084 18840 8090
rect 18788 8026 18840 8032
rect 18604 7812 18656 7818
rect 18524 7772 18604 7800
rect 18420 6792 18472 6798
rect 18420 6734 18472 6740
rect 18420 6656 18472 6662
rect 18418 6624 18420 6633
rect 18472 6624 18474 6633
rect 18418 6559 18474 6568
rect 18328 5908 18380 5914
rect 18328 5850 18380 5856
rect 18420 5908 18472 5914
rect 18420 5850 18472 5856
rect 18328 5704 18380 5710
rect 18328 5646 18380 5652
rect 17992 5468 18300 5477
rect 17992 5466 17998 5468
rect 18054 5466 18078 5468
rect 18134 5466 18158 5468
rect 18214 5466 18238 5468
rect 18294 5466 18300 5468
rect 18054 5414 18056 5466
rect 18236 5414 18238 5466
rect 17992 5412 17998 5414
rect 18054 5412 18078 5414
rect 18134 5412 18158 5414
rect 18214 5412 18238 5414
rect 18294 5412 18300 5414
rect 17992 5403 18300 5412
rect 18340 4826 18368 5646
rect 18432 5370 18460 5850
rect 18420 5364 18472 5370
rect 18420 5306 18472 5312
rect 18328 4820 18380 4826
rect 18328 4762 18380 4768
rect 18524 4758 18552 7772
rect 18604 7754 18656 7760
rect 18800 7478 18828 8026
rect 18604 7472 18656 7478
rect 18604 7414 18656 7420
rect 18788 7472 18840 7478
rect 18788 7414 18840 7420
rect 18616 5234 18644 7414
rect 18788 7336 18840 7342
rect 18892 7290 18920 9551
rect 18984 8956 19012 10934
rect 19168 9586 19196 10950
rect 19352 10810 19380 12786
rect 19432 12640 19484 12646
rect 19432 12582 19484 12588
rect 19444 12345 19472 12582
rect 19430 12336 19486 12345
rect 19430 12271 19486 12280
rect 19432 12232 19484 12238
rect 19432 12174 19484 12180
rect 19444 11150 19472 12174
rect 19616 11620 19668 11626
rect 19616 11562 19668 11568
rect 19628 11286 19656 11562
rect 19812 11506 19840 13466
rect 19892 13456 19944 13462
rect 19892 13398 19944 13404
rect 19904 12238 19932 13398
rect 19892 12232 19944 12238
rect 19892 12174 19944 12180
rect 19720 11478 19840 11506
rect 19616 11280 19668 11286
rect 19616 11222 19668 11228
rect 19524 11212 19576 11218
rect 19524 11154 19576 11160
rect 19432 11144 19484 11150
rect 19432 11086 19484 11092
rect 19340 10804 19392 10810
rect 19340 10746 19392 10752
rect 19432 10736 19484 10742
rect 19432 10678 19484 10684
rect 19340 10668 19392 10674
rect 19340 10610 19392 10616
rect 19352 10130 19380 10610
rect 19444 10470 19472 10678
rect 19432 10464 19484 10470
rect 19432 10406 19484 10412
rect 19340 10124 19392 10130
rect 19340 10066 19392 10072
rect 19156 9580 19208 9586
rect 19156 9522 19208 9528
rect 19248 9512 19300 9518
rect 19248 9454 19300 9460
rect 19260 9382 19288 9454
rect 19352 9450 19380 10066
rect 19432 9920 19484 9926
rect 19432 9862 19484 9868
rect 19444 9722 19472 9862
rect 19432 9716 19484 9722
rect 19432 9658 19484 9664
rect 19340 9444 19392 9450
rect 19340 9386 19392 9392
rect 19248 9376 19300 9382
rect 19248 9318 19300 9324
rect 18984 8928 19104 8956
rect 18972 8832 19024 8838
rect 18972 8774 19024 8780
rect 18984 8430 19012 8774
rect 18972 8424 19024 8430
rect 19076 8401 19104 8928
rect 19352 8838 19380 9386
rect 19340 8832 19392 8838
rect 19340 8774 19392 8780
rect 18972 8366 19024 8372
rect 19062 8392 19118 8401
rect 19062 8327 19118 8336
rect 18970 7440 19026 7449
rect 18970 7375 18972 7384
rect 19024 7375 19026 7384
rect 18972 7346 19024 7352
rect 18840 7284 18920 7290
rect 18788 7278 18920 7284
rect 18800 7262 18920 7278
rect 18696 7200 18748 7206
rect 18696 7142 18748 7148
rect 18708 6798 18736 7142
rect 18696 6792 18748 6798
rect 18694 6760 18696 6769
rect 18748 6760 18750 6769
rect 18800 6746 18828 7262
rect 18972 7200 19024 7206
rect 18972 7142 19024 7148
rect 18984 7018 19012 7142
rect 18892 6990 19012 7018
rect 18892 6866 18920 6990
rect 18972 6928 19024 6934
rect 18972 6870 19024 6876
rect 18880 6860 18932 6866
rect 18880 6802 18932 6808
rect 18800 6730 18920 6746
rect 18800 6724 18932 6730
rect 18800 6718 18880 6724
rect 18694 6695 18750 6704
rect 18880 6666 18932 6672
rect 18788 6656 18840 6662
rect 18788 6598 18840 6604
rect 18800 6497 18828 6598
rect 18786 6488 18842 6497
rect 18786 6423 18842 6432
rect 18800 6322 18828 6423
rect 18984 6322 19012 6870
rect 19076 6361 19104 8327
rect 19340 8288 19392 8294
rect 19340 8230 19392 8236
rect 19352 7954 19380 8230
rect 19340 7948 19392 7954
rect 19340 7890 19392 7896
rect 19340 7744 19392 7750
rect 19444 7732 19472 9658
rect 19536 8498 19564 11154
rect 19628 10266 19656 11222
rect 19720 11121 19748 11478
rect 19904 11370 19932 12174
rect 19812 11342 19932 11370
rect 19706 11112 19762 11121
rect 19706 11047 19708 11056
rect 19760 11047 19762 11056
rect 19708 11018 19760 11024
rect 19720 10987 19748 11018
rect 19708 10600 19760 10606
rect 19708 10542 19760 10548
rect 19616 10260 19668 10266
rect 19616 10202 19668 10208
rect 19720 9994 19748 10542
rect 19708 9988 19760 9994
rect 19708 9930 19760 9936
rect 19616 9376 19668 9382
rect 19616 9318 19668 9324
rect 19628 8974 19656 9318
rect 19616 8968 19668 8974
rect 19616 8910 19668 8916
rect 19524 8492 19576 8498
rect 19524 8434 19576 8440
rect 19392 7704 19472 7732
rect 19340 7686 19392 7692
rect 19352 7410 19380 7686
rect 19340 7404 19392 7410
rect 19340 7346 19392 7352
rect 19432 7268 19484 7274
rect 19432 7210 19484 7216
rect 19340 6792 19392 6798
rect 19154 6760 19210 6769
rect 19154 6695 19210 6704
rect 19338 6760 19340 6769
rect 19392 6760 19394 6769
rect 19338 6695 19394 6704
rect 19062 6352 19118 6361
rect 18788 6316 18840 6322
rect 18788 6258 18840 6264
rect 18972 6316 19024 6322
rect 19168 6322 19196 6695
rect 19340 6656 19392 6662
rect 19340 6598 19392 6604
rect 19352 6390 19380 6598
rect 19340 6384 19392 6390
rect 19340 6326 19392 6332
rect 19062 6287 19118 6296
rect 19156 6316 19208 6322
rect 18972 6258 19024 6264
rect 19156 6258 19208 6264
rect 18696 6112 18748 6118
rect 18696 6054 18748 6060
rect 19340 6112 19392 6118
rect 19340 6054 19392 6060
rect 18708 5778 18736 6054
rect 19352 5846 19380 6054
rect 18972 5840 19024 5846
rect 19340 5840 19392 5846
rect 18972 5782 19024 5788
rect 19154 5808 19210 5817
rect 18696 5772 18748 5778
rect 18696 5714 18748 5720
rect 18696 5636 18748 5642
rect 18696 5578 18748 5584
rect 18604 5228 18656 5234
rect 18604 5170 18656 5176
rect 18708 5098 18736 5578
rect 18984 5370 19012 5782
rect 19340 5782 19392 5788
rect 19154 5743 19156 5752
rect 19208 5743 19210 5752
rect 19156 5714 19208 5720
rect 19352 5574 19380 5782
rect 19444 5642 19472 7210
rect 19536 6458 19564 8434
rect 19628 7546 19656 8910
rect 19616 7540 19668 7546
rect 19616 7482 19668 7488
rect 19616 7404 19668 7410
rect 19616 7346 19668 7352
rect 19628 6474 19656 7346
rect 19720 6662 19748 9930
rect 19812 7970 19840 11342
rect 19892 11280 19944 11286
rect 19892 11222 19944 11228
rect 19904 11150 19932 11222
rect 19892 11144 19944 11150
rect 19892 11086 19944 11092
rect 19904 10742 19932 11086
rect 19892 10736 19944 10742
rect 19892 10678 19944 10684
rect 19890 9752 19946 9761
rect 19890 9687 19946 9696
rect 19904 9586 19932 9687
rect 19892 9580 19944 9586
rect 19892 9522 19944 9528
rect 19892 8900 19944 8906
rect 19996 8888 20024 13874
rect 20260 13320 20312 13326
rect 20260 13262 20312 13268
rect 20272 13190 20300 13262
rect 20260 13184 20312 13190
rect 20260 13126 20312 13132
rect 20168 12844 20220 12850
rect 20168 12786 20220 12792
rect 20180 12442 20208 12786
rect 20168 12436 20220 12442
rect 20168 12378 20220 12384
rect 20076 12232 20128 12238
rect 20074 12200 20076 12209
rect 20128 12200 20130 12209
rect 20074 12135 20130 12144
rect 20180 11830 20208 12378
rect 20076 11824 20128 11830
rect 20076 11766 20128 11772
rect 20168 11824 20220 11830
rect 20168 11766 20220 11772
rect 20088 10130 20116 11766
rect 20272 11762 20300 13126
rect 20260 11756 20312 11762
rect 20260 11698 20312 11704
rect 20168 11688 20220 11694
rect 20168 11630 20220 11636
rect 20076 10124 20128 10130
rect 20076 10066 20128 10072
rect 20076 9512 20128 9518
rect 20074 9480 20076 9489
rect 20128 9480 20130 9489
rect 20074 9415 20130 9424
rect 20180 8906 20208 11630
rect 20364 11354 20392 13874
rect 20456 11762 20484 14350
rect 21640 14340 21692 14346
rect 21640 14282 21692 14288
rect 20833 13628 21141 13637
rect 20833 13626 20839 13628
rect 20895 13626 20919 13628
rect 20975 13626 20999 13628
rect 21055 13626 21079 13628
rect 21135 13626 21141 13628
rect 20895 13574 20897 13626
rect 21077 13574 21079 13626
rect 20833 13572 20839 13574
rect 20895 13572 20919 13574
rect 20975 13572 20999 13574
rect 21055 13572 21079 13574
rect 21135 13572 21141 13574
rect 20833 13563 21141 13572
rect 21652 13326 21680 14282
rect 23673 14172 23981 14181
rect 23673 14170 23679 14172
rect 23735 14170 23759 14172
rect 23815 14170 23839 14172
rect 23895 14170 23919 14172
rect 23975 14170 23981 14172
rect 23735 14118 23737 14170
rect 23917 14118 23919 14170
rect 23673 14116 23679 14118
rect 23735 14116 23759 14118
rect 23815 14116 23839 14118
rect 23895 14116 23919 14118
rect 23975 14116 23981 14118
rect 23673 14107 23981 14116
rect 21272 13320 21324 13326
rect 21272 13262 21324 13268
rect 21640 13320 21692 13326
rect 21640 13262 21692 13268
rect 20536 13252 20588 13258
rect 20536 13194 20588 13200
rect 20548 12714 20576 13194
rect 20626 12880 20682 12889
rect 20626 12815 20682 12824
rect 20812 12844 20864 12850
rect 20536 12708 20588 12714
rect 20536 12650 20588 12656
rect 20444 11756 20496 11762
rect 20444 11698 20496 11704
rect 20444 11620 20496 11626
rect 20444 11562 20496 11568
rect 20352 11348 20404 11354
rect 20352 11290 20404 11296
rect 20352 11076 20404 11082
rect 20352 11018 20404 11024
rect 20364 10169 20392 11018
rect 20456 10810 20484 11562
rect 20536 11008 20588 11014
rect 20534 10976 20536 10985
rect 20588 10976 20590 10985
rect 20534 10911 20590 10920
rect 20444 10804 20496 10810
rect 20444 10746 20496 10752
rect 20536 10804 20588 10810
rect 20536 10746 20588 10752
rect 20350 10160 20406 10169
rect 20350 10095 20406 10104
rect 20260 9988 20312 9994
rect 20260 9930 20312 9936
rect 19944 8860 20024 8888
rect 19892 8842 19944 8848
rect 19892 8492 19944 8498
rect 19996 8480 20024 8860
rect 20168 8900 20220 8906
rect 20168 8842 20220 8848
rect 20076 8492 20128 8498
rect 19996 8452 20076 8480
rect 19892 8434 19944 8440
rect 20076 8434 20128 8440
rect 19904 8090 19932 8434
rect 19892 8084 19944 8090
rect 19892 8026 19944 8032
rect 19812 7942 19932 7970
rect 19800 7472 19852 7478
rect 19800 7414 19852 7420
rect 19812 7313 19840 7414
rect 19798 7304 19854 7313
rect 19798 7239 19854 7248
rect 19812 6866 19840 7239
rect 19800 6860 19852 6866
rect 19800 6802 19852 6808
rect 19904 6798 19932 7942
rect 20180 7886 20208 8842
rect 20272 8514 20300 9930
rect 20444 9920 20496 9926
rect 20444 9862 20496 9868
rect 20456 9654 20484 9862
rect 20444 9648 20496 9654
rect 20548 9625 20576 10746
rect 20640 10674 20668 12815
rect 20812 12786 20864 12792
rect 20824 12646 20852 12786
rect 20812 12640 20864 12646
rect 20812 12582 20864 12588
rect 20833 12540 21141 12549
rect 20833 12538 20839 12540
rect 20895 12538 20919 12540
rect 20975 12538 20999 12540
rect 21055 12538 21079 12540
rect 21135 12538 21141 12540
rect 20895 12486 20897 12538
rect 21077 12486 21079 12538
rect 20833 12484 20839 12486
rect 20895 12484 20919 12486
rect 20975 12484 20999 12486
rect 21055 12484 21079 12486
rect 21135 12484 21141 12486
rect 20833 12475 21141 12484
rect 21088 12232 21140 12238
rect 21088 12174 21140 12180
rect 20720 12164 20772 12170
rect 20720 12106 20772 12112
rect 20732 11354 20760 12106
rect 21100 11642 21128 12174
rect 21180 12164 21232 12170
rect 21180 12106 21232 12112
rect 21192 11762 21220 12106
rect 21180 11756 21232 11762
rect 21180 11698 21232 11704
rect 21100 11614 21220 11642
rect 20833 11452 21141 11461
rect 20833 11450 20839 11452
rect 20895 11450 20919 11452
rect 20975 11450 20999 11452
rect 21055 11450 21079 11452
rect 21135 11450 21141 11452
rect 20895 11398 20897 11450
rect 21077 11398 21079 11450
rect 20833 11396 20839 11398
rect 20895 11396 20919 11398
rect 20975 11396 20999 11398
rect 21055 11396 21079 11398
rect 21135 11396 21141 11398
rect 20833 11387 21141 11396
rect 20720 11348 20772 11354
rect 20720 11290 20772 11296
rect 21192 11218 21220 11614
rect 21180 11212 21232 11218
rect 21180 11154 21232 11160
rect 20996 11144 21048 11150
rect 20812 11138 20864 11144
rect 20720 11122 20772 11128
rect 20718 11112 20720 11121
rect 20772 11112 20774 11121
rect 20996 11086 21048 11092
rect 20812 11080 20864 11086
rect 20718 11047 20774 11056
rect 20628 10668 20680 10674
rect 20628 10610 20680 10616
rect 20444 9590 20496 9596
rect 20534 9616 20590 9625
rect 20352 9580 20404 9586
rect 20534 9551 20536 9560
rect 20352 9522 20404 9528
rect 20588 9551 20590 9560
rect 20536 9522 20588 9528
rect 20364 9353 20392 9522
rect 20444 9444 20496 9450
rect 20444 9386 20496 9392
rect 20350 9344 20406 9353
rect 20350 9279 20406 9288
rect 20352 9172 20404 9178
rect 20352 9114 20404 9120
rect 20364 8634 20392 9114
rect 20456 9042 20484 9386
rect 20534 9344 20590 9353
rect 20640 9330 20668 10610
rect 20824 10452 20852 11080
rect 21008 10985 21036 11086
rect 20994 10976 21050 10985
rect 20994 10911 21050 10920
rect 21008 10810 21036 10911
rect 20996 10804 21048 10810
rect 20996 10746 21048 10752
rect 21284 10713 21312 13262
rect 21652 12238 21680 13262
rect 23673 13084 23981 13093
rect 23673 13082 23679 13084
rect 23735 13082 23759 13084
rect 23815 13082 23839 13084
rect 23895 13082 23919 13084
rect 23975 13082 23981 13084
rect 23735 13030 23737 13082
rect 23917 13030 23919 13082
rect 23673 13028 23679 13030
rect 23735 13028 23759 13030
rect 23815 13028 23839 13030
rect 23895 13028 23919 13030
rect 23975 13028 23981 13030
rect 23673 13019 23981 13028
rect 21732 12640 21784 12646
rect 21732 12582 21784 12588
rect 22100 12640 22152 12646
rect 22100 12582 22152 12588
rect 21640 12232 21692 12238
rect 21640 12174 21692 12180
rect 21364 12096 21416 12102
rect 21364 12038 21416 12044
rect 21270 10704 21326 10713
rect 21270 10639 21326 10648
rect 20732 10424 20852 10452
rect 20732 9450 20760 10424
rect 20833 10364 21141 10373
rect 20833 10362 20839 10364
rect 20895 10362 20919 10364
rect 20975 10362 20999 10364
rect 21055 10362 21079 10364
rect 21135 10362 21141 10364
rect 20895 10310 20897 10362
rect 21077 10310 21079 10362
rect 20833 10308 20839 10310
rect 20895 10308 20919 10310
rect 20975 10308 20999 10310
rect 21055 10308 21079 10310
rect 21135 10308 21141 10310
rect 20833 10299 21141 10308
rect 20904 10260 20956 10266
rect 20904 10202 20956 10208
rect 21180 10260 21232 10266
rect 21180 10202 21232 10208
rect 20916 10169 20944 10202
rect 20902 10160 20958 10169
rect 20902 10095 20958 10104
rect 21192 9586 21220 10202
rect 21284 10198 21312 10639
rect 21376 10606 21404 12038
rect 21640 11756 21692 11762
rect 21640 11698 21692 11704
rect 21652 11082 21680 11698
rect 21744 11354 21772 12582
rect 22112 12170 22140 12582
rect 22100 12164 22152 12170
rect 22100 12106 22152 12112
rect 23112 12164 23164 12170
rect 23112 12106 23164 12112
rect 22560 12096 22612 12102
rect 22560 12038 22612 12044
rect 21824 11824 21876 11830
rect 21824 11766 21876 11772
rect 21732 11348 21784 11354
rect 21732 11290 21784 11296
rect 21640 11076 21692 11082
rect 21640 11018 21692 11024
rect 21364 10600 21416 10606
rect 21364 10542 21416 10548
rect 21272 10192 21324 10198
rect 21272 10134 21324 10140
rect 21180 9580 21232 9586
rect 21180 9522 21232 9528
rect 20720 9444 20772 9450
rect 20720 9386 20772 9392
rect 21180 9376 21232 9382
rect 20640 9302 20760 9330
rect 21180 9318 21232 9324
rect 20534 9279 20590 9288
rect 20548 9178 20576 9279
rect 20536 9172 20588 9178
rect 20536 9114 20588 9120
rect 20444 9036 20496 9042
rect 20444 8978 20496 8984
rect 20732 8974 20760 9302
rect 20833 9276 21141 9285
rect 20833 9274 20839 9276
rect 20895 9274 20919 9276
rect 20975 9274 20999 9276
rect 21055 9274 21079 9276
rect 21135 9274 21141 9276
rect 20895 9222 20897 9274
rect 21077 9222 21079 9274
rect 20833 9220 20839 9222
rect 20895 9220 20919 9222
rect 20975 9220 20999 9222
rect 21055 9220 21079 9222
rect 21135 9220 21141 9222
rect 20833 9211 21141 9220
rect 21192 9160 21220 9318
rect 21100 9132 21220 9160
rect 20996 9104 21048 9110
rect 20996 9046 21048 9052
rect 20536 8968 20588 8974
rect 20720 8968 20772 8974
rect 20588 8916 20668 8922
rect 20536 8910 20668 8916
rect 20720 8910 20772 8916
rect 20548 8894 20668 8910
rect 20536 8832 20588 8838
rect 20536 8774 20588 8780
rect 20352 8628 20404 8634
rect 20352 8570 20404 8576
rect 20272 8486 20484 8514
rect 20258 8120 20314 8129
rect 20258 8055 20260 8064
rect 20312 8055 20314 8064
rect 20260 8026 20312 8032
rect 20168 7880 20220 7886
rect 20168 7822 20220 7828
rect 20352 7744 20404 7750
rect 20352 7686 20404 7692
rect 19982 7440 20038 7449
rect 19982 7375 19984 7384
rect 20036 7375 20038 7384
rect 19984 7346 20036 7352
rect 20364 6866 20392 7686
rect 20456 7002 20484 8486
rect 20548 7886 20576 8774
rect 20640 8634 20668 8894
rect 20732 8838 20760 8910
rect 20720 8832 20772 8838
rect 20720 8774 20772 8780
rect 20628 8628 20680 8634
rect 20628 8570 20680 8576
rect 20640 8430 20668 8570
rect 21008 8498 21036 9046
rect 20720 8492 20772 8498
rect 20720 8434 20772 8440
rect 20996 8492 21048 8498
rect 20996 8434 21048 8440
rect 20628 8424 20680 8430
rect 20628 8366 20680 8372
rect 20732 7970 20760 8434
rect 20810 8392 20866 8401
rect 20810 8327 20812 8336
rect 20864 8327 20866 8336
rect 20812 8298 20864 8304
rect 21100 8294 21128 9132
rect 21180 8832 21232 8838
rect 21180 8774 21232 8780
rect 21088 8288 21140 8294
rect 21088 8230 21140 8236
rect 20833 8188 21141 8197
rect 20833 8186 20839 8188
rect 20895 8186 20919 8188
rect 20975 8186 20999 8188
rect 21055 8186 21079 8188
rect 21135 8186 21141 8188
rect 20895 8134 20897 8186
rect 21077 8134 21079 8186
rect 20833 8132 20839 8134
rect 20895 8132 20919 8134
rect 20975 8132 20999 8134
rect 21055 8132 21079 8134
rect 21135 8132 21141 8134
rect 20833 8123 21141 8132
rect 20640 7942 20760 7970
rect 20536 7880 20588 7886
rect 20536 7822 20588 7828
rect 20444 6996 20496 7002
rect 20444 6938 20496 6944
rect 20352 6860 20404 6866
rect 20352 6802 20404 6808
rect 19892 6792 19944 6798
rect 19892 6734 19944 6740
rect 20076 6792 20128 6798
rect 20076 6734 20128 6740
rect 19800 6724 19852 6730
rect 19800 6666 19852 6672
rect 19708 6656 19760 6662
rect 19708 6598 19760 6604
rect 19812 6474 19840 6666
rect 19524 6452 19576 6458
rect 19524 6394 19576 6400
rect 19628 6446 19840 6474
rect 19628 6118 19656 6446
rect 19904 6186 19932 6734
rect 19984 6248 20036 6254
rect 20088 6236 20116 6734
rect 20260 6316 20312 6322
rect 20260 6258 20312 6264
rect 20036 6208 20116 6236
rect 19984 6190 20036 6196
rect 20272 6186 20300 6258
rect 20456 6186 20484 6938
rect 20536 6860 20588 6866
rect 20536 6802 20588 6808
rect 20548 6458 20576 6802
rect 20640 6798 20668 7942
rect 20720 7812 20772 7818
rect 20720 7754 20772 7760
rect 20732 6866 20760 7754
rect 20812 7404 20864 7410
rect 20812 7346 20864 7352
rect 20824 7313 20852 7346
rect 20810 7304 20866 7313
rect 20810 7239 20866 7248
rect 20833 7100 21141 7109
rect 20833 7098 20839 7100
rect 20895 7098 20919 7100
rect 20975 7098 20999 7100
rect 21055 7098 21079 7100
rect 21135 7098 21141 7100
rect 20895 7046 20897 7098
rect 21077 7046 21079 7098
rect 20833 7044 20839 7046
rect 20895 7044 20919 7046
rect 20975 7044 20999 7046
rect 21055 7044 21079 7046
rect 21135 7044 21141 7046
rect 20833 7035 21141 7044
rect 20720 6860 20772 6866
rect 20720 6802 20772 6808
rect 20628 6792 20680 6798
rect 20628 6734 20680 6740
rect 20536 6452 20588 6458
rect 20536 6394 20588 6400
rect 19892 6180 19944 6186
rect 19892 6122 19944 6128
rect 20260 6180 20312 6186
rect 20260 6122 20312 6128
rect 20444 6180 20496 6186
rect 20444 6122 20496 6128
rect 19616 6112 19668 6118
rect 19616 6054 19668 6060
rect 20456 5914 20484 6122
rect 19616 5908 19668 5914
rect 19616 5850 19668 5856
rect 20444 5908 20496 5914
rect 20444 5850 20496 5856
rect 19432 5636 19484 5642
rect 19432 5578 19484 5584
rect 19340 5568 19392 5574
rect 19340 5510 19392 5516
rect 18972 5364 19024 5370
rect 18972 5306 19024 5312
rect 19444 5166 19472 5578
rect 19628 5234 19656 5850
rect 20548 5642 20576 6394
rect 20640 5914 20668 6734
rect 21192 6497 21220 8774
rect 21284 7478 21312 10134
rect 21376 8430 21404 10542
rect 21548 10532 21600 10538
rect 21548 10474 21600 10480
rect 21456 10464 21508 10470
rect 21456 10406 21508 10412
rect 21468 9926 21496 10406
rect 21456 9920 21508 9926
rect 21456 9862 21508 9868
rect 21468 9382 21496 9862
rect 21456 9376 21508 9382
rect 21456 9318 21508 9324
rect 21364 8424 21416 8430
rect 21364 8366 21416 8372
rect 21376 7886 21404 8366
rect 21364 7880 21416 7886
rect 21364 7822 21416 7828
rect 21272 7472 21324 7478
rect 21272 7414 21324 7420
rect 21454 7304 21510 7313
rect 21272 7268 21324 7274
rect 21560 7274 21588 10474
rect 21652 9042 21680 11018
rect 21744 10554 21772 11290
rect 21836 11150 21864 11766
rect 22572 11762 22600 12038
rect 22192 11756 22244 11762
rect 22192 11698 22244 11704
rect 22560 11756 22612 11762
rect 22560 11698 22612 11704
rect 21916 11688 21968 11694
rect 22204 11665 22232 11698
rect 21916 11630 21968 11636
rect 22190 11656 22246 11665
rect 21824 11144 21876 11150
rect 21824 11086 21876 11092
rect 21744 10526 21864 10554
rect 21732 9512 21784 9518
rect 21732 9454 21784 9460
rect 21640 9036 21692 9042
rect 21640 8978 21692 8984
rect 21640 8832 21692 8838
rect 21640 8774 21692 8780
rect 21652 8498 21680 8774
rect 21744 8498 21772 9454
rect 21640 8492 21692 8498
rect 21640 8434 21692 8440
rect 21732 8492 21784 8498
rect 21732 8434 21784 8440
rect 21744 7886 21772 8434
rect 21732 7880 21784 7886
rect 21732 7822 21784 7828
rect 21640 7744 21692 7750
rect 21640 7686 21692 7692
rect 21652 7546 21680 7686
rect 21640 7540 21692 7546
rect 21640 7482 21692 7488
rect 21744 7410 21772 7822
rect 21732 7404 21784 7410
rect 21732 7346 21784 7352
rect 21454 7239 21510 7248
rect 21548 7268 21600 7274
rect 21272 7210 21324 7216
rect 21284 6934 21312 7210
rect 21272 6928 21324 6934
rect 21272 6870 21324 6876
rect 21468 6798 21496 7239
rect 21548 7210 21600 7216
rect 21456 6792 21508 6798
rect 21456 6734 21508 6740
rect 21744 6633 21772 7346
rect 21730 6624 21786 6633
rect 21730 6559 21786 6568
rect 21178 6488 21234 6497
rect 21836 6458 21864 10526
rect 21928 7546 21956 11630
rect 22190 11591 22246 11600
rect 22008 11552 22060 11558
rect 22008 11494 22060 11500
rect 22192 11552 22244 11558
rect 22192 11494 22244 11500
rect 22020 9178 22048 11494
rect 22204 9586 22232 11494
rect 22192 9580 22244 9586
rect 22192 9522 22244 9528
rect 22468 9512 22520 9518
rect 22468 9454 22520 9460
rect 22376 9444 22428 9450
rect 22376 9386 22428 9392
rect 22192 9376 22244 9382
rect 22192 9318 22244 9324
rect 22008 9172 22060 9178
rect 22008 9114 22060 9120
rect 22204 9081 22232 9318
rect 22190 9072 22246 9081
rect 22190 9007 22246 9016
rect 22284 8968 22336 8974
rect 22284 8910 22336 8916
rect 22100 8832 22152 8838
rect 22100 8774 22152 8780
rect 22008 8628 22060 8634
rect 22008 8570 22060 8576
rect 22020 8362 22048 8570
rect 22008 8356 22060 8362
rect 22008 8298 22060 8304
rect 22112 7818 22140 8774
rect 22296 8634 22324 8910
rect 22284 8628 22336 8634
rect 22284 8570 22336 8576
rect 22192 8356 22244 8362
rect 22192 8298 22244 8304
rect 22100 7812 22152 7818
rect 22100 7754 22152 7760
rect 21916 7540 21968 7546
rect 21916 7482 21968 7488
rect 21178 6423 21234 6432
rect 21824 6452 21876 6458
rect 21824 6394 21876 6400
rect 20720 6316 20772 6322
rect 20720 6258 20772 6264
rect 20628 5908 20680 5914
rect 20628 5850 20680 5856
rect 20536 5636 20588 5642
rect 20536 5578 20588 5584
rect 20350 5536 20406 5545
rect 20350 5471 20406 5480
rect 20364 5234 20392 5471
rect 19616 5228 19668 5234
rect 19616 5170 19668 5176
rect 20352 5228 20404 5234
rect 20352 5170 20404 5176
rect 19432 5160 19484 5166
rect 19432 5102 19484 5108
rect 20364 5098 20392 5170
rect 18696 5092 18748 5098
rect 18696 5034 18748 5040
rect 20352 5092 20404 5098
rect 20352 5034 20404 5040
rect 18512 4752 18564 4758
rect 18512 4694 18564 4700
rect 17592 4684 17644 4690
rect 17592 4626 17644 4632
rect 20364 4622 20392 5034
rect 20548 5030 20576 5578
rect 20640 5370 20668 5850
rect 20628 5364 20680 5370
rect 20628 5306 20680 5312
rect 20732 5234 20760 6258
rect 21180 6248 21232 6254
rect 21180 6190 21232 6196
rect 20833 6012 21141 6021
rect 20833 6010 20839 6012
rect 20895 6010 20919 6012
rect 20975 6010 20999 6012
rect 21055 6010 21079 6012
rect 21135 6010 21141 6012
rect 20895 5958 20897 6010
rect 21077 5958 21079 6010
rect 20833 5956 20839 5958
rect 20895 5956 20919 5958
rect 20975 5956 20999 5958
rect 21055 5956 21079 5958
rect 21135 5956 21141 5958
rect 20833 5947 21141 5956
rect 20720 5228 20772 5234
rect 20720 5170 20772 5176
rect 21192 5098 21220 6190
rect 22112 6118 22140 7754
rect 22204 7750 22232 8298
rect 22296 8022 22324 8570
rect 22388 8498 22416 9386
rect 22480 8634 22508 9454
rect 22572 8838 22600 11698
rect 23124 11558 23152 12106
rect 23673 11996 23981 12005
rect 23673 11994 23679 11996
rect 23735 11994 23759 11996
rect 23815 11994 23839 11996
rect 23895 11994 23919 11996
rect 23975 11994 23981 11996
rect 23735 11942 23737 11994
rect 23917 11942 23919 11994
rect 23673 11940 23679 11942
rect 23735 11940 23759 11942
rect 23815 11940 23839 11942
rect 23895 11940 23919 11942
rect 23975 11940 23981 11942
rect 23673 11931 23981 11940
rect 23112 11552 23164 11558
rect 23112 11494 23164 11500
rect 23124 9926 23152 11494
rect 23673 10908 23981 10917
rect 23673 10906 23679 10908
rect 23735 10906 23759 10908
rect 23815 10906 23839 10908
rect 23895 10906 23919 10908
rect 23975 10906 23981 10908
rect 23735 10854 23737 10906
rect 23917 10854 23919 10906
rect 23673 10852 23679 10854
rect 23735 10852 23759 10854
rect 23815 10852 23839 10854
rect 23895 10852 23919 10854
rect 23975 10852 23981 10854
rect 23673 10843 23981 10852
rect 23112 9920 23164 9926
rect 23112 9862 23164 9868
rect 23020 9580 23072 9586
rect 23020 9522 23072 9528
rect 23032 8974 23060 9522
rect 23020 8968 23072 8974
rect 23020 8910 23072 8916
rect 22560 8832 22612 8838
rect 22560 8774 22612 8780
rect 22836 8832 22888 8838
rect 22836 8774 22888 8780
rect 22468 8628 22520 8634
rect 22468 8570 22520 8576
rect 22848 8566 22876 8774
rect 23032 8634 23060 8910
rect 23020 8628 23072 8634
rect 23020 8570 23072 8576
rect 22836 8560 22888 8566
rect 22836 8502 22888 8508
rect 22376 8492 22428 8498
rect 22376 8434 22428 8440
rect 23032 8294 23060 8570
rect 22560 8288 22612 8294
rect 22560 8230 22612 8236
rect 23020 8288 23072 8294
rect 23020 8230 23072 8236
rect 22284 8016 22336 8022
rect 22284 7958 22336 7964
rect 22192 7744 22244 7750
rect 22192 7686 22244 7692
rect 22296 7410 22324 7958
rect 22572 7410 22600 8230
rect 23020 7744 23072 7750
rect 23124 7732 23152 9862
rect 23673 9820 23981 9829
rect 23673 9818 23679 9820
rect 23735 9818 23759 9820
rect 23815 9818 23839 9820
rect 23895 9818 23919 9820
rect 23975 9818 23981 9820
rect 23735 9766 23737 9818
rect 23917 9766 23919 9818
rect 23673 9764 23679 9766
rect 23735 9764 23759 9766
rect 23815 9764 23839 9766
rect 23895 9764 23919 9766
rect 23975 9764 23981 9766
rect 23673 9755 23981 9764
rect 23673 8732 23981 8741
rect 23673 8730 23679 8732
rect 23735 8730 23759 8732
rect 23815 8730 23839 8732
rect 23895 8730 23919 8732
rect 23975 8730 23981 8732
rect 23735 8678 23737 8730
rect 23917 8678 23919 8730
rect 23673 8676 23679 8678
rect 23735 8676 23759 8678
rect 23815 8676 23839 8678
rect 23895 8676 23919 8678
rect 23975 8676 23981 8678
rect 23673 8667 23981 8676
rect 23072 7704 23152 7732
rect 23020 7686 23072 7692
rect 23032 7546 23060 7686
rect 23673 7644 23981 7653
rect 23673 7642 23679 7644
rect 23735 7642 23759 7644
rect 23815 7642 23839 7644
rect 23895 7642 23919 7644
rect 23975 7642 23981 7644
rect 23735 7590 23737 7642
rect 23917 7590 23919 7642
rect 23673 7588 23679 7590
rect 23735 7588 23759 7590
rect 23815 7588 23839 7590
rect 23895 7588 23919 7590
rect 23975 7588 23981 7590
rect 23673 7579 23981 7588
rect 23020 7540 23072 7546
rect 23020 7482 23072 7488
rect 22284 7404 22336 7410
rect 22284 7346 22336 7352
rect 22560 7404 22612 7410
rect 22560 7346 22612 7352
rect 23673 6556 23981 6565
rect 23673 6554 23679 6556
rect 23735 6554 23759 6556
rect 23815 6554 23839 6556
rect 23895 6554 23919 6556
rect 23975 6554 23981 6556
rect 23735 6502 23737 6554
rect 23917 6502 23919 6554
rect 23673 6500 23679 6502
rect 23735 6500 23759 6502
rect 23815 6500 23839 6502
rect 23895 6500 23919 6502
rect 23975 6500 23981 6502
rect 23673 6491 23981 6500
rect 22100 6112 22152 6118
rect 22100 6054 22152 6060
rect 21180 5092 21232 5098
rect 21180 5034 21232 5040
rect 20536 5024 20588 5030
rect 20536 4966 20588 4972
rect 20833 4924 21141 4933
rect 20833 4922 20839 4924
rect 20895 4922 20919 4924
rect 20975 4922 20999 4924
rect 21055 4922 21079 4924
rect 21135 4922 21141 4924
rect 20895 4870 20897 4922
rect 21077 4870 21079 4922
rect 20833 4868 20839 4870
rect 20895 4868 20919 4870
rect 20975 4868 20999 4870
rect 21055 4868 21079 4870
rect 21135 4868 21141 4870
rect 20833 4859 21141 4868
rect 22112 4826 22140 6054
rect 23673 5468 23981 5477
rect 23673 5466 23679 5468
rect 23735 5466 23759 5468
rect 23815 5466 23839 5468
rect 23895 5466 23919 5468
rect 23975 5466 23981 5468
rect 23735 5414 23737 5466
rect 23917 5414 23919 5466
rect 23673 5412 23679 5414
rect 23735 5412 23759 5414
rect 23815 5412 23839 5414
rect 23895 5412 23919 5414
rect 23975 5412 23981 5414
rect 23673 5403 23981 5412
rect 22100 4820 22152 4826
rect 22100 4762 22152 4768
rect 20352 4616 20404 4622
rect 20352 4558 20404 4564
rect 17992 4380 18300 4389
rect 17992 4378 17998 4380
rect 18054 4378 18078 4380
rect 18134 4378 18158 4380
rect 18214 4378 18238 4380
rect 18294 4378 18300 4380
rect 18054 4326 18056 4378
rect 18236 4326 18238 4378
rect 17992 4324 17998 4326
rect 18054 4324 18078 4326
rect 18134 4324 18158 4326
rect 18214 4324 18238 4326
rect 18294 4324 18300 4326
rect 17992 4315 18300 4324
rect 23673 4380 23981 4389
rect 23673 4378 23679 4380
rect 23735 4378 23759 4380
rect 23815 4378 23839 4380
rect 23895 4378 23919 4380
rect 23975 4378 23981 4380
rect 23735 4326 23737 4378
rect 23917 4326 23919 4378
rect 23673 4324 23679 4326
rect 23735 4324 23759 4326
rect 23815 4324 23839 4326
rect 23895 4324 23919 4326
rect 23975 4324 23981 4326
rect 23673 4315 23981 4324
rect 17132 4276 17184 4282
rect 17132 4218 17184 4224
rect 16672 4208 16724 4214
rect 16672 4150 16724 4156
rect 15752 4140 15804 4146
rect 15752 4082 15804 4088
rect 15152 3836 15460 3845
rect 15152 3834 15158 3836
rect 15214 3834 15238 3836
rect 15294 3834 15318 3836
rect 15374 3834 15398 3836
rect 15454 3834 15460 3836
rect 15214 3782 15216 3834
rect 15396 3782 15398 3834
rect 15152 3780 15158 3782
rect 15214 3780 15238 3782
rect 15294 3780 15318 3782
rect 15374 3780 15398 3782
rect 15454 3780 15460 3782
rect 15152 3771 15460 3780
rect 15016 3664 15068 3670
rect 15016 3606 15068 3612
rect 15764 3534 15792 4082
rect 16684 3738 16712 4150
rect 17406 4040 17462 4049
rect 17406 3975 17462 3984
rect 16672 3732 16724 3738
rect 16672 3674 16724 3680
rect 12348 3528 12400 3534
rect 12348 3470 12400 3476
rect 13912 3528 13964 3534
rect 13912 3470 13964 3476
rect 15752 3528 15804 3534
rect 15752 3470 15804 3476
rect 12311 3292 12619 3301
rect 12311 3290 12317 3292
rect 12373 3290 12397 3292
rect 12453 3290 12477 3292
rect 12533 3290 12557 3292
rect 12613 3290 12619 3292
rect 12373 3238 12375 3290
rect 12555 3238 12557 3290
rect 12311 3236 12317 3238
rect 12373 3236 12397 3238
rect 12453 3236 12477 3238
rect 12533 3236 12557 3238
rect 12613 3236 12619 3238
rect 12311 3227 12619 3236
rect 13924 3194 13952 3470
rect 14372 3460 14424 3466
rect 14372 3402 14424 3408
rect 14384 3194 14412 3402
rect 17316 3392 17368 3398
rect 17316 3334 17368 3340
rect 13912 3188 13964 3194
rect 13912 3130 13964 3136
rect 14372 3188 14424 3194
rect 14372 3130 14424 3136
rect 12164 3120 12216 3126
rect 12164 3062 12216 3068
rect 15660 2848 15712 2854
rect 15660 2790 15712 2796
rect 16856 2848 16908 2854
rect 16856 2790 16908 2796
rect 15152 2748 15460 2757
rect 15152 2746 15158 2748
rect 15214 2746 15238 2748
rect 15294 2746 15318 2748
rect 15374 2746 15398 2748
rect 15454 2746 15460 2748
rect 15214 2694 15216 2746
rect 15396 2694 15398 2746
rect 15152 2692 15158 2694
rect 15214 2692 15238 2694
rect 15294 2692 15318 2694
rect 15374 2692 15398 2694
rect 15454 2692 15460 2694
rect 15152 2683 15460 2692
rect 11980 2644 12032 2650
rect 11980 2586 12032 2592
rect 11612 2440 11664 2446
rect 11612 2382 11664 2388
rect 11888 2440 11940 2446
rect 11888 2382 11940 2388
rect 12716 2440 12768 2446
rect 12716 2382 12768 2388
rect 13084 2440 13136 2446
rect 13084 2382 13136 2388
rect 13728 2440 13780 2446
rect 13728 2382 13780 2388
rect 14372 2440 14424 2446
rect 14372 2382 14424 2388
rect 15016 2440 15068 2446
rect 15016 2382 15068 2388
rect 11796 2372 11848 2378
rect 11796 2314 11848 2320
rect 11808 800 11836 2314
rect 12311 2204 12619 2213
rect 12311 2202 12317 2204
rect 12373 2202 12397 2204
rect 12453 2202 12477 2204
rect 12533 2202 12557 2204
rect 12613 2202 12619 2204
rect 12373 2150 12375 2202
rect 12555 2150 12557 2202
rect 12311 2148 12317 2150
rect 12373 2148 12397 2150
rect 12453 2148 12477 2150
rect 12533 2148 12557 2150
rect 12613 2148 12619 2150
rect 12311 2139 12619 2148
rect 12452 870 12572 898
rect 12452 800 12480 870
rect 1490 0 1546 800
rect 2134 0 2190 800
rect 2778 0 2834 800
rect 3422 0 3478 800
rect 4066 0 4122 800
rect 4710 0 4766 800
rect 5354 0 5410 800
rect 5998 0 6054 800
rect 6642 0 6698 800
rect 7286 0 7342 800
rect 7930 0 7986 800
rect 8574 0 8630 800
rect 9218 0 9274 800
rect 9862 0 9918 800
rect 10506 0 10562 800
rect 11150 0 11206 800
rect 11794 0 11850 800
rect 12438 0 12494 800
rect 12544 762 12572 870
rect 12728 762 12756 2382
rect 13096 800 13124 2382
rect 13740 800 13768 2382
rect 14384 800 14412 2382
rect 15028 800 15056 2382
rect 15672 800 15700 2790
rect 16868 2650 16896 2790
rect 16856 2644 16908 2650
rect 16856 2586 16908 2592
rect 17328 2582 17356 3334
rect 17420 3194 17448 3975
rect 20833 3836 21141 3845
rect 20833 3834 20839 3836
rect 20895 3834 20919 3836
rect 20975 3834 20999 3836
rect 21055 3834 21079 3836
rect 21135 3834 21141 3836
rect 20895 3782 20897 3834
rect 21077 3782 21079 3834
rect 20833 3780 20839 3782
rect 20895 3780 20919 3782
rect 20975 3780 20999 3782
rect 21055 3780 21079 3782
rect 21135 3780 21141 3782
rect 20833 3771 21141 3780
rect 23388 3528 23440 3534
rect 17958 3496 18014 3505
rect 23388 3470 23440 3476
rect 17958 3431 17960 3440
rect 18012 3431 18014 3440
rect 17960 3402 18012 3408
rect 17992 3292 18300 3301
rect 17992 3290 17998 3292
rect 18054 3290 18078 3292
rect 18134 3290 18158 3292
rect 18214 3290 18238 3292
rect 18294 3290 18300 3292
rect 18054 3238 18056 3290
rect 18236 3238 18238 3290
rect 17992 3236 17998 3238
rect 18054 3236 18078 3238
rect 18134 3236 18158 3238
rect 18214 3236 18238 3238
rect 18294 3236 18300 3238
rect 17992 3227 18300 3236
rect 17408 3188 17460 3194
rect 17408 3130 17460 3136
rect 18328 2848 18380 2854
rect 18328 2790 18380 2796
rect 20720 2848 20772 2854
rect 20720 2790 20772 2796
rect 22744 2848 22796 2854
rect 22744 2790 22796 2796
rect 17316 2576 17368 2582
rect 17316 2518 17368 2524
rect 16304 2440 16356 2446
rect 16304 2382 16356 2388
rect 16948 2440 17000 2446
rect 16948 2382 17000 2388
rect 17592 2440 17644 2446
rect 17592 2382 17644 2388
rect 16316 800 16344 2382
rect 16396 2372 16448 2378
rect 16396 2314 16448 2320
rect 16408 2106 16436 2314
rect 16396 2100 16448 2106
rect 16396 2042 16448 2048
rect 16960 800 16988 2382
rect 17604 800 17632 2382
rect 17992 2204 18300 2213
rect 17992 2202 17998 2204
rect 18054 2202 18078 2204
rect 18134 2202 18158 2204
rect 18214 2202 18238 2204
rect 18294 2202 18300 2204
rect 18054 2150 18056 2202
rect 18236 2150 18238 2202
rect 17992 2148 17998 2150
rect 18054 2148 18078 2150
rect 18134 2148 18158 2150
rect 18214 2148 18238 2150
rect 18294 2148 18300 2150
rect 17992 2139 18300 2148
rect 18340 1442 18368 2790
rect 18880 2440 18932 2446
rect 18880 2382 18932 2388
rect 19524 2440 19576 2446
rect 19524 2382 19576 2388
rect 20168 2440 20220 2446
rect 20168 2382 20220 2388
rect 18248 1414 18368 1442
rect 18248 800 18276 1414
rect 18892 800 18920 2382
rect 19536 800 19564 2382
rect 20180 800 20208 2382
rect 20732 1442 20760 2790
rect 20833 2748 21141 2757
rect 20833 2746 20839 2748
rect 20895 2746 20919 2748
rect 20975 2746 20999 2748
rect 21055 2746 21079 2748
rect 21135 2746 21141 2748
rect 20895 2694 20897 2746
rect 21077 2694 21079 2746
rect 20833 2692 20839 2694
rect 20895 2692 20919 2694
rect 20975 2692 20999 2694
rect 21055 2692 21079 2694
rect 21135 2692 21141 2694
rect 20833 2683 21141 2692
rect 21456 2440 21508 2446
rect 21456 2382 21508 2388
rect 22100 2440 22152 2446
rect 22100 2382 22152 2388
rect 20732 1414 20852 1442
rect 20824 800 20852 1414
rect 21468 800 21496 2382
rect 22112 800 22140 2382
rect 22756 800 22784 2790
rect 23400 800 23428 3470
rect 23673 3292 23981 3301
rect 23673 3290 23679 3292
rect 23735 3290 23759 3292
rect 23815 3290 23839 3292
rect 23895 3290 23919 3292
rect 23975 3290 23981 3292
rect 23735 3238 23737 3290
rect 23917 3238 23919 3290
rect 23673 3236 23679 3238
rect 23735 3236 23759 3238
rect 23815 3236 23839 3238
rect 23895 3236 23919 3238
rect 23975 3236 23981 3238
rect 23673 3227 23981 3236
rect 23673 2204 23981 2213
rect 23673 2202 23679 2204
rect 23735 2202 23759 2204
rect 23815 2202 23839 2204
rect 23895 2202 23919 2204
rect 23975 2202 23981 2204
rect 23735 2150 23737 2202
rect 23917 2150 23919 2202
rect 23673 2148 23679 2150
rect 23735 2148 23759 2150
rect 23815 2148 23839 2150
rect 23895 2148 23919 2150
rect 23975 2148 23981 2150
rect 23673 2139 23981 2148
rect 12544 734 12756 762
rect 13082 0 13138 800
rect 13726 0 13782 800
rect 14370 0 14426 800
rect 15014 0 15070 800
rect 15658 0 15714 800
rect 16302 0 16358 800
rect 16946 0 17002 800
rect 17590 0 17646 800
rect 18234 0 18290 800
rect 18878 0 18934 800
rect 19522 0 19578 800
rect 20166 0 20222 800
rect 20810 0 20866 800
rect 21454 0 21510 800
rect 22098 0 22154 800
rect 22742 0 22798 800
rect 23386 0 23442 800
<< via2 >>
rect 3796 22330 3852 22332
rect 3876 22330 3932 22332
rect 3956 22330 4012 22332
rect 4036 22330 4092 22332
rect 3796 22278 3842 22330
rect 3842 22278 3852 22330
rect 3876 22278 3906 22330
rect 3906 22278 3918 22330
rect 3918 22278 3932 22330
rect 3956 22278 3970 22330
rect 3970 22278 3982 22330
rect 3982 22278 4012 22330
rect 4036 22278 4046 22330
rect 4046 22278 4092 22330
rect 3796 22276 3852 22278
rect 3876 22276 3932 22278
rect 3956 22276 4012 22278
rect 4036 22276 4092 22278
rect 9477 22330 9533 22332
rect 9557 22330 9613 22332
rect 9637 22330 9693 22332
rect 9717 22330 9773 22332
rect 9477 22278 9523 22330
rect 9523 22278 9533 22330
rect 9557 22278 9587 22330
rect 9587 22278 9599 22330
rect 9599 22278 9613 22330
rect 9637 22278 9651 22330
rect 9651 22278 9663 22330
rect 9663 22278 9693 22330
rect 9717 22278 9727 22330
rect 9727 22278 9773 22330
rect 9477 22276 9533 22278
rect 9557 22276 9613 22278
rect 9637 22276 9693 22278
rect 9717 22276 9773 22278
rect 15158 22330 15214 22332
rect 15238 22330 15294 22332
rect 15318 22330 15374 22332
rect 15398 22330 15454 22332
rect 15158 22278 15204 22330
rect 15204 22278 15214 22330
rect 15238 22278 15268 22330
rect 15268 22278 15280 22330
rect 15280 22278 15294 22330
rect 15318 22278 15332 22330
rect 15332 22278 15344 22330
rect 15344 22278 15374 22330
rect 15398 22278 15408 22330
rect 15408 22278 15454 22330
rect 15158 22276 15214 22278
rect 15238 22276 15294 22278
rect 15318 22276 15374 22278
rect 15398 22276 15454 22278
rect 20839 22330 20895 22332
rect 20919 22330 20975 22332
rect 20999 22330 21055 22332
rect 21079 22330 21135 22332
rect 20839 22278 20885 22330
rect 20885 22278 20895 22330
rect 20919 22278 20949 22330
rect 20949 22278 20961 22330
rect 20961 22278 20975 22330
rect 20999 22278 21013 22330
rect 21013 22278 21025 22330
rect 21025 22278 21055 22330
rect 21079 22278 21089 22330
rect 21089 22278 21135 22330
rect 20839 22276 20895 22278
rect 20919 22276 20975 22278
rect 20999 22276 21055 22278
rect 21079 22276 21135 22278
rect 6636 21786 6692 21788
rect 6716 21786 6772 21788
rect 6796 21786 6852 21788
rect 6876 21786 6932 21788
rect 6636 21734 6682 21786
rect 6682 21734 6692 21786
rect 6716 21734 6746 21786
rect 6746 21734 6758 21786
rect 6758 21734 6772 21786
rect 6796 21734 6810 21786
rect 6810 21734 6822 21786
rect 6822 21734 6852 21786
rect 6876 21734 6886 21786
rect 6886 21734 6932 21786
rect 6636 21732 6692 21734
rect 6716 21732 6772 21734
rect 6796 21732 6852 21734
rect 6876 21732 6932 21734
rect 3796 21242 3852 21244
rect 3876 21242 3932 21244
rect 3956 21242 4012 21244
rect 4036 21242 4092 21244
rect 3796 21190 3842 21242
rect 3842 21190 3852 21242
rect 3876 21190 3906 21242
rect 3906 21190 3918 21242
rect 3918 21190 3932 21242
rect 3956 21190 3970 21242
rect 3970 21190 3982 21242
rect 3982 21190 4012 21242
rect 4036 21190 4046 21242
rect 4046 21190 4092 21242
rect 3796 21188 3852 21190
rect 3876 21188 3932 21190
rect 3956 21188 4012 21190
rect 4036 21188 4092 21190
rect 4894 20748 4896 20768
rect 4896 20748 4948 20768
rect 4948 20748 4950 20768
rect 4894 20712 4950 20748
rect 3796 20154 3852 20156
rect 3876 20154 3932 20156
rect 3956 20154 4012 20156
rect 4036 20154 4092 20156
rect 3796 20102 3842 20154
rect 3842 20102 3852 20154
rect 3876 20102 3906 20154
rect 3906 20102 3918 20154
rect 3918 20102 3932 20154
rect 3956 20102 3970 20154
rect 3970 20102 3982 20154
rect 3982 20102 4012 20154
rect 4036 20102 4046 20154
rect 4046 20102 4092 20154
rect 3796 20100 3852 20102
rect 3876 20100 3932 20102
rect 3956 20100 4012 20102
rect 4036 20100 4092 20102
rect 3698 19352 3754 19408
rect 3796 19066 3852 19068
rect 3876 19066 3932 19068
rect 3956 19066 4012 19068
rect 4036 19066 4092 19068
rect 3796 19014 3842 19066
rect 3842 19014 3852 19066
rect 3876 19014 3906 19066
rect 3906 19014 3918 19066
rect 3918 19014 3932 19066
rect 3956 19014 3970 19066
rect 3970 19014 3982 19066
rect 3982 19014 4012 19066
rect 4036 19014 4046 19066
rect 4046 19014 4092 19066
rect 3796 19012 3852 19014
rect 3876 19012 3932 19014
rect 3956 19012 4012 19014
rect 4036 19012 4092 19014
rect 3422 16632 3478 16688
rect 3796 17978 3852 17980
rect 3876 17978 3932 17980
rect 3956 17978 4012 17980
rect 4036 17978 4092 17980
rect 3796 17926 3842 17978
rect 3842 17926 3852 17978
rect 3876 17926 3906 17978
rect 3906 17926 3918 17978
rect 3918 17926 3932 17978
rect 3956 17926 3970 17978
rect 3970 17926 3982 17978
rect 3982 17926 4012 17978
rect 4036 17926 4046 17978
rect 4046 17926 4092 17978
rect 3796 17924 3852 17926
rect 3876 17924 3932 17926
rect 3956 17924 4012 17926
rect 4036 17924 4092 17926
rect 3796 16890 3852 16892
rect 3876 16890 3932 16892
rect 3956 16890 4012 16892
rect 4036 16890 4092 16892
rect 3796 16838 3842 16890
rect 3842 16838 3852 16890
rect 3876 16838 3906 16890
rect 3906 16838 3918 16890
rect 3918 16838 3932 16890
rect 3956 16838 3970 16890
rect 3970 16838 3982 16890
rect 3982 16838 4012 16890
rect 4036 16838 4046 16890
rect 4046 16838 4092 16890
rect 3796 16836 3852 16838
rect 3876 16836 3932 16838
rect 3956 16836 4012 16838
rect 4036 16836 4092 16838
rect 3238 10532 3294 10568
rect 3238 10512 3240 10532
rect 3240 10512 3292 10532
rect 3292 10512 3294 10532
rect 3796 15802 3852 15804
rect 3876 15802 3932 15804
rect 3956 15802 4012 15804
rect 4036 15802 4092 15804
rect 3796 15750 3842 15802
rect 3842 15750 3852 15802
rect 3876 15750 3906 15802
rect 3906 15750 3918 15802
rect 3918 15750 3932 15802
rect 3956 15750 3970 15802
rect 3970 15750 3982 15802
rect 3982 15750 4012 15802
rect 4036 15750 4046 15802
rect 4046 15750 4092 15802
rect 3796 15748 3852 15750
rect 3876 15748 3932 15750
rect 3956 15748 4012 15750
rect 4036 15748 4092 15750
rect 3796 14714 3852 14716
rect 3876 14714 3932 14716
rect 3956 14714 4012 14716
rect 4036 14714 4092 14716
rect 3796 14662 3842 14714
rect 3842 14662 3852 14714
rect 3876 14662 3906 14714
rect 3906 14662 3918 14714
rect 3918 14662 3932 14714
rect 3956 14662 3970 14714
rect 3970 14662 3982 14714
rect 3982 14662 4012 14714
rect 4036 14662 4046 14714
rect 4046 14662 4092 14714
rect 3796 14660 3852 14662
rect 3876 14660 3932 14662
rect 3956 14660 4012 14662
rect 4036 14660 4092 14662
rect 4434 15000 4490 15056
rect 2870 4140 2926 4176
rect 2870 4120 2872 4140
rect 2872 4120 2924 4140
rect 2924 4120 2926 4140
rect 2502 3984 2558 4040
rect 3796 13626 3852 13628
rect 3876 13626 3932 13628
rect 3956 13626 4012 13628
rect 4036 13626 4092 13628
rect 3796 13574 3842 13626
rect 3842 13574 3852 13626
rect 3876 13574 3906 13626
rect 3906 13574 3918 13626
rect 3918 13574 3932 13626
rect 3956 13574 3970 13626
rect 3970 13574 3982 13626
rect 3982 13574 4012 13626
rect 4036 13574 4046 13626
rect 4046 13574 4092 13626
rect 3796 13572 3852 13574
rect 3876 13572 3932 13574
rect 3956 13572 4012 13574
rect 4036 13572 4092 13574
rect 4526 13776 4582 13832
rect 3796 12538 3852 12540
rect 3876 12538 3932 12540
rect 3956 12538 4012 12540
rect 4036 12538 4092 12540
rect 3796 12486 3842 12538
rect 3842 12486 3852 12538
rect 3876 12486 3906 12538
rect 3906 12486 3918 12538
rect 3918 12486 3932 12538
rect 3956 12486 3970 12538
rect 3970 12486 3982 12538
rect 3982 12486 4012 12538
rect 4036 12486 4046 12538
rect 4046 12486 4092 12538
rect 3796 12484 3852 12486
rect 3876 12484 3932 12486
rect 3956 12484 4012 12486
rect 4036 12484 4092 12486
rect 5078 14048 5134 14104
rect 4526 12552 4582 12608
rect 4250 11892 4306 11928
rect 4250 11872 4252 11892
rect 4252 11872 4304 11892
rect 4304 11872 4306 11892
rect 3796 11450 3852 11452
rect 3876 11450 3932 11452
rect 3956 11450 4012 11452
rect 4036 11450 4092 11452
rect 3796 11398 3842 11450
rect 3842 11398 3852 11450
rect 3876 11398 3906 11450
rect 3906 11398 3918 11450
rect 3918 11398 3932 11450
rect 3956 11398 3970 11450
rect 3970 11398 3982 11450
rect 3982 11398 4012 11450
rect 4036 11398 4046 11450
rect 4046 11398 4092 11450
rect 3796 11396 3852 11398
rect 3876 11396 3932 11398
rect 3956 11396 4012 11398
rect 4036 11396 4092 11398
rect 3796 10362 3852 10364
rect 3876 10362 3932 10364
rect 3956 10362 4012 10364
rect 4036 10362 4092 10364
rect 3796 10310 3842 10362
rect 3842 10310 3852 10362
rect 3876 10310 3906 10362
rect 3906 10310 3918 10362
rect 3918 10310 3932 10362
rect 3956 10310 3970 10362
rect 3970 10310 3982 10362
rect 3982 10310 4012 10362
rect 4036 10310 4046 10362
rect 4046 10310 4092 10362
rect 3796 10308 3852 10310
rect 3876 10308 3932 10310
rect 3956 10308 4012 10310
rect 4036 10308 4092 10310
rect 3796 9274 3852 9276
rect 3876 9274 3932 9276
rect 3956 9274 4012 9276
rect 4036 9274 4092 9276
rect 3796 9222 3842 9274
rect 3842 9222 3852 9274
rect 3876 9222 3906 9274
rect 3906 9222 3918 9274
rect 3918 9222 3932 9274
rect 3956 9222 3970 9274
rect 3970 9222 3982 9274
rect 3982 9222 4012 9274
rect 4036 9222 4046 9274
rect 4046 9222 4092 9274
rect 3796 9220 3852 9222
rect 3876 9220 3932 9222
rect 3956 9220 4012 9222
rect 4036 9220 4092 9222
rect 3796 8186 3852 8188
rect 3876 8186 3932 8188
rect 3956 8186 4012 8188
rect 4036 8186 4092 8188
rect 3796 8134 3842 8186
rect 3842 8134 3852 8186
rect 3876 8134 3906 8186
rect 3906 8134 3918 8186
rect 3918 8134 3932 8186
rect 3956 8134 3970 8186
rect 3970 8134 3982 8186
rect 3982 8134 4012 8186
rect 4036 8134 4046 8186
rect 4046 8134 4092 8186
rect 3796 8132 3852 8134
rect 3876 8132 3932 8134
rect 3956 8132 4012 8134
rect 4036 8132 4092 8134
rect 3796 7098 3852 7100
rect 3876 7098 3932 7100
rect 3956 7098 4012 7100
rect 4036 7098 4092 7100
rect 3796 7046 3842 7098
rect 3842 7046 3852 7098
rect 3876 7046 3906 7098
rect 3906 7046 3918 7098
rect 3918 7046 3932 7098
rect 3956 7046 3970 7098
rect 3970 7046 3982 7098
rect 3982 7046 4012 7098
rect 4036 7046 4046 7098
rect 4046 7046 4092 7098
rect 3796 7044 3852 7046
rect 3876 7044 3932 7046
rect 3956 7044 4012 7046
rect 4036 7044 4092 7046
rect 3796 6010 3852 6012
rect 3876 6010 3932 6012
rect 3956 6010 4012 6012
rect 4036 6010 4092 6012
rect 3796 5958 3842 6010
rect 3842 5958 3852 6010
rect 3876 5958 3906 6010
rect 3906 5958 3918 6010
rect 3918 5958 3932 6010
rect 3956 5958 3970 6010
rect 3970 5958 3982 6010
rect 3982 5958 4012 6010
rect 4036 5958 4046 6010
rect 4046 5958 4092 6010
rect 3796 5956 3852 5958
rect 3876 5956 3932 5958
rect 3956 5956 4012 5958
rect 4036 5956 4092 5958
rect 3796 4922 3852 4924
rect 3876 4922 3932 4924
rect 3956 4922 4012 4924
rect 4036 4922 4092 4924
rect 3796 4870 3842 4922
rect 3842 4870 3852 4922
rect 3876 4870 3906 4922
rect 3906 4870 3918 4922
rect 3918 4870 3932 4922
rect 3956 4870 3970 4922
rect 3970 4870 3982 4922
rect 3982 4870 4012 4922
rect 4036 4870 4046 4922
rect 4046 4870 4092 4922
rect 3796 4868 3852 4870
rect 3876 4868 3932 4870
rect 3956 4868 4012 4870
rect 4036 4868 4092 4870
rect 4066 4664 4122 4720
rect 5170 13252 5226 13288
rect 5170 13232 5172 13252
rect 5172 13232 5224 13252
rect 5224 13232 5226 13252
rect 4342 9424 4398 9480
rect 4894 8880 4950 8936
rect 4802 7404 4858 7440
rect 4802 7384 4804 7404
rect 4804 7384 4856 7404
rect 4856 7384 4858 7404
rect 4802 6724 4858 6760
rect 4802 6704 4804 6724
rect 4804 6704 4856 6724
rect 4856 6704 4858 6724
rect 3796 3834 3852 3836
rect 3876 3834 3932 3836
rect 3956 3834 4012 3836
rect 4036 3834 4092 3836
rect 3796 3782 3842 3834
rect 3842 3782 3852 3834
rect 3876 3782 3906 3834
rect 3906 3782 3918 3834
rect 3918 3782 3932 3834
rect 3956 3782 3970 3834
rect 3970 3782 3982 3834
rect 3982 3782 4012 3834
rect 4036 3782 4046 3834
rect 4046 3782 4092 3834
rect 3796 3780 3852 3782
rect 3876 3780 3932 3782
rect 3956 3780 4012 3782
rect 4036 3780 4092 3782
rect 3422 3476 3424 3496
rect 3424 3476 3476 3496
rect 3476 3476 3478 3496
rect 3422 3440 3478 3476
rect 2686 2896 2742 2952
rect 1858 1944 1914 2000
rect 6636 20698 6692 20700
rect 6716 20698 6772 20700
rect 6796 20698 6852 20700
rect 6876 20698 6932 20700
rect 6636 20646 6682 20698
rect 6682 20646 6692 20698
rect 6716 20646 6746 20698
rect 6746 20646 6758 20698
rect 6758 20646 6772 20698
rect 6796 20646 6810 20698
rect 6810 20646 6822 20698
rect 6822 20646 6852 20698
rect 6876 20646 6886 20698
rect 6886 20646 6932 20698
rect 6636 20644 6692 20646
rect 6716 20644 6772 20646
rect 6796 20644 6852 20646
rect 6876 20644 6932 20646
rect 6636 19610 6692 19612
rect 6716 19610 6772 19612
rect 6796 19610 6852 19612
rect 6876 19610 6932 19612
rect 6636 19558 6682 19610
rect 6682 19558 6692 19610
rect 6716 19558 6746 19610
rect 6746 19558 6758 19610
rect 6758 19558 6772 19610
rect 6796 19558 6810 19610
rect 6810 19558 6822 19610
rect 6822 19558 6852 19610
rect 6876 19558 6886 19610
rect 6886 19558 6932 19610
rect 6636 19556 6692 19558
rect 6716 19556 6772 19558
rect 6796 19556 6852 19558
rect 6876 19556 6932 19558
rect 6366 19352 6422 19408
rect 6636 18522 6692 18524
rect 6716 18522 6772 18524
rect 6796 18522 6852 18524
rect 6876 18522 6932 18524
rect 6636 18470 6682 18522
rect 6682 18470 6692 18522
rect 6716 18470 6746 18522
rect 6746 18470 6758 18522
rect 6758 18470 6772 18522
rect 6796 18470 6810 18522
rect 6810 18470 6822 18522
rect 6822 18470 6852 18522
rect 6876 18470 6886 18522
rect 6886 18470 6932 18522
rect 6636 18468 6692 18470
rect 6716 18468 6772 18470
rect 6796 18468 6852 18470
rect 6876 18468 6932 18470
rect 6636 17434 6692 17436
rect 6716 17434 6772 17436
rect 6796 17434 6852 17436
rect 6876 17434 6932 17436
rect 6636 17382 6682 17434
rect 6682 17382 6692 17434
rect 6716 17382 6746 17434
rect 6746 17382 6758 17434
rect 6758 17382 6772 17434
rect 6796 17382 6810 17434
rect 6810 17382 6822 17434
rect 6822 17382 6852 17434
rect 6876 17382 6886 17434
rect 6886 17382 6932 17434
rect 6636 17380 6692 17382
rect 6716 17380 6772 17382
rect 6796 17380 6852 17382
rect 6876 17380 6932 17382
rect 6636 16346 6692 16348
rect 6716 16346 6772 16348
rect 6796 16346 6852 16348
rect 6876 16346 6932 16348
rect 6636 16294 6682 16346
rect 6682 16294 6692 16346
rect 6716 16294 6746 16346
rect 6746 16294 6758 16346
rect 6758 16294 6772 16346
rect 6796 16294 6810 16346
rect 6810 16294 6822 16346
rect 6822 16294 6852 16346
rect 6876 16294 6886 16346
rect 6886 16294 6932 16346
rect 6636 16292 6692 16294
rect 6716 16292 6772 16294
rect 6796 16292 6852 16294
rect 6876 16292 6932 16294
rect 6636 15258 6692 15260
rect 6716 15258 6772 15260
rect 6796 15258 6852 15260
rect 6876 15258 6932 15260
rect 6636 15206 6682 15258
rect 6682 15206 6692 15258
rect 6716 15206 6746 15258
rect 6746 15206 6758 15258
rect 6758 15206 6772 15258
rect 6796 15206 6810 15258
rect 6810 15206 6822 15258
rect 6822 15206 6852 15258
rect 6876 15206 6886 15258
rect 6886 15206 6932 15258
rect 6636 15204 6692 15206
rect 6716 15204 6772 15206
rect 6796 15204 6852 15206
rect 6876 15204 6932 15206
rect 6642 15036 6644 15056
rect 6644 15036 6696 15056
rect 6696 15036 6698 15056
rect 6642 15000 6698 15036
rect 6636 14170 6692 14172
rect 6716 14170 6772 14172
rect 6796 14170 6852 14172
rect 6876 14170 6932 14172
rect 6636 14118 6682 14170
rect 6682 14118 6692 14170
rect 6716 14118 6746 14170
rect 6746 14118 6758 14170
rect 6758 14118 6772 14170
rect 6796 14118 6810 14170
rect 6810 14118 6822 14170
rect 6822 14118 6852 14170
rect 6876 14118 6886 14170
rect 6886 14118 6932 14170
rect 6636 14116 6692 14118
rect 6716 14116 6772 14118
rect 6796 14116 6852 14118
rect 6876 14116 6932 14118
rect 6642 13268 6644 13288
rect 6644 13268 6696 13288
rect 6696 13268 6698 13288
rect 6642 13232 6698 13268
rect 7378 17992 7434 18048
rect 9477 21242 9533 21244
rect 9557 21242 9613 21244
rect 9637 21242 9693 21244
rect 9717 21242 9773 21244
rect 9477 21190 9523 21242
rect 9523 21190 9533 21242
rect 9557 21190 9587 21242
rect 9587 21190 9599 21242
rect 9599 21190 9613 21242
rect 9637 21190 9651 21242
rect 9651 21190 9663 21242
rect 9663 21190 9693 21242
rect 9717 21190 9727 21242
rect 9727 21190 9773 21242
rect 9477 21188 9533 21190
rect 9557 21188 9613 21190
rect 9637 21188 9693 21190
rect 9717 21188 9773 21190
rect 6636 13082 6692 13084
rect 6716 13082 6772 13084
rect 6796 13082 6852 13084
rect 6876 13082 6932 13084
rect 6636 13030 6682 13082
rect 6682 13030 6692 13082
rect 6716 13030 6746 13082
rect 6746 13030 6758 13082
rect 6758 13030 6772 13082
rect 6796 13030 6810 13082
rect 6810 13030 6822 13082
rect 6822 13030 6852 13082
rect 6876 13030 6886 13082
rect 6886 13030 6932 13082
rect 6636 13028 6692 13030
rect 6716 13028 6772 13030
rect 6796 13028 6852 13030
rect 6876 13028 6932 13030
rect 5538 10648 5594 10704
rect 5446 8880 5502 8936
rect 6826 12280 6882 12336
rect 6636 11994 6692 11996
rect 6716 11994 6772 11996
rect 6796 11994 6852 11996
rect 6876 11994 6932 11996
rect 6636 11942 6682 11994
rect 6682 11942 6692 11994
rect 6716 11942 6746 11994
rect 6746 11942 6758 11994
rect 6758 11942 6772 11994
rect 6796 11942 6810 11994
rect 6810 11942 6822 11994
rect 6822 11942 6852 11994
rect 6876 11942 6886 11994
rect 6886 11942 6932 11994
rect 6636 11940 6692 11942
rect 6716 11940 6772 11942
rect 6796 11940 6852 11942
rect 6876 11940 6932 11942
rect 6636 10906 6692 10908
rect 6716 10906 6772 10908
rect 6796 10906 6852 10908
rect 6876 10906 6932 10908
rect 6636 10854 6682 10906
rect 6682 10854 6692 10906
rect 6716 10854 6746 10906
rect 6746 10854 6758 10906
rect 6758 10854 6772 10906
rect 6796 10854 6810 10906
rect 6810 10854 6822 10906
rect 6822 10854 6852 10906
rect 6876 10854 6886 10906
rect 6886 10854 6932 10906
rect 6636 10852 6692 10854
rect 6716 10852 6772 10854
rect 6796 10852 6852 10854
rect 6876 10852 6932 10854
rect 6734 10004 6736 10024
rect 6736 10004 6788 10024
rect 6788 10004 6790 10024
rect 6734 9968 6790 10004
rect 6636 9818 6692 9820
rect 6716 9818 6772 9820
rect 6796 9818 6852 9820
rect 6876 9818 6932 9820
rect 6636 9766 6682 9818
rect 6682 9766 6692 9818
rect 6716 9766 6746 9818
rect 6746 9766 6758 9818
rect 6758 9766 6772 9818
rect 6796 9766 6810 9818
rect 6810 9766 6822 9818
rect 6822 9766 6852 9818
rect 6876 9766 6886 9818
rect 6886 9766 6932 9818
rect 6636 9764 6692 9766
rect 6716 9764 6772 9766
rect 6796 9764 6852 9766
rect 6876 9764 6932 9766
rect 6366 8916 6368 8936
rect 6368 8916 6420 8936
rect 6420 8916 6422 8936
rect 6366 8880 6422 8916
rect 7010 9444 7066 9480
rect 7010 9424 7012 9444
rect 7012 9424 7064 9444
rect 7064 9424 7066 9444
rect 6636 8730 6692 8732
rect 6716 8730 6772 8732
rect 6796 8730 6852 8732
rect 6876 8730 6932 8732
rect 6636 8678 6682 8730
rect 6682 8678 6692 8730
rect 6716 8678 6746 8730
rect 6746 8678 6758 8730
rect 6758 8678 6772 8730
rect 6796 8678 6810 8730
rect 6810 8678 6822 8730
rect 6822 8678 6852 8730
rect 6876 8678 6886 8730
rect 6886 8678 6932 8730
rect 6636 8676 6692 8678
rect 6716 8676 6772 8678
rect 6796 8676 6852 8678
rect 6876 8676 6932 8678
rect 8114 20748 8116 20768
rect 8116 20748 8168 20768
rect 8168 20748 8170 20768
rect 8114 20712 8170 20748
rect 9477 20154 9533 20156
rect 9557 20154 9613 20156
rect 9637 20154 9693 20156
rect 9717 20154 9773 20156
rect 9477 20102 9523 20154
rect 9523 20102 9533 20154
rect 9557 20102 9587 20154
rect 9587 20102 9599 20154
rect 9599 20102 9613 20154
rect 9637 20102 9651 20154
rect 9651 20102 9663 20154
rect 9663 20102 9693 20154
rect 9717 20102 9727 20154
rect 9727 20102 9773 20154
rect 9477 20100 9533 20102
rect 9557 20100 9613 20102
rect 9637 20100 9693 20102
rect 9717 20100 9773 20102
rect 9477 19066 9533 19068
rect 9557 19066 9613 19068
rect 9637 19066 9693 19068
rect 9717 19066 9773 19068
rect 9477 19014 9523 19066
rect 9523 19014 9533 19066
rect 9557 19014 9587 19066
rect 9587 19014 9599 19066
rect 9599 19014 9613 19066
rect 9637 19014 9651 19066
rect 9651 19014 9663 19066
rect 9663 19014 9693 19066
rect 9717 19014 9727 19066
rect 9727 19014 9773 19066
rect 9477 19012 9533 19014
rect 9557 19012 9613 19014
rect 9637 19012 9693 19014
rect 9717 19012 9773 19014
rect 9477 17978 9533 17980
rect 9557 17978 9613 17980
rect 9637 17978 9693 17980
rect 9717 17978 9773 17980
rect 9477 17926 9523 17978
rect 9523 17926 9533 17978
rect 9557 17926 9587 17978
rect 9587 17926 9599 17978
rect 9599 17926 9613 17978
rect 9637 17926 9651 17978
rect 9651 17926 9663 17978
rect 9663 17926 9693 17978
rect 9717 17926 9727 17978
rect 9727 17926 9773 17978
rect 9477 17924 9533 17926
rect 9557 17924 9613 17926
rect 9637 17924 9693 17926
rect 9717 17924 9773 17926
rect 9477 16890 9533 16892
rect 9557 16890 9613 16892
rect 9637 16890 9693 16892
rect 9717 16890 9773 16892
rect 9477 16838 9523 16890
rect 9523 16838 9533 16890
rect 9557 16838 9587 16890
rect 9587 16838 9599 16890
rect 9599 16838 9613 16890
rect 9637 16838 9651 16890
rect 9651 16838 9663 16890
rect 9663 16838 9693 16890
rect 9717 16838 9727 16890
rect 9727 16838 9773 16890
rect 9477 16836 9533 16838
rect 9557 16836 9613 16838
rect 9637 16836 9693 16838
rect 9717 16836 9773 16838
rect 9477 15802 9533 15804
rect 9557 15802 9613 15804
rect 9637 15802 9693 15804
rect 9717 15802 9773 15804
rect 9477 15750 9523 15802
rect 9523 15750 9533 15802
rect 9557 15750 9587 15802
rect 9587 15750 9599 15802
rect 9599 15750 9613 15802
rect 9637 15750 9651 15802
rect 9651 15750 9663 15802
rect 9663 15750 9693 15802
rect 9717 15750 9727 15802
rect 9727 15750 9773 15802
rect 9477 15748 9533 15750
rect 9557 15748 9613 15750
rect 9637 15748 9693 15750
rect 9717 15748 9773 15750
rect 8114 11892 8170 11928
rect 8114 11872 8116 11892
rect 8116 11872 8168 11892
rect 8168 11872 8170 11892
rect 8482 12008 8538 12064
rect 7562 11192 7618 11248
rect 6636 7642 6692 7644
rect 6716 7642 6772 7644
rect 6796 7642 6852 7644
rect 6876 7642 6932 7644
rect 6636 7590 6682 7642
rect 6682 7590 6692 7642
rect 6716 7590 6746 7642
rect 6746 7590 6758 7642
rect 6758 7590 6772 7642
rect 6796 7590 6810 7642
rect 6810 7590 6822 7642
rect 6822 7590 6852 7642
rect 6876 7590 6886 7642
rect 6886 7590 6932 7642
rect 6636 7588 6692 7590
rect 6716 7588 6772 7590
rect 6796 7588 6852 7590
rect 6876 7588 6932 7590
rect 7194 7828 7196 7848
rect 7196 7828 7248 7848
rect 7248 7828 7250 7848
rect 7194 7792 7250 7828
rect 8022 10512 8078 10568
rect 5998 6724 6054 6760
rect 5998 6704 6000 6724
rect 6000 6704 6052 6724
rect 6052 6704 6054 6724
rect 4894 3712 4950 3768
rect 6636 6554 6692 6556
rect 6716 6554 6772 6556
rect 6796 6554 6852 6556
rect 6876 6554 6932 6556
rect 6636 6502 6682 6554
rect 6682 6502 6692 6554
rect 6716 6502 6746 6554
rect 6746 6502 6758 6554
rect 6758 6502 6772 6554
rect 6796 6502 6810 6554
rect 6810 6502 6822 6554
rect 6822 6502 6852 6554
rect 6876 6502 6886 6554
rect 6886 6502 6932 6554
rect 6636 6500 6692 6502
rect 6716 6500 6772 6502
rect 6796 6500 6852 6502
rect 6876 6500 6932 6502
rect 5906 4120 5962 4176
rect 5814 3440 5870 3496
rect 3796 2746 3852 2748
rect 3876 2746 3932 2748
rect 3956 2746 4012 2748
rect 4036 2746 4092 2748
rect 3796 2694 3842 2746
rect 3842 2694 3852 2746
rect 3876 2694 3906 2746
rect 3906 2694 3918 2746
rect 3918 2694 3932 2746
rect 3956 2694 3970 2746
rect 3970 2694 3982 2746
rect 3982 2694 4012 2746
rect 4036 2694 4046 2746
rect 4046 2694 4092 2746
rect 3796 2692 3852 2694
rect 3876 2692 3932 2694
rect 3956 2692 4012 2694
rect 4036 2692 4092 2694
rect 5078 2624 5134 2680
rect 4250 2488 4306 2544
rect 6636 5466 6692 5468
rect 6716 5466 6772 5468
rect 6796 5466 6852 5468
rect 6876 5466 6932 5468
rect 6636 5414 6682 5466
rect 6682 5414 6692 5466
rect 6716 5414 6746 5466
rect 6746 5414 6758 5466
rect 6758 5414 6772 5466
rect 6796 5414 6810 5466
rect 6810 5414 6822 5466
rect 6822 5414 6852 5466
rect 6876 5414 6886 5466
rect 6886 5414 6932 5466
rect 6636 5412 6692 5414
rect 6716 5412 6772 5414
rect 6796 5412 6852 5414
rect 6876 5412 6932 5414
rect 7654 8336 7710 8392
rect 7838 9324 7840 9344
rect 7840 9324 7892 9344
rect 7892 9324 7894 9344
rect 7838 9288 7894 9324
rect 6636 4378 6692 4380
rect 6716 4378 6772 4380
rect 6796 4378 6852 4380
rect 6876 4378 6932 4380
rect 6636 4326 6682 4378
rect 6682 4326 6692 4378
rect 6716 4326 6746 4378
rect 6746 4326 6758 4378
rect 6758 4326 6772 4378
rect 6796 4326 6810 4378
rect 6810 4326 6822 4378
rect 6822 4326 6852 4378
rect 6876 4326 6886 4378
rect 6886 4326 6932 4378
rect 6636 4324 6692 4326
rect 6716 4324 6772 4326
rect 6796 4324 6852 4326
rect 6876 4324 6932 4326
rect 7286 3712 7342 3768
rect 6636 3290 6692 3292
rect 6716 3290 6772 3292
rect 6796 3290 6852 3292
rect 6876 3290 6932 3292
rect 6636 3238 6682 3290
rect 6682 3238 6692 3290
rect 6716 3238 6746 3290
rect 6746 3238 6758 3290
rect 6758 3238 6772 3290
rect 6796 3238 6810 3290
rect 6810 3238 6822 3290
rect 6822 3238 6852 3290
rect 6876 3238 6886 3290
rect 6886 3238 6932 3290
rect 6636 3236 6692 3238
rect 6716 3236 6772 3238
rect 6796 3236 6852 3238
rect 6876 3236 6932 3238
rect 8482 10004 8484 10024
rect 8484 10004 8536 10024
rect 8536 10004 8538 10024
rect 8482 9968 8538 10004
rect 8390 9696 8446 9752
rect 8390 7828 8392 7848
rect 8392 7828 8444 7848
rect 8444 7828 8446 7848
rect 8390 7792 8446 7828
rect 9477 14714 9533 14716
rect 9557 14714 9613 14716
rect 9637 14714 9693 14716
rect 9717 14714 9773 14716
rect 9477 14662 9523 14714
rect 9523 14662 9533 14714
rect 9557 14662 9587 14714
rect 9587 14662 9599 14714
rect 9599 14662 9613 14714
rect 9637 14662 9651 14714
rect 9651 14662 9663 14714
rect 9663 14662 9693 14714
rect 9717 14662 9727 14714
rect 9727 14662 9773 14714
rect 9477 14660 9533 14662
rect 9557 14660 9613 14662
rect 9637 14660 9693 14662
rect 9717 14660 9773 14662
rect 9477 13626 9533 13628
rect 9557 13626 9613 13628
rect 9637 13626 9693 13628
rect 9717 13626 9773 13628
rect 9477 13574 9523 13626
rect 9523 13574 9533 13626
rect 9557 13574 9587 13626
rect 9587 13574 9599 13626
rect 9599 13574 9613 13626
rect 9637 13574 9651 13626
rect 9651 13574 9663 13626
rect 9663 13574 9693 13626
rect 9717 13574 9727 13626
rect 9727 13574 9773 13626
rect 9477 13572 9533 13574
rect 9557 13572 9613 13574
rect 9637 13572 9693 13574
rect 9717 13572 9773 13574
rect 9477 12538 9533 12540
rect 9557 12538 9613 12540
rect 9637 12538 9693 12540
rect 9717 12538 9773 12540
rect 9477 12486 9523 12538
rect 9523 12486 9533 12538
rect 9557 12486 9587 12538
rect 9587 12486 9599 12538
rect 9599 12486 9613 12538
rect 9637 12486 9651 12538
rect 9651 12486 9663 12538
rect 9663 12486 9693 12538
rect 9717 12486 9727 12538
rect 9727 12486 9773 12538
rect 9477 12484 9533 12486
rect 9557 12484 9613 12486
rect 9637 12484 9693 12486
rect 9717 12484 9773 12486
rect 8758 10668 8814 10704
rect 8758 10648 8760 10668
rect 8760 10648 8812 10668
rect 8812 10648 8814 10668
rect 3422 2388 3424 2408
rect 3424 2388 3476 2408
rect 3476 2388 3478 2408
rect 3422 2352 3478 2388
rect 6636 2202 6692 2204
rect 6716 2202 6772 2204
rect 6796 2202 6852 2204
rect 6876 2202 6932 2204
rect 6636 2150 6682 2202
rect 6682 2150 6692 2202
rect 6716 2150 6746 2202
rect 6746 2150 6758 2202
rect 6758 2150 6772 2202
rect 6796 2150 6810 2202
rect 6810 2150 6822 2202
rect 6822 2150 6852 2202
rect 6876 2150 6886 2202
rect 6886 2150 6932 2202
rect 6636 2148 6692 2150
rect 6716 2148 6772 2150
rect 6796 2148 6852 2150
rect 6876 2148 6932 2150
rect 7654 2896 7710 2952
rect 7838 2644 7894 2680
rect 7838 2624 7840 2644
rect 7840 2624 7892 2644
rect 7892 2624 7894 2644
rect 8298 2896 8354 2952
rect 9770 12008 9826 12064
rect 9477 11450 9533 11452
rect 9557 11450 9613 11452
rect 9637 11450 9693 11452
rect 9717 11450 9773 11452
rect 9477 11398 9523 11450
rect 9523 11398 9533 11450
rect 9557 11398 9587 11450
rect 9587 11398 9599 11450
rect 9599 11398 9613 11450
rect 9637 11398 9651 11450
rect 9651 11398 9663 11450
rect 9663 11398 9693 11450
rect 9717 11398 9727 11450
rect 9727 11398 9773 11450
rect 9477 11396 9533 11398
rect 9557 11396 9613 11398
rect 9637 11396 9693 11398
rect 9717 11396 9773 11398
rect 9402 10668 9458 10704
rect 9402 10648 9404 10668
rect 9404 10648 9456 10668
rect 9456 10648 9458 10668
rect 9477 10362 9533 10364
rect 9557 10362 9613 10364
rect 9637 10362 9693 10364
rect 9717 10362 9773 10364
rect 9477 10310 9523 10362
rect 9523 10310 9533 10362
rect 9557 10310 9587 10362
rect 9587 10310 9599 10362
rect 9599 10310 9613 10362
rect 9637 10310 9651 10362
rect 9651 10310 9663 10362
rect 9663 10310 9693 10362
rect 9717 10310 9727 10362
rect 9727 10310 9773 10362
rect 9477 10308 9533 10310
rect 9557 10308 9613 10310
rect 9637 10308 9693 10310
rect 9717 10308 9773 10310
rect 9494 10104 9550 10160
rect 9310 9696 9366 9752
rect 9477 9274 9533 9276
rect 9557 9274 9613 9276
rect 9637 9274 9693 9276
rect 9717 9274 9773 9276
rect 9477 9222 9523 9274
rect 9523 9222 9533 9274
rect 9557 9222 9587 9274
rect 9587 9222 9599 9274
rect 9599 9222 9613 9274
rect 9637 9222 9651 9274
rect 9651 9222 9663 9274
rect 9663 9222 9693 9274
rect 9717 9222 9727 9274
rect 9727 9222 9773 9274
rect 9477 9220 9533 9222
rect 9557 9220 9613 9222
rect 9637 9220 9693 9222
rect 9717 9220 9773 9222
rect 10138 9152 10194 9208
rect 9862 8744 9918 8800
rect 9477 8186 9533 8188
rect 9557 8186 9613 8188
rect 9637 8186 9693 8188
rect 9717 8186 9773 8188
rect 9477 8134 9523 8186
rect 9523 8134 9533 8186
rect 9557 8134 9587 8186
rect 9587 8134 9599 8186
rect 9599 8134 9613 8186
rect 9637 8134 9651 8186
rect 9651 8134 9663 8186
rect 9663 8134 9693 8186
rect 9717 8134 9727 8186
rect 9727 8134 9773 8186
rect 9477 8132 9533 8134
rect 9557 8132 9613 8134
rect 9637 8132 9693 8134
rect 9717 8132 9773 8134
rect 9477 7098 9533 7100
rect 9557 7098 9613 7100
rect 9637 7098 9693 7100
rect 9717 7098 9773 7100
rect 9477 7046 9523 7098
rect 9523 7046 9533 7098
rect 9557 7046 9587 7098
rect 9587 7046 9599 7098
rect 9599 7046 9613 7098
rect 9637 7046 9651 7098
rect 9651 7046 9663 7098
rect 9663 7046 9693 7098
rect 9717 7046 9727 7098
rect 9727 7046 9773 7098
rect 9477 7044 9533 7046
rect 9557 7044 9613 7046
rect 9637 7044 9693 7046
rect 9717 7044 9773 7046
rect 9477 6010 9533 6012
rect 9557 6010 9613 6012
rect 9637 6010 9693 6012
rect 9717 6010 9773 6012
rect 9477 5958 9523 6010
rect 9523 5958 9533 6010
rect 9557 5958 9587 6010
rect 9587 5958 9599 6010
rect 9599 5958 9613 6010
rect 9637 5958 9651 6010
rect 9651 5958 9663 6010
rect 9663 5958 9693 6010
rect 9717 5958 9727 6010
rect 9727 5958 9773 6010
rect 9477 5956 9533 5958
rect 9557 5956 9613 5958
rect 9637 5956 9693 5958
rect 9717 5956 9773 5958
rect 9494 5752 9550 5808
rect 8206 2352 8262 2408
rect 9477 4922 9533 4924
rect 9557 4922 9613 4924
rect 9637 4922 9693 4924
rect 9717 4922 9773 4924
rect 9477 4870 9523 4922
rect 9523 4870 9533 4922
rect 9557 4870 9587 4922
rect 9587 4870 9599 4922
rect 9599 4870 9613 4922
rect 9637 4870 9651 4922
rect 9651 4870 9663 4922
rect 9663 4870 9693 4922
rect 9717 4870 9727 4922
rect 9727 4870 9773 4922
rect 9477 4868 9533 4870
rect 9557 4868 9613 4870
rect 9637 4868 9693 4870
rect 9717 4868 9773 4870
rect 10322 8744 10378 8800
rect 12317 21786 12373 21788
rect 12397 21786 12453 21788
rect 12477 21786 12533 21788
rect 12557 21786 12613 21788
rect 12317 21734 12363 21786
rect 12363 21734 12373 21786
rect 12397 21734 12427 21786
rect 12427 21734 12439 21786
rect 12439 21734 12453 21786
rect 12477 21734 12491 21786
rect 12491 21734 12503 21786
rect 12503 21734 12533 21786
rect 12557 21734 12567 21786
rect 12567 21734 12613 21786
rect 12317 21732 12373 21734
rect 12397 21732 12453 21734
rect 12477 21732 12533 21734
rect 12557 21732 12613 21734
rect 12317 20698 12373 20700
rect 12397 20698 12453 20700
rect 12477 20698 12533 20700
rect 12557 20698 12613 20700
rect 12317 20646 12363 20698
rect 12363 20646 12373 20698
rect 12397 20646 12427 20698
rect 12427 20646 12439 20698
rect 12439 20646 12453 20698
rect 12477 20646 12491 20698
rect 12491 20646 12503 20698
rect 12503 20646 12533 20698
rect 12557 20646 12567 20698
rect 12567 20646 12613 20698
rect 12317 20644 12373 20646
rect 12397 20644 12453 20646
rect 12477 20644 12533 20646
rect 12557 20644 12613 20646
rect 12317 19610 12373 19612
rect 12397 19610 12453 19612
rect 12477 19610 12533 19612
rect 12557 19610 12613 19612
rect 12317 19558 12363 19610
rect 12363 19558 12373 19610
rect 12397 19558 12427 19610
rect 12427 19558 12439 19610
rect 12439 19558 12453 19610
rect 12477 19558 12491 19610
rect 12491 19558 12503 19610
rect 12503 19558 12533 19610
rect 12557 19558 12567 19610
rect 12567 19558 12613 19610
rect 12317 19556 12373 19558
rect 12397 19556 12453 19558
rect 12477 19556 12533 19558
rect 12557 19556 12613 19558
rect 10966 9696 11022 9752
rect 12317 18522 12373 18524
rect 12397 18522 12453 18524
rect 12477 18522 12533 18524
rect 12557 18522 12613 18524
rect 12317 18470 12363 18522
rect 12363 18470 12373 18522
rect 12397 18470 12427 18522
rect 12427 18470 12439 18522
rect 12439 18470 12453 18522
rect 12477 18470 12491 18522
rect 12491 18470 12503 18522
rect 12503 18470 12533 18522
rect 12557 18470 12567 18522
rect 12567 18470 12613 18522
rect 12317 18468 12373 18470
rect 12397 18468 12453 18470
rect 12477 18468 12533 18470
rect 12557 18468 12613 18470
rect 12317 17434 12373 17436
rect 12397 17434 12453 17436
rect 12477 17434 12533 17436
rect 12557 17434 12613 17436
rect 12317 17382 12363 17434
rect 12363 17382 12373 17434
rect 12397 17382 12427 17434
rect 12427 17382 12439 17434
rect 12439 17382 12453 17434
rect 12477 17382 12491 17434
rect 12491 17382 12503 17434
rect 12503 17382 12533 17434
rect 12557 17382 12567 17434
rect 12567 17382 12613 17434
rect 12317 17380 12373 17382
rect 12397 17380 12453 17382
rect 12477 17380 12533 17382
rect 12557 17380 12613 17382
rect 12317 16346 12373 16348
rect 12397 16346 12453 16348
rect 12477 16346 12533 16348
rect 12557 16346 12613 16348
rect 12317 16294 12363 16346
rect 12363 16294 12373 16346
rect 12397 16294 12427 16346
rect 12427 16294 12439 16346
rect 12439 16294 12453 16346
rect 12477 16294 12491 16346
rect 12491 16294 12503 16346
rect 12503 16294 12533 16346
rect 12557 16294 12567 16346
rect 12567 16294 12613 16346
rect 12317 16292 12373 16294
rect 12397 16292 12453 16294
rect 12477 16292 12533 16294
rect 12557 16292 12613 16294
rect 12317 15258 12373 15260
rect 12397 15258 12453 15260
rect 12477 15258 12533 15260
rect 12557 15258 12613 15260
rect 12317 15206 12363 15258
rect 12363 15206 12373 15258
rect 12397 15206 12427 15258
rect 12427 15206 12439 15258
rect 12439 15206 12453 15258
rect 12477 15206 12491 15258
rect 12491 15206 12503 15258
rect 12503 15206 12533 15258
rect 12557 15206 12567 15258
rect 12567 15206 12613 15258
rect 12317 15204 12373 15206
rect 12397 15204 12453 15206
rect 12477 15204 12533 15206
rect 12557 15204 12613 15206
rect 12317 14170 12373 14172
rect 12397 14170 12453 14172
rect 12477 14170 12533 14172
rect 12557 14170 12613 14172
rect 12317 14118 12363 14170
rect 12363 14118 12373 14170
rect 12397 14118 12427 14170
rect 12427 14118 12439 14170
rect 12439 14118 12453 14170
rect 12477 14118 12491 14170
rect 12491 14118 12503 14170
rect 12503 14118 12533 14170
rect 12557 14118 12567 14170
rect 12567 14118 12613 14170
rect 12317 14116 12373 14118
rect 12397 14116 12453 14118
rect 12477 14116 12533 14118
rect 12557 14116 12613 14118
rect 17998 21786 18054 21788
rect 18078 21786 18134 21788
rect 18158 21786 18214 21788
rect 18238 21786 18294 21788
rect 17998 21734 18044 21786
rect 18044 21734 18054 21786
rect 18078 21734 18108 21786
rect 18108 21734 18120 21786
rect 18120 21734 18134 21786
rect 18158 21734 18172 21786
rect 18172 21734 18184 21786
rect 18184 21734 18214 21786
rect 18238 21734 18248 21786
rect 18248 21734 18294 21786
rect 17998 21732 18054 21734
rect 18078 21732 18134 21734
rect 18158 21732 18214 21734
rect 18238 21732 18294 21734
rect 23679 21786 23735 21788
rect 23759 21786 23815 21788
rect 23839 21786 23895 21788
rect 23919 21786 23975 21788
rect 23679 21734 23725 21786
rect 23725 21734 23735 21786
rect 23759 21734 23789 21786
rect 23789 21734 23801 21786
rect 23801 21734 23815 21786
rect 23839 21734 23853 21786
rect 23853 21734 23865 21786
rect 23865 21734 23895 21786
rect 23919 21734 23929 21786
rect 23929 21734 23975 21786
rect 23679 21732 23735 21734
rect 23759 21732 23815 21734
rect 23839 21732 23895 21734
rect 23919 21732 23975 21734
rect 15158 21242 15214 21244
rect 15238 21242 15294 21244
rect 15318 21242 15374 21244
rect 15398 21242 15454 21244
rect 15158 21190 15204 21242
rect 15204 21190 15214 21242
rect 15238 21190 15268 21242
rect 15268 21190 15280 21242
rect 15280 21190 15294 21242
rect 15318 21190 15332 21242
rect 15332 21190 15344 21242
rect 15344 21190 15374 21242
rect 15398 21190 15408 21242
rect 15408 21190 15454 21242
rect 15158 21188 15214 21190
rect 15238 21188 15294 21190
rect 15318 21188 15374 21190
rect 15398 21188 15454 21190
rect 20839 21242 20895 21244
rect 20919 21242 20975 21244
rect 20999 21242 21055 21244
rect 21079 21242 21135 21244
rect 20839 21190 20885 21242
rect 20885 21190 20895 21242
rect 20919 21190 20949 21242
rect 20949 21190 20961 21242
rect 20961 21190 20975 21242
rect 20999 21190 21013 21242
rect 21013 21190 21025 21242
rect 21025 21190 21055 21242
rect 21079 21190 21089 21242
rect 21089 21190 21135 21242
rect 20839 21188 20895 21190
rect 20919 21188 20975 21190
rect 20999 21188 21055 21190
rect 21079 21188 21135 21190
rect 17998 20698 18054 20700
rect 18078 20698 18134 20700
rect 18158 20698 18214 20700
rect 18238 20698 18294 20700
rect 17998 20646 18044 20698
rect 18044 20646 18054 20698
rect 18078 20646 18108 20698
rect 18108 20646 18120 20698
rect 18120 20646 18134 20698
rect 18158 20646 18172 20698
rect 18172 20646 18184 20698
rect 18184 20646 18214 20698
rect 18238 20646 18248 20698
rect 18248 20646 18294 20698
rect 17998 20644 18054 20646
rect 18078 20644 18134 20646
rect 18158 20644 18214 20646
rect 18238 20644 18294 20646
rect 23679 20698 23735 20700
rect 23759 20698 23815 20700
rect 23839 20698 23895 20700
rect 23919 20698 23975 20700
rect 23679 20646 23725 20698
rect 23725 20646 23735 20698
rect 23759 20646 23789 20698
rect 23789 20646 23801 20698
rect 23801 20646 23815 20698
rect 23839 20646 23853 20698
rect 23853 20646 23865 20698
rect 23865 20646 23895 20698
rect 23919 20646 23929 20698
rect 23929 20646 23975 20698
rect 23679 20644 23735 20646
rect 23759 20644 23815 20646
rect 23839 20644 23895 20646
rect 23919 20644 23975 20646
rect 15158 20154 15214 20156
rect 15238 20154 15294 20156
rect 15318 20154 15374 20156
rect 15398 20154 15454 20156
rect 15158 20102 15204 20154
rect 15204 20102 15214 20154
rect 15238 20102 15268 20154
rect 15268 20102 15280 20154
rect 15280 20102 15294 20154
rect 15318 20102 15332 20154
rect 15332 20102 15344 20154
rect 15344 20102 15374 20154
rect 15398 20102 15408 20154
rect 15408 20102 15454 20154
rect 15158 20100 15214 20102
rect 15238 20100 15294 20102
rect 15318 20100 15374 20102
rect 15398 20100 15454 20102
rect 20839 20154 20895 20156
rect 20919 20154 20975 20156
rect 20999 20154 21055 20156
rect 21079 20154 21135 20156
rect 20839 20102 20885 20154
rect 20885 20102 20895 20154
rect 20919 20102 20949 20154
rect 20949 20102 20961 20154
rect 20961 20102 20975 20154
rect 20999 20102 21013 20154
rect 21013 20102 21025 20154
rect 21025 20102 21055 20154
rect 21079 20102 21089 20154
rect 21089 20102 21135 20154
rect 20839 20100 20895 20102
rect 20919 20100 20975 20102
rect 20999 20100 21055 20102
rect 21079 20100 21135 20102
rect 17998 19610 18054 19612
rect 18078 19610 18134 19612
rect 18158 19610 18214 19612
rect 18238 19610 18294 19612
rect 17998 19558 18044 19610
rect 18044 19558 18054 19610
rect 18078 19558 18108 19610
rect 18108 19558 18120 19610
rect 18120 19558 18134 19610
rect 18158 19558 18172 19610
rect 18172 19558 18184 19610
rect 18184 19558 18214 19610
rect 18238 19558 18248 19610
rect 18248 19558 18294 19610
rect 17998 19556 18054 19558
rect 18078 19556 18134 19558
rect 18158 19556 18214 19558
rect 18238 19556 18294 19558
rect 15158 19066 15214 19068
rect 15238 19066 15294 19068
rect 15318 19066 15374 19068
rect 15398 19066 15454 19068
rect 15158 19014 15204 19066
rect 15204 19014 15214 19066
rect 15238 19014 15268 19066
rect 15268 19014 15280 19066
rect 15280 19014 15294 19066
rect 15318 19014 15332 19066
rect 15332 19014 15344 19066
rect 15344 19014 15374 19066
rect 15398 19014 15408 19066
rect 15408 19014 15454 19066
rect 15158 19012 15214 19014
rect 15238 19012 15294 19014
rect 15318 19012 15374 19014
rect 15398 19012 15454 19014
rect 23679 19610 23735 19612
rect 23759 19610 23815 19612
rect 23839 19610 23895 19612
rect 23919 19610 23975 19612
rect 23679 19558 23725 19610
rect 23725 19558 23735 19610
rect 23759 19558 23789 19610
rect 23789 19558 23801 19610
rect 23801 19558 23815 19610
rect 23839 19558 23853 19610
rect 23853 19558 23865 19610
rect 23865 19558 23895 19610
rect 23919 19558 23929 19610
rect 23929 19558 23975 19610
rect 23679 19556 23735 19558
rect 23759 19556 23815 19558
rect 23839 19556 23895 19558
rect 23919 19556 23975 19558
rect 20839 19066 20895 19068
rect 20919 19066 20975 19068
rect 20999 19066 21055 19068
rect 21079 19066 21135 19068
rect 20839 19014 20885 19066
rect 20885 19014 20895 19066
rect 20919 19014 20949 19066
rect 20949 19014 20961 19066
rect 20961 19014 20975 19066
rect 20999 19014 21013 19066
rect 21013 19014 21025 19066
rect 21025 19014 21055 19066
rect 21079 19014 21089 19066
rect 21089 19014 21135 19066
rect 20839 19012 20895 19014
rect 20919 19012 20975 19014
rect 20999 19012 21055 19014
rect 21079 19012 21135 19014
rect 17998 18522 18054 18524
rect 18078 18522 18134 18524
rect 18158 18522 18214 18524
rect 18238 18522 18294 18524
rect 17998 18470 18044 18522
rect 18044 18470 18054 18522
rect 18078 18470 18108 18522
rect 18108 18470 18120 18522
rect 18120 18470 18134 18522
rect 18158 18470 18172 18522
rect 18172 18470 18184 18522
rect 18184 18470 18214 18522
rect 18238 18470 18248 18522
rect 18248 18470 18294 18522
rect 17998 18468 18054 18470
rect 18078 18468 18134 18470
rect 18158 18468 18214 18470
rect 18238 18468 18294 18470
rect 15158 17978 15214 17980
rect 15238 17978 15294 17980
rect 15318 17978 15374 17980
rect 15398 17978 15454 17980
rect 15158 17926 15204 17978
rect 15204 17926 15214 17978
rect 15238 17926 15268 17978
rect 15268 17926 15280 17978
rect 15280 17926 15294 17978
rect 15318 17926 15332 17978
rect 15332 17926 15344 17978
rect 15344 17926 15374 17978
rect 15398 17926 15408 17978
rect 15408 17926 15454 17978
rect 15158 17924 15214 17926
rect 15238 17924 15294 17926
rect 15318 17924 15374 17926
rect 15398 17924 15454 17926
rect 9477 3834 9533 3836
rect 9557 3834 9613 3836
rect 9637 3834 9693 3836
rect 9717 3834 9773 3836
rect 9477 3782 9523 3834
rect 9523 3782 9533 3834
rect 9557 3782 9587 3834
rect 9587 3782 9599 3834
rect 9599 3782 9613 3834
rect 9637 3782 9651 3834
rect 9651 3782 9663 3834
rect 9663 3782 9693 3834
rect 9717 3782 9727 3834
rect 9727 3782 9773 3834
rect 9477 3780 9533 3782
rect 9557 3780 9613 3782
rect 9637 3780 9693 3782
rect 9717 3780 9773 3782
rect 11242 9424 11298 9480
rect 11426 8916 11428 8936
rect 11428 8916 11480 8936
rect 11480 8916 11482 8936
rect 11426 8880 11482 8916
rect 12070 12180 12072 12200
rect 12072 12180 12124 12200
rect 12124 12180 12126 12200
rect 12070 12144 12126 12180
rect 12317 13082 12373 13084
rect 12397 13082 12453 13084
rect 12477 13082 12533 13084
rect 12557 13082 12613 13084
rect 12317 13030 12363 13082
rect 12363 13030 12373 13082
rect 12397 13030 12427 13082
rect 12427 13030 12439 13082
rect 12439 13030 12453 13082
rect 12477 13030 12491 13082
rect 12491 13030 12503 13082
rect 12503 13030 12533 13082
rect 12557 13030 12567 13082
rect 12567 13030 12613 13082
rect 12317 13028 12373 13030
rect 12397 13028 12453 13030
rect 12477 13028 12533 13030
rect 12557 13028 12613 13030
rect 12898 12416 12954 12472
rect 12317 11994 12373 11996
rect 12397 11994 12453 11996
rect 12477 11994 12533 11996
rect 12557 11994 12613 11996
rect 12317 11942 12363 11994
rect 12363 11942 12373 11994
rect 12397 11942 12427 11994
rect 12427 11942 12439 11994
rect 12439 11942 12453 11994
rect 12477 11942 12491 11994
rect 12491 11942 12503 11994
rect 12503 11942 12533 11994
rect 12557 11942 12567 11994
rect 12567 11942 12613 11994
rect 12317 11940 12373 11942
rect 12397 11940 12453 11942
rect 12477 11940 12533 11942
rect 12557 11940 12613 11942
rect 12317 10906 12373 10908
rect 12397 10906 12453 10908
rect 12477 10906 12533 10908
rect 12557 10906 12613 10908
rect 12317 10854 12363 10906
rect 12363 10854 12373 10906
rect 12397 10854 12427 10906
rect 12427 10854 12439 10906
rect 12439 10854 12453 10906
rect 12477 10854 12491 10906
rect 12491 10854 12503 10906
rect 12503 10854 12533 10906
rect 12557 10854 12567 10906
rect 12567 10854 12613 10906
rect 12317 10852 12373 10854
rect 12397 10852 12453 10854
rect 12477 10852 12533 10854
rect 12557 10852 12613 10854
rect 12622 10124 12678 10160
rect 12622 10104 12624 10124
rect 12624 10104 12676 10124
rect 12676 10104 12678 10124
rect 12317 9818 12373 9820
rect 12397 9818 12453 9820
rect 12477 9818 12533 9820
rect 12557 9818 12613 9820
rect 12317 9766 12363 9818
rect 12363 9766 12373 9818
rect 12397 9766 12427 9818
rect 12427 9766 12439 9818
rect 12439 9766 12453 9818
rect 12477 9766 12491 9818
rect 12491 9766 12503 9818
rect 12503 9766 12533 9818
rect 12557 9766 12567 9818
rect 12567 9766 12613 9818
rect 12317 9764 12373 9766
rect 12397 9764 12453 9766
rect 12477 9764 12533 9766
rect 12557 9764 12613 9766
rect 12070 9424 12126 9480
rect 12438 9580 12494 9616
rect 12438 9560 12440 9580
rect 12440 9560 12492 9580
rect 12492 9560 12494 9580
rect 12898 9832 12954 9888
rect 12317 8730 12373 8732
rect 12397 8730 12453 8732
rect 12477 8730 12533 8732
rect 12557 8730 12613 8732
rect 12317 8678 12363 8730
rect 12363 8678 12373 8730
rect 12397 8678 12427 8730
rect 12427 8678 12439 8730
rect 12439 8678 12453 8730
rect 12477 8678 12491 8730
rect 12491 8678 12503 8730
rect 12503 8678 12533 8730
rect 12557 8678 12567 8730
rect 12567 8678 12613 8730
rect 12317 8676 12373 8678
rect 12397 8676 12453 8678
rect 12477 8676 12533 8678
rect 12557 8676 12613 8678
rect 11886 8508 11888 8528
rect 11888 8508 11940 8528
rect 11940 8508 11942 8528
rect 11886 8472 11942 8508
rect 9477 2746 9533 2748
rect 9557 2746 9613 2748
rect 9637 2746 9693 2748
rect 9717 2746 9773 2748
rect 9477 2694 9523 2746
rect 9523 2694 9533 2746
rect 9557 2694 9587 2746
rect 9587 2694 9599 2746
rect 9599 2694 9613 2746
rect 9637 2694 9651 2746
rect 9651 2694 9663 2746
rect 9663 2694 9693 2746
rect 9717 2694 9727 2746
rect 9727 2694 9773 2746
rect 9477 2692 9533 2694
rect 9557 2692 9613 2694
rect 9637 2692 9693 2694
rect 9717 2692 9773 2694
rect 12317 7642 12373 7644
rect 12397 7642 12453 7644
rect 12477 7642 12533 7644
rect 12557 7642 12613 7644
rect 12317 7590 12363 7642
rect 12363 7590 12373 7642
rect 12397 7590 12427 7642
rect 12427 7590 12439 7642
rect 12439 7590 12453 7642
rect 12477 7590 12491 7642
rect 12491 7590 12503 7642
rect 12503 7590 12533 7642
rect 12557 7590 12567 7642
rect 12567 7590 12613 7642
rect 12317 7588 12373 7590
rect 12397 7588 12453 7590
rect 12477 7588 12533 7590
rect 12557 7588 12613 7590
rect 15158 16890 15214 16892
rect 15238 16890 15294 16892
rect 15318 16890 15374 16892
rect 15398 16890 15454 16892
rect 15158 16838 15204 16890
rect 15204 16838 15214 16890
rect 15238 16838 15268 16890
rect 15268 16838 15280 16890
rect 15280 16838 15294 16890
rect 15318 16838 15332 16890
rect 15332 16838 15344 16890
rect 15344 16838 15374 16890
rect 15398 16838 15408 16890
rect 15408 16838 15454 16890
rect 15158 16836 15214 16838
rect 15238 16836 15294 16838
rect 15318 16836 15374 16838
rect 15398 16836 15454 16838
rect 15158 15802 15214 15804
rect 15238 15802 15294 15804
rect 15318 15802 15374 15804
rect 15398 15802 15454 15804
rect 15158 15750 15204 15802
rect 15204 15750 15214 15802
rect 15238 15750 15268 15802
rect 15268 15750 15280 15802
rect 15280 15750 15294 15802
rect 15318 15750 15332 15802
rect 15332 15750 15344 15802
rect 15344 15750 15374 15802
rect 15398 15750 15408 15802
rect 15408 15750 15454 15802
rect 15158 15748 15214 15750
rect 15238 15748 15294 15750
rect 15318 15748 15374 15750
rect 15398 15748 15454 15750
rect 13082 7656 13138 7712
rect 12317 6554 12373 6556
rect 12397 6554 12453 6556
rect 12477 6554 12533 6556
rect 12557 6554 12613 6556
rect 12317 6502 12363 6554
rect 12363 6502 12373 6554
rect 12397 6502 12427 6554
rect 12427 6502 12439 6554
rect 12439 6502 12453 6554
rect 12477 6502 12491 6554
rect 12491 6502 12503 6554
rect 12503 6502 12533 6554
rect 12557 6502 12567 6554
rect 12567 6502 12613 6554
rect 12317 6500 12373 6502
rect 12397 6500 12453 6502
rect 12477 6500 12533 6502
rect 12557 6500 12613 6502
rect 13634 8608 13690 8664
rect 14002 8608 14058 8664
rect 13910 8472 13966 8528
rect 15158 14714 15214 14716
rect 15238 14714 15294 14716
rect 15318 14714 15374 14716
rect 15398 14714 15454 14716
rect 15158 14662 15204 14714
rect 15204 14662 15214 14714
rect 15238 14662 15268 14714
rect 15268 14662 15280 14714
rect 15280 14662 15294 14714
rect 15318 14662 15332 14714
rect 15332 14662 15344 14714
rect 15344 14662 15374 14714
rect 15398 14662 15408 14714
rect 15408 14662 15454 14714
rect 15158 14660 15214 14662
rect 15238 14660 15294 14662
rect 15318 14660 15374 14662
rect 15398 14660 15454 14662
rect 15382 13812 15384 13832
rect 15384 13812 15436 13832
rect 15436 13812 15438 13832
rect 15382 13776 15438 13812
rect 15158 13626 15214 13628
rect 15238 13626 15294 13628
rect 15318 13626 15374 13628
rect 15398 13626 15454 13628
rect 15158 13574 15204 13626
rect 15204 13574 15214 13626
rect 15238 13574 15268 13626
rect 15268 13574 15280 13626
rect 15280 13574 15294 13626
rect 15318 13574 15332 13626
rect 15332 13574 15344 13626
rect 15344 13574 15374 13626
rect 15398 13574 15408 13626
rect 15408 13574 15454 13626
rect 15158 13572 15214 13574
rect 15238 13572 15294 13574
rect 15318 13572 15374 13574
rect 15398 13572 15454 13574
rect 14554 12280 14610 12336
rect 14646 12008 14702 12064
rect 14830 11636 14832 11656
rect 14832 11636 14884 11656
rect 14884 11636 14886 11656
rect 14830 11600 14886 11636
rect 14738 11192 14794 11248
rect 14462 9832 14518 9888
rect 14370 9560 14426 9616
rect 14278 8472 14334 8528
rect 14830 11092 14832 11112
rect 14832 11092 14884 11112
rect 14884 11092 14886 11112
rect 14830 11056 14886 11092
rect 14462 9424 14518 9480
rect 14554 9016 14610 9072
rect 14830 9152 14886 9208
rect 15158 12538 15214 12540
rect 15238 12538 15294 12540
rect 15318 12538 15374 12540
rect 15398 12538 15454 12540
rect 15158 12486 15204 12538
rect 15204 12486 15214 12538
rect 15238 12486 15268 12538
rect 15268 12486 15280 12538
rect 15280 12486 15294 12538
rect 15318 12486 15332 12538
rect 15332 12486 15344 12538
rect 15344 12486 15374 12538
rect 15398 12486 15408 12538
rect 15408 12486 15454 12538
rect 15158 12484 15214 12486
rect 15238 12484 15294 12486
rect 15318 12484 15374 12486
rect 15398 12484 15454 12486
rect 15014 12416 15070 12472
rect 15658 12180 15660 12200
rect 15660 12180 15712 12200
rect 15712 12180 15714 12200
rect 15158 11450 15214 11452
rect 15238 11450 15294 11452
rect 15318 11450 15374 11452
rect 15398 11450 15454 11452
rect 15158 11398 15204 11450
rect 15204 11398 15214 11450
rect 15238 11398 15268 11450
rect 15268 11398 15280 11450
rect 15280 11398 15294 11450
rect 15318 11398 15332 11450
rect 15332 11398 15344 11450
rect 15344 11398 15374 11450
rect 15398 11398 15408 11450
rect 15408 11398 15454 11450
rect 15158 11396 15214 11398
rect 15238 11396 15294 11398
rect 15318 11396 15374 11398
rect 15398 11396 15454 11398
rect 15658 12144 15714 12180
rect 15290 10784 15346 10840
rect 15158 10362 15214 10364
rect 15238 10362 15294 10364
rect 15318 10362 15374 10364
rect 15398 10362 15454 10364
rect 15158 10310 15204 10362
rect 15204 10310 15214 10362
rect 15238 10310 15268 10362
rect 15268 10310 15280 10362
rect 15280 10310 15294 10362
rect 15318 10310 15332 10362
rect 15332 10310 15344 10362
rect 15344 10310 15374 10362
rect 15398 10310 15408 10362
rect 15408 10310 15454 10362
rect 15158 10308 15214 10310
rect 15238 10308 15294 10310
rect 15318 10308 15374 10310
rect 15398 10308 15454 10310
rect 15290 9988 15346 10024
rect 15290 9968 15292 9988
rect 15292 9968 15344 9988
rect 15344 9968 15346 9988
rect 15382 9424 15438 9480
rect 15158 9274 15214 9276
rect 15238 9274 15294 9276
rect 15318 9274 15374 9276
rect 15398 9274 15454 9276
rect 15158 9222 15204 9274
rect 15204 9222 15214 9274
rect 15238 9222 15268 9274
rect 15268 9222 15280 9274
rect 15280 9222 15294 9274
rect 15318 9222 15332 9274
rect 15332 9222 15344 9274
rect 15344 9222 15374 9274
rect 15398 9222 15408 9274
rect 15408 9222 15454 9274
rect 15158 9220 15214 9222
rect 15238 9220 15294 9222
rect 15318 9220 15374 9222
rect 15398 9220 15454 9222
rect 14462 8492 14518 8528
rect 14462 8472 14464 8492
rect 14464 8472 14516 8492
rect 14516 8472 14518 8492
rect 14646 7384 14702 7440
rect 13910 6432 13966 6488
rect 12317 5466 12373 5468
rect 12397 5466 12453 5468
rect 12477 5466 12533 5468
rect 12557 5466 12613 5468
rect 12317 5414 12363 5466
rect 12363 5414 12373 5466
rect 12397 5414 12427 5466
rect 12427 5414 12439 5466
rect 12439 5414 12453 5466
rect 12477 5414 12491 5466
rect 12491 5414 12503 5466
rect 12503 5414 12533 5466
rect 12557 5414 12567 5466
rect 12567 5414 12613 5466
rect 12317 5412 12373 5414
rect 12397 5412 12453 5414
rect 12477 5412 12533 5414
rect 12557 5412 12613 5414
rect 11886 4564 11888 4584
rect 11888 4564 11940 4584
rect 11940 4564 11942 4584
rect 11886 4528 11942 4564
rect 12714 4528 12770 4584
rect 12317 4378 12373 4380
rect 12397 4378 12453 4380
rect 12477 4378 12533 4380
rect 12557 4378 12613 4380
rect 12317 4326 12363 4378
rect 12363 4326 12373 4378
rect 12397 4326 12427 4378
rect 12427 4326 12439 4378
rect 12439 4326 12453 4378
rect 12477 4326 12491 4378
rect 12491 4326 12503 4378
rect 12503 4326 12533 4378
rect 12557 4326 12567 4378
rect 12567 4326 12613 4378
rect 12317 4324 12373 4326
rect 12397 4324 12453 4326
rect 12477 4324 12533 4326
rect 12557 4324 12613 4326
rect 17998 17434 18054 17436
rect 18078 17434 18134 17436
rect 18158 17434 18214 17436
rect 18238 17434 18294 17436
rect 17998 17382 18044 17434
rect 18044 17382 18054 17434
rect 18078 17382 18108 17434
rect 18108 17382 18120 17434
rect 18120 17382 18134 17434
rect 18158 17382 18172 17434
rect 18172 17382 18184 17434
rect 18184 17382 18214 17434
rect 18238 17382 18248 17434
rect 18248 17382 18294 17434
rect 17998 17380 18054 17382
rect 18078 17380 18134 17382
rect 18158 17380 18214 17382
rect 18238 17380 18294 17382
rect 17998 16346 18054 16348
rect 18078 16346 18134 16348
rect 18158 16346 18214 16348
rect 18238 16346 18294 16348
rect 17998 16294 18044 16346
rect 18044 16294 18054 16346
rect 18078 16294 18108 16346
rect 18108 16294 18120 16346
rect 18120 16294 18134 16346
rect 18158 16294 18172 16346
rect 18172 16294 18184 16346
rect 18184 16294 18214 16346
rect 18238 16294 18248 16346
rect 18248 16294 18294 16346
rect 17998 16292 18054 16294
rect 18078 16292 18134 16294
rect 18158 16292 18214 16294
rect 18238 16292 18294 16294
rect 16762 15036 16764 15056
rect 16764 15036 16816 15056
rect 16816 15036 16818 15056
rect 16762 15000 16818 15036
rect 15158 8186 15214 8188
rect 15238 8186 15294 8188
rect 15318 8186 15374 8188
rect 15398 8186 15454 8188
rect 15158 8134 15204 8186
rect 15204 8134 15214 8186
rect 15238 8134 15268 8186
rect 15268 8134 15280 8186
rect 15280 8134 15294 8186
rect 15318 8134 15332 8186
rect 15332 8134 15344 8186
rect 15344 8134 15374 8186
rect 15398 8134 15408 8186
rect 15408 8134 15454 8186
rect 15158 8132 15214 8134
rect 15238 8132 15294 8134
rect 15318 8132 15374 8134
rect 15398 8132 15454 8134
rect 15158 7098 15214 7100
rect 15238 7098 15294 7100
rect 15318 7098 15374 7100
rect 15398 7098 15454 7100
rect 15158 7046 15204 7098
rect 15204 7046 15214 7098
rect 15238 7046 15268 7098
rect 15268 7046 15280 7098
rect 15280 7046 15294 7098
rect 15318 7046 15332 7098
rect 15332 7046 15344 7098
rect 15344 7046 15374 7098
rect 15398 7046 15408 7098
rect 15408 7046 15454 7098
rect 15158 7044 15214 7046
rect 15238 7044 15294 7046
rect 15318 7044 15374 7046
rect 15398 7044 15454 7046
rect 15934 12008 15990 12064
rect 17998 15258 18054 15260
rect 18078 15258 18134 15260
rect 18158 15258 18214 15260
rect 18238 15258 18294 15260
rect 17998 15206 18044 15258
rect 18044 15206 18054 15258
rect 18078 15206 18108 15258
rect 18108 15206 18120 15258
rect 18120 15206 18134 15258
rect 18158 15206 18172 15258
rect 18172 15206 18184 15258
rect 18184 15206 18214 15258
rect 18238 15206 18248 15258
rect 18248 15206 18294 15258
rect 17998 15204 18054 15206
rect 18078 15204 18134 15206
rect 18158 15204 18214 15206
rect 18238 15204 18294 15206
rect 16026 11192 16082 11248
rect 16394 10784 16450 10840
rect 16486 10104 16542 10160
rect 16486 9988 16542 10024
rect 16486 9968 16488 9988
rect 16488 9968 16540 9988
rect 16540 9968 16542 9988
rect 16486 9560 16542 9616
rect 15158 6010 15214 6012
rect 15238 6010 15294 6012
rect 15318 6010 15374 6012
rect 15398 6010 15454 6012
rect 15158 5958 15204 6010
rect 15204 5958 15214 6010
rect 15238 5958 15268 6010
rect 15268 5958 15280 6010
rect 15280 5958 15294 6010
rect 15318 5958 15332 6010
rect 15332 5958 15344 6010
rect 15344 5958 15374 6010
rect 15398 5958 15408 6010
rect 15408 5958 15454 6010
rect 15158 5956 15214 5958
rect 15238 5956 15294 5958
rect 15318 5956 15374 5958
rect 15398 5956 15454 5958
rect 15158 4922 15214 4924
rect 15238 4922 15294 4924
rect 15318 4922 15374 4924
rect 15398 4922 15454 4924
rect 15158 4870 15204 4922
rect 15204 4870 15214 4922
rect 15238 4870 15268 4922
rect 15268 4870 15280 4922
rect 15280 4870 15294 4922
rect 15318 4870 15332 4922
rect 15332 4870 15344 4922
rect 15344 4870 15374 4922
rect 15398 4870 15408 4922
rect 15408 4870 15454 4922
rect 15158 4868 15214 4870
rect 15238 4868 15294 4870
rect 15318 4868 15374 4870
rect 15398 4868 15454 4870
rect 16026 6840 16082 6896
rect 14922 4528 14978 4584
rect 16302 7656 16358 7712
rect 16486 9152 16542 9208
rect 17998 14170 18054 14172
rect 18078 14170 18134 14172
rect 18158 14170 18214 14172
rect 18238 14170 18294 14172
rect 17998 14118 18044 14170
rect 18044 14118 18054 14170
rect 18078 14118 18108 14170
rect 18108 14118 18120 14170
rect 18120 14118 18134 14170
rect 18158 14118 18172 14170
rect 18172 14118 18184 14170
rect 18184 14118 18214 14170
rect 18238 14118 18248 14170
rect 18248 14118 18294 14170
rect 17998 14116 18054 14118
rect 18078 14116 18134 14118
rect 18158 14116 18214 14118
rect 18238 14116 18294 14118
rect 23679 18522 23735 18524
rect 23759 18522 23815 18524
rect 23839 18522 23895 18524
rect 23919 18522 23975 18524
rect 23679 18470 23725 18522
rect 23725 18470 23735 18522
rect 23759 18470 23789 18522
rect 23789 18470 23801 18522
rect 23801 18470 23815 18522
rect 23839 18470 23853 18522
rect 23853 18470 23865 18522
rect 23865 18470 23895 18522
rect 23919 18470 23929 18522
rect 23929 18470 23975 18522
rect 23679 18468 23735 18470
rect 23759 18468 23815 18470
rect 23839 18468 23895 18470
rect 23919 18468 23975 18470
rect 20839 17978 20895 17980
rect 20919 17978 20975 17980
rect 20999 17978 21055 17980
rect 21079 17978 21135 17980
rect 20839 17926 20885 17978
rect 20885 17926 20895 17978
rect 20919 17926 20949 17978
rect 20949 17926 20961 17978
rect 20961 17926 20975 17978
rect 20999 17926 21013 17978
rect 21013 17926 21025 17978
rect 21025 17926 21055 17978
rect 21079 17926 21089 17978
rect 21089 17926 21135 17978
rect 20839 17924 20895 17926
rect 20919 17924 20975 17926
rect 20999 17924 21055 17926
rect 21079 17924 21135 17926
rect 23679 17434 23735 17436
rect 23759 17434 23815 17436
rect 23839 17434 23895 17436
rect 23919 17434 23975 17436
rect 23679 17382 23725 17434
rect 23725 17382 23735 17434
rect 23759 17382 23789 17434
rect 23789 17382 23801 17434
rect 23801 17382 23815 17434
rect 23839 17382 23853 17434
rect 23853 17382 23865 17434
rect 23865 17382 23895 17434
rect 23919 17382 23929 17434
rect 23929 17382 23975 17434
rect 23679 17380 23735 17382
rect 23759 17380 23815 17382
rect 23839 17380 23895 17382
rect 23919 17380 23975 17382
rect 20839 16890 20895 16892
rect 20919 16890 20975 16892
rect 20999 16890 21055 16892
rect 21079 16890 21135 16892
rect 20839 16838 20885 16890
rect 20885 16838 20895 16890
rect 20919 16838 20949 16890
rect 20949 16838 20961 16890
rect 20961 16838 20975 16890
rect 20999 16838 21013 16890
rect 21013 16838 21025 16890
rect 21025 16838 21055 16890
rect 21079 16838 21089 16890
rect 21089 16838 21135 16890
rect 20839 16836 20895 16838
rect 20919 16836 20975 16838
rect 20999 16836 21055 16838
rect 21079 16836 21135 16838
rect 23679 16346 23735 16348
rect 23759 16346 23815 16348
rect 23839 16346 23895 16348
rect 23919 16346 23975 16348
rect 23679 16294 23725 16346
rect 23725 16294 23735 16346
rect 23759 16294 23789 16346
rect 23789 16294 23801 16346
rect 23801 16294 23815 16346
rect 23839 16294 23853 16346
rect 23853 16294 23865 16346
rect 23865 16294 23895 16346
rect 23919 16294 23929 16346
rect 23929 16294 23975 16346
rect 23679 16292 23735 16294
rect 23759 16292 23815 16294
rect 23839 16292 23895 16294
rect 23919 16292 23975 16294
rect 20839 15802 20895 15804
rect 20919 15802 20975 15804
rect 20999 15802 21055 15804
rect 21079 15802 21135 15804
rect 20839 15750 20885 15802
rect 20885 15750 20895 15802
rect 20919 15750 20949 15802
rect 20949 15750 20961 15802
rect 20961 15750 20975 15802
rect 20999 15750 21013 15802
rect 21013 15750 21025 15802
rect 21025 15750 21055 15802
rect 21079 15750 21089 15802
rect 21089 15750 21135 15802
rect 20839 15748 20895 15750
rect 20919 15748 20975 15750
rect 20999 15748 21055 15750
rect 21079 15748 21135 15750
rect 17774 13232 17830 13288
rect 16946 11772 16948 11792
rect 16948 11772 17000 11792
rect 17000 11772 17002 11792
rect 16946 11736 17002 11772
rect 17038 11600 17094 11656
rect 16854 7964 16856 7984
rect 16856 7964 16908 7984
rect 16908 7964 16910 7984
rect 16854 7928 16910 7964
rect 16946 7656 17002 7712
rect 16762 5752 16818 5808
rect 17130 10784 17186 10840
rect 17314 10648 17370 10704
rect 17130 9832 17186 9888
rect 17130 9424 17186 9480
rect 17222 9152 17278 9208
rect 17222 7656 17278 7712
rect 18234 13268 18236 13288
rect 18236 13268 18288 13288
rect 18288 13268 18290 13288
rect 18234 13232 18290 13268
rect 17998 13082 18054 13084
rect 18078 13082 18134 13084
rect 18158 13082 18214 13084
rect 18238 13082 18294 13084
rect 17998 13030 18044 13082
rect 18044 13030 18054 13082
rect 18078 13030 18108 13082
rect 18108 13030 18120 13082
rect 18120 13030 18134 13082
rect 18158 13030 18172 13082
rect 18172 13030 18184 13082
rect 18184 13030 18214 13082
rect 18238 13030 18248 13082
rect 18248 13030 18294 13082
rect 17998 13028 18054 13030
rect 18078 13028 18134 13030
rect 18158 13028 18214 13030
rect 18238 13028 18294 13030
rect 17998 11994 18054 11996
rect 18078 11994 18134 11996
rect 18158 11994 18214 11996
rect 18238 11994 18294 11996
rect 17998 11942 18044 11994
rect 18044 11942 18054 11994
rect 18078 11942 18108 11994
rect 18108 11942 18120 11994
rect 18120 11942 18134 11994
rect 18158 11942 18172 11994
rect 18172 11942 18184 11994
rect 18184 11942 18214 11994
rect 18238 11942 18248 11994
rect 18248 11942 18294 11994
rect 17998 11940 18054 11942
rect 18078 11940 18134 11942
rect 18158 11940 18214 11942
rect 18238 11940 18294 11942
rect 17998 10906 18054 10908
rect 18078 10906 18134 10908
rect 18158 10906 18214 10908
rect 18238 10906 18294 10908
rect 17998 10854 18044 10906
rect 18044 10854 18054 10906
rect 18078 10854 18108 10906
rect 18108 10854 18120 10906
rect 18120 10854 18134 10906
rect 18158 10854 18172 10906
rect 18172 10854 18184 10906
rect 18184 10854 18214 10906
rect 18238 10854 18248 10906
rect 18248 10854 18294 10906
rect 17998 10852 18054 10854
rect 18078 10852 18134 10854
rect 18158 10852 18214 10854
rect 18238 10852 18294 10854
rect 17998 9818 18054 9820
rect 18078 9818 18134 9820
rect 18158 9818 18214 9820
rect 18238 9818 18294 9820
rect 17998 9766 18044 9818
rect 18044 9766 18054 9818
rect 18078 9766 18108 9818
rect 18108 9766 18120 9818
rect 18120 9766 18134 9818
rect 18158 9766 18172 9818
rect 18172 9766 18184 9818
rect 18184 9766 18214 9818
rect 18238 9766 18248 9818
rect 18248 9766 18294 9818
rect 17998 9764 18054 9766
rect 18078 9764 18134 9766
rect 18158 9764 18214 9766
rect 18238 9764 18294 9766
rect 17682 9424 17738 9480
rect 17958 9288 18014 9344
rect 17590 7792 17646 7848
rect 23679 15258 23735 15260
rect 23759 15258 23815 15260
rect 23839 15258 23895 15260
rect 23919 15258 23975 15260
rect 23679 15206 23725 15258
rect 23725 15206 23735 15258
rect 23759 15206 23789 15258
rect 23789 15206 23801 15258
rect 23801 15206 23815 15258
rect 23839 15206 23853 15258
rect 23853 15206 23865 15258
rect 23865 15206 23895 15258
rect 23919 15206 23929 15258
rect 23929 15206 23975 15258
rect 23679 15204 23735 15206
rect 23759 15204 23815 15206
rect 23839 15204 23895 15206
rect 23919 15204 23975 15206
rect 18878 11736 18934 11792
rect 18786 11600 18842 11656
rect 19062 11600 19118 11656
rect 20839 14714 20895 14716
rect 20919 14714 20975 14716
rect 20999 14714 21055 14716
rect 21079 14714 21135 14716
rect 20839 14662 20885 14714
rect 20885 14662 20895 14714
rect 20919 14662 20949 14714
rect 20949 14662 20961 14714
rect 20961 14662 20975 14714
rect 20999 14662 21013 14714
rect 21013 14662 21025 14714
rect 21025 14662 21055 14714
rect 21079 14662 21089 14714
rect 21089 14662 21135 14714
rect 20839 14660 20895 14662
rect 20919 14660 20975 14662
rect 20999 14660 21055 14662
rect 21079 14660 21135 14662
rect 19522 13776 19578 13832
rect 19706 12824 19762 12880
rect 19246 11076 19302 11112
rect 19246 11056 19248 11076
rect 19248 11056 19300 11076
rect 19300 11056 19302 11076
rect 17998 8730 18054 8732
rect 18078 8730 18134 8732
rect 18158 8730 18214 8732
rect 18238 8730 18294 8732
rect 17998 8678 18044 8730
rect 18044 8678 18054 8730
rect 18078 8678 18108 8730
rect 18108 8678 18120 8730
rect 18120 8678 18134 8730
rect 18158 8678 18172 8730
rect 18172 8678 18184 8730
rect 18184 8678 18214 8730
rect 18238 8678 18248 8730
rect 18248 8678 18294 8730
rect 17998 8676 18054 8678
rect 18078 8676 18134 8678
rect 18158 8676 18214 8678
rect 18238 8676 18294 8678
rect 18602 9716 18658 9752
rect 18602 9696 18604 9716
rect 18604 9696 18656 9716
rect 18656 9696 18658 9716
rect 18510 8880 18566 8936
rect 18050 7828 18052 7848
rect 18052 7828 18104 7848
rect 18104 7828 18106 7848
rect 18050 7792 18106 7828
rect 17998 7642 18054 7644
rect 18078 7642 18134 7644
rect 18158 7642 18214 7644
rect 18238 7642 18294 7644
rect 17998 7590 18044 7642
rect 18044 7590 18054 7642
rect 18078 7590 18108 7642
rect 18108 7590 18120 7642
rect 18120 7590 18134 7642
rect 18158 7590 18172 7642
rect 18172 7590 18184 7642
rect 18184 7590 18214 7642
rect 18238 7590 18248 7642
rect 18248 7590 18294 7642
rect 17998 7588 18054 7590
rect 18078 7588 18134 7590
rect 18158 7588 18214 7590
rect 18238 7588 18294 7590
rect 17682 6840 17738 6896
rect 17682 6432 17738 6488
rect 17998 6554 18054 6556
rect 18078 6554 18134 6556
rect 18158 6554 18214 6556
rect 18238 6554 18294 6556
rect 17998 6502 18044 6554
rect 18044 6502 18054 6554
rect 18078 6502 18108 6554
rect 18108 6502 18120 6554
rect 18120 6502 18134 6554
rect 18158 6502 18172 6554
rect 18172 6502 18184 6554
rect 18184 6502 18214 6554
rect 18238 6502 18248 6554
rect 18248 6502 18294 6554
rect 17998 6500 18054 6502
rect 18078 6500 18134 6502
rect 18158 6500 18214 6502
rect 18238 6500 18294 6502
rect 18050 6296 18106 6352
rect 18694 9152 18750 9208
rect 18878 9560 18934 9616
rect 18418 6604 18420 6624
rect 18420 6604 18472 6624
rect 18472 6604 18474 6624
rect 18418 6568 18474 6604
rect 17998 5466 18054 5468
rect 18078 5466 18134 5468
rect 18158 5466 18214 5468
rect 18238 5466 18294 5468
rect 17998 5414 18044 5466
rect 18044 5414 18054 5466
rect 18078 5414 18108 5466
rect 18108 5414 18120 5466
rect 18120 5414 18134 5466
rect 18158 5414 18172 5466
rect 18172 5414 18184 5466
rect 18184 5414 18214 5466
rect 18238 5414 18248 5466
rect 18248 5414 18294 5466
rect 17998 5412 18054 5414
rect 18078 5412 18134 5414
rect 18158 5412 18214 5414
rect 18238 5412 18294 5414
rect 19430 12280 19486 12336
rect 19062 8336 19118 8392
rect 18970 7404 19026 7440
rect 18970 7384 18972 7404
rect 18972 7384 19024 7404
rect 19024 7384 19026 7404
rect 18694 6740 18696 6760
rect 18696 6740 18748 6760
rect 18748 6740 18750 6760
rect 18694 6704 18750 6740
rect 18786 6432 18842 6488
rect 19706 11076 19762 11112
rect 19706 11056 19708 11076
rect 19708 11056 19760 11076
rect 19760 11056 19762 11076
rect 19154 6704 19210 6760
rect 19338 6740 19340 6760
rect 19340 6740 19392 6760
rect 19392 6740 19394 6760
rect 19338 6704 19394 6740
rect 19062 6296 19118 6352
rect 19154 5772 19210 5808
rect 19154 5752 19156 5772
rect 19156 5752 19208 5772
rect 19208 5752 19210 5772
rect 19890 9696 19946 9752
rect 20074 12180 20076 12200
rect 20076 12180 20128 12200
rect 20128 12180 20130 12200
rect 20074 12144 20130 12180
rect 20074 9460 20076 9480
rect 20076 9460 20128 9480
rect 20128 9460 20130 9480
rect 20074 9424 20130 9460
rect 20839 13626 20895 13628
rect 20919 13626 20975 13628
rect 20999 13626 21055 13628
rect 21079 13626 21135 13628
rect 20839 13574 20885 13626
rect 20885 13574 20895 13626
rect 20919 13574 20949 13626
rect 20949 13574 20961 13626
rect 20961 13574 20975 13626
rect 20999 13574 21013 13626
rect 21013 13574 21025 13626
rect 21025 13574 21055 13626
rect 21079 13574 21089 13626
rect 21089 13574 21135 13626
rect 20839 13572 20895 13574
rect 20919 13572 20975 13574
rect 20999 13572 21055 13574
rect 21079 13572 21135 13574
rect 23679 14170 23735 14172
rect 23759 14170 23815 14172
rect 23839 14170 23895 14172
rect 23919 14170 23975 14172
rect 23679 14118 23725 14170
rect 23725 14118 23735 14170
rect 23759 14118 23789 14170
rect 23789 14118 23801 14170
rect 23801 14118 23815 14170
rect 23839 14118 23853 14170
rect 23853 14118 23865 14170
rect 23865 14118 23895 14170
rect 23919 14118 23929 14170
rect 23929 14118 23975 14170
rect 23679 14116 23735 14118
rect 23759 14116 23815 14118
rect 23839 14116 23895 14118
rect 23919 14116 23975 14118
rect 20626 12824 20682 12880
rect 20534 10956 20536 10976
rect 20536 10956 20588 10976
rect 20588 10956 20590 10976
rect 20534 10920 20590 10956
rect 20350 10104 20406 10160
rect 19798 7248 19854 7304
rect 20839 12538 20895 12540
rect 20919 12538 20975 12540
rect 20999 12538 21055 12540
rect 21079 12538 21135 12540
rect 20839 12486 20885 12538
rect 20885 12486 20895 12538
rect 20919 12486 20949 12538
rect 20949 12486 20961 12538
rect 20961 12486 20975 12538
rect 20999 12486 21013 12538
rect 21013 12486 21025 12538
rect 21025 12486 21055 12538
rect 21079 12486 21089 12538
rect 21089 12486 21135 12538
rect 20839 12484 20895 12486
rect 20919 12484 20975 12486
rect 20999 12484 21055 12486
rect 21079 12484 21135 12486
rect 20839 11450 20895 11452
rect 20919 11450 20975 11452
rect 20999 11450 21055 11452
rect 21079 11450 21135 11452
rect 20839 11398 20885 11450
rect 20885 11398 20895 11450
rect 20919 11398 20949 11450
rect 20949 11398 20961 11450
rect 20961 11398 20975 11450
rect 20999 11398 21013 11450
rect 21013 11398 21025 11450
rect 21025 11398 21055 11450
rect 21079 11398 21089 11450
rect 21089 11398 21135 11450
rect 20839 11396 20895 11398
rect 20919 11396 20975 11398
rect 20999 11396 21055 11398
rect 21079 11396 21135 11398
rect 20718 11070 20720 11112
rect 20720 11070 20772 11112
rect 20772 11070 20774 11112
rect 20718 11056 20774 11070
rect 20534 9580 20590 9616
rect 20534 9560 20536 9580
rect 20536 9560 20588 9580
rect 20588 9560 20590 9580
rect 20350 9288 20406 9344
rect 20534 9288 20590 9344
rect 20994 10920 21050 10976
rect 23679 13082 23735 13084
rect 23759 13082 23815 13084
rect 23839 13082 23895 13084
rect 23919 13082 23975 13084
rect 23679 13030 23725 13082
rect 23725 13030 23735 13082
rect 23759 13030 23789 13082
rect 23789 13030 23801 13082
rect 23801 13030 23815 13082
rect 23839 13030 23853 13082
rect 23853 13030 23865 13082
rect 23865 13030 23895 13082
rect 23919 13030 23929 13082
rect 23929 13030 23975 13082
rect 23679 13028 23735 13030
rect 23759 13028 23815 13030
rect 23839 13028 23895 13030
rect 23919 13028 23975 13030
rect 21270 10648 21326 10704
rect 20839 10362 20895 10364
rect 20919 10362 20975 10364
rect 20999 10362 21055 10364
rect 21079 10362 21135 10364
rect 20839 10310 20885 10362
rect 20885 10310 20895 10362
rect 20919 10310 20949 10362
rect 20949 10310 20961 10362
rect 20961 10310 20975 10362
rect 20999 10310 21013 10362
rect 21013 10310 21025 10362
rect 21025 10310 21055 10362
rect 21079 10310 21089 10362
rect 21089 10310 21135 10362
rect 20839 10308 20895 10310
rect 20919 10308 20975 10310
rect 20999 10308 21055 10310
rect 21079 10308 21135 10310
rect 20902 10104 20958 10160
rect 20839 9274 20895 9276
rect 20919 9274 20975 9276
rect 20999 9274 21055 9276
rect 21079 9274 21135 9276
rect 20839 9222 20885 9274
rect 20885 9222 20895 9274
rect 20919 9222 20949 9274
rect 20949 9222 20961 9274
rect 20961 9222 20975 9274
rect 20999 9222 21013 9274
rect 21013 9222 21025 9274
rect 21025 9222 21055 9274
rect 21079 9222 21089 9274
rect 21089 9222 21135 9274
rect 20839 9220 20895 9222
rect 20919 9220 20975 9222
rect 20999 9220 21055 9222
rect 21079 9220 21135 9222
rect 20258 8084 20314 8120
rect 20258 8064 20260 8084
rect 20260 8064 20312 8084
rect 20312 8064 20314 8084
rect 19982 7404 20038 7440
rect 19982 7384 19984 7404
rect 19984 7384 20036 7404
rect 20036 7384 20038 7404
rect 20810 8356 20866 8392
rect 20810 8336 20812 8356
rect 20812 8336 20864 8356
rect 20864 8336 20866 8356
rect 20839 8186 20895 8188
rect 20919 8186 20975 8188
rect 20999 8186 21055 8188
rect 21079 8186 21135 8188
rect 20839 8134 20885 8186
rect 20885 8134 20895 8186
rect 20919 8134 20949 8186
rect 20949 8134 20961 8186
rect 20961 8134 20975 8186
rect 20999 8134 21013 8186
rect 21013 8134 21025 8186
rect 21025 8134 21055 8186
rect 21079 8134 21089 8186
rect 21089 8134 21135 8186
rect 20839 8132 20895 8134
rect 20919 8132 20975 8134
rect 20999 8132 21055 8134
rect 21079 8132 21135 8134
rect 20810 7248 20866 7304
rect 20839 7098 20895 7100
rect 20919 7098 20975 7100
rect 20999 7098 21055 7100
rect 21079 7098 21135 7100
rect 20839 7046 20885 7098
rect 20885 7046 20895 7098
rect 20919 7046 20949 7098
rect 20949 7046 20961 7098
rect 20961 7046 20975 7098
rect 20999 7046 21013 7098
rect 21013 7046 21025 7098
rect 21025 7046 21055 7098
rect 21079 7046 21089 7098
rect 21089 7046 21135 7098
rect 20839 7044 20895 7046
rect 20919 7044 20975 7046
rect 20999 7044 21055 7046
rect 21079 7044 21135 7046
rect 21454 7248 21510 7304
rect 21730 6568 21786 6624
rect 21178 6432 21234 6488
rect 22190 11600 22246 11656
rect 22190 9016 22246 9072
rect 20350 5480 20406 5536
rect 20839 6010 20895 6012
rect 20919 6010 20975 6012
rect 20999 6010 21055 6012
rect 21079 6010 21135 6012
rect 20839 5958 20885 6010
rect 20885 5958 20895 6010
rect 20919 5958 20949 6010
rect 20949 5958 20961 6010
rect 20961 5958 20975 6010
rect 20999 5958 21013 6010
rect 21013 5958 21025 6010
rect 21025 5958 21055 6010
rect 21079 5958 21089 6010
rect 21089 5958 21135 6010
rect 20839 5956 20895 5958
rect 20919 5956 20975 5958
rect 20999 5956 21055 5958
rect 21079 5956 21135 5958
rect 23679 11994 23735 11996
rect 23759 11994 23815 11996
rect 23839 11994 23895 11996
rect 23919 11994 23975 11996
rect 23679 11942 23725 11994
rect 23725 11942 23735 11994
rect 23759 11942 23789 11994
rect 23789 11942 23801 11994
rect 23801 11942 23815 11994
rect 23839 11942 23853 11994
rect 23853 11942 23865 11994
rect 23865 11942 23895 11994
rect 23919 11942 23929 11994
rect 23929 11942 23975 11994
rect 23679 11940 23735 11942
rect 23759 11940 23815 11942
rect 23839 11940 23895 11942
rect 23919 11940 23975 11942
rect 23679 10906 23735 10908
rect 23759 10906 23815 10908
rect 23839 10906 23895 10908
rect 23919 10906 23975 10908
rect 23679 10854 23725 10906
rect 23725 10854 23735 10906
rect 23759 10854 23789 10906
rect 23789 10854 23801 10906
rect 23801 10854 23815 10906
rect 23839 10854 23853 10906
rect 23853 10854 23865 10906
rect 23865 10854 23895 10906
rect 23919 10854 23929 10906
rect 23929 10854 23975 10906
rect 23679 10852 23735 10854
rect 23759 10852 23815 10854
rect 23839 10852 23895 10854
rect 23919 10852 23975 10854
rect 23679 9818 23735 9820
rect 23759 9818 23815 9820
rect 23839 9818 23895 9820
rect 23919 9818 23975 9820
rect 23679 9766 23725 9818
rect 23725 9766 23735 9818
rect 23759 9766 23789 9818
rect 23789 9766 23801 9818
rect 23801 9766 23815 9818
rect 23839 9766 23853 9818
rect 23853 9766 23865 9818
rect 23865 9766 23895 9818
rect 23919 9766 23929 9818
rect 23929 9766 23975 9818
rect 23679 9764 23735 9766
rect 23759 9764 23815 9766
rect 23839 9764 23895 9766
rect 23919 9764 23975 9766
rect 23679 8730 23735 8732
rect 23759 8730 23815 8732
rect 23839 8730 23895 8732
rect 23919 8730 23975 8732
rect 23679 8678 23725 8730
rect 23725 8678 23735 8730
rect 23759 8678 23789 8730
rect 23789 8678 23801 8730
rect 23801 8678 23815 8730
rect 23839 8678 23853 8730
rect 23853 8678 23865 8730
rect 23865 8678 23895 8730
rect 23919 8678 23929 8730
rect 23929 8678 23975 8730
rect 23679 8676 23735 8678
rect 23759 8676 23815 8678
rect 23839 8676 23895 8678
rect 23919 8676 23975 8678
rect 23679 7642 23735 7644
rect 23759 7642 23815 7644
rect 23839 7642 23895 7644
rect 23919 7642 23975 7644
rect 23679 7590 23725 7642
rect 23725 7590 23735 7642
rect 23759 7590 23789 7642
rect 23789 7590 23801 7642
rect 23801 7590 23815 7642
rect 23839 7590 23853 7642
rect 23853 7590 23865 7642
rect 23865 7590 23895 7642
rect 23919 7590 23929 7642
rect 23929 7590 23975 7642
rect 23679 7588 23735 7590
rect 23759 7588 23815 7590
rect 23839 7588 23895 7590
rect 23919 7588 23975 7590
rect 23679 6554 23735 6556
rect 23759 6554 23815 6556
rect 23839 6554 23895 6556
rect 23919 6554 23975 6556
rect 23679 6502 23725 6554
rect 23725 6502 23735 6554
rect 23759 6502 23789 6554
rect 23789 6502 23801 6554
rect 23801 6502 23815 6554
rect 23839 6502 23853 6554
rect 23853 6502 23865 6554
rect 23865 6502 23895 6554
rect 23919 6502 23929 6554
rect 23929 6502 23975 6554
rect 23679 6500 23735 6502
rect 23759 6500 23815 6502
rect 23839 6500 23895 6502
rect 23919 6500 23975 6502
rect 20839 4922 20895 4924
rect 20919 4922 20975 4924
rect 20999 4922 21055 4924
rect 21079 4922 21135 4924
rect 20839 4870 20885 4922
rect 20885 4870 20895 4922
rect 20919 4870 20949 4922
rect 20949 4870 20961 4922
rect 20961 4870 20975 4922
rect 20999 4870 21013 4922
rect 21013 4870 21025 4922
rect 21025 4870 21055 4922
rect 21079 4870 21089 4922
rect 21089 4870 21135 4922
rect 20839 4868 20895 4870
rect 20919 4868 20975 4870
rect 20999 4868 21055 4870
rect 21079 4868 21135 4870
rect 23679 5466 23735 5468
rect 23759 5466 23815 5468
rect 23839 5466 23895 5468
rect 23919 5466 23975 5468
rect 23679 5414 23725 5466
rect 23725 5414 23735 5466
rect 23759 5414 23789 5466
rect 23789 5414 23801 5466
rect 23801 5414 23815 5466
rect 23839 5414 23853 5466
rect 23853 5414 23865 5466
rect 23865 5414 23895 5466
rect 23919 5414 23929 5466
rect 23929 5414 23975 5466
rect 23679 5412 23735 5414
rect 23759 5412 23815 5414
rect 23839 5412 23895 5414
rect 23919 5412 23975 5414
rect 17998 4378 18054 4380
rect 18078 4378 18134 4380
rect 18158 4378 18214 4380
rect 18238 4378 18294 4380
rect 17998 4326 18044 4378
rect 18044 4326 18054 4378
rect 18078 4326 18108 4378
rect 18108 4326 18120 4378
rect 18120 4326 18134 4378
rect 18158 4326 18172 4378
rect 18172 4326 18184 4378
rect 18184 4326 18214 4378
rect 18238 4326 18248 4378
rect 18248 4326 18294 4378
rect 17998 4324 18054 4326
rect 18078 4324 18134 4326
rect 18158 4324 18214 4326
rect 18238 4324 18294 4326
rect 23679 4378 23735 4380
rect 23759 4378 23815 4380
rect 23839 4378 23895 4380
rect 23919 4378 23975 4380
rect 23679 4326 23725 4378
rect 23725 4326 23735 4378
rect 23759 4326 23789 4378
rect 23789 4326 23801 4378
rect 23801 4326 23815 4378
rect 23839 4326 23853 4378
rect 23853 4326 23865 4378
rect 23865 4326 23895 4378
rect 23919 4326 23929 4378
rect 23929 4326 23975 4378
rect 23679 4324 23735 4326
rect 23759 4324 23815 4326
rect 23839 4324 23895 4326
rect 23919 4324 23975 4326
rect 15158 3834 15214 3836
rect 15238 3834 15294 3836
rect 15318 3834 15374 3836
rect 15398 3834 15454 3836
rect 15158 3782 15204 3834
rect 15204 3782 15214 3834
rect 15238 3782 15268 3834
rect 15268 3782 15280 3834
rect 15280 3782 15294 3834
rect 15318 3782 15332 3834
rect 15332 3782 15344 3834
rect 15344 3782 15374 3834
rect 15398 3782 15408 3834
rect 15408 3782 15454 3834
rect 15158 3780 15214 3782
rect 15238 3780 15294 3782
rect 15318 3780 15374 3782
rect 15398 3780 15454 3782
rect 17406 3984 17462 4040
rect 12317 3290 12373 3292
rect 12397 3290 12453 3292
rect 12477 3290 12533 3292
rect 12557 3290 12613 3292
rect 12317 3238 12363 3290
rect 12363 3238 12373 3290
rect 12397 3238 12427 3290
rect 12427 3238 12439 3290
rect 12439 3238 12453 3290
rect 12477 3238 12491 3290
rect 12491 3238 12503 3290
rect 12503 3238 12533 3290
rect 12557 3238 12567 3290
rect 12567 3238 12613 3290
rect 12317 3236 12373 3238
rect 12397 3236 12453 3238
rect 12477 3236 12533 3238
rect 12557 3236 12613 3238
rect 15158 2746 15214 2748
rect 15238 2746 15294 2748
rect 15318 2746 15374 2748
rect 15398 2746 15454 2748
rect 15158 2694 15204 2746
rect 15204 2694 15214 2746
rect 15238 2694 15268 2746
rect 15268 2694 15280 2746
rect 15280 2694 15294 2746
rect 15318 2694 15332 2746
rect 15332 2694 15344 2746
rect 15344 2694 15374 2746
rect 15398 2694 15408 2746
rect 15408 2694 15454 2746
rect 15158 2692 15214 2694
rect 15238 2692 15294 2694
rect 15318 2692 15374 2694
rect 15398 2692 15454 2694
rect 12317 2202 12373 2204
rect 12397 2202 12453 2204
rect 12477 2202 12533 2204
rect 12557 2202 12613 2204
rect 12317 2150 12363 2202
rect 12363 2150 12373 2202
rect 12397 2150 12427 2202
rect 12427 2150 12439 2202
rect 12439 2150 12453 2202
rect 12477 2150 12491 2202
rect 12491 2150 12503 2202
rect 12503 2150 12533 2202
rect 12557 2150 12567 2202
rect 12567 2150 12613 2202
rect 12317 2148 12373 2150
rect 12397 2148 12453 2150
rect 12477 2148 12533 2150
rect 12557 2148 12613 2150
rect 20839 3834 20895 3836
rect 20919 3834 20975 3836
rect 20999 3834 21055 3836
rect 21079 3834 21135 3836
rect 20839 3782 20885 3834
rect 20885 3782 20895 3834
rect 20919 3782 20949 3834
rect 20949 3782 20961 3834
rect 20961 3782 20975 3834
rect 20999 3782 21013 3834
rect 21013 3782 21025 3834
rect 21025 3782 21055 3834
rect 21079 3782 21089 3834
rect 21089 3782 21135 3834
rect 20839 3780 20895 3782
rect 20919 3780 20975 3782
rect 20999 3780 21055 3782
rect 21079 3780 21135 3782
rect 17958 3460 18014 3496
rect 17958 3440 17960 3460
rect 17960 3440 18012 3460
rect 18012 3440 18014 3460
rect 17998 3290 18054 3292
rect 18078 3290 18134 3292
rect 18158 3290 18214 3292
rect 18238 3290 18294 3292
rect 17998 3238 18044 3290
rect 18044 3238 18054 3290
rect 18078 3238 18108 3290
rect 18108 3238 18120 3290
rect 18120 3238 18134 3290
rect 18158 3238 18172 3290
rect 18172 3238 18184 3290
rect 18184 3238 18214 3290
rect 18238 3238 18248 3290
rect 18248 3238 18294 3290
rect 17998 3236 18054 3238
rect 18078 3236 18134 3238
rect 18158 3236 18214 3238
rect 18238 3236 18294 3238
rect 17998 2202 18054 2204
rect 18078 2202 18134 2204
rect 18158 2202 18214 2204
rect 18238 2202 18294 2204
rect 17998 2150 18044 2202
rect 18044 2150 18054 2202
rect 18078 2150 18108 2202
rect 18108 2150 18120 2202
rect 18120 2150 18134 2202
rect 18158 2150 18172 2202
rect 18172 2150 18184 2202
rect 18184 2150 18214 2202
rect 18238 2150 18248 2202
rect 18248 2150 18294 2202
rect 17998 2148 18054 2150
rect 18078 2148 18134 2150
rect 18158 2148 18214 2150
rect 18238 2148 18294 2150
rect 20839 2746 20895 2748
rect 20919 2746 20975 2748
rect 20999 2746 21055 2748
rect 21079 2746 21135 2748
rect 20839 2694 20885 2746
rect 20885 2694 20895 2746
rect 20919 2694 20949 2746
rect 20949 2694 20961 2746
rect 20961 2694 20975 2746
rect 20999 2694 21013 2746
rect 21013 2694 21025 2746
rect 21025 2694 21055 2746
rect 21079 2694 21089 2746
rect 21089 2694 21135 2746
rect 20839 2692 20895 2694
rect 20919 2692 20975 2694
rect 20999 2692 21055 2694
rect 21079 2692 21135 2694
rect 23679 3290 23735 3292
rect 23759 3290 23815 3292
rect 23839 3290 23895 3292
rect 23919 3290 23975 3292
rect 23679 3238 23725 3290
rect 23725 3238 23735 3290
rect 23759 3238 23789 3290
rect 23789 3238 23801 3290
rect 23801 3238 23815 3290
rect 23839 3238 23853 3290
rect 23853 3238 23865 3290
rect 23865 3238 23895 3290
rect 23919 3238 23929 3290
rect 23929 3238 23975 3290
rect 23679 3236 23735 3238
rect 23759 3236 23815 3238
rect 23839 3236 23895 3238
rect 23919 3236 23975 3238
rect 23679 2202 23735 2204
rect 23759 2202 23815 2204
rect 23839 2202 23895 2204
rect 23919 2202 23975 2204
rect 23679 2150 23725 2202
rect 23725 2150 23735 2202
rect 23759 2150 23789 2202
rect 23789 2150 23801 2202
rect 23801 2150 23815 2202
rect 23839 2150 23853 2202
rect 23853 2150 23865 2202
rect 23865 2150 23895 2202
rect 23919 2150 23929 2202
rect 23929 2150 23975 2202
rect 23679 2148 23735 2150
rect 23759 2148 23815 2150
rect 23839 2148 23895 2150
rect 23919 2148 23975 2150
<< metal3 >>
rect 3786 22336 4102 22337
rect 3786 22272 3792 22336
rect 3856 22272 3872 22336
rect 3936 22272 3952 22336
rect 4016 22272 4032 22336
rect 4096 22272 4102 22336
rect 3786 22271 4102 22272
rect 9467 22336 9783 22337
rect 9467 22272 9473 22336
rect 9537 22272 9553 22336
rect 9617 22272 9633 22336
rect 9697 22272 9713 22336
rect 9777 22272 9783 22336
rect 9467 22271 9783 22272
rect 15148 22336 15464 22337
rect 15148 22272 15154 22336
rect 15218 22272 15234 22336
rect 15298 22272 15314 22336
rect 15378 22272 15394 22336
rect 15458 22272 15464 22336
rect 15148 22271 15464 22272
rect 20829 22336 21145 22337
rect 20829 22272 20835 22336
rect 20899 22272 20915 22336
rect 20979 22272 20995 22336
rect 21059 22272 21075 22336
rect 21139 22272 21145 22336
rect 20829 22271 21145 22272
rect 6626 21792 6942 21793
rect 6626 21728 6632 21792
rect 6696 21728 6712 21792
rect 6776 21728 6792 21792
rect 6856 21728 6872 21792
rect 6936 21728 6942 21792
rect 6626 21727 6942 21728
rect 12307 21792 12623 21793
rect 12307 21728 12313 21792
rect 12377 21728 12393 21792
rect 12457 21728 12473 21792
rect 12537 21728 12553 21792
rect 12617 21728 12623 21792
rect 12307 21727 12623 21728
rect 17988 21792 18304 21793
rect 17988 21728 17994 21792
rect 18058 21728 18074 21792
rect 18138 21728 18154 21792
rect 18218 21728 18234 21792
rect 18298 21728 18304 21792
rect 17988 21727 18304 21728
rect 23669 21792 23985 21793
rect 23669 21728 23675 21792
rect 23739 21728 23755 21792
rect 23819 21728 23835 21792
rect 23899 21728 23915 21792
rect 23979 21728 23985 21792
rect 23669 21727 23985 21728
rect 3786 21248 4102 21249
rect 3786 21184 3792 21248
rect 3856 21184 3872 21248
rect 3936 21184 3952 21248
rect 4016 21184 4032 21248
rect 4096 21184 4102 21248
rect 3786 21183 4102 21184
rect 9467 21248 9783 21249
rect 9467 21184 9473 21248
rect 9537 21184 9553 21248
rect 9617 21184 9633 21248
rect 9697 21184 9713 21248
rect 9777 21184 9783 21248
rect 9467 21183 9783 21184
rect 15148 21248 15464 21249
rect 15148 21184 15154 21248
rect 15218 21184 15234 21248
rect 15298 21184 15314 21248
rect 15378 21184 15394 21248
rect 15458 21184 15464 21248
rect 15148 21183 15464 21184
rect 20829 21248 21145 21249
rect 20829 21184 20835 21248
rect 20899 21184 20915 21248
rect 20979 21184 20995 21248
rect 21059 21184 21075 21248
rect 21139 21184 21145 21248
rect 20829 21183 21145 21184
rect 4286 20708 4292 20772
rect 4356 20770 4362 20772
rect 4889 20770 4955 20773
rect 4356 20768 4955 20770
rect 4356 20712 4894 20768
rect 4950 20712 4955 20768
rect 4356 20710 4955 20712
rect 4356 20708 4362 20710
rect 4889 20707 4955 20710
rect 7598 20708 7604 20772
rect 7668 20770 7674 20772
rect 8109 20770 8175 20773
rect 7668 20768 8175 20770
rect 7668 20712 8114 20768
rect 8170 20712 8175 20768
rect 7668 20710 8175 20712
rect 7668 20708 7674 20710
rect 8109 20707 8175 20710
rect 6626 20704 6942 20705
rect 6626 20640 6632 20704
rect 6696 20640 6712 20704
rect 6776 20640 6792 20704
rect 6856 20640 6872 20704
rect 6936 20640 6942 20704
rect 6626 20639 6942 20640
rect 12307 20704 12623 20705
rect 12307 20640 12313 20704
rect 12377 20640 12393 20704
rect 12457 20640 12473 20704
rect 12537 20640 12553 20704
rect 12617 20640 12623 20704
rect 12307 20639 12623 20640
rect 17988 20704 18304 20705
rect 17988 20640 17994 20704
rect 18058 20640 18074 20704
rect 18138 20640 18154 20704
rect 18218 20640 18234 20704
rect 18298 20640 18304 20704
rect 17988 20639 18304 20640
rect 23669 20704 23985 20705
rect 23669 20640 23675 20704
rect 23739 20640 23755 20704
rect 23819 20640 23835 20704
rect 23899 20640 23915 20704
rect 23979 20640 23985 20704
rect 23669 20639 23985 20640
rect 3786 20160 4102 20161
rect 3786 20096 3792 20160
rect 3856 20096 3872 20160
rect 3936 20096 3952 20160
rect 4016 20096 4032 20160
rect 4096 20096 4102 20160
rect 3786 20095 4102 20096
rect 9467 20160 9783 20161
rect 9467 20096 9473 20160
rect 9537 20096 9553 20160
rect 9617 20096 9633 20160
rect 9697 20096 9713 20160
rect 9777 20096 9783 20160
rect 9467 20095 9783 20096
rect 15148 20160 15464 20161
rect 15148 20096 15154 20160
rect 15218 20096 15234 20160
rect 15298 20096 15314 20160
rect 15378 20096 15394 20160
rect 15458 20096 15464 20160
rect 15148 20095 15464 20096
rect 20829 20160 21145 20161
rect 20829 20096 20835 20160
rect 20899 20096 20915 20160
rect 20979 20096 20995 20160
rect 21059 20096 21075 20160
rect 21139 20096 21145 20160
rect 20829 20095 21145 20096
rect 6626 19616 6942 19617
rect 6626 19552 6632 19616
rect 6696 19552 6712 19616
rect 6776 19552 6792 19616
rect 6856 19552 6872 19616
rect 6936 19552 6942 19616
rect 6626 19551 6942 19552
rect 12307 19616 12623 19617
rect 12307 19552 12313 19616
rect 12377 19552 12393 19616
rect 12457 19552 12473 19616
rect 12537 19552 12553 19616
rect 12617 19552 12623 19616
rect 12307 19551 12623 19552
rect 17988 19616 18304 19617
rect 17988 19552 17994 19616
rect 18058 19552 18074 19616
rect 18138 19552 18154 19616
rect 18218 19552 18234 19616
rect 18298 19552 18304 19616
rect 17988 19551 18304 19552
rect 23669 19616 23985 19617
rect 23669 19552 23675 19616
rect 23739 19552 23755 19616
rect 23819 19552 23835 19616
rect 23899 19552 23915 19616
rect 23979 19552 23985 19616
rect 23669 19551 23985 19552
rect 3550 19348 3556 19412
rect 3620 19410 3626 19412
rect 3693 19410 3759 19413
rect 6361 19412 6427 19413
rect 6310 19410 6316 19412
rect 3620 19408 3759 19410
rect 3620 19352 3698 19408
rect 3754 19352 3759 19408
rect 3620 19350 3759 19352
rect 6270 19350 6316 19410
rect 6380 19408 6427 19412
rect 6422 19352 6427 19408
rect 3620 19348 3626 19350
rect 3693 19347 3759 19350
rect 6310 19348 6316 19350
rect 6380 19348 6427 19352
rect 6361 19347 6427 19348
rect 3786 19072 4102 19073
rect 3786 19008 3792 19072
rect 3856 19008 3872 19072
rect 3936 19008 3952 19072
rect 4016 19008 4032 19072
rect 4096 19008 4102 19072
rect 3786 19007 4102 19008
rect 9467 19072 9783 19073
rect 9467 19008 9473 19072
rect 9537 19008 9553 19072
rect 9617 19008 9633 19072
rect 9697 19008 9713 19072
rect 9777 19008 9783 19072
rect 9467 19007 9783 19008
rect 15148 19072 15464 19073
rect 15148 19008 15154 19072
rect 15218 19008 15234 19072
rect 15298 19008 15314 19072
rect 15378 19008 15394 19072
rect 15458 19008 15464 19072
rect 15148 19007 15464 19008
rect 20829 19072 21145 19073
rect 20829 19008 20835 19072
rect 20899 19008 20915 19072
rect 20979 19008 20995 19072
rect 21059 19008 21075 19072
rect 21139 19008 21145 19072
rect 20829 19007 21145 19008
rect 6626 18528 6942 18529
rect 6626 18464 6632 18528
rect 6696 18464 6712 18528
rect 6776 18464 6792 18528
rect 6856 18464 6872 18528
rect 6936 18464 6942 18528
rect 6626 18463 6942 18464
rect 12307 18528 12623 18529
rect 12307 18464 12313 18528
rect 12377 18464 12393 18528
rect 12457 18464 12473 18528
rect 12537 18464 12553 18528
rect 12617 18464 12623 18528
rect 12307 18463 12623 18464
rect 17988 18528 18304 18529
rect 17988 18464 17994 18528
rect 18058 18464 18074 18528
rect 18138 18464 18154 18528
rect 18218 18464 18234 18528
rect 18298 18464 18304 18528
rect 17988 18463 18304 18464
rect 23669 18528 23985 18529
rect 23669 18464 23675 18528
rect 23739 18464 23755 18528
rect 23819 18464 23835 18528
rect 23899 18464 23915 18528
rect 23979 18464 23985 18528
rect 23669 18463 23985 18464
rect 7373 18052 7439 18053
rect 7373 18048 7420 18052
rect 7484 18050 7490 18052
rect 7373 17992 7378 18048
rect 7373 17988 7420 17992
rect 7484 17990 7530 18050
rect 7484 17988 7490 17990
rect 7373 17987 7439 17988
rect 3786 17984 4102 17985
rect 3786 17920 3792 17984
rect 3856 17920 3872 17984
rect 3936 17920 3952 17984
rect 4016 17920 4032 17984
rect 4096 17920 4102 17984
rect 3786 17919 4102 17920
rect 9467 17984 9783 17985
rect 9467 17920 9473 17984
rect 9537 17920 9553 17984
rect 9617 17920 9633 17984
rect 9697 17920 9713 17984
rect 9777 17920 9783 17984
rect 9467 17919 9783 17920
rect 15148 17984 15464 17985
rect 15148 17920 15154 17984
rect 15218 17920 15234 17984
rect 15298 17920 15314 17984
rect 15378 17920 15394 17984
rect 15458 17920 15464 17984
rect 15148 17919 15464 17920
rect 20829 17984 21145 17985
rect 20829 17920 20835 17984
rect 20899 17920 20915 17984
rect 20979 17920 20995 17984
rect 21059 17920 21075 17984
rect 21139 17920 21145 17984
rect 20829 17919 21145 17920
rect 6626 17440 6942 17441
rect 6626 17376 6632 17440
rect 6696 17376 6712 17440
rect 6776 17376 6792 17440
rect 6856 17376 6872 17440
rect 6936 17376 6942 17440
rect 6626 17375 6942 17376
rect 12307 17440 12623 17441
rect 12307 17376 12313 17440
rect 12377 17376 12393 17440
rect 12457 17376 12473 17440
rect 12537 17376 12553 17440
rect 12617 17376 12623 17440
rect 12307 17375 12623 17376
rect 17988 17440 18304 17441
rect 17988 17376 17994 17440
rect 18058 17376 18074 17440
rect 18138 17376 18154 17440
rect 18218 17376 18234 17440
rect 18298 17376 18304 17440
rect 17988 17375 18304 17376
rect 23669 17440 23985 17441
rect 23669 17376 23675 17440
rect 23739 17376 23755 17440
rect 23819 17376 23835 17440
rect 23899 17376 23915 17440
rect 23979 17376 23985 17440
rect 23669 17375 23985 17376
rect 3786 16896 4102 16897
rect 3786 16832 3792 16896
rect 3856 16832 3872 16896
rect 3936 16832 3952 16896
rect 4016 16832 4032 16896
rect 4096 16832 4102 16896
rect 3786 16831 4102 16832
rect 9467 16896 9783 16897
rect 9467 16832 9473 16896
rect 9537 16832 9553 16896
rect 9617 16832 9633 16896
rect 9697 16832 9713 16896
rect 9777 16832 9783 16896
rect 9467 16831 9783 16832
rect 15148 16896 15464 16897
rect 15148 16832 15154 16896
rect 15218 16832 15234 16896
rect 15298 16832 15314 16896
rect 15378 16832 15394 16896
rect 15458 16832 15464 16896
rect 15148 16831 15464 16832
rect 20829 16896 21145 16897
rect 20829 16832 20835 16896
rect 20899 16832 20915 16896
rect 20979 16832 20995 16896
rect 21059 16832 21075 16896
rect 21139 16832 21145 16896
rect 20829 16831 21145 16832
rect 3417 16692 3483 16693
rect 3366 16690 3372 16692
rect 3326 16630 3372 16690
rect 3436 16688 3483 16692
rect 3478 16632 3483 16688
rect 3366 16628 3372 16630
rect 3436 16628 3483 16632
rect 3417 16627 3483 16628
rect 6626 16352 6942 16353
rect 6626 16288 6632 16352
rect 6696 16288 6712 16352
rect 6776 16288 6792 16352
rect 6856 16288 6872 16352
rect 6936 16288 6942 16352
rect 6626 16287 6942 16288
rect 12307 16352 12623 16353
rect 12307 16288 12313 16352
rect 12377 16288 12393 16352
rect 12457 16288 12473 16352
rect 12537 16288 12553 16352
rect 12617 16288 12623 16352
rect 12307 16287 12623 16288
rect 17988 16352 18304 16353
rect 17988 16288 17994 16352
rect 18058 16288 18074 16352
rect 18138 16288 18154 16352
rect 18218 16288 18234 16352
rect 18298 16288 18304 16352
rect 17988 16287 18304 16288
rect 23669 16352 23985 16353
rect 23669 16288 23675 16352
rect 23739 16288 23755 16352
rect 23819 16288 23835 16352
rect 23899 16288 23915 16352
rect 23979 16288 23985 16352
rect 23669 16287 23985 16288
rect 3786 15808 4102 15809
rect 3786 15744 3792 15808
rect 3856 15744 3872 15808
rect 3936 15744 3952 15808
rect 4016 15744 4032 15808
rect 4096 15744 4102 15808
rect 3786 15743 4102 15744
rect 9467 15808 9783 15809
rect 9467 15744 9473 15808
rect 9537 15744 9553 15808
rect 9617 15744 9633 15808
rect 9697 15744 9713 15808
rect 9777 15744 9783 15808
rect 9467 15743 9783 15744
rect 15148 15808 15464 15809
rect 15148 15744 15154 15808
rect 15218 15744 15234 15808
rect 15298 15744 15314 15808
rect 15378 15744 15394 15808
rect 15458 15744 15464 15808
rect 15148 15743 15464 15744
rect 20829 15808 21145 15809
rect 20829 15744 20835 15808
rect 20899 15744 20915 15808
rect 20979 15744 20995 15808
rect 21059 15744 21075 15808
rect 21139 15744 21145 15808
rect 20829 15743 21145 15744
rect 6626 15264 6942 15265
rect 6626 15200 6632 15264
rect 6696 15200 6712 15264
rect 6776 15200 6792 15264
rect 6856 15200 6872 15264
rect 6936 15200 6942 15264
rect 6626 15199 6942 15200
rect 12307 15264 12623 15265
rect 12307 15200 12313 15264
rect 12377 15200 12393 15264
rect 12457 15200 12473 15264
rect 12537 15200 12553 15264
rect 12617 15200 12623 15264
rect 12307 15199 12623 15200
rect 17988 15264 18304 15265
rect 17988 15200 17994 15264
rect 18058 15200 18074 15264
rect 18138 15200 18154 15264
rect 18218 15200 18234 15264
rect 18298 15200 18304 15264
rect 17988 15199 18304 15200
rect 23669 15264 23985 15265
rect 23669 15200 23675 15264
rect 23739 15200 23755 15264
rect 23819 15200 23835 15264
rect 23899 15200 23915 15264
rect 23979 15200 23985 15264
rect 23669 15199 23985 15200
rect 4429 15058 4495 15061
rect 6637 15058 6703 15061
rect 4429 15056 6703 15058
rect 4429 15000 4434 15056
rect 4490 15000 6642 15056
rect 6698 15000 6703 15056
rect 4429 14998 6703 15000
rect 4429 14995 4495 14998
rect 6637 14995 6703 14998
rect 16430 14996 16436 15060
rect 16500 15058 16506 15060
rect 16757 15058 16823 15061
rect 16500 15056 16823 15058
rect 16500 15000 16762 15056
rect 16818 15000 16823 15056
rect 16500 14998 16823 15000
rect 16500 14996 16506 14998
rect 16757 14995 16823 14998
rect 3786 14720 4102 14721
rect 3786 14656 3792 14720
rect 3856 14656 3872 14720
rect 3936 14656 3952 14720
rect 4016 14656 4032 14720
rect 4096 14656 4102 14720
rect 3786 14655 4102 14656
rect 9467 14720 9783 14721
rect 9467 14656 9473 14720
rect 9537 14656 9553 14720
rect 9617 14656 9633 14720
rect 9697 14656 9713 14720
rect 9777 14656 9783 14720
rect 9467 14655 9783 14656
rect 15148 14720 15464 14721
rect 15148 14656 15154 14720
rect 15218 14656 15234 14720
rect 15298 14656 15314 14720
rect 15378 14656 15394 14720
rect 15458 14656 15464 14720
rect 15148 14655 15464 14656
rect 20829 14720 21145 14721
rect 20829 14656 20835 14720
rect 20899 14656 20915 14720
rect 20979 14656 20995 14720
rect 21059 14656 21075 14720
rect 21139 14656 21145 14720
rect 20829 14655 21145 14656
rect 6626 14176 6942 14177
rect 6626 14112 6632 14176
rect 6696 14112 6712 14176
rect 6776 14112 6792 14176
rect 6856 14112 6872 14176
rect 6936 14112 6942 14176
rect 6626 14111 6942 14112
rect 12307 14176 12623 14177
rect 12307 14112 12313 14176
rect 12377 14112 12393 14176
rect 12457 14112 12473 14176
rect 12537 14112 12553 14176
rect 12617 14112 12623 14176
rect 12307 14111 12623 14112
rect 17988 14176 18304 14177
rect 17988 14112 17994 14176
rect 18058 14112 18074 14176
rect 18138 14112 18154 14176
rect 18218 14112 18234 14176
rect 18298 14112 18304 14176
rect 17988 14111 18304 14112
rect 23669 14176 23985 14177
rect 23669 14112 23675 14176
rect 23739 14112 23755 14176
rect 23819 14112 23835 14176
rect 23899 14112 23915 14176
rect 23979 14112 23985 14176
rect 23669 14111 23985 14112
rect 5073 14106 5139 14109
rect 4662 14104 5139 14106
rect 4662 14048 5078 14104
rect 5134 14048 5139 14104
rect 4662 14046 5139 14048
rect 4521 13834 4587 13837
rect 4662 13834 4722 14046
rect 5073 14043 5139 14046
rect 4521 13832 4722 13834
rect 4521 13776 4526 13832
rect 4582 13776 4722 13832
rect 4521 13774 4722 13776
rect 15377 13834 15443 13837
rect 15694 13834 15700 13836
rect 15377 13832 15700 13834
rect 15377 13776 15382 13832
rect 15438 13776 15700 13832
rect 15377 13774 15700 13776
rect 4521 13771 4587 13774
rect 15377 13771 15443 13774
rect 15694 13772 15700 13774
rect 15764 13772 15770 13836
rect 19517 13834 19583 13837
rect 20110 13834 20116 13836
rect 19517 13832 20116 13834
rect 19517 13776 19522 13832
rect 19578 13776 20116 13832
rect 19517 13774 20116 13776
rect 19517 13771 19583 13774
rect 20110 13772 20116 13774
rect 20180 13772 20186 13836
rect 3786 13632 4102 13633
rect 3786 13568 3792 13632
rect 3856 13568 3872 13632
rect 3936 13568 3952 13632
rect 4016 13568 4032 13632
rect 4096 13568 4102 13632
rect 3786 13567 4102 13568
rect 9467 13632 9783 13633
rect 9467 13568 9473 13632
rect 9537 13568 9553 13632
rect 9617 13568 9633 13632
rect 9697 13568 9713 13632
rect 9777 13568 9783 13632
rect 9467 13567 9783 13568
rect 15148 13632 15464 13633
rect 15148 13568 15154 13632
rect 15218 13568 15234 13632
rect 15298 13568 15314 13632
rect 15378 13568 15394 13632
rect 15458 13568 15464 13632
rect 15148 13567 15464 13568
rect 20829 13632 21145 13633
rect 20829 13568 20835 13632
rect 20899 13568 20915 13632
rect 20979 13568 20995 13632
rect 21059 13568 21075 13632
rect 21139 13568 21145 13632
rect 20829 13567 21145 13568
rect 5165 13290 5231 13293
rect 6637 13290 6703 13293
rect 5165 13288 6703 13290
rect 5165 13232 5170 13288
rect 5226 13232 6642 13288
rect 6698 13232 6703 13288
rect 5165 13230 6703 13232
rect 5165 13227 5231 13230
rect 6637 13227 6703 13230
rect 17769 13290 17835 13293
rect 18229 13290 18295 13293
rect 17769 13288 18295 13290
rect 17769 13232 17774 13288
rect 17830 13232 18234 13288
rect 18290 13232 18295 13288
rect 17769 13230 18295 13232
rect 17769 13227 17835 13230
rect 18229 13227 18295 13230
rect 6626 13088 6942 13089
rect 6626 13024 6632 13088
rect 6696 13024 6712 13088
rect 6776 13024 6792 13088
rect 6856 13024 6872 13088
rect 6936 13024 6942 13088
rect 6626 13023 6942 13024
rect 12307 13088 12623 13089
rect 12307 13024 12313 13088
rect 12377 13024 12393 13088
rect 12457 13024 12473 13088
rect 12537 13024 12553 13088
rect 12617 13024 12623 13088
rect 12307 13023 12623 13024
rect 17988 13088 18304 13089
rect 17988 13024 17994 13088
rect 18058 13024 18074 13088
rect 18138 13024 18154 13088
rect 18218 13024 18234 13088
rect 18298 13024 18304 13088
rect 17988 13023 18304 13024
rect 23669 13088 23985 13089
rect 23669 13024 23675 13088
rect 23739 13024 23755 13088
rect 23819 13024 23835 13088
rect 23899 13024 23915 13088
rect 23979 13024 23985 13088
rect 23669 13023 23985 13024
rect 19701 12882 19767 12885
rect 20621 12882 20687 12885
rect 19701 12880 20687 12882
rect 19701 12824 19706 12880
rect 19762 12824 20626 12880
rect 20682 12824 20687 12880
rect 19701 12822 20687 12824
rect 19701 12819 19767 12822
rect 20621 12819 20687 12822
rect 4521 12610 4587 12613
rect 5022 12610 5028 12612
rect 4521 12608 5028 12610
rect 4521 12552 4526 12608
rect 4582 12552 5028 12608
rect 4521 12550 5028 12552
rect 4521 12547 4587 12550
rect 5022 12548 5028 12550
rect 5092 12548 5098 12612
rect 3786 12544 4102 12545
rect 3786 12480 3792 12544
rect 3856 12480 3872 12544
rect 3936 12480 3952 12544
rect 4016 12480 4032 12544
rect 4096 12480 4102 12544
rect 3786 12479 4102 12480
rect 9467 12544 9783 12545
rect 9467 12480 9473 12544
rect 9537 12480 9553 12544
rect 9617 12480 9633 12544
rect 9697 12480 9713 12544
rect 9777 12480 9783 12544
rect 9467 12479 9783 12480
rect 15148 12544 15464 12545
rect 15148 12480 15154 12544
rect 15218 12480 15234 12544
rect 15298 12480 15314 12544
rect 15378 12480 15394 12544
rect 15458 12480 15464 12544
rect 15148 12479 15464 12480
rect 20829 12544 21145 12545
rect 20829 12480 20835 12544
rect 20899 12480 20915 12544
rect 20979 12480 20995 12544
rect 21059 12480 21075 12544
rect 21139 12480 21145 12544
rect 20829 12479 21145 12480
rect 12893 12474 12959 12477
rect 15009 12474 15075 12477
rect 12893 12472 15075 12474
rect 12893 12416 12898 12472
rect 12954 12416 15014 12472
rect 15070 12416 15075 12472
rect 12893 12414 15075 12416
rect 12893 12411 12959 12414
rect 15009 12411 15075 12414
rect 4286 12276 4292 12340
rect 4356 12338 4362 12340
rect 6821 12338 6887 12341
rect 4356 12336 6887 12338
rect 4356 12280 6826 12336
rect 6882 12280 6887 12336
rect 4356 12278 6887 12280
rect 4356 12276 4362 12278
rect 6821 12275 6887 12278
rect 14549 12338 14615 12341
rect 19425 12338 19491 12341
rect 14549 12336 19491 12338
rect 14549 12280 14554 12336
rect 14610 12280 19430 12336
rect 19486 12280 19491 12336
rect 14549 12278 19491 12280
rect 14549 12275 14615 12278
rect 19425 12275 19491 12278
rect 6310 12140 6316 12204
rect 6380 12202 6386 12204
rect 12065 12202 12131 12205
rect 12934 12202 12940 12204
rect 6380 12142 7114 12202
rect 6380 12140 6386 12142
rect 7054 12066 7114 12142
rect 12065 12200 12940 12202
rect 12065 12144 12070 12200
rect 12126 12144 12940 12200
rect 12065 12142 12940 12144
rect 12065 12139 12131 12142
rect 12934 12140 12940 12142
rect 13004 12202 13010 12204
rect 15653 12202 15719 12205
rect 20069 12202 20135 12205
rect 13004 12200 20135 12202
rect 13004 12144 15658 12200
rect 15714 12144 20074 12200
rect 20130 12144 20135 12200
rect 13004 12142 20135 12144
rect 13004 12140 13010 12142
rect 15653 12139 15719 12142
rect 20069 12139 20135 12142
rect 8477 12068 8543 12069
rect 8477 12066 8524 12068
rect 7054 12064 8524 12066
rect 8588 12066 8594 12068
rect 9765 12066 9831 12069
rect 8588 12064 9831 12066
rect 7054 12008 8482 12064
rect 8588 12008 9770 12064
rect 9826 12008 9831 12064
rect 7054 12006 8524 12008
rect 8477 12004 8524 12006
rect 8588 12006 9831 12008
rect 8588 12004 8594 12006
rect 8477 12003 8543 12004
rect 9765 12003 9831 12006
rect 14641 12066 14707 12069
rect 15929 12066 15995 12069
rect 14641 12064 15995 12066
rect 14641 12008 14646 12064
rect 14702 12008 15934 12064
rect 15990 12008 15995 12064
rect 14641 12006 15995 12008
rect 14641 12003 14707 12006
rect 15929 12003 15995 12006
rect 6626 12000 6942 12001
rect 6626 11936 6632 12000
rect 6696 11936 6712 12000
rect 6776 11936 6792 12000
rect 6856 11936 6872 12000
rect 6936 11936 6942 12000
rect 6626 11935 6942 11936
rect 12307 12000 12623 12001
rect 12307 11936 12313 12000
rect 12377 11936 12393 12000
rect 12457 11936 12473 12000
rect 12537 11936 12553 12000
rect 12617 11936 12623 12000
rect 12307 11935 12623 11936
rect 17988 12000 18304 12001
rect 17988 11936 17994 12000
rect 18058 11936 18074 12000
rect 18138 11936 18154 12000
rect 18218 11936 18234 12000
rect 18298 11936 18304 12000
rect 17988 11935 18304 11936
rect 23669 12000 23985 12001
rect 23669 11936 23675 12000
rect 23739 11936 23755 12000
rect 23819 11936 23835 12000
rect 23899 11936 23915 12000
rect 23979 11936 23985 12000
rect 23669 11935 23985 11936
rect 4245 11932 4311 11933
rect 8109 11932 8175 11933
rect 4245 11930 4292 11932
rect 4200 11928 4292 11930
rect 4200 11872 4250 11928
rect 4200 11870 4292 11872
rect 4245 11868 4292 11870
rect 4356 11868 4362 11932
rect 8109 11928 8156 11932
rect 8220 11930 8226 11932
rect 8109 11872 8114 11928
rect 8109 11868 8156 11872
rect 8220 11870 8266 11930
rect 8220 11868 8226 11870
rect 4245 11867 4311 11868
rect 8109 11867 8175 11868
rect 16941 11794 17007 11797
rect 18873 11794 18939 11797
rect 16941 11792 18939 11794
rect 16941 11736 16946 11792
rect 17002 11736 18878 11792
rect 18934 11736 18939 11792
rect 16941 11734 18939 11736
rect 16941 11731 17007 11734
rect 18873 11731 18939 11734
rect 14825 11658 14891 11661
rect 17033 11658 17099 11661
rect 18781 11658 18847 11661
rect 14825 11656 18847 11658
rect 14825 11600 14830 11656
rect 14886 11600 17038 11656
rect 17094 11600 18786 11656
rect 18842 11600 18847 11656
rect 14825 11598 18847 11600
rect 14825 11595 14891 11598
rect 17033 11595 17099 11598
rect 18781 11595 18847 11598
rect 19057 11658 19123 11661
rect 22185 11658 22251 11661
rect 19057 11656 22251 11658
rect 19057 11600 19062 11656
rect 19118 11600 22190 11656
rect 22246 11600 22251 11656
rect 19057 11598 22251 11600
rect 19057 11595 19123 11598
rect 22185 11595 22251 11598
rect 3786 11456 4102 11457
rect 3786 11392 3792 11456
rect 3856 11392 3872 11456
rect 3936 11392 3952 11456
rect 4016 11392 4032 11456
rect 4096 11392 4102 11456
rect 3786 11391 4102 11392
rect 9467 11456 9783 11457
rect 9467 11392 9473 11456
rect 9537 11392 9553 11456
rect 9617 11392 9633 11456
rect 9697 11392 9713 11456
rect 9777 11392 9783 11456
rect 9467 11391 9783 11392
rect 15148 11456 15464 11457
rect 15148 11392 15154 11456
rect 15218 11392 15234 11456
rect 15298 11392 15314 11456
rect 15378 11392 15394 11456
rect 15458 11392 15464 11456
rect 15148 11391 15464 11392
rect 20829 11456 21145 11457
rect 20829 11392 20835 11456
rect 20899 11392 20915 11456
rect 20979 11392 20995 11456
rect 21059 11392 21075 11456
rect 21139 11392 21145 11456
rect 20829 11391 21145 11392
rect 7557 11252 7623 11253
rect 7557 11248 7604 11252
rect 7668 11250 7674 11252
rect 14733 11250 14799 11253
rect 16021 11250 16087 11253
rect 7557 11192 7562 11248
rect 7557 11188 7604 11192
rect 7668 11190 7714 11250
rect 14733 11248 16087 11250
rect 14733 11192 14738 11248
rect 14794 11192 16026 11248
rect 16082 11192 16087 11248
rect 14733 11190 16087 11192
rect 7668 11188 7674 11190
rect 7557 11187 7623 11188
rect 14733 11187 14799 11190
rect 16021 11187 16087 11190
rect 14825 11114 14891 11117
rect 19241 11114 19307 11117
rect 14825 11112 19307 11114
rect 14825 11056 14830 11112
rect 14886 11056 19246 11112
rect 19302 11056 19307 11112
rect 14825 11054 19307 11056
rect 14825 11051 14891 11054
rect 19241 11051 19307 11054
rect 19701 11114 19767 11117
rect 20713 11114 20779 11117
rect 19701 11112 20779 11114
rect 19701 11056 19706 11112
rect 19762 11056 20718 11112
rect 20774 11056 20779 11112
rect 19701 11054 20779 11056
rect 19701 11051 19767 11054
rect 20713 11051 20779 11054
rect 20529 10978 20595 10981
rect 20989 10978 21055 10981
rect 20529 10976 21055 10978
rect 20529 10920 20534 10976
rect 20590 10920 20994 10976
rect 21050 10920 21055 10976
rect 20529 10918 21055 10920
rect 20529 10915 20595 10918
rect 20989 10915 21055 10918
rect 6626 10912 6942 10913
rect 6626 10848 6632 10912
rect 6696 10848 6712 10912
rect 6776 10848 6792 10912
rect 6856 10848 6872 10912
rect 6936 10848 6942 10912
rect 6626 10847 6942 10848
rect 12307 10912 12623 10913
rect 12307 10848 12313 10912
rect 12377 10848 12393 10912
rect 12457 10848 12473 10912
rect 12537 10848 12553 10912
rect 12617 10848 12623 10912
rect 12307 10847 12623 10848
rect 17988 10912 18304 10913
rect 17988 10848 17994 10912
rect 18058 10848 18074 10912
rect 18138 10848 18154 10912
rect 18218 10848 18234 10912
rect 18298 10848 18304 10912
rect 17988 10847 18304 10848
rect 23669 10912 23985 10913
rect 23669 10848 23675 10912
rect 23739 10848 23755 10912
rect 23819 10848 23835 10912
rect 23899 10848 23915 10912
rect 23979 10848 23985 10912
rect 23669 10847 23985 10848
rect 15285 10842 15351 10845
rect 16389 10842 16455 10845
rect 17125 10842 17191 10845
rect 15285 10840 17191 10842
rect 15285 10784 15290 10840
rect 15346 10784 16394 10840
rect 16450 10784 17130 10840
rect 17186 10784 17191 10840
rect 15285 10782 17191 10784
rect 15285 10779 15351 10782
rect 16389 10779 16455 10782
rect 17125 10779 17191 10782
rect 5533 10706 5599 10709
rect 8753 10706 8819 10709
rect 9397 10706 9463 10709
rect 5533 10704 8819 10706
rect 5533 10648 5538 10704
rect 5594 10648 8758 10704
rect 8814 10648 8819 10704
rect 5533 10646 8819 10648
rect 5533 10643 5599 10646
rect 8753 10643 8819 10646
rect 9262 10704 9463 10706
rect 9262 10648 9402 10704
rect 9458 10648 9463 10704
rect 9262 10646 9463 10648
rect 3233 10570 3299 10573
rect 8017 10570 8083 10573
rect 9262 10570 9322 10646
rect 9397 10643 9463 10646
rect 17309 10706 17375 10709
rect 21265 10706 21331 10709
rect 17309 10704 21331 10706
rect 17309 10648 17314 10704
rect 17370 10648 21270 10704
rect 21326 10648 21331 10704
rect 17309 10646 21331 10648
rect 17309 10643 17375 10646
rect 21265 10643 21331 10646
rect 3233 10568 9322 10570
rect 3233 10512 3238 10568
rect 3294 10512 8022 10568
rect 8078 10512 9322 10568
rect 3233 10510 9322 10512
rect 3233 10507 3299 10510
rect 8017 10507 8083 10510
rect 3786 10368 4102 10369
rect 3786 10304 3792 10368
rect 3856 10304 3872 10368
rect 3936 10304 3952 10368
rect 4016 10304 4032 10368
rect 4096 10304 4102 10368
rect 3786 10303 4102 10304
rect 9262 10162 9322 10510
rect 9467 10368 9783 10369
rect 9467 10304 9473 10368
rect 9537 10304 9553 10368
rect 9617 10304 9633 10368
rect 9697 10304 9713 10368
rect 9777 10304 9783 10368
rect 9467 10303 9783 10304
rect 15148 10368 15464 10369
rect 15148 10304 15154 10368
rect 15218 10304 15234 10368
rect 15298 10304 15314 10368
rect 15378 10304 15394 10368
rect 15458 10304 15464 10368
rect 15148 10303 15464 10304
rect 20829 10368 21145 10369
rect 20829 10304 20835 10368
rect 20899 10304 20915 10368
rect 20979 10304 20995 10368
rect 21059 10304 21075 10368
rect 21139 10304 21145 10368
rect 20829 10303 21145 10304
rect 9489 10162 9555 10165
rect 9262 10160 9555 10162
rect 9262 10104 9494 10160
rect 9550 10104 9555 10160
rect 9262 10102 9555 10104
rect 9489 10099 9555 10102
rect 12617 10162 12683 10165
rect 16481 10162 16547 10165
rect 12617 10160 16547 10162
rect 12617 10104 12622 10160
rect 12678 10104 16486 10160
rect 16542 10104 16547 10160
rect 12617 10102 16547 10104
rect 12617 10099 12683 10102
rect 16481 10099 16547 10102
rect 20345 10162 20411 10165
rect 20897 10162 20963 10165
rect 20345 10160 20963 10162
rect 20345 10104 20350 10160
rect 20406 10104 20902 10160
rect 20958 10104 20963 10160
rect 20345 10102 20963 10104
rect 20345 10099 20411 10102
rect 20897 10099 20963 10102
rect 6729 10026 6795 10029
rect 8477 10026 8543 10029
rect 6729 10024 8543 10026
rect 6729 9968 6734 10024
rect 6790 9968 8482 10024
rect 8538 9968 8543 10024
rect 6729 9966 8543 9968
rect 6729 9963 6795 9966
rect 8477 9963 8543 9966
rect 15285 10026 15351 10029
rect 16481 10026 16547 10029
rect 15285 10024 16547 10026
rect 15285 9968 15290 10024
rect 15346 9968 16486 10024
rect 16542 9968 16547 10024
rect 15285 9966 16547 9968
rect 15285 9963 15351 9966
rect 16481 9963 16547 9966
rect 12893 9892 12959 9893
rect 12893 9890 12940 9892
rect 12848 9888 12940 9890
rect 12848 9832 12898 9888
rect 12848 9830 12940 9832
rect 12893 9828 12940 9830
rect 13004 9828 13010 9892
rect 14457 9890 14523 9893
rect 17125 9890 17191 9893
rect 14457 9888 17191 9890
rect 14457 9832 14462 9888
rect 14518 9832 17130 9888
rect 17186 9832 17191 9888
rect 14457 9830 17191 9832
rect 12893 9827 12959 9828
rect 14457 9827 14523 9830
rect 17125 9827 17191 9830
rect 6626 9824 6942 9825
rect 6626 9760 6632 9824
rect 6696 9760 6712 9824
rect 6776 9760 6792 9824
rect 6856 9760 6872 9824
rect 6936 9760 6942 9824
rect 6626 9759 6942 9760
rect 12307 9824 12623 9825
rect 12307 9760 12313 9824
rect 12377 9760 12393 9824
rect 12457 9760 12473 9824
rect 12537 9760 12553 9824
rect 12617 9760 12623 9824
rect 12307 9759 12623 9760
rect 17988 9824 18304 9825
rect 17988 9760 17994 9824
rect 18058 9760 18074 9824
rect 18138 9760 18154 9824
rect 18218 9760 18234 9824
rect 18298 9760 18304 9824
rect 17988 9759 18304 9760
rect 23669 9824 23985 9825
rect 23669 9760 23675 9824
rect 23739 9760 23755 9824
rect 23819 9760 23835 9824
rect 23899 9760 23915 9824
rect 23979 9760 23985 9824
rect 23669 9759 23985 9760
rect 8385 9756 8451 9757
rect 9305 9756 9371 9757
rect 10961 9756 11027 9757
rect 8334 9754 8340 9756
rect 8294 9694 8340 9754
rect 8404 9752 8451 9756
rect 9254 9754 9260 9756
rect 8446 9696 8451 9752
rect 8334 9692 8340 9694
rect 8404 9692 8451 9696
rect 9214 9694 9260 9754
rect 9324 9752 9371 9756
rect 10910 9754 10916 9756
rect 9366 9696 9371 9752
rect 9254 9692 9260 9694
rect 9324 9692 9371 9696
rect 10870 9694 10916 9754
rect 10980 9752 11027 9756
rect 11022 9696 11027 9752
rect 10910 9692 10916 9694
rect 10980 9692 11027 9696
rect 8385 9691 8451 9692
rect 9305 9691 9371 9692
rect 10961 9691 11027 9692
rect 18597 9754 18663 9757
rect 19885 9754 19951 9757
rect 18597 9752 19951 9754
rect 18597 9696 18602 9752
rect 18658 9696 19890 9752
rect 19946 9696 19951 9752
rect 18597 9694 19951 9696
rect 18597 9691 18663 9694
rect 19885 9691 19951 9694
rect 12433 9618 12499 9621
rect 14365 9618 14431 9621
rect 16481 9618 16547 9621
rect 12433 9616 16547 9618
rect 12433 9560 12438 9616
rect 12494 9560 14370 9616
rect 14426 9560 16486 9616
rect 16542 9560 16547 9616
rect 12433 9558 16547 9560
rect 12433 9555 12499 9558
rect 14365 9555 14431 9558
rect 16481 9555 16547 9558
rect 18873 9618 18939 9621
rect 20529 9618 20595 9621
rect 18873 9616 20595 9618
rect 18873 9560 18878 9616
rect 18934 9560 20534 9616
rect 20590 9560 20595 9616
rect 18873 9558 20595 9560
rect 18873 9555 18939 9558
rect 20529 9555 20595 9558
rect 4337 9482 4403 9485
rect 7005 9482 7071 9485
rect 4337 9480 7071 9482
rect 4337 9424 4342 9480
rect 4398 9424 7010 9480
rect 7066 9424 7071 9480
rect 4337 9422 7071 9424
rect 4337 9419 4403 9422
rect 7005 9419 7071 9422
rect 7414 9420 7420 9484
rect 7484 9482 7490 9484
rect 11237 9482 11303 9485
rect 7484 9480 11303 9482
rect 7484 9424 11242 9480
rect 11298 9424 11303 9480
rect 7484 9422 11303 9424
rect 7484 9420 7490 9422
rect 11237 9419 11303 9422
rect 12065 9482 12131 9485
rect 14457 9482 14523 9485
rect 12065 9480 14523 9482
rect 12065 9424 12070 9480
rect 12126 9424 14462 9480
rect 14518 9424 14523 9480
rect 12065 9422 14523 9424
rect 12065 9419 12131 9422
rect 14457 9419 14523 9422
rect 15377 9482 15443 9485
rect 17125 9482 17191 9485
rect 17677 9482 17743 9485
rect 15377 9480 17743 9482
rect 15377 9424 15382 9480
rect 15438 9424 17130 9480
rect 17186 9424 17682 9480
rect 17738 9424 17743 9480
rect 15377 9422 17743 9424
rect 15377 9419 15443 9422
rect 17125 9419 17191 9422
rect 17677 9419 17743 9422
rect 20069 9482 20135 9485
rect 20294 9482 20300 9484
rect 20069 9480 20300 9482
rect 20069 9424 20074 9480
rect 20130 9424 20300 9480
rect 20069 9422 20300 9424
rect 20069 9419 20135 9422
rect 20294 9420 20300 9422
rect 20364 9420 20370 9484
rect 7833 9346 7899 9349
rect 7966 9346 7972 9348
rect 7833 9344 7972 9346
rect 7833 9288 7838 9344
rect 7894 9288 7972 9344
rect 7833 9286 7972 9288
rect 7833 9283 7899 9286
rect 7966 9284 7972 9286
rect 8036 9284 8042 9348
rect 17953 9346 18019 9349
rect 20345 9346 20411 9349
rect 20529 9346 20595 9349
rect 17953 9344 20595 9346
rect 17953 9288 17958 9344
rect 18014 9288 20350 9344
rect 20406 9288 20534 9344
rect 20590 9288 20595 9344
rect 17953 9286 20595 9288
rect 17953 9283 18019 9286
rect 20345 9283 20411 9286
rect 20529 9283 20595 9286
rect 3786 9280 4102 9281
rect 3786 9216 3792 9280
rect 3856 9216 3872 9280
rect 3936 9216 3952 9280
rect 4016 9216 4032 9280
rect 4096 9216 4102 9280
rect 3786 9215 4102 9216
rect 9467 9280 9783 9281
rect 9467 9216 9473 9280
rect 9537 9216 9553 9280
rect 9617 9216 9633 9280
rect 9697 9216 9713 9280
rect 9777 9216 9783 9280
rect 9467 9215 9783 9216
rect 15148 9280 15464 9281
rect 15148 9216 15154 9280
rect 15218 9216 15234 9280
rect 15298 9216 15314 9280
rect 15378 9216 15394 9280
rect 15458 9216 15464 9280
rect 15148 9215 15464 9216
rect 20829 9280 21145 9281
rect 20829 9216 20835 9280
rect 20899 9216 20915 9280
rect 20979 9216 20995 9280
rect 21059 9216 21075 9280
rect 21139 9216 21145 9280
rect 20829 9215 21145 9216
rect 10133 9210 10199 9213
rect 14825 9210 14891 9213
rect 16481 9212 16547 9213
rect 16430 9210 16436 9212
rect 10133 9208 14891 9210
rect 10133 9152 10138 9208
rect 10194 9152 14830 9208
rect 14886 9152 14891 9208
rect 10133 9150 14891 9152
rect 16390 9150 16436 9210
rect 16500 9208 16547 9212
rect 16542 9152 16547 9208
rect 10133 9147 10199 9150
rect 14825 9147 14891 9150
rect 16430 9148 16436 9150
rect 16500 9148 16547 9152
rect 16481 9147 16547 9148
rect 17217 9210 17283 9213
rect 18689 9210 18755 9213
rect 17217 9208 18755 9210
rect 17217 9152 17222 9208
rect 17278 9152 18694 9208
rect 18750 9152 18755 9208
rect 17217 9150 18755 9152
rect 17217 9147 17283 9150
rect 18689 9147 18755 9150
rect 14549 9074 14615 9077
rect 22185 9074 22251 9077
rect 14549 9072 22251 9074
rect 14549 9016 14554 9072
rect 14610 9016 22190 9072
rect 22246 9016 22251 9072
rect 14549 9014 22251 9016
rect 14549 9011 14615 9014
rect 22185 9011 22251 9014
rect 4889 8938 4955 8941
rect 5441 8938 5507 8941
rect 6361 8938 6427 8941
rect 4889 8936 6427 8938
rect 4889 8880 4894 8936
rect 4950 8880 5446 8936
rect 5502 8880 6366 8936
rect 6422 8880 6427 8936
rect 4889 8878 6427 8880
rect 4889 8875 4955 8878
rect 5441 8875 5507 8878
rect 6361 8875 6427 8878
rect 11421 8938 11487 8941
rect 18505 8938 18571 8941
rect 11421 8936 18571 8938
rect 11421 8880 11426 8936
rect 11482 8880 18510 8936
rect 18566 8880 18571 8936
rect 11421 8878 18571 8880
rect 11421 8875 11487 8878
rect 18505 8875 18571 8878
rect 9857 8802 9923 8805
rect 10317 8802 10383 8805
rect 9857 8800 10383 8802
rect 9857 8744 9862 8800
rect 9918 8744 10322 8800
rect 10378 8744 10383 8800
rect 9857 8742 10383 8744
rect 9857 8739 9923 8742
rect 10317 8739 10383 8742
rect 6626 8736 6942 8737
rect 6626 8672 6632 8736
rect 6696 8672 6712 8736
rect 6776 8672 6792 8736
rect 6856 8672 6872 8736
rect 6936 8672 6942 8736
rect 6626 8671 6942 8672
rect 12307 8736 12623 8737
rect 12307 8672 12313 8736
rect 12377 8672 12393 8736
rect 12457 8672 12473 8736
rect 12537 8672 12553 8736
rect 12617 8672 12623 8736
rect 12307 8671 12623 8672
rect 17988 8736 18304 8737
rect 17988 8672 17994 8736
rect 18058 8672 18074 8736
rect 18138 8672 18154 8736
rect 18218 8672 18234 8736
rect 18298 8672 18304 8736
rect 17988 8671 18304 8672
rect 23669 8736 23985 8737
rect 23669 8672 23675 8736
rect 23739 8672 23755 8736
rect 23819 8672 23835 8736
rect 23899 8672 23915 8736
rect 23979 8672 23985 8736
rect 23669 8671 23985 8672
rect 13629 8666 13695 8669
rect 13997 8666 14063 8669
rect 13629 8664 14063 8666
rect 13629 8608 13634 8664
rect 13690 8608 14002 8664
rect 14058 8608 14063 8664
rect 13629 8606 14063 8608
rect 13629 8603 13695 8606
rect 13997 8603 14063 8606
rect 11881 8530 11947 8533
rect 13905 8530 13971 8533
rect 11881 8528 13971 8530
rect 11881 8472 11886 8528
rect 11942 8472 13910 8528
rect 13966 8472 13971 8528
rect 11881 8470 13971 8472
rect 11881 8467 11947 8470
rect 13905 8467 13971 8470
rect 14273 8530 14339 8533
rect 14457 8530 14523 8533
rect 14273 8528 14523 8530
rect 14273 8472 14278 8528
rect 14334 8472 14462 8528
rect 14518 8472 14523 8528
rect 14273 8470 14523 8472
rect 14273 8467 14339 8470
rect 14457 8467 14523 8470
rect 7649 8394 7715 8397
rect 7782 8394 7788 8396
rect 7649 8392 7788 8394
rect 7649 8336 7654 8392
rect 7710 8336 7788 8392
rect 7649 8334 7788 8336
rect 7649 8331 7715 8334
rect 7782 8332 7788 8334
rect 7852 8332 7858 8396
rect 19057 8394 19123 8397
rect 20805 8394 20871 8397
rect 19057 8392 20871 8394
rect 19057 8336 19062 8392
rect 19118 8336 20810 8392
rect 20866 8336 20871 8392
rect 19057 8334 20871 8336
rect 19057 8331 19123 8334
rect 20805 8331 20871 8334
rect 3786 8192 4102 8193
rect 3786 8128 3792 8192
rect 3856 8128 3872 8192
rect 3936 8128 3952 8192
rect 4016 8128 4032 8192
rect 4096 8128 4102 8192
rect 3786 8127 4102 8128
rect 9467 8192 9783 8193
rect 9467 8128 9473 8192
rect 9537 8128 9553 8192
rect 9617 8128 9633 8192
rect 9697 8128 9713 8192
rect 9777 8128 9783 8192
rect 9467 8127 9783 8128
rect 15148 8192 15464 8193
rect 15148 8128 15154 8192
rect 15218 8128 15234 8192
rect 15298 8128 15314 8192
rect 15378 8128 15394 8192
rect 15458 8128 15464 8192
rect 15148 8127 15464 8128
rect 20829 8192 21145 8193
rect 20829 8128 20835 8192
rect 20899 8128 20915 8192
rect 20979 8128 20995 8192
rect 21059 8128 21075 8192
rect 21139 8128 21145 8192
rect 20829 8127 21145 8128
rect 20110 8060 20116 8124
rect 20180 8122 20186 8124
rect 20253 8122 20319 8125
rect 20180 8120 20319 8122
rect 20180 8064 20258 8120
rect 20314 8064 20319 8120
rect 20180 8062 20319 8064
rect 20180 8060 20186 8062
rect 20253 8059 20319 8062
rect 10910 7924 10916 7988
rect 10980 7986 10986 7988
rect 16849 7986 16915 7989
rect 10980 7984 16915 7986
rect 10980 7928 16854 7984
rect 16910 7928 16915 7984
rect 10980 7926 16915 7928
rect 10980 7924 10986 7926
rect 16849 7923 16915 7926
rect 7189 7850 7255 7853
rect 8385 7850 8451 7853
rect 7189 7848 8451 7850
rect 7189 7792 7194 7848
rect 7250 7792 8390 7848
rect 8446 7792 8451 7848
rect 7189 7790 8451 7792
rect 7189 7787 7255 7790
rect 8385 7787 8451 7790
rect 17585 7850 17651 7853
rect 18045 7850 18111 7853
rect 17585 7848 18111 7850
rect 17585 7792 17590 7848
rect 17646 7792 18050 7848
rect 18106 7792 18111 7848
rect 17585 7790 18111 7792
rect 17585 7787 17651 7790
rect 18045 7787 18111 7790
rect 13077 7714 13143 7717
rect 16297 7714 16363 7717
rect 16941 7714 17007 7717
rect 17217 7714 17283 7717
rect 13077 7712 17283 7714
rect 13077 7656 13082 7712
rect 13138 7656 16302 7712
rect 16358 7656 16946 7712
rect 17002 7656 17222 7712
rect 17278 7656 17283 7712
rect 13077 7654 17283 7656
rect 13077 7651 13143 7654
rect 16297 7651 16363 7654
rect 16941 7651 17007 7654
rect 17217 7651 17283 7654
rect 6626 7648 6942 7649
rect 6626 7584 6632 7648
rect 6696 7584 6712 7648
rect 6776 7584 6792 7648
rect 6856 7584 6872 7648
rect 6936 7584 6942 7648
rect 6626 7583 6942 7584
rect 12307 7648 12623 7649
rect 12307 7584 12313 7648
rect 12377 7584 12393 7648
rect 12457 7584 12473 7648
rect 12537 7584 12553 7648
rect 12617 7584 12623 7648
rect 12307 7583 12623 7584
rect 17988 7648 18304 7649
rect 17988 7584 17994 7648
rect 18058 7584 18074 7648
rect 18138 7584 18154 7648
rect 18218 7584 18234 7648
rect 18298 7584 18304 7648
rect 17988 7583 18304 7584
rect 23669 7648 23985 7649
rect 23669 7584 23675 7648
rect 23739 7584 23755 7648
rect 23819 7584 23835 7648
rect 23899 7584 23915 7648
rect 23979 7584 23985 7648
rect 23669 7583 23985 7584
rect 3366 7380 3372 7444
rect 3436 7442 3442 7444
rect 4797 7442 4863 7445
rect 3436 7440 4863 7442
rect 3436 7384 4802 7440
rect 4858 7384 4863 7440
rect 3436 7382 4863 7384
rect 3436 7380 3442 7382
rect 4797 7379 4863 7382
rect 14641 7442 14707 7445
rect 18965 7442 19031 7445
rect 19977 7442 20043 7445
rect 14641 7440 20043 7442
rect 14641 7384 14646 7440
rect 14702 7384 18970 7440
rect 19026 7384 19982 7440
rect 20038 7384 20043 7440
rect 14641 7382 20043 7384
rect 14641 7379 14707 7382
rect 18965 7379 19031 7382
rect 19977 7379 20043 7382
rect 19793 7306 19859 7309
rect 20805 7306 20871 7309
rect 21449 7306 21515 7309
rect 19793 7304 21515 7306
rect 19793 7248 19798 7304
rect 19854 7248 20810 7304
rect 20866 7248 21454 7304
rect 21510 7248 21515 7304
rect 19793 7246 21515 7248
rect 19793 7243 19859 7246
rect 20805 7243 20871 7246
rect 21449 7243 21515 7246
rect 3786 7104 4102 7105
rect 3786 7040 3792 7104
rect 3856 7040 3872 7104
rect 3936 7040 3952 7104
rect 4016 7040 4032 7104
rect 4096 7040 4102 7104
rect 3786 7039 4102 7040
rect 9467 7104 9783 7105
rect 9467 7040 9473 7104
rect 9537 7040 9553 7104
rect 9617 7040 9633 7104
rect 9697 7040 9713 7104
rect 9777 7040 9783 7104
rect 9467 7039 9783 7040
rect 15148 7104 15464 7105
rect 15148 7040 15154 7104
rect 15218 7040 15234 7104
rect 15298 7040 15314 7104
rect 15378 7040 15394 7104
rect 15458 7040 15464 7104
rect 15148 7039 15464 7040
rect 20829 7104 21145 7105
rect 20829 7040 20835 7104
rect 20899 7040 20915 7104
rect 20979 7040 20995 7104
rect 21059 7040 21075 7104
rect 21139 7040 21145 7104
rect 20829 7039 21145 7040
rect 16021 6898 16087 6901
rect 17677 6898 17743 6901
rect 16021 6896 17743 6898
rect 16021 6840 16026 6896
rect 16082 6840 17682 6896
rect 17738 6840 17743 6896
rect 16021 6838 17743 6840
rect 16021 6835 16087 6838
rect 17677 6835 17743 6838
rect 4797 6762 4863 6765
rect 5993 6762 6059 6765
rect 4797 6760 6059 6762
rect 4797 6704 4802 6760
rect 4858 6704 5998 6760
rect 6054 6704 6059 6760
rect 4797 6702 6059 6704
rect 4797 6699 4863 6702
rect 5993 6699 6059 6702
rect 18689 6762 18755 6765
rect 19149 6762 19215 6765
rect 19333 6762 19399 6765
rect 18689 6760 19399 6762
rect 18689 6704 18694 6760
rect 18750 6704 19154 6760
rect 19210 6704 19338 6760
rect 19394 6704 19399 6760
rect 18689 6702 19399 6704
rect 18689 6699 18755 6702
rect 19149 6699 19215 6702
rect 19333 6699 19399 6702
rect 18413 6626 18479 6629
rect 21725 6626 21791 6629
rect 18413 6624 21791 6626
rect 18413 6568 18418 6624
rect 18474 6568 21730 6624
rect 21786 6568 21791 6624
rect 18413 6566 21791 6568
rect 18413 6563 18479 6566
rect 21725 6563 21791 6566
rect 6626 6560 6942 6561
rect 6626 6496 6632 6560
rect 6696 6496 6712 6560
rect 6776 6496 6792 6560
rect 6856 6496 6872 6560
rect 6936 6496 6942 6560
rect 6626 6495 6942 6496
rect 12307 6560 12623 6561
rect 12307 6496 12313 6560
rect 12377 6496 12393 6560
rect 12457 6496 12473 6560
rect 12537 6496 12553 6560
rect 12617 6496 12623 6560
rect 12307 6495 12623 6496
rect 17988 6560 18304 6561
rect 17988 6496 17994 6560
rect 18058 6496 18074 6560
rect 18138 6496 18154 6560
rect 18218 6496 18234 6560
rect 18298 6496 18304 6560
rect 17988 6495 18304 6496
rect 23669 6560 23985 6561
rect 23669 6496 23675 6560
rect 23739 6496 23755 6560
rect 23819 6496 23835 6560
rect 23899 6496 23915 6560
rect 23979 6496 23985 6560
rect 23669 6495 23985 6496
rect 13905 6490 13971 6493
rect 15694 6490 15700 6492
rect 13905 6488 15700 6490
rect 13905 6432 13910 6488
rect 13966 6432 15700 6488
rect 13905 6430 15700 6432
rect 13905 6427 13971 6430
rect 15694 6428 15700 6430
rect 15764 6490 15770 6492
rect 17677 6490 17743 6493
rect 15764 6488 17743 6490
rect 15764 6432 17682 6488
rect 17738 6432 17743 6488
rect 15764 6430 17743 6432
rect 15764 6428 15770 6430
rect 17677 6427 17743 6430
rect 18781 6490 18847 6493
rect 21173 6490 21239 6493
rect 18781 6488 21239 6490
rect 18781 6432 18786 6488
rect 18842 6432 21178 6488
rect 21234 6432 21239 6488
rect 18781 6430 21239 6432
rect 18781 6427 18847 6430
rect 21173 6427 21239 6430
rect 18045 6354 18111 6357
rect 19057 6354 19123 6357
rect 18045 6352 19123 6354
rect 18045 6296 18050 6352
rect 18106 6296 19062 6352
rect 19118 6296 19123 6352
rect 18045 6294 19123 6296
rect 18045 6291 18111 6294
rect 19057 6291 19123 6294
rect 3786 6016 4102 6017
rect 3786 5952 3792 6016
rect 3856 5952 3872 6016
rect 3936 5952 3952 6016
rect 4016 5952 4032 6016
rect 4096 5952 4102 6016
rect 3786 5951 4102 5952
rect 9467 6016 9783 6017
rect 9467 5952 9473 6016
rect 9537 5952 9553 6016
rect 9617 5952 9633 6016
rect 9697 5952 9713 6016
rect 9777 5952 9783 6016
rect 9467 5951 9783 5952
rect 15148 6016 15464 6017
rect 15148 5952 15154 6016
rect 15218 5952 15234 6016
rect 15298 5952 15314 6016
rect 15378 5952 15394 6016
rect 15458 5952 15464 6016
rect 15148 5951 15464 5952
rect 20829 6016 21145 6017
rect 20829 5952 20835 6016
rect 20899 5952 20915 6016
rect 20979 5952 20995 6016
rect 21059 5952 21075 6016
rect 21139 5952 21145 6016
rect 20829 5951 21145 5952
rect 9254 5748 9260 5812
rect 9324 5810 9330 5812
rect 9489 5810 9555 5813
rect 9324 5808 9555 5810
rect 9324 5752 9494 5808
rect 9550 5752 9555 5808
rect 9324 5750 9555 5752
rect 9324 5748 9330 5750
rect 9489 5747 9555 5750
rect 16757 5810 16823 5813
rect 19149 5810 19215 5813
rect 16757 5808 19215 5810
rect 16757 5752 16762 5808
rect 16818 5752 19154 5808
rect 19210 5752 19215 5808
rect 16757 5750 19215 5752
rect 16757 5747 16823 5750
rect 19149 5747 19215 5750
rect 20345 5540 20411 5541
rect 20294 5538 20300 5540
rect 20254 5478 20300 5538
rect 20364 5536 20411 5540
rect 20406 5480 20411 5536
rect 20294 5476 20300 5478
rect 20364 5476 20411 5480
rect 20345 5475 20411 5476
rect 6626 5472 6942 5473
rect 6626 5408 6632 5472
rect 6696 5408 6712 5472
rect 6776 5408 6792 5472
rect 6856 5408 6872 5472
rect 6936 5408 6942 5472
rect 6626 5407 6942 5408
rect 12307 5472 12623 5473
rect 12307 5408 12313 5472
rect 12377 5408 12393 5472
rect 12457 5408 12473 5472
rect 12537 5408 12553 5472
rect 12617 5408 12623 5472
rect 12307 5407 12623 5408
rect 17988 5472 18304 5473
rect 17988 5408 17994 5472
rect 18058 5408 18074 5472
rect 18138 5408 18154 5472
rect 18218 5408 18234 5472
rect 18298 5408 18304 5472
rect 17988 5407 18304 5408
rect 23669 5472 23985 5473
rect 23669 5408 23675 5472
rect 23739 5408 23755 5472
rect 23819 5408 23835 5472
rect 23899 5408 23915 5472
rect 23979 5408 23985 5472
rect 23669 5407 23985 5408
rect 3786 4928 4102 4929
rect 3786 4864 3792 4928
rect 3856 4864 3872 4928
rect 3936 4864 3952 4928
rect 4016 4864 4032 4928
rect 4096 4864 4102 4928
rect 3786 4863 4102 4864
rect 9467 4928 9783 4929
rect 9467 4864 9473 4928
rect 9537 4864 9553 4928
rect 9617 4864 9633 4928
rect 9697 4864 9713 4928
rect 9777 4864 9783 4928
rect 9467 4863 9783 4864
rect 15148 4928 15464 4929
rect 15148 4864 15154 4928
rect 15218 4864 15234 4928
rect 15298 4864 15314 4928
rect 15378 4864 15394 4928
rect 15458 4864 15464 4928
rect 15148 4863 15464 4864
rect 20829 4928 21145 4929
rect 20829 4864 20835 4928
rect 20899 4864 20915 4928
rect 20979 4864 20995 4928
rect 21059 4864 21075 4928
rect 21139 4864 21145 4928
rect 20829 4863 21145 4864
rect 4061 4722 4127 4725
rect 8334 4722 8340 4724
rect 4061 4720 8340 4722
rect 4061 4664 4066 4720
rect 4122 4664 8340 4720
rect 4061 4662 8340 4664
rect 4061 4659 4127 4662
rect 8334 4660 8340 4662
rect 8404 4660 8410 4724
rect 11881 4586 11947 4589
rect 12709 4586 12775 4589
rect 14917 4586 14983 4589
rect 11881 4584 14983 4586
rect 11881 4528 11886 4584
rect 11942 4528 12714 4584
rect 12770 4528 14922 4584
rect 14978 4528 14983 4584
rect 11881 4526 14983 4528
rect 11881 4523 11947 4526
rect 12709 4523 12775 4526
rect 14917 4523 14983 4526
rect 6626 4384 6942 4385
rect 6626 4320 6632 4384
rect 6696 4320 6712 4384
rect 6776 4320 6792 4384
rect 6856 4320 6872 4384
rect 6936 4320 6942 4384
rect 6626 4319 6942 4320
rect 12307 4384 12623 4385
rect 12307 4320 12313 4384
rect 12377 4320 12393 4384
rect 12457 4320 12473 4384
rect 12537 4320 12553 4384
rect 12617 4320 12623 4384
rect 12307 4319 12623 4320
rect 17988 4384 18304 4385
rect 17988 4320 17994 4384
rect 18058 4320 18074 4384
rect 18138 4320 18154 4384
rect 18218 4320 18234 4384
rect 18298 4320 18304 4384
rect 17988 4319 18304 4320
rect 23669 4384 23985 4385
rect 23669 4320 23675 4384
rect 23739 4320 23755 4384
rect 23819 4320 23835 4384
rect 23899 4320 23915 4384
rect 23979 4320 23985 4384
rect 23669 4319 23985 4320
rect 2865 4178 2931 4181
rect 5901 4178 5967 4181
rect 2865 4176 5967 4178
rect 2865 4120 2870 4176
rect 2926 4120 5906 4176
rect 5962 4120 5967 4176
rect 2865 4118 5967 4120
rect 2865 4115 2931 4118
rect 5901 4115 5967 4118
rect 2497 4042 2563 4045
rect 3550 4042 3556 4044
rect 2497 4040 3556 4042
rect 2497 3984 2502 4040
rect 2558 3984 3556 4040
rect 2497 3982 3556 3984
rect 2497 3979 2563 3982
rect 3550 3980 3556 3982
rect 3620 3980 3626 4044
rect 8518 3980 8524 4044
rect 8588 4042 8594 4044
rect 17401 4042 17467 4045
rect 8588 4040 17467 4042
rect 8588 3984 17406 4040
rect 17462 3984 17467 4040
rect 8588 3982 17467 3984
rect 8588 3980 8594 3982
rect 17401 3979 17467 3982
rect 3786 3840 4102 3841
rect 3786 3776 3792 3840
rect 3856 3776 3872 3840
rect 3936 3776 3952 3840
rect 4016 3776 4032 3840
rect 4096 3776 4102 3840
rect 3786 3775 4102 3776
rect 9467 3840 9783 3841
rect 9467 3776 9473 3840
rect 9537 3776 9553 3840
rect 9617 3776 9633 3840
rect 9697 3776 9713 3840
rect 9777 3776 9783 3840
rect 9467 3775 9783 3776
rect 15148 3840 15464 3841
rect 15148 3776 15154 3840
rect 15218 3776 15234 3840
rect 15298 3776 15314 3840
rect 15378 3776 15394 3840
rect 15458 3776 15464 3840
rect 15148 3775 15464 3776
rect 20829 3840 21145 3841
rect 20829 3776 20835 3840
rect 20899 3776 20915 3840
rect 20979 3776 20995 3840
rect 21059 3776 21075 3840
rect 21139 3776 21145 3840
rect 20829 3775 21145 3776
rect 4889 3770 4955 3773
rect 7281 3770 7347 3773
rect 4889 3768 7347 3770
rect 4889 3712 4894 3768
rect 4950 3712 7286 3768
rect 7342 3712 7347 3768
rect 4889 3710 7347 3712
rect 4889 3707 4955 3710
rect 7281 3707 7347 3710
rect 3417 3498 3483 3501
rect 4286 3498 4292 3500
rect 3417 3496 4292 3498
rect 3417 3440 3422 3496
rect 3478 3440 4292 3496
rect 3417 3438 4292 3440
rect 3417 3435 3483 3438
rect 4286 3436 4292 3438
rect 4356 3498 4362 3500
rect 5809 3498 5875 3501
rect 4356 3496 5875 3498
rect 4356 3440 5814 3496
rect 5870 3440 5875 3496
rect 4356 3438 5875 3440
rect 4356 3436 4362 3438
rect 5809 3435 5875 3438
rect 7966 3436 7972 3500
rect 8036 3498 8042 3500
rect 17953 3498 18019 3501
rect 8036 3496 18019 3498
rect 8036 3440 17958 3496
rect 18014 3440 18019 3496
rect 8036 3438 18019 3440
rect 8036 3436 8042 3438
rect 17953 3435 18019 3438
rect 6626 3296 6942 3297
rect 6626 3232 6632 3296
rect 6696 3232 6712 3296
rect 6776 3232 6792 3296
rect 6856 3232 6872 3296
rect 6936 3232 6942 3296
rect 6626 3231 6942 3232
rect 12307 3296 12623 3297
rect 12307 3232 12313 3296
rect 12377 3232 12393 3296
rect 12457 3232 12473 3296
rect 12537 3232 12553 3296
rect 12617 3232 12623 3296
rect 12307 3231 12623 3232
rect 17988 3296 18304 3297
rect 17988 3232 17994 3296
rect 18058 3232 18074 3296
rect 18138 3232 18154 3296
rect 18218 3232 18234 3296
rect 18298 3232 18304 3296
rect 17988 3231 18304 3232
rect 23669 3296 23985 3297
rect 23669 3232 23675 3296
rect 23739 3232 23755 3296
rect 23819 3232 23835 3296
rect 23899 3232 23915 3296
rect 23979 3232 23985 3296
rect 23669 3231 23985 3232
rect 2681 2954 2747 2957
rect 7649 2954 7715 2957
rect 8293 2954 8359 2957
rect 2681 2952 8359 2954
rect 2681 2896 2686 2952
rect 2742 2896 7654 2952
rect 7710 2896 8298 2952
rect 8354 2896 8359 2952
rect 2681 2894 8359 2896
rect 2681 2891 2747 2894
rect 7649 2891 7715 2894
rect 8293 2891 8359 2894
rect 3786 2752 4102 2753
rect 3786 2688 3792 2752
rect 3856 2688 3872 2752
rect 3936 2688 3952 2752
rect 4016 2688 4032 2752
rect 4096 2688 4102 2752
rect 3786 2687 4102 2688
rect 9467 2752 9783 2753
rect 9467 2688 9473 2752
rect 9537 2688 9553 2752
rect 9617 2688 9633 2752
rect 9697 2688 9713 2752
rect 9777 2688 9783 2752
rect 9467 2687 9783 2688
rect 15148 2752 15464 2753
rect 15148 2688 15154 2752
rect 15218 2688 15234 2752
rect 15298 2688 15314 2752
rect 15378 2688 15394 2752
rect 15458 2688 15464 2752
rect 15148 2687 15464 2688
rect 20829 2752 21145 2753
rect 20829 2688 20835 2752
rect 20899 2688 20915 2752
rect 20979 2688 20995 2752
rect 21059 2688 21075 2752
rect 21139 2688 21145 2752
rect 20829 2687 21145 2688
rect 5073 2684 5139 2685
rect 7833 2684 7899 2685
rect 5022 2682 5028 2684
rect 4982 2622 5028 2682
rect 5092 2680 5139 2684
rect 5134 2624 5139 2680
rect 5022 2620 5028 2622
rect 5092 2620 5139 2624
rect 7782 2620 7788 2684
rect 7852 2682 7899 2684
rect 7852 2680 7944 2682
rect 7894 2624 7944 2680
rect 7852 2622 7944 2624
rect 7852 2620 7899 2622
rect 5073 2619 5139 2620
rect 7833 2619 7899 2620
rect 4245 2546 4311 2549
rect 8518 2546 8524 2548
rect 4245 2544 8524 2546
rect 4245 2488 4250 2544
rect 4306 2488 8524 2544
rect 4245 2486 8524 2488
rect 4245 2483 4311 2486
rect 8518 2484 8524 2486
rect 8588 2484 8594 2548
rect 3417 2410 3483 2413
rect 8201 2412 8267 2413
rect 8150 2410 8156 2412
rect 3417 2408 8156 2410
rect 8220 2410 8267 2412
rect 8220 2408 8348 2410
rect 3417 2352 3422 2408
rect 3478 2352 8156 2408
rect 8262 2352 8348 2408
rect 3417 2350 8156 2352
rect 3417 2347 3483 2350
rect 8150 2348 8156 2350
rect 8220 2350 8348 2352
rect 8220 2348 8267 2350
rect 8201 2347 8267 2348
rect 6626 2208 6942 2209
rect 6626 2144 6632 2208
rect 6696 2144 6712 2208
rect 6776 2144 6792 2208
rect 6856 2144 6872 2208
rect 6936 2144 6942 2208
rect 6626 2143 6942 2144
rect 12307 2208 12623 2209
rect 12307 2144 12313 2208
rect 12377 2144 12393 2208
rect 12457 2144 12473 2208
rect 12537 2144 12553 2208
rect 12617 2144 12623 2208
rect 12307 2143 12623 2144
rect 17988 2208 18304 2209
rect 17988 2144 17994 2208
rect 18058 2144 18074 2208
rect 18138 2144 18154 2208
rect 18218 2144 18234 2208
rect 18298 2144 18304 2208
rect 17988 2143 18304 2144
rect 23669 2208 23985 2209
rect 23669 2144 23675 2208
rect 23739 2144 23755 2208
rect 23819 2144 23835 2208
rect 23899 2144 23915 2208
rect 23979 2144 23985 2208
rect 23669 2143 23985 2144
rect 1853 2002 1919 2005
rect 7966 2002 7972 2004
rect 1853 2000 7972 2002
rect 1853 1944 1858 2000
rect 1914 1944 7972 2000
rect 1853 1942 7972 1944
rect 1853 1939 1919 1942
rect 7966 1940 7972 1942
rect 8036 1940 8042 2004
<< via3 >>
rect 3792 22332 3856 22336
rect 3792 22276 3796 22332
rect 3796 22276 3852 22332
rect 3852 22276 3856 22332
rect 3792 22272 3856 22276
rect 3872 22332 3936 22336
rect 3872 22276 3876 22332
rect 3876 22276 3932 22332
rect 3932 22276 3936 22332
rect 3872 22272 3936 22276
rect 3952 22332 4016 22336
rect 3952 22276 3956 22332
rect 3956 22276 4012 22332
rect 4012 22276 4016 22332
rect 3952 22272 4016 22276
rect 4032 22332 4096 22336
rect 4032 22276 4036 22332
rect 4036 22276 4092 22332
rect 4092 22276 4096 22332
rect 4032 22272 4096 22276
rect 9473 22332 9537 22336
rect 9473 22276 9477 22332
rect 9477 22276 9533 22332
rect 9533 22276 9537 22332
rect 9473 22272 9537 22276
rect 9553 22332 9617 22336
rect 9553 22276 9557 22332
rect 9557 22276 9613 22332
rect 9613 22276 9617 22332
rect 9553 22272 9617 22276
rect 9633 22332 9697 22336
rect 9633 22276 9637 22332
rect 9637 22276 9693 22332
rect 9693 22276 9697 22332
rect 9633 22272 9697 22276
rect 9713 22332 9777 22336
rect 9713 22276 9717 22332
rect 9717 22276 9773 22332
rect 9773 22276 9777 22332
rect 9713 22272 9777 22276
rect 15154 22332 15218 22336
rect 15154 22276 15158 22332
rect 15158 22276 15214 22332
rect 15214 22276 15218 22332
rect 15154 22272 15218 22276
rect 15234 22332 15298 22336
rect 15234 22276 15238 22332
rect 15238 22276 15294 22332
rect 15294 22276 15298 22332
rect 15234 22272 15298 22276
rect 15314 22332 15378 22336
rect 15314 22276 15318 22332
rect 15318 22276 15374 22332
rect 15374 22276 15378 22332
rect 15314 22272 15378 22276
rect 15394 22332 15458 22336
rect 15394 22276 15398 22332
rect 15398 22276 15454 22332
rect 15454 22276 15458 22332
rect 15394 22272 15458 22276
rect 20835 22332 20899 22336
rect 20835 22276 20839 22332
rect 20839 22276 20895 22332
rect 20895 22276 20899 22332
rect 20835 22272 20899 22276
rect 20915 22332 20979 22336
rect 20915 22276 20919 22332
rect 20919 22276 20975 22332
rect 20975 22276 20979 22332
rect 20915 22272 20979 22276
rect 20995 22332 21059 22336
rect 20995 22276 20999 22332
rect 20999 22276 21055 22332
rect 21055 22276 21059 22332
rect 20995 22272 21059 22276
rect 21075 22332 21139 22336
rect 21075 22276 21079 22332
rect 21079 22276 21135 22332
rect 21135 22276 21139 22332
rect 21075 22272 21139 22276
rect 6632 21788 6696 21792
rect 6632 21732 6636 21788
rect 6636 21732 6692 21788
rect 6692 21732 6696 21788
rect 6632 21728 6696 21732
rect 6712 21788 6776 21792
rect 6712 21732 6716 21788
rect 6716 21732 6772 21788
rect 6772 21732 6776 21788
rect 6712 21728 6776 21732
rect 6792 21788 6856 21792
rect 6792 21732 6796 21788
rect 6796 21732 6852 21788
rect 6852 21732 6856 21788
rect 6792 21728 6856 21732
rect 6872 21788 6936 21792
rect 6872 21732 6876 21788
rect 6876 21732 6932 21788
rect 6932 21732 6936 21788
rect 6872 21728 6936 21732
rect 12313 21788 12377 21792
rect 12313 21732 12317 21788
rect 12317 21732 12373 21788
rect 12373 21732 12377 21788
rect 12313 21728 12377 21732
rect 12393 21788 12457 21792
rect 12393 21732 12397 21788
rect 12397 21732 12453 21788
rect 12453 21732 12457 21788
rect 12393 21728 12457 21732
rect 12473 21788 12537 21792
rect 12473 21732 12477 21788
rect 12477 21732 12533 21788
rect 12533 21732 12537 21788
rect 12473 21728 12537 21732
rect 12553 21788 12617 21792
rect 12553 21732 12557 21788
rect 12557 21732 12613 21788
rect 12613 21732 12617 21788
rect 12553 21728 12617 21732
rect 17994 21788 18058 21792
rect 17994 21732 17998 21788
rect 17998 21732 18054 21788
rect 18054 21732 18058 21788
rect 17994 21728 18058 21732
rect 18074 21788 18138 21792
rect 18074 21732 18078 21788
rect 18078 21732 18134 21788
rect 18134 21732 18138 21788
rect 18074 21728 18138 21732
rect 18154 21788 18218 21792
rect 18154 21732 18158 21788
rect 18158 21732 18214 21788
rect 18214 21732 18218 21788
rect 18154 21728 18218 21732
rect 18234 21788 18298 21792
rect 18234 21732 18238 21788
rect 18238 21732 18294 21788
rect 18294 21732 18298 21788
rect 18234 21728 18298 21732
rect 23675 21788 23739 21792
rect 23675 21732 23679 21788
rect 23679 21732 23735 21788
rect 23735 21732 23739 21788
rect 23675 21728 23739 21732
rect 23755 21788 23819 21792
rect 23755 21732 23759 21788
rect 23759 21732 23815 21788
rect 23815 21732 23819 21788
rect 23755 21728 23819 21732
rect 23835 21788 23899 21792
rect 23835 21732 23839 21788
rect 23839 21732 23895 21788
rect 23895 21732 23899 21788
rect 23835 21728 23899 21732
rect 23915 21788 23979 21792
rect 23915 21732 23919 21788
rect 23919 21732 23975 21788
rect 23975 21732 23979 21788
rect 23915 21728 23979 21732
rect 3792 21244 3856 21248
rect 3792 21188 3796 21244
rect 3796 21188 3852 21244
rect 3852 21188 3856 21244
rect 3792 21184 3856 21188
rect 3872 21244 3936 21248
rect 3872 21188 3876 21244
rect 3876 21188 3932 21244
rect 3932 21188 3936 21244
rect 3872 21184 3936 21188
rect 3952 21244 4016 21248
rect 3952 21188 3956 21244
rect 3956 21188 4012 21244
rect 4012 21188 4016 21244
rect 3952 21184 4016 21188
rect 4032 21244 4096 21248
rect 4032 21188 4036 21244
rect 4036 21188 4092 21244
rect 4092 21188 4096 21244
rect 4032 21184 4096 21188
rect 9473 21244 9537 21248
rect 9473 21188 9477 21244
rect 9477 21188 9533 21244
rect 9533 21188 9537 21244
rect 9473 21184 9537 21188
rect 9553 21244 9617 21248
rect 9553 21188 9557 21244
rect 9557 21188 9613 21244
rect 9613 21188 9617 21244
rect 9553 21184 9617 21188
rect 9633 21244 9697 21248
rect 9633 21188 9637 21244
rect 9637 21188 9693 21244
rect 9693 21188 9697 21244
rect 9633 21184 9697 21188
rect 9713 21244 9777 21248
rect 9713 21188 9717 21244
rect 9717 21188 9773 21244
rect 9773 21188 9777 21244
rect 9713 21184 9777 21188
rect 15154 21244 15218 21248
rect 15154 21188 15158 21244
rect 15158 21188 15214 21244
rect 15214 21188 15218 21244
rect 15154 21184 15218 21188
rect 15234 21244 15298 21248
rect 15234 21188 15238 21244
rect 15238 21188 15294 21244
rect 15294 21188 15298 21244
rect 15234 21184 15298 21188
rect 15314 21244 15378 21248
rect 15314 21188 15318 21244
rect 15318 21188 15374 21244
rect 15374 21188 15378 21244
rect 15314 21184 15378 21188
rect 15394 21244 15458 21248
rect 15394 21188 15398 21244
rect 15398 21188 15454 21244
rect 15454 21188 15458 21244
rect 15394 21184 15458 21188
rect 20835 21244 20899 21248
rect 20835 21188 20839 21244
rect 20839 21188 20895 21244
rect 20895 21188 20899 21244
rect 20835 21184 20899 21188
rect 20915 21244 20979 21248
rect 20915 21188 20919 21244
rect 20919 21188 20975 21244
rect 20975 21188 20979 21244
rect 20915 21184 20979 21188
rect 20995 21244 21059 21248
rect 20995 21188 20999 21244
rect 20999 21188 21055 21244
rect 21055 21188 21059 21244
rect 20995 21184 21059 21188
rect 21075 21244 21139 21248
rect 21075 21188 21079 21244
rect 21079 21188 21135 21244
rect 21135 21188 21139 21244
rect 21075 21184 21139 21188
rect 4292 20708 4356 20772
rect 7604 20708 7668 20772
rect 6632 20700 6696 20704
rect 6632 20644 6636 20700
rect 6636 20644 6692 20700
rect 6692 20644 6696 20700
rect 6632 20640 6696 20644
rect 6712 20700 6776 20704
rect 6712 20644 6716 20700
rect 6716 20644 6772 20700
rect 6772 20644 6776 20700
rect 6712 20640 6776 20644
rect 6792 20700 6856 20704
rect 6792 20644 6796 20700
rect 6796 20644 6852 20700
rect 6852 20644 6856 20700
rect 6792 20640 6856 20644
rect 6872 20700 6936 20704
rect 6872 20644 6876 20700
rect 6876 20644 6932 20700
rect 6932 20644 6936 20700
rect 6872 20640 6936 20644
rect 12313 20700 12377 20704
rect 12313 20644 12317 20700
rect 12317 20644 12373 20700
rect 12373 20644 12377 20700
rect 12313 20640 12377 20644
rect 12393 20700 12457 20704
rect 12393 20644 12397 20700
rect 12397 20644 12453 20700
rect 12453 20644 12457 20700
rect 12393 20640 12457 20644
rect 12473 20700 12537 20704
rect 12473 20644 12477 20700
rect 12477 20644 12533 20700
rect 12533 20644 12537 20700
rect 12473 20640 12537 20644
rect 12553 20700 12617 20704
rect 12553 20644 12557 20700
rect 12557 20644 12613 20700
rect 12613 20644 12617 20700
rect 12553 20640 12617 20644
rect 17994 20700 18058 20704
rect 17994 20644 17998 20700
rect 17998 20644 18054 20700
rect 18054 20644 18058 20700
rect 17994 20640 18058 20644
rect 18074 20700 18138 20704
rect 18074 20644 18078 20700
rect 18078 20644 18134 20700
rect 18134 20644 18138 20700
rect 18074 20640 18138 20644
rect 18154 20700 18218 20704
rect 18154 20644 18158 20700
rect 18158 20644 18214 20700
rect 18214 20644 18218 20700
rect 18154 20640 18218 20644
rect 18234 20700 18298 20704
rect 18234 20644 18238 20700
rect 18238 20644 18294 20700
rect 18294 20644 18298 20700
rect 18234 20640 18298 20644
rect 23675 20700 23739 20704
rect 23675 20644 23679 20700
rect 23679 20644 23735 20700
rect 23735 20644 23739 20700
rect 23675 20640 23739 20644
rect 23755 20700 23819 20704
rect 23755 20644 23759 20700
rect 23759 20644 23815 20700
rect 23815 20644 23819 20700
rect 23755 20640 23819 20644
rect 23835 20700 23899 20704
rect 23835 20644 23839 20700
rect 23839 20644 23895 20700
rect 23895 20644 23899 20700
rect 23835 20640 23899 20644
rect 23915 20700 23979 20704
rect 23915 20644 23919 20700
rect 23919 20644 23975 20700
rect 23975 20644 23979 20700
rect 23915 20640 23979 20644
rect 3792 20156 3856 20160
rect 3792 20100 3796 20156
rect 3796 20100 3852 20156
rect 3852 20100 3856 20156
rect 3792 20096 3856 20100
rect 3872 20156 3936 20160
rect 3872 20100 3876 20156
rect 3876 20100 3932 20156
rect 3932 20100 3936 20156
rect 3872 20096 3936 20100
rect 3952 20156 4016 20160
rect 3952 20100 3956 20156
rect 3956 20100 4012 20156
rect 4012 20100 4016 20156
rect 3952 20096 4016 20100
rect 4032 20156 4096 20160
rect 4032 20100 4036 20156
rect 4036 20100 4092 20156
rect 4092 20100 4096 20156
rect 4032 20096 4096 20100
rect 9473 20156 9537 20160
rect 9473 20100 9477 20156
rect 9477 20100 9533 20156
rect 9533 20100 9537 20156
rect 9473 20096 9537 20100
rect 9553 20156 9617 20160
rect 9553 20100 9557 20156
rect 9557 20100 9613 20156
rect 9613 20100 9617 20156
rect 9553 20096 9617 20100
rect 9633 20156 9697 20160
rect 9633 20100 9637 20156
rect 9637 20100 9693 20156
rect 9693 20100 9697 20156
rect 9633 20096 9697 20100
rect 9713 20156 9777 20160
rect 9713 20100 9717 20156
rect 9717 20100 9773 20156
rect 9773 20100 9777 20156
rect 9713 20096 9777 20100
rect 15154 20156 15218 20160
rect 15154 20100 15158 20156
rect 15158 20100 15214 20156
rect 15214 20100 15218 20156
rect 15154 20096 15218 20100
rect 15234 20156 15298 20160
rect 15234 20100 15238 20156
rect 15238 20100 15294 20156
rect 15294 20100 15298 20156
rect 15234 20096 15298 20100
rect 15314 20156 15378 20160
rect 15314 20100 15318 20156
rect 15318 20100 15374 20156
rect 15374 20100 15378 20156
rect 15314 20096 15378 20100
rect 15394 20156 15458 20160
rect 15394 20100 15398 20156
rect 15398 20100 15454 20156
rect 15454 20100 15458 20156
rect 15394 20096 15458 20100
rect 20835 20156 20899 20160
rect 20835 20100 20839 20156
rect 20839 20100 20895 20156
rect 20895 20100 20899 20156
rect 20835 20096 20899 20100
rect 20915 20156 20979 20160
rect 20915 20100 20919 20156
rect 20919 20100 20975 20156
rect 20975 20100 20979 20156
rect 20915 20096 20979 20100
rect 20995 20156 21059 20160
rect 20995 20100 20999 20156
rect 20999 20100 21055 20156
rect 21055 20100 21059 20156
rect 20995 20096 21059 20100
rect 21075 20156 21139 20160
rect 21075 20100 21079 20156
rect 21079 20100 21135 20156
rect 21135 20100 21139 20156
rect 21075 20096 21139 20100
rect 6632 19612 6696 19616
rect 6632 19556 6636 19612
rect 6636 19556 6692 19612
rect 6692 19556 6696 19612
rect 6632 19552 6696 19556
rect 6712 19612 6776 19616
rect 6712 19556 6716 19612
rect 6716 19556 6772 19612
rect 6772 19556 6776 19612
rect 6712 19552 6776 19556
rect 6792 19612 6856 19616
rect 6792 19556 6796 19612
rect 6796 19556 6852 19612
rect 6852 19556 6856 19612
rect 6792 19552 6856 19556
rect 6872 19612 6936 19616
rect 6872 19556 6876 19612
rect 6876 19556 6932 19612
rect 6932 19556 6936 19612
rect 6872 19552 6936 19556
rect 12313 19612 12377 19616
rect 12313 19556 12317 19612
rect 12317 19556 12373 19612
rect 12373 19556 12377 19612
rect 12313 19552 12377 19556
rect 12393 19612 12457 19616
rect 12393 19556 12397 19612
rect 12397 19556 12453 19612
rect 12453 19556 12457 19612
rect 12393 19552 12457 19556
rect 12473 19612 12537 19616
rect 12473 19556 12477 19612
rect 12477 19556 12533 19612
rect 12533 19556 12537 19612
rect 12473 19552 12537 19556
rect 12553 19612 12617 19616
rect 12553 19556 12557 19612
rect 12557 19556 12613 19612
rect 12613 19556 12617 19612
rect 12553 19552 12617 19556
rect 17994 19612 18058 19616
rect 17994 19556 17998 19612
rect 17998 19556 18054 19612
rect 18054 19556 18058 19612
rect 17994 19552 18058 19556
rect 18074 19612 18138 19616
rect 18074 19556 18078 19612
rect 18078 19556 18134 19612
rect 18134 19556 18138 19612
rect 18074 19552 18138 19556
rect 18154 19612 18218 19616
rect 18154 19556 18158 19612
rect 18158 19556 18214 19612
rect 18214 19556 18218 19612
rect 18154 19552 18218 19556
rect 18234 19612 18298 19616
rect 18234 19556 18238 19612
rect 18238 19556 18294 19612
rect 18294 19556 18298 19612
rect 18234 19552 18298 19556
rect 23675 19612 23739 19616
rect 23675 19556 23679 19612
rect 23679 19556 23735 19612
rect 23735 19556 23739 19612
rect 23675 19552 23739 19556
rect 23755 19612 23819 19616
rect 23755 19556 23759 19612
rect 23759 19556 23815 19612
rect 23815 19556 23819 19612
rect 23755 19552 23819 19556
rect 23835 19612 23899 19616
rect 23835 19556 23839 19612
rect 23839 19556 23895 19612
rect 23895 19556 23899 19612
rect 23835 19552 23899 19556
rect 23915 19612 23979 19616
rect 23915 19556 23919 19612
rect 23919 19556 23975 19612
rect 23975 19556 23979 19612
rect 23915 19552 23979 19556
rect 3556 19348 3620 19412
rect 6316 19408 6380 19412
rect 6316 19352 6366 19408
rect 6366 19352 6380 19408
rect 6316 19348 6380 19352
rect 3792 19068 3856 19072
rect 3792 19012 3796 19068
rect 3796 19012 3852 19068
rect 3852 19012 3856 19068
rect 3792 19008 3856 19012
rect 3872 19068 3936 19072
rect 3872 19012 3876 19068
rect 3876 19012 3932 19068
rect 3932 19012 3936 19068
rect 3872 19008 3936 19012
rect 3952 19068 4016 19072
rect 3952 19012 3956 19068
rect 3956 19012 4012 19068
rect 4012 19012 4016 19068
rect 3952 19008 4016 19012
rect 4032 19068 4096 19072
rect 4032 19012 4036 19068
rect 4036 19012 4092 19068
rect 4092 19012 4096 19068
rect 4032 19008 4096 19012
rect 9473 19068 9537 19072
rect 9473 19012 9477 19068
rect 9477 19012 9533 19068
rect 9533 19012 9537 19068
rect 9473 19008 9537 19012
rect 9553 19068 9617 19072
rect 9553 19012 9557 19068
rect 9557 19012 9613 19068
rect 9613 19012 9617 19068
rect 9553 19008 9617 19012
rect 9633 19068 9697 19072
rect 9633 19012 9637 19068
rect 9637 19012 9693 19068
rect 9693 19012 9697 19068
rect 9633 19008 9697 19012
rect 9713 19068 9777 19072
rect 9713 19012 9717 19068
rect 9717 19012 9773 19068
rect 9773 19012 9777 19068
rect 9713 19008 9777 19012
rect 15154 19068 15218 19072
rect 15154 19012 15158 19068
rect 15158 19012 15214 19068
rect 15214 19012 15218 19068
rect 15154 19008 15218 19012
rect 15234 19068 15298 19072
rect 15234 19012 15238 19068
rect 15238 19012 15294 19068
rect 15294 19012 15298 19068
rect 15234 19008 15298 19012
rect 15314 19068 15378 19072
rect 15314 19012 15318 19068
rect 15318 19012 15374 19068
rect 15374 19012 15378 19068
rect 15314 19008 15378 19012
rect 15394 19068 15458 19072
rect 15394 19012 15398 19068
rect 15398 19012 15454 19068
rect 15454 19012 15458 19068
rect 15394 19008 15458 19012
rect 20835 19068 20899 19072
rect 20835 19012 20839 19068
rect 20839 19012 20895 19068
rect 20895 19012 20899 19068
rect 20835 19008 20899 19012
rect 20915 19068 20979 19072
rect 20915 19012 20919 19068
rect 20919 19012 20975 19068
rect 20975 19012 20979 19068
rect 20915 19008 20979 19012
rect 20995 19068 21059 19072
rect 20995 19012 20999 19068
rect 20999 19012 21055 19068
rect 21055 19012 21059 19068
rect 20995 19008 21059 19012
rect 21075 19068 21139 19072
rect 21075 19012 21079 19068
rect 21079 19012 21135 19068
rect 21135 19012 21139 19068
rect 21075 19008 21139 19012
rect 6632 18524 6696 18528
rect 6632 18468 6636 18524
rect 6636 18468 6692 18524
rect 6692 18468 6696 18524
rect 6632 18464 6696 18468
rect 6712 18524 6776 18528
rect 6712 18468 6716 18524
rect 6716 18468 6772 18524
rect 6772 18468 6776 18524
rect 6712 18464 6776 18468
rect 6792 18524 6856 18528
rect 6792 18468 6796 18524
rect 6796 18468 6852 18524
rect 6852 18468 6856 18524
rect 6792 18464 6856 18468
rect 6872 18524 6936 18528
rect 6872 18468 6876 18524
rect 6876 18468 6932 18524
rect 6932 18468 6936 18524
rect 6872 18464 6936 18468
rect 12313 18524 12377 18528
rect 12313 18468 12317 18524
rect 12317 18468 12373 18524
rect 12373 18468 12377 18524
rect 12313 18464 12377 18468
rect 12393 18524 12457 18528
rect 12393 18468 12397 18524
rect 12397 18468 12453 18524
rect 12453 18468 12457 18524
rect 12393 18464 12457 18468
rect 12473 18524 12537 18528
rect 12473 18468 12477 18524
rect 12477 18468 12533 18524
rect 12533 18468 12537 18524
rect 12473 18464 12537 18468
rect 12553 18524 12617 18528
rect 12553 18468 12557 18524
rect 12557 18468 12613 18524
rect 12613 18468 12617 18524
rect 12553 18464 12617 18468
rect 17994 18524 18058 18528
rect 17994 18468 17998 18524
rect 17998 18468 18054 18524
rect 18054 18468 18058 18524
rect 17994 18464 18058 18468
rect 18074 18524 18138 18528
rect 18074 18468 18078 18524
rect 18078 18468 18134 18524
rect 18134 18468 18138 18524
rect 18074 18464 18138 18468
rect 18154 18524 18218 18528
rect 18154 18468 18158 18524
rect 18158 18468 18214 18524
rect 18214 18468 18218 18524
rect 18154 18464 18218 18468
rect 18234 18524 18298 18528
rect 18234 18468 18238 18524
rect 18238 18468 18294 18524
rect 18294 18468 18298 18524
rect 18234 18464 18298 18468
rect 23675 18524 23739 18528
rect 23675 18468 23679 18524
rect 23679 18468 23735 18524
rect 23735 18468 23739 18524
rect 23675 18464 23739 18468
rect 23755 18524 23819 18528
rect 23755 18468 23759 18524
rect 23759 18468 23815 18524
rect 23815 18468 23819 18524
rect 23755 18464 23819 18468
rect 23835 18524 23899 18528
rect 23835 18468 23839 18524
rect 23839 18468 23895 18524
rect 23895 18468 23899 18524
rect 23835 18464 23899 18468
rect 23915 18524 23979 18528
rect 23915 18468 23919 18524
rect 23919 18468 23975 18524
rect 23975 18468 23979 18524
rect 23915 18464 23979 18468
rect 7420 18048 7484 18052
rect 7420 17992 7434 18048
rect 7434 17992 7484 18048
rect 7420 17988 7484 17992
rect 3792 17980 3856 17984
rect 3792 17924 3796 17980
rect 3796 17924 3852 17980
rect 3852 17924 3856 17980
rect 3792 17920 3856 17924
rect 3872 17980 3936 17984
rect 3872 17924 3876 17980
rect 3876 17924 3932 17980
rect 3932 17924 3936 17980
rect 3872 17920 3936 17924
rect 3952 17980 4016 17984
rect 3952 17924 3956 17980
rect 3956 17924 4012 17980
rect 4012 17924 4016 17980
rect 3952 17920 4016 17924
rect 4032 17980 4096 17984
rect 4032 17924 4036 17980
rect 4036 17924 4092 17980
rect 4092 17924 4096 17980
rect 4032 17920 4096 17924
rect 9473 17980 9537 17984
rect 9473 17924 9477 17980
rect 9477 17924 9533 17980
rect 9533 17924 9537 17980
rect 9473 17920 9537 17924
rect 9553 17980 9617 17984
rect 9553 17924 9557 17980
rect 9557 17924 9613 17980
rect 9613 17924 9617 17980
rect 9553 17920 9617 17924
rect 9633 17980 9697 17984
rect 9633 17924 9637 17980
rect 9637 17924 9693 17980
rect 9693 17924 9697 17980
rect 9633 17920 9697 17924
rect 9713 17980 9777 17984
rect 9713 17924 9717 17980
rect 9717 17924 9773 17980
rect 9773 17924 9777 17980
rect 9713 17920 9777 17924
rect 15154 17980 15218 17984
rect 15154 17924 15158 17980
rect 15158 17924 15214 17980
rect 15214 17924 15218 17980
rect 15154 17920 15218 17924
rect 15234 17980 15298 17984
rect 15234 17924 15238 17980
rect 15238 17924 15294 17980
rect 15294 17924 15298 17980
rect 15234 17920 15298 17924
rect 15314 17980 15378 17984
rect 15314 17924 15318 17980
rect 15318 17924 15374 17980
rect 15374 17924 15378 17980
rect 15314 17920 15378 17924
rect 15394 17980 15458 17984
rect 15394 17924 15398 17980
rect 15398 17924 15454 17980
rect 15454 17924 15458 17980
rect 15394 17920 15458 17924
rect 20835 17980 20899 17984
rect 20835 17924 20839 17980
rect 20839 17924 20895 17980
rect 20895 17924 20899 17980
rect 20835 17920 20899 17924
rect 20915 17980 20979 17984
rect 20915 17924 20919 17980
rect 20919 17924 20975 17980
rect 20975 17924 20979 17980
rect 20915 17920 20979 17924
rect 20995 17980 21059 17984
rect 20995 17924 20999 17980
rect 20999 17924 21055 17980
rect 21055 17924 21059 17980
rect 20995 17920 21059 17924
rect 21075 17980 21139 17984
rect 21075 17924 21079 17980
rect 21079 17924 21135 17980
rect 21135 17924 21139 17980
rect 21075 17920 21139 17924
rect 6632 17436 6696 17440
rect 6632 17380 6636 17436
rect 6636 17380 6692 17436
rect 6692 17380 6696 17436
rect 6632 17376 6696 17380
rect 6712 17436 6776 17440
rect 6712 17380 6716 17436
rect 6716 17380 6772 17436
rect 6772 17380 6776 17436
rect 6712 17376 6776 17380
rect 6792 17436 6856 17440
rect 6792 17380 6796 17436
rect 6796 17380 6852 17436
rect 6852 17380 6856 17436
rect 6792 17376 6856 17380
rect 6872 17436 6936 17440
rect 6872 17380 6876 17436
rect 6876 17380 6932 17436
rect 6932 17380 6936 17436
rect 6872 17376 6936 17380
rect 12313 17436 12377 17440
rect 12313 17380 12317 17436
rect 12317 17380 12373 17436
rect 12373 17380 12377 17436
rect 12313 17376 12377 17380
rect 12393 17436 12457 17440
rect 12393 17380 12397 17436
rect 12397 17380 12453 17436
rect 12453 17380 12457 17436
rect 12393 17376 12457 17380
rect 12473 17436 12537 17440
rect 12473 17380 12477 17436
rect 12477 17380 12533 17436
rect 12533 17380 12537 17436
rect 12473 17376 12537 17380
rect 12553 17436 12617 17440
rect 12553 17380 12557 17436
rect 12557 17380 12613 17436
rect 12613 17380 12617 17436
rect 12553 17376 12617 17380
rect 17994 17436 18058 17440
rect 17994 17380 17998 17436
rect 17998 17380 18054 17436
rect 18054 17380 18058 17436
rect 17994 17376 18058 17380
rect 18074 17436 18138 17440
rect 18074 17380 18078 17436
rect 18078 17380 18134 17436
rect 18134 17380 18138 17436
rect 18074 17376 18138 17380
rect 18154 17436 18218 17440
rect 18154 17380 18158 17436
rect 18158 17380 18214 17436
rect 18214 17380 18218 17436
rect 18154 17376 18218 17380
rect 18234 17436 18298 17440
rect 18234 17380 18238 17436
rect 18238 17380 18294 17436
rect 18294 17380 18298 17436
rect 18234 17376 18298 17380
rect 23675 17436 23739 17440
rect 23675 17380 23679 17436
rect 23679 17380 23735 17436
rect 23735 17380 23739 17436
rect 23675 17376 23739 17380
rect 23755 17436 23819 17440
rect 23755 17380 23759 17436
rect 23759 17380 23815 17436
rect 23815 17380 23819 17436
rect 23755 17376 23819 17380
rect 23835 17436 23899 17440
rect 23835 17380 23839 17436
rect 23839 17380 23895 17436
rect 23895 17380 23899 17436
rect 23835 17376 23899 17380
rect 23915 17436 23979 17440
rect 23915 17380 23919 17436
rect 23919 17380 23975 17436
rect 23975 17380 23979 17436
rect 23915 17376 23979 17380
rect 3792 16892 3856 16896
rect 3792 16836 3796 16892
rect 3796 16836 3852 16892
rect 3852 16836 3856 16892
rect 3792 16832 3856 16836
rect 3872 16892 3936 16896
rect 3872 16836 3876 16892
rect 3876 16836 3932 16892
rect 3932 16836 3936 16892
rect 3872 16832 3936 16836
rect 3952 16892 4016 16896
rect 3952 16836 3956 16892
rect 3956 16836 4012 16892
rect 4012 16836 4016 16892
rect 3952 16832 4016 16836
rect 4032 16892 4096 16896
rect 4032 16836 4036 16892
rect 4036 16836 4092 16892
rect 4092 16836 4096 16892
rect 4032 16832 4096 16836
rect 9473 16892 9537 16896
rect 9473 16836 9477 16892
rect 9477 16836 9533 16892
rect 9533 16836 9537 16892
rect 9473 16832 9537 16836
rect 9553 16892 9617 16896
rect 9553 16836 9557 16892
rect 9557 16836 9613 16892
rect 9613 16836 9617 16892
rect 9553 16832 9617 16836
rect 9633 16892 9697 16896
rect 9633 16836 9637 16892
rect 9637 16836 9693 16892
rect 9693 16836 9697 16892
rect 9633 16832 9697 16836
rect 9713 16892 9777 16896
rect 9713 16836 9717 16892
rect 9717 16836 9773 16892
rect 9773 16836 9777 16892
rect 9713 16832 9777 16836
rect 15154 16892 15218 16896
rect 15154 16836 15158 16892
rect 15158 16836 15214 16892
rect 15214 16836 15218 16892
rect 15154 16832 15218 16836
rect 15234 16892 15298 16896
rect 15234 16836 15238 16892
rect 15238 16836 15294 16892
rect 15294 16836 15298 16892
rect 15234 16832 15298 16836
rect 15314 16892 15378 16896
rect 15314 16836 15318 16892
rect 15318 16836 15374 16892
rect 15374 16836 15378 16892
rect 15314 16832 15378 16836
rect 15394 16892 15458 16896
rect 15394 16836 15398 16892
rect 15398 16836 15454 16892
rect 15454 16836 15458 16892
rect 15394 16832 15458 16836
rect 20835 16892 20899 16896
rect 20835 16836 20839 16892
rect 20839 16836 20895 16892
rect 20895 16836 20899 16892
rect 20835 16832 20899 16836
rect 20915 16892 20979 16896
rect 20915 16836 20919 16892
rect 20919 16836 20975 16892
rect 20975 16836 20979 16892
rect 20915 16832 20979 16836
rect 20995 16892 21059 16896
rect 20995 16836 20999 16892
rect 20999 16836 21055 16892
rect 21055 16836 21059 16892
rect 20995 16832 21059 16836
rect 21075 16892 21139 16896
rect 21075 16836 21079 16892
rect 21079 16836 21135 16892
rect 21135 16836 21139 16892
rect 21075 16832 21139 16836
rect 3372 16688 3436 16692
rect 3372 16632 3422 16688
rect 3422 16632 3436 16688
rect 3372 16628 3436 16632
rect 6632 16348 6696 16352
rect 6632 16292 6636 16348
rect 6636 16292 6692 16348
rect 6692 16292 6696 16348
rect 6632 16288 6696 16292
rect 6712 16348 6776 16352
rect 6712 16292 6716 16348
rect 6716 16292 6772 16348
rect 6772 16292 6776 16348
rect 6712 16288 6776 16292
rect 6792 16348 6856 16352
rect 6792 16292 6796 16348
rect 6796 16292 6852 16348
rect 6852 16292 6856 16348
rect 6792 16288 6856 16292
rect 6872 16348 6936 16352
rect 6872 16292 6876 16348
rect 6876 16292 6932 16348
rect 6932 16292 6936 16348
rect 6872 16288 6936 16292
rect 12313 16348 12377 16352
rect 12313 16292 12317 16348
rect 12317 16292 12373 16348
rect 12373 16292 12377 16348
rect 12313 16288 12377 16292
rect 12393 16348 12457 16352
rect 12393 16292 12397 16348
rect 12397 16292 12453 16348
rect 12453 16292 12457 16348
rect 12393 16288 12457 16292
rect 12473 16348 12537 16352
rect 12473 16292 12477 16348
rect 12477 16292 12533 16348
rect 12533 16292 12537 16348
rect 12473 16288 12537 16292
rect 12553 16348 12617 16352
rect 12553 16292 12557 16348
rect 12557 16292 12613 16348
rect 12613 16292 12617 16348
rect 12553 16288 12617 16292
rect 17994 16348 18058 16352
rect 17994 16292 17998 16348
rect 17998 16292 18054 16348
rect 18054 16292 18058 16348
rect 17994 16288 18058 16292
rect 18074 16348 18138 16352
rect 18074 16292 18078 16348
rect 18078 16292 18134 16348
rect 18134 16292 18138 16348
rect 18074 16288 18138 16292
rect 18154 16348 18218 16352
rect 18154 16292 18158 16348
rect 18158 16292 18214 16348
rect 18214 16292 18218 16348
rect 18154 16288 18218 16292
rect 18234 16348 18298 16352
rect 18234 16292 18238 16348
rect 18238 16292 18294 16348
rect 18294 16292 18298 16348
rect 18234 16288 18298 16292
rect 23675 16348 23739 16352
rect 23675 16292 23679 16348
rect 23679 16292 23735 16348
rect 23735 16292 23739 16348
rect 23675 16288 23739 16292
rect 23755 16348 23819 16352
rect 23755 16292 23759 16348
rect 23759 16292 23815 16348
rect 23815 16292 23819 16348
rect 23755 16288 23819 16292
rect 23835 16348 23899 16352
rect 23835 16292 23839 16348
rect 23839 16292 23895 16348
rect 23895 16292 23899 16348
rect 23835 16288 23899 16292
rect 23915 16348 23979 16352
rect 23915 16292 23919 16348
rect 23919 16292 23975 16348
rect 23975 16292 23979 16348
rect 23915 16288 23979 16292
rect 3792 15804 3856 15808
rect 3792 15748 3796 15804
rect 3796 15748 3852 15804
rect 3852 15748 3856 15804
rect 3792 15744 3856 15748
rect 3872 15804 3936 15808
rect 3872 15748 3876 15804
rect 3876 15748 3932 15804
rect 3932 15748 3936 15804
rect 3872 15744 3936 15748
rect 3952 15804 4016 15808
rect 3952 15748 3956 15804
rect 3956 15748 4012 15804
rect 4012 15748 4016 15804
rect 3952 15744 4016 15748
rect 4032 15804 4096 15808
rect 4032 15748 4036 15804
rect 4036 15748 4092 15804
rect 4092 15748 4096 15804
rect 4032 15744 4096 15748
rect 9473 15804 9537 15808
rect 9473 15748 9477 15804
rect 9477 15748 9533 15804
rect 9533 15748 9537 15804
rect 9473 15744 9537 15748
rect 9553 15804 9617 15808
rect 9553 15748 9557 15804
rect 9557 15748 9613 15804
rect 9613 15748 9617 15804
rect 9553 15744 9617 15748
rect 9633 15804 9697 15808
rect 9633 15748 9637 15804
rect 9637 15748 9693 15804
rect 9693 15748 9697 15804
rect 9633 15744 9697 15748
rect 9713 15804 9777 15808
rect 9713 15748 9717 15804
rect 9717 15748 9773 15804
rect 9773 15748 9777 15804
rect 9713 15744 9777 15748
rect 15154 15804 15218 15808
rect 15154 15748 15158 15804
rect 15158 15748 15214 15804
rect 15214 15748 15218 15804
rect 15154 15744 15218 15748
rect 15234 15804 15298 15808
rect 15234 15748 15238 15804
rect 15238 15748 15294 15804
rect 15294 15748 15298 15804
rect 15234 15744 15298 15748
rect 15314 15804 15378 15808
rect 15314 15748 15318 15804
rect 15318 15748 15374 15804
rect 15374 15748 15378 15804
rect 15314 15744 15378 15748
rect 15394 15804 15458 15808
rect 15394 15748 15398 15804
rect 15398 15748 15454 15804
rect 15454 15748 15458 15804
rect 15394 15744 15458 15748
rect 20835 15804 20899 15808
rect 20835 15748 20839 15804
rect 20839 15748 20895 15804
rect 20895 15748 20899 15804
rect 20835 15744 20899 15748
rect 20915 15804 20979 15808
rect 20915 15748 20919 15804
rect 20919 15748 20975 15804
rect 20975 15748 20979 15804
rect 20915 15744 20979 15748
rect 20995 15804 21059 15808
rect 20995 15748 20999 15804
rect 20999 15748 21055 15804
rect 21055 15748 21059 15804
rect 20995 15744 21059 15748
rect 21075 15804 21139 15808
rect 21075 15748 21079 15804
rect 21079 15748 21135 15804
rect 21135 15748 21139 15804
rect 21075 15744 21139 15748
rect 6632 15260 6696 15264
rect 6632 15204 6636 15260
rect 6636 15204 6692 15260
rect 6692 15204 6696 15260
rect 6632 15200 6696 15204
rect 6712 15260 6776 15264
rect 6712 15204 6716 15260
rect 6716 15204 6772 15260
rect 6772 15204 6776 15260
rect 6712 15200 6776 15204
rect 6792 15260 6856 15264
rect 6792 15204 6796 15260
rect 6796 15204 6852 15260
rect 6852 15204 6856 15260
rect 6792 15200 6856 15204
rect 6872 15260 6936 15264
rect 6872 15204 6876 15260
rect 6876 15204 6932 15260
rect 6932 15204 6936 15260
rect 6872 15200 6936 15204
rect 12313 15260 12377 15264
rect 12313 15204 12317 15260
rect 12317 15204 12373 15260
rect 12373 15204 12377 15260
rect 12313 15200 12377 15204
rect 12393 15260 12457 15264
rect 12393 15204 12397 15260
rect 12397 15204 12453 15260
rect 12453 15204 12457 15260
rect 12393 15200 12457 15204
rect 12473 15260 12537 15264
rect 12473 15204 12477 15260
rect 12477 15204 12533 15260
rect 12533 15204 12537 15260
rect 12473 15200 12537 15204
rect 12553 15260 12617 15264
rect 12553 15204 12557 15260
rect 12557 15204 12613 15260
rect 12613 15204 12617 15260
rect 12553 15200 12617 15204
rect 17994 15260 18058 15264
rect 17994 15204 17998 15260
rect 17998 15204 18054 15260
rect 18054 15204 18058 15260
rect 17994 15200 18058 15204
rect 18074 15260 18138 15264
rect 18074 15204 18078 15260
rect 18078 15204 18134 15260
rect 18134 15204 18138 15260
rect 18074 15200 18138 15204
rect 18154 15260 18218 15264
rect 18154 15204 18158 15260
rect 18158 15204 18214 15260
rect 18214 15204 18218 15260
rect 18154 15200 18218 15204
rect 18234 15260 18298 15264
rect 18234 15204 18238 15260
rect 18238 15204 18294 15260
rect 18294 15204 18298 15260
rect 18234 15200 18298 15204
rect 23675 15260 23739 15264
rect 23675 15204 23679 15260
rect 23679 15204 23735 15260
rect 23735 15204 23739 15260
rect 23675 15200 23739 15204
rect 23755 15260 23819 15264
rect 23755 15204 23759 15260
rect 23759 15204 23815 15260
rect 23815 15204 23819 15260
rect 23755 15200 23819 15204
rect 23835 15260 23899 15264
rect 23835 15204 23839 15260
rect 23839 15204 23895 15260
rect 23895 15204 23899 15260
rect 23835 15200 23899 15204
rect 23915 15260 23979 15264
rect 23915 15204 23919 15260
rect 23919 15204 23975 15260
rect 23975 15204 23979 15260
rect 23915 15200 23979 15204
rect 16436 14996 16500 15060
rect 3792 14716 3856 14720
rect 3792 14660 3796 14716
rect 3796 14660 3852 14716
rect 3852 14660 3856 14716
rect 3792 14656 3856 14660
rect 3872 14716 3936 14720
rect 3872 14660 3876 14716
rect 3876 14660 3932 14716
rect 3932 14660 3936 14716
rect 3872 14656 3936 14660
rect 3952 14716 4016 14720
rect 3952 14660 3956 14716
rect 3956 14660 4012 14716
rect 4012 14660 4016 14716
rect 3952 14656 4016 14660
rect 4032 14716 4096 14720
rect 4032 14660 4036 14716
rect 4036 14660 4092 14716
rect 4092 14660 4096 14716
rect 4032 14656 4096 14660
rect 9473 14716 9537 14720
rect 9473 14660 9477 14716
rect 9477 14660 9533 14716
rect 9533 14660 9537 14716
rect 9473 14656 9537 14660
rect 9553 14716 9617 14720
rect 9553 14660 9557 14716
rect 9557 14660 9613 14716
rect 9613 14660 9617 14716
rect 9553 14656 9617 14660
rect 9633 14716 9697 14720
rect 9633 14660 9637 14716
rect 9637 14660 9693 14716
rect 9693 14660 9697 14716
rect 9633 14656 9697 14660
rect 9713 14716 9777 14720
rect 9713 14660 9717 14716
rect 9717 14660 9773 14716
rect 9773 14660 9777 14716
rect 9713 14656 9777 14660
rect 15154 14716 15218 14720
rect 15154 14660 15158 14716
rect 15158 14660 15214 14716
rect 15214 14660 15218 14716
rect 15154 14656 15218 14660
rect 15234 14716 15298 14720
rect 15234 14660 15238 14716
rect 15238 14660 15294 14716
rect 15294 14660 15298 14716
rect 15234 14656 15298 14660
rect 15314 14716 15378 14720
rect 15314 14660 15318 14716
rect 15318 14660 15374 14716
rect 15374 14660 15378 14716
rect 15314 14656 15378 14660
rect 15394 14716 15458 14720
rect 15394 14660 15398 14716
rect 15398 14660 15454 14716
rect 15454 14660 15458 14716
rect 15394 14656 15458 14660
rect 20835 14716 20899 14720
rect 20835 14660 20839 14716
rect 20839 14660 20895 14716
rect 20895 14660 20899 14716
rect 20835 14656 20899 14660
rect 20915 14716 20979 14720
rect 20915 14660 20919 14716
rect 20919 14660 20975 14716
rect 20975 14660 20979 14716
rect 20915 14656 20979 14660
rect 20995 14716 21059 14720
rect 20995 14660 20999 14716
rect 20999 14660 21055 14716
rect 21055 14660 21059 14716
rect 20995 14656 21059 14660
rect 21075 14716 21139 14720
rect 21075 14660 21079 14716
rect 21079 14660 21135 14716
rect 21135 14660 21139 14716
rect 21075 14656 21139 14660
rect 6632 14172 6696 14176
rect 6632 14116 6636 14172
rect 6636 14116 6692 14172
rect 6692 14116 6696 14172
rect 6632 14112 6696 14116
rect 6712 14172 6776 14176
rect 6712 14116 6716 14172
rect 6716 14116 6772 14172
rect 6772 14116 6776 14172
rect 6712 14112 6776 14116
rect 6792 14172 6856 14176
rect 6792 14116 6796 14172
rect 6796 14116 6852 14172
rect 6852 14116 6856 14172
rect 6792 14112 6856 14116
rect 6872 14172 6936 14176
rect 6872 14116 6876 14172
rect 6876 14116 6932 14172
rect 6932 14116 6936 14172
rect 6872 14112 6936 14116
rect 12313 14172 12377 14176
rect 12313 14116 12317 14172
rect 12317 14116 12373 14172
rect 12373 14116 12377 14172
rect 12313 14112 12377 14116
rect 12393 14172 12457 14176
rect 12393 14116 12397 14172
rect 12397 14116 12453 14172
rect 12453 14116 12457 14172
rect 12393 14112 12457 14116
rect 12473 14172 12537 14176
rect 12473 14116 12477 14172
rect 12477 14116 12533 14172
rect 12533 14116 12537 14172
rect 12473 14112 12537 14116
rect 12553 14172 12617 14176
rect 12553 14116 12557 14172
rect 12557 14116 12613 14172
rect 12613 14116 12617 14172
rect 12553 14112 12617 14116
rect 17994 14172 18058 14176
rect 17994 14116 17998 14172
rect 17998 14116 18054 14172
rect 18054 14116 18058 14172
rect 17994 14112 18058 14116
rect 18074 14172 18138 14176
rect 18074 14116 18078 14172
rect 18078 14116 18134 14172
rect 18134 14116 18138 14172
rect 18074 14112 18138 14116
rect 18154 14172 18218 14176
rect 18154 14116 18158 14172
rect 18158 14116 18214 14172
rect 18214 14116 18218 14172
rect 18154 14112 18218 14116
rect 18234 14172 18298 14176
rect 18234 14116 18238 14172
rect 18238 14116 18294 14172
rect 18294 14116 18298 14172
rect 18234 14112 18298 14116
rect 23675 14172 23739 14176
rect 23675 14116 23679 14172
rect 23679 14116 23735 14172
rect 23735 14116 23739 14172
rect 23675 14112 23739 14116
rect 23755 14172 23819 14176
rect 23755 14116 23759 14172
rect 23759 14116 23815 14172
rect 23815 14116 23819 14172
rect 23755 14112 23819 14116
rect 23835 14172 23899 14176
rect 23835 14116 23839 14172
rect 23839 14116 23895 14172
rect 23895 14116 23899 14172
rect 23835 14112 23899 14116
rect 23915 14172 23979 14176
rect 23915 14116 23919 14172
rect 23919 14116 23975 14172
rect 23975 14116 23979 14172
rect 23915 14112 23979 14116
rect 15700 13772 15764 13836
rect 20116 13772 20180 13836
rect 3792 13628 3856 13632
rect 3792 13572 3796 13628
rect 3796 13572 3852 13628
rect 3852 13572 3856 13628
rect 3792 13568 3856 13572
rect 3872 13628 3936 13632
rect 3872 13572 3876 13628
rect 3876 13572 3932 13628
rect 3932 13572 3936 13628
rect 3872 13568 3936 13572
rect 3952 13628 4016 13632
rect 3952 13572 3956 13628
rect 3956 13572 4012 13628
rect 4012 13572 4016 13628
rect 3952 13568 4016 13572
rect 4032 13628 4096 13632
rect 4032 13572 4036 13628
rect 4036 13572 4092 13628
rect 4092 13572 4096 13628
rect 4032 13568 4096 13572
rect 9473 13628 9537 13632
rect 9473 13572 9477 13628
rect 9477 13572 9533 13628
rect 9533 13572 9537 13628
rect 9473 13568 9537 13572
rect 9553 13628 9617 13632
rect 9553 13572 9557 13628
rect 9557 13572 9613 13628
rect 9613 13572 9617 13628
rect 9553 13568 9617 13572
rect 9633 13628 9697 13632
rect 9633 13572 9637 13628
rect 9637 13572 9693 13628
rect 9693 13572 9697 13628
rect 9633 13568 9697 13572
rect 9713 13628 9777 13632
rect 9713 13572 9717 13628
rect 9717 13572 9773 13628
rect 9773 13572 9777 13628
rect 9713 13568 9777 13572
rect 15154 13628 15218 13632
rect 15154 13572 15158 13628
rect 15158 13572 15214 13628
rect 15214 13572 15218 13628
rect 15154 13568 15218 13572
rect 15234 13628 15298 13632
rect 15234 13572 15238 13628
rect 15238 13572 15294 13628
rect 15294 13572 15298 13628
rect 15234 13568 15298 13572
rect 15314 13628 15378 13632
rect 15314 13572 15318 13628
rect 15318 13572 15374 13628
rect 15374 13572 15378 13628
rect 15314 13568 15378 13572
rect 15394 13628 15458 13632
rect 15394 13572 15398 13628
rect 15398 13572 15454 13628
rect 15454 13572 15458 13628
rect 15394 13568 15458 13572
rect 20835 13628 20899 13632
rect 20835 13572 20839 13628
rect 20839 13572 20895 13628
rect 20895 13572 20899 13628
rect 20835 13568 20899 13572
rect 20915 13628 20979 13632
rect 20915 13572 20919 13628
rect 20919 13572 20975 13628
rect 20975 13572 20979 13628
rect 20915 13568 20979 13572
rect 20995 13628 21059 13632
rect 20995 13572 20999 13628
rect 20999 13572 21055 13628
rect 21055 13572 21059 13628
rect 20995 13568 21059 13572
rect 21075 13628 21139 13632
rect 21075 13572 21079 13628
rect 21079 13572 21135 13628
rect 21135 13572 21139 13628
rect 21075 13568 21139 13572
rect 6632 13084 6696 13088
rect 6632 13028 6636 13084
rect 6636 13028 6692 13084
rect 6692 13028 6696 13084
rect 6632 13024 6696 13028
rect 6712 13084 6776 13088
rect 6712 13028 6716 13084
rect 6716 13028 6772 13084
rect 6772 13028 6776 13084
rect 6712 13024 6776 13028
rect 6792 13084 6856 13088
rect 6792 13028 6796 13084
rect 6796 13028 6852 13084
rect 6852 13028 6856 13084
rect 6792 13024 6856 13028
rect 6872 13084 6936 13088
rect 6872 13028 6876 13084
rect 6876 13028 6932 13084
rect 6932 13028 6936 13084
rect 6872 13024 6936 13028
rect 12313 13084 12377 13088
rect 12313 13028 12317 13084
rect 12317 13028 12373 13084
rect 12373 13028 12377 13084
rect 12313 13024 12377 13028
rect 12393 13084 12457 13088
rect 12393 13028 12397 13084
rect 12397 13028 12453 13084
rect 12453 13028 12457 13084
rect 12393 13024 12457 13028
rect 12473 13084 12537 13088
rect 12473 13028 12477 13084
rect 12477 13028 12533 13084
rect 12533 13028 12537 13084
rect 12473 13024 12537 13028
rect 12553 13084 12617 13088
rect 12553 13028 12557 13084
rect 12557 13028 12613 13084
rect 12613 13028 12617 13084
rect 12553 13024 12617 13028
rect 17994 13084 18058 13088
rect 17994 13028 17998 13084
rect 17998 13028 18054 13084
rect 18054 13028 18058 13084
rect 17994 13024 18058 13028
rect 18074 13084 18138 13088
rect 18074 13028 18078 13084
rect 18078 13028 18134 13084
rect 18134 13028 18138 13084
rect 18074 13024 18138 13028
rect 18154 13084 18218 13088
rect 18154 13028 18158 13084
rect 18158 13028 18214 13084
rect 18214 13028 18218 13084
rect 18154 13024 18218 13028
rect 18234 13084 18298 13088
rect 18234 13028 18238 13084
rect 18238 13028 18294 13084
rect 18294 13028 18298 13084
rect 18234 13024 18298 13028
rect 23675 13084 23739 13088
rect 23675 13028 23679 13084
rect 23679 13028 23735 13084
rect 23735 13028 23739 13084
rect 23675 13024 23739 13028
rect 23755 13084 23819 13088
rect 23755 13028 23759 13084
rect 23759 13028 23815 13084
rect 23815 13028 23819 13084
rect 23755 13024 23819 13028
rect 23835 13084 23899 13088
rect 23835 13028 23839 13084
rect 23839 13028 23895 13084
rect 23895 13028 23899 13084
rect 23835 13024 23899 13028
rect 23915 13084 23979 13088
rect 23915 13028 23919 13084
rect 23919 13028 23975 13084
rect 23975 13028 23979 13084
rect 23915 13024 23979 13028
rect 5028 12548 5092 12612
rect 3792 12540 3856 12544
rect 3792 12484 3796 12540
rect 3796 12484 3852 12540
rect 3852 12484 3856 12540
rect 3792 12480 3856 12484
rect 3872 12540 3936 12544
rect 3872 12484 3876 12540
rect 3876 12484 3932 12540
rect 3932 12484 3936 12540
rect 3872 12480 3936 12484
rect 3952 12540 4016 12544
rect 3952 12484 3956 12540
rect 3956 12484 4012 12540
rect 4012 12484 4016 12540
rect 3952 12480 4016 12484
rect 4032 12540 4096 12544
rect 4032 12484 4036 12540
rect 4036 12484 4092 12540
rect 4092 12484 4096 12540
rect 4032 12480 4096 12484
rect 9473 12540 9537 12544
rect 9473 12484 9477 12540
rect 9477 12484 9533 12540
rect 9533 12484 9537 12540
rect 9473 12480 9537 12484
rect 9553 12540 9617 12544
rect 9553 12484 9557 12540
rect 9557 12484 9613 12540
rect 9613 12484 9617 12540
rect 9553 12480 9617 12484
rect 9633 12540 9697 12544
rect 9633 12484 9637 12540
rect 9637 12484 9693 12540
rect 9693 12484 9697 12540
rect 9633 12480 9697 12484
rect 9713 12540 9777 12544
rect 9713 12484 9717 12540
rect 9717 12484 9773 12540
rect 9773 12484 9777 12540
rect 9713 12480 9777 12484
rect 15154 12540 15218 12544
rect 15154 12484 15158 12540
rect 15158 12484 15214 12540
rect 15214 12484 15218 12540
rect 15154 12480 15218 12484
rect 15234 12540 15298 12544
rect 15234 12484 15238 12540
rect 15238 12484 15294 12540
rect 15294 12484 15298 12540
rect 15234 12480 15298 12484
rect 15314 12540 15378 12544
rect 15314 12484 15318 12540
rect 15318 12484 15374 12540
rect 15374 12484 15378 12540
rect 15314 12480 15378 12484
rect 15394 12540 15458 12544
rect 15394 12484 15398 12540
rect 15398 12484 15454 12540
rect 15454 12484 15458 12540
rect 15394 12480 15458 12484
rect 20835 12540 20899 12544
rect 20835 12484 20839 12540
rect 20839 12484 20895 12540
rect 20895 12484 20899 12540
rect 20835 12480 20899 12484
rect 20915 12540 20979 12544
rect 20915 12484 20919 12540
rect 20919 12484 20975 12540
rect 20975 12484 20979 12540
rect 20915 12480 20979 12484
rect 20995 12540 21059 12544
rect 20995 12484 20999 12540
rect 20999 12484 21055 12540
rect 21055 12484 21059 12540
rect 20995 12480 21059 12484
rect 21075 12540 21139 12544
rect 21075 12484 21079 12540
rect 21079 12484 21135 12540
rect 21135 12484 21139 12540
rect 21075 12480 21139 12484
rect 4292 12276 4356 12340
rect 6316 12140 6380 12204
rect 12940 12140 13004 12204
rect 8524 12064 8588 12068
rect 8524 12008 8538 12064
rect 8538 12008 8588 12064
rect 8524 12004 8588 12008
rect 6632 11996 6696 12000
rect 6632 11940 6636 11996
rect 6636 11940 6692 11996
rect 6692 11940 6696 11996
rect 6632 11936 6696 11940
rect 6712 11996 6776 12000
rect 6712 11940 6716 11996
rect 6716 11940 6772 11996
rect 6772 11940 6776 11996
rect 6712 11936 6776 11940
rect 6792 11996 6856 12000
rect 6792 11940 6796 11996
rect 6796 11940 6852 11996
rect 6852 11940 6856 11996
rect 6792 11936 6856 11940
rect 6872 11996 6936 12000
rect 6872 11940 6876 11996
rect 6876 11940 6932 11996
rect 6932 11940 6936 11996
rect 6872 11936 6936 11940
rect 12313 11996 12377 12000
rect 12313 11940 12317 11996
rect 12317 11940 12373 11996
rect 12373 11940 12377 11996
rect 12313 11936 12377 11940
rect 12393 11996 12457 12000
rect 12393 11940 12397 11996
rect 12397 11940 12453 11996
rect 12453 11940 12457 11996
rect 12393 11936 12457 11940
rect 12473 11996 12537 12000
rect 12473 11940 12477 11996
rect 12477 11940 12533 11996
rect 12533 11940 12537 11996
rect 12473 11936 12537 11940
rect 12553 11996 12617 12000
rect 12553 11940 12557 11996
rect 12557 11940 12613 11996
rect 12613 11940 12617 11996
rect 12553 11936 12617 11940
rect 17994 11996 18058 12000
rect 17994 11940 17998 11996
rect 17998 11940 18054 11996
rect 18054 11940 18058 11996
rect 17994 11936 18058 11940
rect 18074 11996 18138 12000
rect 18074 11940 18078 11996
rect 18078 11940 18134 11996
rect 18134 11940 18138 11996
rect 18074 11936 18138 11940
rect 18154 11996 18218 12000
rect 18154 11940 18158 11996
rect 18158 11940 18214 11996
rect 18214 11940 18218 11996
rect 18154 11936 18218 11940
rect 18234 11996 18298 12000
rect 18234 11940 18238 11996
rect 18238 11940 18294 11996
rect 18294 11940 18298 11996
rect 18234 11936 18298 11940
rect 23675 11996 23739 12000
rect 23675 11940 23679 11996
rect 23679 11940 23735 11996
rect 23735 11940 23739 11996
rect 23675 11936 23739 11940
rect 23755 11996 23819 12000
rect 23755 11940 23759 11996
rect 23759 11940 23815 11996
rect 23815 11940 23819 11996
rect 23755 11936 23819 11940
rect 23835 11996 23899 12000
rect 23835 11940 23839 11996
rect 23839 11940 23895 11996
rect 23895 11940 23899 11996
rect 23835 11936 23899 11940
rect 23915 11996 23979 12000
rect 23915 11940 23919 11996
rect 23919 11940 23975 11996
rect 23975 11940 23979 11996
rect 23915 11936 23979 11940
rect 4292 11928 4356 11932
rect 4292 11872 4306 11928
rect 4306 11872 4356 11928
rect 4292 11868 4356 11872
rect 8156 11928 8220 11932
rect 8156 11872 8170 11928
rect 8170 11872 8220 11928
rect 8156 11868 8220 11872
rect 3792 11452 3856 11456
rect 3792 11396 3796 11452
rect 3796 11396 3852 11452
rect 3852 11396 3856 11452
rect 3792 11392 3856 11396
rect 3872 11452 3936 11456
rect 3872 11396 3876 11452
rect 3876 11396 3932 11452
rect 3932 11396 3936 11452
rect 3872 11392 3936 11396
rect 3952 11452 4016 11456
rect 3952 11396 3956 11452
rect 3956 11396 4012 11452
rect 4012 11396 4016 11452
rect 3952 11392 4016 11396
rect 4032 11452 4096 11456
rect 4032 11396 4036 11452
rect 4036 11396 4092 11452
rect 4092 11396 4096 11452
rect 4032 11392 4096 11396
rect 9473 11452 9537 11456
rect 9473 11396 9477 11452
rect 9477 11396 9533 11452
rect 9533 11396 9537 11452
rect 9473 11392 9537 11396
rect 9553 11452 9617 11456
rect 9553 11396 9557 11452
rect 9557 11396 9613 11452
rect 9613 11396 9617 11452
rect 9553 11392 9617 11396
rect 9633 11452 9697 11456
rect 9633 11396 9637 11452
rect 9637 11396 9693 11452
rect 9693 11396 9697 11452
rect 9633 11392 9697 11396
rect 9713 11452 9777 11456
rect 9713 11396 9717 11452
rect 9717 11396 9773 11452
rect 9773 11396 9777 11452
rect 9713 11392 9777 11396
rect 15154 11452 15218 11456
rect 15154 11396 15158 11452
rect 15158 11396 15214 11452
rect 15214 11396 15218 11452
rect 15154 11392 15218 11396
rect 15234 11452 15298 11456
rect 15234 11396 15238 11452
rect 15238 11396 15294 11452
rect 15294 11396 15298 11452
rect 15234 11392 15298 11396
rect 15314 11452 15378 11456
rect 15314 11396 15318 11452
rect 15318 11396 15374 11452
rect 15374 11396 15378 11452
rect 15314 11392 15378 11396
rect 15394 11452 15458 11456
rect 15394 11396 15398 11452
rect 15398 11396 15454 11452
rect 15454 11396 15458 11452
rect 15394 11392 15458 11396
rect 20835 11452 20899 11456
rect 20835 11396 20839 11452
rect 20839 11396 20895 11452
rect 20895 11396 20899 11452
rect 20835 11392 20899 11396
rect 20915 11452 20979 11456
rect 20915 11396 20919 11452
rect 20919 11396 20975 11452
rect 20975 11396 20979 11452
rect 20915 11392 20979 11396
rect 20995 11452 21059 11456
rect 20995 11396 20999 11452
rect 20999 11396 21055 11452
rect 21055 11396 21059 11452
rect 20995 11392 21059 11396
rect 21075 11452 21139 11456
rect 21075 11396 21079 11452
rect 21079 11396 21135 11452
rect 21135 11396 21139 11452
rect 21075 11392 21139 11396
rect 7604 11248 7668 11252
rect 7604 11192 7618 11248
rect 7618 11192 7668 11248
rect 7604 11188 7668 11192
rect 6632 10908 6696 10912
rect 6632 10852 6636 10908
rect 6636 10852 6692 10908
rect 6692 10852 6696 10908
rect 6632 10848 6696 10852
rect 6712 10908 6776 10912
rect 6712 10852 6716 10908
rect 6716 10852 6772 10908
rect 6772 10852 6776 10908
rect 6712 10848 6776 10852
rect 6792 10908 6856 10912
rect 6792 10852 6796 10908
rect 6796 10852 6852 10908
rect 6852 10852 6856 10908
rect 6792 10848 6856 10852
rect 6872 10908 6936 10912
rect 6872 10852 6876 10908
rect 6876 10852 6932 10908
rect 6932 10852 6936 10908
rect 6872 10848 6936 10852
rect 12313 10908 12377 10912
rect 12313 10852 12317 10908
rect 12317 10852 12373 10908
rect 12373 10852 12377 10908
rect 12313 10848 12377 10852
rect 12393 10908 12457 10912
rect 12393 10852 12397 10908
rect 12397 10852 12453 10908
rect 12453 10852 12457 10908
rect 12393 10848 12457 10852
rect 12473 10908 12537 10912
rect 12473 10852 12477 10908
rect 12477 10852 12533 10908
rect 12533 10852 12537 10908
rect 12473 10848 12537 10852
rect 12553 10908 12617 10912
rect 12553 10852 12557 10908
rect 12557 10852 12613 10908
rect 12613 10852 12617 10908
rect 12553 10848 12617 10852
rect 17994 10908 18058 10912
rect 17994 10852 17998 10908
rect 17998 10852 18054 10908
rect 18054 10852 18058 10908
rect 17994 10848 18058 10852
rect 18074 10908 18138 10912
rect 18074 10852 18078 10908
rect 18078 10852 18134 10908
rect 18134 10852 18138 10908
rect 18074 10848 18138 10852
rect 18154 10908 18218 10912
rect 18154 10852 18158 10908
rect 18158 10852 18214 10908
rect 18214 10852 18218 10908
rect 18154 10848 18218 10852
rect 18234 10908 18298 10912
rect 18234 10852 18238 10908
rect 18238 10852 18294 10908
rect 18294 10852 18298 10908
rect 18234 10848 18298 10852
rect 23675 10908 23739 10912
rect 23675 10852 23679 10908
rect 23679 10852 23735 10908
rect 23735 10852 23739 10908
rect 23675 10848 23739 10852
rect 23755 10908 23819 10912
rect 23755 10852 23759 10908
rect 23759 10852 23815 10908
rect 23815 10852 23819 10908
rect 23755 10848 23819 10852
rect 23835 10908 23899 10912
rect 23835 10852 23839 10908
rect 23839 10852 23895 10908
rect 23895 10852 23899 10908
rect 23835 10848 23899 10852
rect 23915 10908 23979 10912
rect 23915 10852 23919 10908
rect 23919 10852 23975 10908
rect 23975 10852 23979 10908
rect 23915 10848 23979 10852
rect 3792 10364 3856 10368
rect 3792 10308 3796 10364
rect 3796 10308 3852 10364
rect 3852 10308 3856 10364
rect 3792 10304 3856 10308
rect 3872 10364 3936 10368
rect 3872 10308 3876 10364
rect 3876 10308 3932 10364
rect 3932 10308 3936 10364
rect 3872 10304 3936 10308
rect 3952 10364 4016 10368
rect 3952 10308 3956 10364
rect 3956 10308 4012 10364
rect 4012 10308 4016 10364
rect 3952 10304 4016 10308
rect 4032 10364 4096 10368
rect 4032 10308 4036 10364
rect 4036 10308 4092 10364
rect 4092 10308 4096 10364
rect 4032 10304 4096 10308
rect 9473 10364 9537 10368
rect 9473 10308 9477 10364
rect 9477 10308 9533 10364
rect 9533 10308 9537 10364
rect 9473 10304 9537 10308
rect 9553 10364 9617 10368
rect 9553 10308 9557 10364
rect 9557 10308 9613 10364
rect 9613 10308 9617 10364
rect 9553 10304 9617 10308
rect 9633 10364 9697 10368
rect 9633 10308 9637 10364
rect 9637 10308 9693 10364
rect 9693 10308 9697 10364
rect 9633 10304 9697 10308
rect 9713 10364 9777 10368
rect 9713 10308 9717 10364
rect 9717 10308 9773 10364
rect 9773 10308 9777 10364
rect 9713 10304 9777 10308
rect 15154 10364 15218 10368
rect 15154 10308 15158 10364
rect 15158 10308 15214 10364
rect 15214 10308 15218 10364
rect 15154 10304 15218 10308
rect 15234 10364 15298 10368
rect 15234 10308 15238 10364
rect 15238 10308 15294 10364
rect 15294 10308 15298 10364
rect 15234 10304 15298 10308
rect 15314 10364 15378 10368
rect 15314 10308 15318 10364
rect 15318 10308 15374 10364
rect 15374 10308 15378 10364
rect 15314 10304 15378 10308
rect 15394 10364 15458 10368
rect 15394 10308 15398 10364
rect 15398 10308 15454 10364
rect 15454 10308 15458 10364
rect 15394 10304 15458 10308
rect 20835 10364 20899 10368
rect 20835 10308 20839 10364
rect 20839 10308 20895 10364
rect 20895 10308 20899 10364
rect 20835 10304 20899 10308
rect 20915 10364 20979 10368
rect 20915 10308 20919 10364
rect 20919 10308 20975 10364
rect 20975 10308 20979 10364
rect 20915 10304 20979 10308
rect 20995 10364 21059 10368
rect 20995 10308 20999 10364
rect 20999 10308 21055 10364
rect 21055 10308 21059 10364
rect 20995 10304 21059 10308
rect 21075 10364 21139 10368
rect 21075 10308 21079 10364
rect 21079 10308 21135 10364
rect 21135 10308 21139 10364
rect 21075 10304 21139 10308
rect 12940 9888 13004 9892
rect 12940 9832 12954 9888
rect 12954 9832 13004 9888
rect 12940 9828 13004 9832
rect 6632 9820 6696 9824
rect 6632 9764 6636 9820
rect 6636 9764 6692 9820
rect 6692 9764 6696 9820
rect 6632 9760 6696 9764
rect 6712 9820 6776 9824
rect 6712 9764 6716 9820
rect 6716 9764 6772 9820
rect 6772 9764 6776 9820
rect 6712 9760 6776 9764
rect 6792 9820 6856 9824
rect 6792 9764 6796 9820
rect 6796 9764 6852 9820
rect 6852 9764 6856 9820
rect 6792 9760 6856 9764
rect 6872 9820 6936 9824
rect 6872 9764 6876 9820
rect 6876 9764 6932 9820
rect 6932 9764 6936 9820
rect 6872 9760 6936 9764
rect 12313 9820 12377 9824
rect 12313 9764 12317 9820
rect 12317 9764 12373 9820
rect 12373 9764 12377 9820
rect 12313 9760 12377 9764
rect 12393 9820 12457 9824
rect 12393 9764 12397 9820
rect 12397 9764 12453 9820
rect 12453 9764 12457 9820
rect 12393 9760 12457 9764
rect 12473 9820 12537 9824
rect 12473 9764 12477 9820
rect 12477 9764 12533 9820
rect 12533 9764 12537 9820
rect 12473 9760 12537 9764
rect 12553 9820 12617 9824
rect 12553 9764 12557 9820
rect 12557 9764 12613 9820
rect 12613 9764 12617 9820
rect 12553 9760 12617 9764
rect 17994 9820 18058 9824
rect 17994 9764 17998 9820
rect 17998 9764 18054 9820
rect 18054 9764 18058 9820
rect 17994 9760 18058 9764
rect 18074 9820 18138 9824
rect 18074 9764 18078 9820
rect 18078 9764 18134 9820
rect 18134 9764 18138 9820
rect 18074 9760 18138 9764
rect 18154 9820 18218 9824
rect 18154 9764 18158 9820
rect 18158 9764 18214 9820
rect 18214 9764 18218 9820
rect 18154 9760 18218 9764
rect 18234 9820 18298 9824
rect 18234 9764 18238 9820
rect 18238 9764 18294 9820
rect 18294 9764 18298 9820
rect 18234 9760 18298 9764
rect 23675 9820 23739 9824
rect 23675 9764 23679 9820
rect 23679 9764 23735 9820
rect 23735 9764 23739 9820
rect 23675 9760 23739 9764
rect 23755 9820 23819 9824
rect 23755 9764 23759 9820
rect 23759 9764 23815 9820
rect 23815 9764 23819 9820
rect 23755 9760 23819 9764
rect 23835 9820 23899 9824
rect 23835 9764 23839 9820
rect 23839 9764 23895 9820
rect 23895 9764 23899 9820
rect 23835 9760 23899 9764
rect 23915 9820 23979 9824
rect 23915 9764 23919 9820
rect 23919 9764 23975 9820
rect 23975 9764 23979 9820
rect 23915 9760 23979 9764
rect 8340 9752 8404 9756
rect 8340 9696 8390 9752
rect 8390 9696 8404 9752
rect 8340 9692 8404 9696
rect 9260 9752 9324 9756
rect 9260 9696 9310 9752
rect 9310 9696 9324 9752
rect 9260 9692 9324 9696
rect 10916 9752 10980 9756
rect 10916 9696 10966 9752
rect 10966 9696 10980 9752
rect 10916 9692 10980 9696
rect 7420 9420 7484 9484
rect 20300 9420 20364 9484
rect 7972 9284 8036 9348
rect 3792 9276 3856 9280
rect 3792 9220 3796 9276
rect 3796 9220 3852 9276
rect 3852 9220 3856 9276
rect 3792 9216 3856 9220
rect 3872 9276 3936 9280
rect 3872 9220 3876 9276
rect 3876 9220 3932 9276
rect 3932 9220 3936 9276
rect 3872 9216 3936 9220
rect 3952 9276 4016 9280
rect 3952 9220 3956 9276
rect 3956 9220 4012 9276
rect 4012 9220 4016 9276
rect 3952 9216 4016 9220
rect 4032 9276 4096 9280
rect 4032 9220 4036 9276
rect 4036 9220 4092 9276
rect 4092 9220 4096 9276
rect 4032 9216 4096 9220
rect 9473 9276 9537 9280
rect 9473 9220 9477 9276
rect 9477 9220 9533 9276
rect 9533 9220 9537 9276
rect 9473 9216 9537 9220
rect 9553 9276 9617 9280
rect 9553 9220 9557 9276
rect 9557 9220 9613 9276
rect 9613 9220 9617 9276
rect 9553 9216 9617 9220
rect 9633 9276 9697 9280
rect 9633 9220 9637 9276
rect 9637 9220 9693 9276
rect 9693 9220 9697 9276
rect 9633 9216 9697 9220
rect 9713 9276 9777 9280
rect 9713 9220 9717 9276
rect 9717 9220 9773 9276
rect 9773 9220 9777 9276
rect 9713 9216 9777 9220
rect 15154 9276 15218 9280
rect 15154 9220 15158 9276
rect 15158 9220 15214 9276
rect 15214 9220 15218 9276
rect 15154 9216 15218 9220
rect 15234 9276 15298 9280
rect 15234 9220 15238 9276
rect 15238 9220 15294 9276
rect 15294 9220 15298 9276
rect 15234 9216 15298 9220
rect 15314 9276 15378 9280
rect 15314 9220 15318 9276
rect 15318 9220 15374 9276
rect 15374 9220 15378 9276
rect 15314 9216 15378 9220
rect 15394 9276 15458 9280
rect 15394 9220 15398 9276
rect 15398 9220 15454 9276
rect 15454 9220 15458 9276
rect 15394 9216 15458 9220
rect 20835 9276 20899 9280
rect 20835 9220 20839 9276
rect 20839 9220 20895 9276
rect 20895 9220 20899 9276
rect 20835 9216 20899 9220
rect 20915 9276 20979 9280
rect 20915 9220 20919 9276
rect 20919 9220 20975 9276
rect 20975 9220 20979 9276
rect 20915 9216 20979 9220
rect 20995 9276 21059 9280
rect 20995 9220 20999 9276
rect 20999 9220 21055 9276
rect 21055 9220 21059 9276
rect 20995 9216 21059 9220
rect 21075 9276 21139 9280
rect 21075 9220 21079 9276
rect 21079 9220 21135 9276
rect 21135 9220 21139 9276
rect 21075 9216 21139 9220
rect 16436 9208 16500 9212
rect 16436 9152 16486 9208
rect 16486 9152 16500 9208
rect 16436 9148 16500 9152
rect 6632 8732 6696 8736
rect 6632 8676 6636 8732
rect 6636 8676 6692 8732
rect 6692 8676 6696 8732
rect 6632 8672 6696 8676
rect 6712 8732 6776 8736
rect 6712 8676 6716 8732
rect 6716 8676 6772 8732
rect 6772 8676 6776 8732
rect 6712 8672 6776 8676
rect 6792 8732 6856 8736
rect 6792 8676 6796 8732
rect 6796 8676 6852 8732
rect 6852 8676 6856 8732
rect 6792 8672 6856 8676
rect 6872 8732 6936 8736
rect 6872 8676 6876 8732
rect 6876 8676 6932 8732
rect 6932 8676 6936 8732
rect 6872 8672 6936 8676
rect 12313 8732 12377 8736
rect 12313 8676 12317 8732
rect 12317 8676 12373 8732
rect 12373 8676 12377 8732
rect 12313 8672 12377 8676
rect 12393 8732 12457 8736
rect 12393 8676 12397 8732
rect 12397 8676 12453 8732
rect 12453 8676 12457 8732
rect 12393 8672 12457 8676
rect 12473 8732 12537 8736
rect 12473 8676 12477 8732
rect 12477 8676 12533 8732
rect 12533 8676 12537 8732
rect 12473 8672 12537 8676
rect 12553 8732 12617 8736
rect 12553 8676 12557 8732
rect 12557 8676 12613 8732
rect 12613 8676 12617 8732
rect 12553 8672 12617 8676
rect 17994 8732 18058 8736
rect 17994 8676 17998 8732
rect 17998 8676 18054 8732
rect 18054 8676 18058 8732
rect 17994 8672 18058 8676
rect 18074 8732 18138 8736
rect 18074 8676 18078 8732
rect 18078 8676 18134 8732
rect 18134 8676 18138 8732
rect 18074 8672 18138 8676
rect 18154 8732 18218 8736
rect 18154 8676 18158 8732
rect 18158 8676 18214 8732
rect 18214 8676 18218 8732
rect 18154 8672 18218 8676
rect 18234 8732 18298 8736
rect 18234 8676 18238 8732
rect 18238 8676 18294 8732
rect 18294 8676 18298 8732
rect 18234 8672 18298 8676
rect 23675 8732 23739 8736
rect 23675 8676 23679 8732
rect 23679 8676 23735 8732
rect 23735 8676 23739 8732
rect 23675 8672 23739 8676
rect 23755 8732 23819 8736
rect 23755 8676 23759 8732
rect 23759 8676 23815 8732
rect 23815 8676 23819 8732
rect 23755 8672 23819 8676
rect 23835 8732 23899 8736
rect 23835 8676 23839 8732
rect 23839 8676 23895 8732
rect 23895 8676 23899 8732
rect 23835 8672 23899 8676
rect 23915 8732 23979 8736
rect 23915 8676 23919 8732
rect 23919 8676 23975 8732
rect 23975 8676 23979 8732
rect 23915 8672 23979 8676
rect 7788 8332 7852 8396
rect 3792 8188 3856 8192
rect 3792 8132 3796 8188
rect 3796 8132 3852 8188
rect 3852 8132 3856 8188
rect 3792 8128 3856 8132
rect 3872 8188 3936 8192
rect 3872 8132 3876 8188
rect 3876 8132 3932 8188
rect 3932 8132 3936 8188
rect 3872 8128 3936 8132
rect 3952 8188 4016 8192
rect 3952 8132 3956 8188
rect 3956 8132 4012 8188
rect 4012 8132 4016 8188
rect 3952 8128 4016 8132
rect 4032 8188 4096 8192
rect 4032 8132 4036 8188
rect 4036 8132 4092 8188
rect 4092 8132 4096 8188
rect 4032 8128 4096 8132
rect 9473 8188 9537 8192
rect 9473 8132 9477 8188
rect 9477 8132 9533 8188
rect 9533 8132 9537 8188
rect 9473 8128 9537 8132
rect 9553 8188 9617 8192
rect 9553 8132 9557 8188
rect 9557 8132 9613 8188
rect 9613 8132 9617 8188
rect 9553 8128 9617 8132
rect 9633 8188 9697 8192
rect 9633 8132 9637 8188
rect 9637 8132 9693 8188
rect 9693 8132 9697 8188
rect 9633 8128 9697 8132
rect 9713 8188 9777 8192
rect 9713 8132 9717 8188
rect 9717 8132 9773 8188
rect 9773 8132 9777 8188
rect 9713 8128 9777 8132
rect 15154 8188 15218 8192
rect 15154 8132 15158 8188
rect 15158 8132 15214 8188
rect 15214 8132 15218 8188
rect 15154 8128 15218 8132
rect 15234 8188 15298 8192
rect 15234 8132 15238 8188
rect 15238 8132 15294 8188
rect 15294 8132 15298 8188
rect 15234 8128 15298 8132
rect 15314 8188 15378 8192
rect 15314 8132 15318 8188
rect 15318 8132 15374 8188
rect 15374 8132 15378 8188
rect 15314 8128 15378 8132
rect 15394 8188 15458 8192
rect 15394 8132 15398 8188
rect 15398 8132 15454 8188
rect 15454 8132 15458 8188
rect 15394 8128 15458 8132
rect 20835 8188 20899 8192
rect 20835 8132 20839 8188
rect 20839 8132 20895 8188
rect 20895 8132 20899 8188
rect 20835 8128 20899 8132
rect 20915 8188 20979 8192
rect 20915 8132 20919 8188
rect 20919 8132 20975 8188
rect 20975 8132 20979 8188
rect 20915 8128 20979 8132
rect 20995 8188 21059 8192
rect 20995 8132 20999 8188
rect 20999 8132 21055 8188
rect 21055 8132 21059 8188
rect 20995 8128 21059 8132
rect 21075 8188 21139 8192
rect 21075 8132 21079 8188
rect 21079 8132 21135 8188
rect 21135 8132 21139 8188
rect 21075 8128 21139 8132
rect 20116 8060 20180 8124
rect 10916 7924 10980 7988
rect 6632 7644 6696 7648
rect 6632 7588 6636 7644
rect 6636 7588 6692 7644
rect 6692 7588 6696 7644
rect 6632 7584 6696 7588
rect 6712 7644 6776 7648
rect 6712 7588 6716 7644
rect 6716 7588 6772 7644
rect 6772 7588 6776 7644
rect 6712 7584 6776 7588
rect 6792 7644 6856 7648
rect 6792 7588 6796 7644
rect 6796 7588 6852 7644
rect 6852 7588 6856 7644
rect 6792 7584 6856 7588
rect 6872 7644 6936 7648
rect 6872 7588 6876 7644
rect 6876 7588 6932 7644
rect 6932 7588 6936 7644
rect 6872 7584 6936 7588
rect 12313 7644 12377 7648
rect 12313 7588 12317 7644
rect 12317 7588 12373 7644
rect 12373 7588 12377 7644
rect 12313 7584 12377 7588
rect 12393 7644 12457 7648
rect 12393 7588 12397 7644
rect 12397 7588 12453 7644
rect 12453 7588 12457 7644
rect 12393 7584 12457 7588
rect 12473 7644 12537 7648
rect 12473 7588 12477 7644
rect 12477 7588 12533 7644
rect 12533 7588 12537 7644
rect 12473 7584 12537 7588
rect 12553 7644 12617 7648
rect 12553 7588 12557 7644
rect 12557 7588 12613 7644
rect 12613 7588 12617 7644
rect 12553 7584 12617 7588
rect 17994 7644 18058 7648
rect 17994 7588 17998 7644
rect 17998 7588 18054 7644
rect 18054 7588 18058 7644
rect 17994 7584 18058 7588
rect 18074 7644 18138 7648
rect 18074 7588 18078 7644
rect 18078 7588 18134 7644
rect 18134 7588 18138 7644
rect 18074 7584 18138 7588
rect 18154 7644 18218 7648
rect 18154 7588 18158 7644
rect 18158 7588 18214 7644
rect 18214 7588 18218 7644
rect 18154 7584 18218 7588
rect 18234 7644 18298 7648
rect 18234 7588 18238 7644
rect 18238 7588 18294 7644
rect 18294 7588 18298 7644
rect 18234 7584 18298 7588
rect 23675 7644 23739 7648
rect 23675 7588 23679 7644
rect 23679 7588 23735 7644
rect 23735 7588 23739 7644
rect 23675 7584 23739 7588
rect 23755 7644 23819 7648
rect 23755 7588 23759 7644
rect 23759 7588 23815 7644
rect 23815 7588 23819 7644
rect 23755 7584 23819 7588
rect 23835 7644 23899 7648
rect 23835 7588 23839 7644
rect 23839 7588 23895 7644
rect 23895 7588 23899 7644
rect 23835 7584 23899 7588
rect 23915 7644 23979 7648
rect 23915 7588 23919 7644
rect 23919 7588 23975 7644
rect 23975 7588 23979 7644
rect 23915 7584 23979 7588
rect 3372 7380 3436 7444
rect 3792 7100 3856 7104
rect 3792 7044 3796 7100
rect 3796 7044 3852 7100
rect 3852 7044 3856 7100
rect 3792 7040 3856 7044
rect 3872 7100 3936 7104
rect 3872 7044 3876 7100
rect 3876 7044 3932 7100
rect 3932 7044 3936 7100
rect 3872 7040 3936 7044
rect 3952 7100 4016 7104
rect 3952 7044 3956 7100
rect 3956 7044 4012 7100
rect 4012 7044 4016 7100
rect 3952 7040 4016 7044
rect 4032 7100 4096 7104
rect 4032 7044 4036 7100
rect 4036 7044 4092 7100
rect 4092 7044 4096 7100
rect 4032 7040 4096 7044
rect 9473 7100 9537 7104
rect 9473 7044 9477 7100
rect 9477 7044 9533 7100
rect 9533 7044 9537 7100
rect 9473 7040 9537 7044
rect 9553 7100 9617 7104
rect 9553 7044 9557 7100
rect 9557 7044 9613 7100
rect 9613 7044 9617 7100
rect 9553 7040 9617 7044
rect 9633 7100 9697 7104
rect 9633 7044 9637 7100
rect 9637 7044 9693 7100
rect 9693 7044 9697 7100
rect 9633 7040 9697 7044
rect 9713 7100 9777 7104
rect 9713 7044 9717 7100
rect 9717 7044 9773 7100
rect 9773 7044 9777 7100
rect 9713 7040 9777 7044
rect 15154 7100 15218 7104
rect 15154 7044 15158 7100
rect 15158 7044 15214 7100
rect 15214 7044 15218 7100
rect 15154 7040 15218 7044
rect 15234 7100 15298 7104
rect 15234 7044 15238 7100
rect 15238 7044 15294 7100
rect 15294 7044 15298 7100
rect 15234 7040 15298 7044
rect 15314 7100 15378 7104
rect 15314 7044 15318 7100
rect 15318 7044 15374 7100
rect 15374 7044 15378 7100
rect 15314 7040 15378 7044
rect 15394 7100 15458 7104
rect 15394 7044 15398 7100
rect 15398 7044 15454 7100
rect 15454 7044 15458 7100
rect 15394 7040 15458 7044
rect 20835 7100 20899 7104
rect 20835 7044 20839 7100
rect 20839 7044 20895 7100
rect 20895 7044 20899 7100
rect 20835 7040 20899 7044
rect 20915 7100 20979 7104
rect 20915 7044 20919 7100
rect 20919 7044 20975 7100
rect 20975 7044 20979 7100
rect 20915 7040 20979 7044
rect 20995 7100 21059 7104
rect 20995 7044 20999 7100
rect 20999 7044 21055 7100
rect 21055 7044 21059 7100
rect 20995 7040 21059 7044
rect 21075 7100 21139 7104
rect 21075 7044 21079 7100
rect 21079 7044 21135 7100
rect 21135 7044 21139 7100
rect 21075 7040 21139 7044
rect 6632 6556 6696 6560
rect 6632 6500 6636 6556
rect 6636 6500 6692 6556
rect 6692 6500 6696 6556
rect 6632 6496 6696 6500
rect 6712 6556 6776 6560
rect 6712 6500 6716 6556
rect 6716 6500 6772 6556
rect 6772 6500 6776 6556
rect 6712 6496 6776 6500
rect 6792 6556 6856 6560
rect 6792 6500 6796 6556
rect 6796 6500 6852 6556
rect 6852 6500 6856 6556
rect 6792 6496 6856 6500
rect 6872 6556 6936 6560
rect 6872 6500 6876 6556
rect 6876 6500 6932 6556
rect 6932 6500 6936 6556
rect 6872 6496 6936 6500
rect 12313 6556 12377 6560
rect 12313 6500 12317 6556
rect 12317 6500 12373 6556
rect 12373 6500 12377 6556
rect 12313 6496 12377 6500
rect 12393 6556 12457 6560
rect 12393 6500 12397 6556
rect 12397 6500 12453 6556
rect 12453 6500 12457 6556
rect 12393 6496 12457 6500
rect 12473 6556 12537 6560
rect 12473 6500 12477 6556
rect 12477 6500 12533 6556
rect 12533 6500 12537 6556
rect 12473 6496 12537 6500
rect 12553 6556 12617 6560
rect 12553 6500 12557 6556
rect 12557 6500 12613 6556
rect 12613 6500 12617 6556
rect 12553 6496 12617 6500
rect 17994 6556 18058 6560
rect 17994 6500 17998 6556
rect 17998 6500 18054 6556
rect 18054 6500 18058 6556
rect 17994 6496 18058 6500
rect 18074 6556 18138 6560
rect 18074 6500 18078 6556
rect 18078 6500 18134 6556
rect 18134 6500 18138 6556
rect 18074 6496 18138 6500
rect 18154 6556 18218 6560
rect 18154 6500 18158 6556
rect 18158 6500 18214 6556
rect 18214 6500 18218 6556
rect 18154 6496 18218 6500
rect 18234 6556 18298 6560
rect 18234 6500 18238 6556
rect 18238 6500 18294 6556
rect 18294 6500 18298 6556
rect 18234 6496 18298 6500
rect 23675 6556 23739 6560
rect 23675 6500 23679 6556
rect 23679 6500 23735 6556
rect 23735 6500 23739 6556
rect 23675 6496 23739 6500
rect 23755 6556 23819 6560
rect 23755 6500 23759 6556
rect 23759 6500 23815 6556
rect 23815 6500 23819 6556
rect 23755 6496 23819 6500
rect 23835 6556 23899 6560
rect 23835 6500 23839 6556
rect 23839 6500 23895 6556
rect 23895 6500 23899 6556
rect 23835 6496 23899 6500
rect 23915 6556 23979 6560
rect 23915 6500 23919 6556
rect 23919 6500 23975 6556
rect 23975 6500 23979 6556
rect 23915 6496 23979 6500
rect 15700 6428 15764 6492
rect 3792 6012 3856 6016
rect 3792 5956 3796 6012
rect 3796 5956 3852 6012
rect 3852 5956 3856 6012
rect 3792 5952 3856 5956
rect 3872 6012 3936 6016
rect 3872 5956 3876 6012
rect 3876 5956 3932 6012
rect 3932 5956 3936 6012
rect 3872 5952 3936 5956
rect 3952 6012 4016 6016
rect 3952 5956 3956 6012
rect 3956 5956 4012 6012
rect 4012 5956 4016 6012
rect 3952 5952 4016 5956
rect 4032 6012 4096 6016
rect 4032 5956 4036 6012
rect 4036 5956 4092 6012
rect 4092 5956 4096 6012
rect 4032 5952 4096 5956
rect 9473 6012 9537 6016
rect 9473 5956 9477 6012
rect 9477 5956 9533 6012
rect 9533 5956 9537 6012
rect 9473 5952 9537 5956
rect 9553 6012 9617 6016
rect 9553 5956 9557 6012
rect 9557 5956 9613 6012
rect 9613 5956 9617 6012
rect 9553 5952 9617 5956
rect 9633 6012 9697 6016
rect 9633 5956 9637 6012
rect 9637 5956 9693 6012
rect 9693 5956 9697 6012
rect 9633 5952 9697 5956
rect 9713 6012 9777 6016
rect 9713 5956 9717 6012
rect 9717 5956 9773 6012
rect 9773 5956 9777 6012
rect 9713 5952 9777 5956
rect 15154 6012 15218 6016
rect 15154 5956 15158 6012
rect 15158 5956 15214 6012
rect 15214 5956 15218 6012
rect 15154 5952 15218 5956
rect 15234 6012 15298 6016
rect 15234 5956 15238 6012
rect 15238 5956 15294 6012
rect 15294 5956 15298 6012
rect 15234 5952 15298 5956
rect 15314 6012 15378 6016
rect 15314 5956 15318 6012
rect 15318 5956 15374 6012
rect 15374 5956 15378 6012
rect 15314 5952 15378 5956
rect 15394 6012 15458 6016
rect 15394 5956 15398 6012
rect 15398 5956 15454 6012
rect 15454 5956 15458 6012
rect 15394 5952 15458 5956
rect 20835 6012 20899 6016
rect 20835 5956 20839 6012
rect 20839 5956 20895 6012
rect 20895 5956 20899 6012
rect 20835 5952 20899 5956
rect 20915 6012 20979 6016
rect 20915 5956 20919 6012
rect 20919 5956 20975 6012
rect 20975 5956 20979 6012
rect 20915 5952 20979 5956
rect 20995 6012 21059 6016
rect 20995 5956 20999 6012
rect 20999 5956 21055 6012
rect 21055 5956 21059 6012
rect 20995 5952 21059 5956
rect 21075 6012 21139 6016
rect 21075 5956 21079 6012
rect 21079 5956 21135 6012
rect 21135 5956 21139 6012
rect 21075 5952 21139 5956
rect 9260 5748 9324 5812
rect 20300 5536 20364 5540
rect 20300 5480 20350 5536
rect 20350 5480 20364 5536
rect 20300 5476 20364 5480
rect 6632 5468 6696 5472
rect 6632 5412 6636 5468
rect 6636 5412 6692 5468
rect 6692 5412 6696 5468
rect 6632 5408 6696 5412
rect 6712 5468 6776 5472
rect 6712 5412 6716 5468
rect 6716 5412 6772 5468
rect 6772 5412 6776 5468
rect 6712 5408 6776 5412
rect 6792 5468 6856 5472
rect 6792 5412 6796 5468
rect 6796 5412 6852 5468
rect 6852 5412 6856 5468
rect 6792 5408 6856 5412
rect 6872 5468 6936 5472
rect 6872 5412 6876 5468
rect 6876 5412 6932 5468
rect 6932 5412 6936 5468
rect 6872 5408 6936 5412
rect 12313 5468 12377 5472
rect 12313 5412 12317 5468
rect 12317 5412 12373 5468
rect 12373 5412 12377 5468
rect 12313 5408 12377 5412
rect 12393 5468 12457 5472
rect 12393 5412 12397 5468
rect 12397 5412 12453 5468
rect 12453 5412 12457 5468
rect 12393 5408 12457 5412
rect 12473 5468 12537 5472
rect 12473 5412 12477 5468
rect 12477 5412 12533 5468
rect 12533 5412 12537 5468
rect 12473 5408 12537 5412
rect 12553 5468 12617 5472
rect 12553 5412 12557 5468
rect 12557 5412 12613 5468
rect 12613 5412 12617 5468
rect 12553 5408 12617 5412
rect 17994 5468 18058 5472
rect 17994 5412 17998 5468
rect 17998 5412 18054 5468
rect 18054 5412 18058 5468
rect 17994 5408 18058 5412
rect 18074 5468 18138 5472
rect 18074 5412 18078 5468
rect 18078 5412 18134 5468
rect 18134 5412 18138 5468
rect 18074 5408 18138 5412
rect 18154 5468 18218 5472
rect 18154 5412 18158 5468
rect 18158 5412 18214 5468
rect 18214 5412 18218 5468
rect 18154 5408 18218 5412
rect 18234 5468 18298 5472
rect 18234 5412 18238 5468
rect 18238 5412 18294 5468
rect 18294 5412 18298 5468
rect 18234 5408 18298 5412
rect 23675 5468 23739 5472
rect 23675 5412 23679 5468
rect 23679 5412 23735 5468
rect 23735 5412 23739 5468
rect 23675 5408 23739 5412
rect 23755 5468 23819 5472
rect 23755 5412 23759 5468
rect 23759 5412 23815 5468
rect 23815 5412 23819 5468
rect 23755 5408 23819 5412
rect 23835 5468 23899 5472
rect 23835 5412 23839 5468
rect 23839 5412 23895 5468
rect 23895 5412 23899 5468
rect 23835 5408 23899 5412
rect 23915 5468 23979 5472
rect 23915 5412 23919 5468
rect 23919 5412 23975 5468
rect 23975 5412 23979 5468
rect 23915 5408 23979 5412
rect 3792 4924 3856 4928
rect 3792 4868 3796 4924
rect 3796 4868 3852 4924
rect 3852 4868 3856 4924
rect 3792 4864 3856 4868
rect 3872 4924 3936 4928
rect 3872 4868 3876 4924
rect 3876 4868 3932 4924
rect 3932 4868 3936 4924
rect 3872 4864 3936 4868
rect 3952 4924 4016 4928
rect 3952 4868 3956 4924
rect 3956 4868 4012 4924
rect 4012 4868 4016 4924
rect 3952 4864 4016 4868
rect 4032 4924 4096 4928
rect 4032 4868 4036 4924
rect 4036 4868 4092 4924
rect 4092 4868 4096 4924
rect 4032 4864 4096 4868
rect 9473 4924 9537 4928
rect 9473 4868 9477 4924
rect 9477 4868 9533 4924
rect 9533 4868 9537 4924
rect 9473 4864 9537 4868
rect 9553 4924 9617 4928
rect 9553 4868 9557 4924
rect 9557 4868 9613 4924
rect 9613 4868 9617 4924
rect 9553 4864 9617 4868
rect 9633 4924 9697 4928
rect 9633 4868 9637 4924
rect 9637 4868 9693 4924
rect 9693 4868 9697 4924
rect 9633 4864 9697 4868
rect 9713 4924 9777 4928
rect 9713 4868 9717 4924
rect 9717 4868 9773 4924
rect 9773 4868 9777 4924
rect 9713 4864 9777 4868
rect 15154 4924 15218 4928
rect 15154 4868 15158 4924
rect 15158 4868 15214 4924
rect 15214 4868 15218 4924
rect 15154 4864 15218 4868
rect 15234 4924 15298 4928
rect 15234 4868 15238 4924
rect 15238 4868 15294 4924
rect 15294 4868 15298 4924
rect 15234 4864 15298 4868
rect 15314 4924 15378 4928
rect 15314 4868 15318 4924
rect 15318 4868 15374 4924
rect 15374 4868 15378 4924
rect 15314 4864 15378 4868
rect 15394 4924 15458 4928
rect 15394 4868 15398 4924
rect 15398 4868 15454 4924
rect 15454 4868 15458 4924
rect 15394 4864 15458 4868
rect 20835 4924 20899 4928
rect 20835 4868 20839 4924
rect 20839 4868 20895 4924
rect 20895 4868 20899 4924
rect 20835 4864 20899 4868
rect 20915 4924 20979 4928
rect 20915 4868 20919 4924
rect 20919 4868 20975 4924
rect 20975 4868 20979 4924
rect 20915 4864 20979 4868
rect 20995 4924 21059 4928
rect 20995 4868 20999 4924
rect 20999 4868 21055 4924
rect 21055 4868 21059 4924
rect 20995 4864 21059 4868
rect 21075 4924 21139 4928
rect 21075 4868 21079 4924
rect 21079 4868 21135 4924
rect 21135 4868 21139 4924
rect 21075 4864 21139 4868
rect 8340 4660 8404 4724
rect 6632 4380 6696 4384
rect 6632 4324 6636 4380
rect 6636 4324 6692 4380
rect 6692 4324 6696 4380
rect 6632 4320 6696 4324
rect 6712 4380 6776 4384
rect 6712 4324 6716 4380
rect 6716 4324 6772 4380
rect 6772 4324 6776 4380
rect 6712 4320 6776 4324
rect 6792 4380 6856 4384
rect 6792 4324 6796 4380
rect 6796 4324 6852 4380
rect 6852 4324 6856 4380
rect 6792 4320 6856 4324
rect 6872 4380 6936 4384
rect 6872 4324 6876 4380
rect 6876 4324 6932 4380
rect 6932 4324 6936 4380
rect 6872 4320 6936 4324
rect 12313 4380 12377 4384
rect 12313 4324 12317 4380
rect 12317 4324 12373 4380
rect 12373 4324 12377 4380
rect 12313 4320 12377 4324
rect 12393 4380 12457 4384
rect 12393 4324 12397 4380
rect 12397 4324 12453 4380
rect 12453 4324 12457 4380
rect 12393 4320 12457 4324
rect 12473 4380 12537 4384
rect 12473 4324 12477 4380
rect 12477 4324 12533 4380
rect 12533 4324 12537 4380
rect 12473 4320 12537 4324
rect 12553 4380 12617 4384
rect 12553 4324 12557 4380
rect 12557 4324 12613 4380
rect 12613 4324 12617 4380
rect 12553 4320 12617 4324
rect 17994 4380 18058 4384
rect 17994 4324 17998 4380
rect 17998 4324 18054 4380
rect 18054 4324 18058 4380
rect 17994 4320 18058 4324
rect 18074 4380 18138 4384
rect 18074 4324 18078 4380
rect 18078 4324 18134 4380
rect 18134 4324 18138 4380
rect 18074 4320 18138 4324
rect 18154 4380 18218 4384
rect 18154 4324 18158 4380
rect 18158 4324 18214 4380
rect 18214 4324 18218 4380
rect 18154 4320 18218 4324
rect 18234 4380 18298 4384
rect 18234 4324 18238 4380
rect 18238 4324 18294 4380
rect 18294 4324 18298 4380
rect 18234 4320 18298 4324
rect 23675 4380 23739 4384
rect 23675 4324 23679 4380
rect 23679 4324 23735 4380
rect 23735 4324 23739 4380
rect 23675 4320 23739 4324
rect 23755 4380 23819 4384
rect 23755 4324 23759 4380
rect 23759 4324 23815 4380
rect 23815 4324 23819 4380
rect 23755 4320 23819 4324
rect 23835 4380 23899 4384
rect 23835 4324 23839 4380
rect 23839 4324 23895 4380
rect 23895 4324 23899 4380
rect 23835 4320 23899 4324
rect 23915 4380 23979 4384
rect 23915 4324 23919 4380
rect 23919 4324 23975 4380
rect 23975 4324 23979 4380
rect 23915 4320 23979 4324
rect 3556 3980 3620 4044
rect 8524 3980 8588 4044
rect 3792 3836 3856 3840
rect 3792 3780 3796 3836
rect 3796 3780 3852 3836
rect 3852 3780 3856 3836
rect 3792 3776 3856 3780
rect 3872 3836 3936 3840
rect 3872 3780 3876 3836
rect 3876 3780 3932 3836
rect 3932 3780 3936 3836
rect 3872 3776 3936 3780
rect 3952 3836 4016 3840
rect 3952 3780 3956 3836
rect 3956 3780 4012 3836
rect 4012 3780 4016 3836
rect 3952 3776 4016 3780
rect 4032 3836 4096 3840
rect 4032 3780 4036 3836
rect 4036 3780 4092 3836
rect 4092 3780 4096 3836
rect 4032 3776 4096 3780
rect 9473 3836 9537 3840
rect 9473 3780 9477 3836
rect 9477 3780 9533 3836
rect 9533 3780 9537 3836
rect 9473 3776 9537 3780
rect 9553 3836 9617 3840
rect 9553 3780 9557 3836
rect 9557 3780 9613 3836
rect 9613 3780 9617 3836
rect 9553 3776 9617 3780
rect 9633 3836 9697 3840
rect 9633 3780 9637 3836
rect 9637 3780 9693 3836
rect 9693 3780 9697 3836
rect 9633 3776 9697 3780
rect 9713 3836 9777 3840
rect 9713 3780 9717 3836
rect 9717 3780 9773 3836
rect 9773 3780 9777 3836
rect 9713 3776 9777 3780
rect 15154 3836 15218 3840
rect 15154 3780 15158 3836
rect 15158 3780 15214 3836
rect 15214 3780 15218 3836
rect 15154 3776 15218 3780
rect 15234 3836 15298 3840
rect 15234 3780 15238 3836
rect 15238 3780 15294 3836
rect 15294 3780 15298 3836
rect 15234 3776 15298 3780
rect 15314 3836 15378 3840
rect 15314 3780 15318 3836
rect 15318 3780 15374 3836
rect 15374 3780 15378 3836
rect 15314 3776 15378 3780
rect 15394 3836 15458 3840
rect 15394 3780 15398 3836
rect 15398 3780 15454 3836
rect 15454 3780 15458 3836
rect 15394 3776 15458 3780
rect 20835 3836 20899 3840
rect 20835 3780 20839 3836
rect 20839 3780 20895 3836
rect 20895 3780 20899 3836
rect 20835 3776 20899 3780
rect 20915 3836 20979 3840
rect 20915 3780 20919 3836
rect 20919 3780 20975 3836
rect 20975 3780 20979 3836
rect 20915 3776 20979 3780
rect 20995 3836 21059 3840
rect 20995 3780 20999 3836
rect 20999 3780 21055 3836
rect 21055 3780 21059 3836
rect 20995 3776 21059 3780
rect 21075 3836 21139 3840
rect 21075 3780 21079 3836
rect 21079 3780 21135 3836
rect 21135 3780 21139 3836
rect 21075 3776 21139 3780
rect 4292 3436 4356 3500
rect 7972 3436 8036 3500
rect 6632 3292 6696 3296
rect 6632 3236 6636 3292
rect 6636 3236 6692 3292
rect 6692 3236 6696 3292
rect 6632 3232 6696 3236
rect 6712 3292 6776 3296
rect 6712 3236 6716 3292
rect 6716 3236 6772 3292
rect 6772 3236 6776 3292
rect 6712 3232 6776 3236
rect 6792 3292 6856 3296
rect 6792 3236 6796 3292
rect 6796 3236 6852 3292
rect 6852 3236 6856 3292
rect 6792 3232 6856 3236
rect 6872 3292 6936 3296
rect 6872 3236 6876 3292
rect 6876 3236 6932 3292
rect 6932 3236 6936 3292
rect 6872 3232 6936 3236
rect 12313 3292 12377 3296
rect 12313 3236 12317 3292
rect 12317 3236 12373 3292
rect 12373 3236 12377 3292
rect 12313 3232 12377 3236
rect 12393 3292 12457 3296
rect 12393 3236 12397 3292
rect 12397 3236 12453 3292
rect 12453 3236 12457 3292
rect 12393 3232 12457 3236
rect 12473 3292 12537 3296
rect 12473 3236 12477 3292
rect 12477 3236 12533 3292
rect 12533 3236 12537 3292
rect 12473 3232 12537 3236
rect 12553 3292 12617 3296
rect 12553 3236 12557 3292
rect 12557 3236 12613 3292
rect 12613 3236 12617 3292
rect 12553 3232 12617 3236
rect 17994 3292 18058 3296
rect 17994 3236 17998 3292
rect 17998 3236 18054 3292
rect 18054 3236 18058 3292
rect 17994 3232 18058 3236
rect 18074 3292 18138 3296
rect 18074 3236 18078 3292
rect 18078 3236 18134 3292
rect 18134 3236 18138 3292
rect 18074 3232 18138 3236
rect 18154 3292 18218 3296
rect 18154 3236 18158 3292
rect 18158 3236 18214 3292
rect 18214 3236 18218 3292
rect 18154 3232 18218 3236
rect 18234 3292 18298 3296
rect 18234 3236 18238 3292
rect 18238 3236 18294 3292
rect 18294 3236 18298 3292
rect 18234 3232 18298 3236
rect 23675 3292 23739 3296
rect 23675 3236 23679 3292
rect 23679 3236 23735 3292
rect 23735 3236 23739 3292
rect 23675 3232 23739 3236
rect 23755 3292 23819 3296
rect 23755 3236 23759 3292
rect 23759 3236 23815 3292
rect 23815 3236 23819 3292
rect 23755 3232 23819 3236
rect 23835 3292 23899 3296
rect 23835 3236 23839 3292
rect 23839 3236 23895 3292
rect 23895 3236 23899 3292
rect 23835 3232 23899 3236
rect 23915 3292 23979 3296
rect 23915 3236 23919 3292
rect 23919 3236 23975 3292
rect 23975 3236 23979 3292
rect 23915 3232 23979 3236
rect 3792 2748 3856 2752
rect 3792 2692 3796 2748
rect 3796 2692 3852 2748
rect 3852 2692 3856 2748
rect 3792 2688 3856 2692
rect 3872 2748 3936 2752
rect 3872 2692 3876 2748
rect 3876 2692 3932 2748
rect 3932 2692 3936 2748
rect 3872 2688 3936 2692
rect 3952 2748 4016 2752
rect 3952 2692 3956 2748
rect 3956 2692 4012 2748
rect 4012 2692 4016 2748
rect 3952 2688 4016 2692
rect 4032 2748 4096 2752
rect 4032 2692 4036 2748
rect 4036 2692 4092 2748
rect 4092 2692 4096 2748
rect 4032 2688 4096 2692
rect 9473 2748 9537 2752
rect 9473 2692 9477 2748
rect 9477 2692 9533 2748
rect 9533 2692 9537 2748
rect 9473 2688 9537 2692
rect 9553 2748 9617 2752
rect 9553 2692 9557 2748
rect 9557 2692 9613 2748
rect 9613 2692 9617 2748
rect 9553 2688 9617 2692
rect 9633 2748 9697 2752
rect 9633 2692 9637 2748
rect 9637 2692 9693 2748
rect 9693 2692 9697 2748
rect 9633 2688 9697 2692
rect 9713 2748 9777 2752
rect 9713 2692 9717 2748
rect 9717 2692 9773 2748
rect 9773 2692 9777 2748
rect 9713 2688 9777 2692
rect 15154 2748 15218 2752
rect 15154 2692 15158 2748
rect 15158 2692 15214 2748
rect 15214 2692 15218 2748
rect 15154 2688 15218 2692
rect 15234 2748 15298 2752
rect 15234 2692 15238 2748
rect 15238 2692 15294 2748
rect 15294 2692 15298 2748
rect 15234 2688 15298 2692
rect 15314 2748 15378 2752
rect 15314 2692 15318 2748
rect 15318 2692 15374 2748
rect 15374 2692 15378 2748
rect 15314 2688 15378 2692
rect 15394 2748 15458 2752
rect 15394 2692 15398 2748
rect 15398 2692 15454 2748
rect 15454 2692 15458 2748
rect 15394 2688 15458 2692
rect 20835 2748 20899 2752
rect 20835 2692 20839 2748
rect 20839 2692 20895 2748
rect 20895 2692 20899 2748
rect 20835 2688 20899 2692
rect 20915 2748 20979 2752
rect 20915 2692 20919 2748
rect 20919 2692 20975 2748
rect 20975 2692 20979 2748
rect 20915 2688 20979 2692
rect 20995 2748 21059 2752
rect 20995 2692 20999 2748
rect 20999 2692 21055 2748
rect 21055 2692 21059 2748
rect 20995 2688 21059 2692
rect 21075 2748 21139 2752
rect 21075 2692 21079 2748
rect 21079 2692 21135 2748
rect 21135 2692 21139 2748
rect 21075 2688 21139 2692
rect 5028 2680 5092 2684
rect 5028 2624 5078 2680
rect 5078 2624 5092 2680
rect 5028 2620 5092 2624
rect 7788 2680 7852 2684
rect 7788 2624 7838 2680
rect 7838 2624 7852 2680
rect 7788 2620 7852 2624
rect 8524 2484 8588 2548
rect 8156 2408 8220 2412
rect 8156 2352 8206 2408
rect 8206 2352 8220 2408
rect 8156 2348 8220 2352
rect 6632 2204 6696 2208
rect 6632 2148 6636 2204
rect 6636 2148 6692 2204
rect 6692 2148 6696 2204
rect 6632 2144 6696 2148
rect 6712 2204 6776 2208
rect 6712 2148 6716 2204
rect 6716 2148 6772 2204
rect 6772 2148 6776 2204
rect 6712 2144 6776 2148
rect 6792 2204 6856 2208
rect 6792 2148 6796 2204
rect 6796 2148 6852 2204
rect 6852 2148 6856 2204
rect 6792 2144 6856 2148
rect 6872 2204 6936 2208
rect 6872 2148 6876 2204
rect 6876 2148 6932 2204
rect 6932 2148 6936 2204
rect 6872 2144 6936 2148
rect 12313 2204 12377 2208
rect 12313 2148 12317 2204
rect 12317 2148 12373 2204
rect 12373 2148 12377 2204
rect 12313 2144 12377 2148
rect 12393 2204 12457 2208
rect 12393 2148 12397 2204
rect 12397 2148 12453 2204
rect 12453 2148 12457 2204
rect 12393 2144 12457 2148
rect 12473 2204 12537 2208
rect 12473 2148 12477 2204
rect 12477 2148 12533 2204
rect 12533 2148 12537 2204
rect 12473 2144 12537 2148
rect 12553 2204 12617 2208
rect 12553 2148 12557 2204
rect 12557 2148 12613 2204
rect 12613 2148 12617 2204
rect 12553 2144 12617 2148
rect 17994 2204 18058 2208
rect 17994 2148 17998 2204
rect 17998 2148 18054 2204
rect 18054 2148 18058 2204
rect 17994 2144 18058 2148
rect 18074 2204 18138 2208
rect 18074 2148 18078 2204
rect 18078 2148 18134 2204
rect 18134 2148 18138 2204
rect 18074 2144 18138 2148
rect 18154 2204 18218 2208
rect 18154 2148 18158 2204
rect 18158 2148 18214 2204
rect 18214 2148 18218 2204
rect 18154 2144 18218 2148
rect 18234 2204 18298 2208
rect 18234 2148 18238 2204
rect 18238 2148 18294 2204
rect 18294 2148 18298 2204
rect 18234 2144 18298 2148
rect 23675 2204 23739 2208
rect 23675 2148 23679 2204
rect 23679 2148 23735 2204
rect 23735 2148 23739 2204
rect 23675 2144 23739 2148
rect 23755 2204 23819 2208
rect 23755 2148 23759 2204
rect 23759 2148 23815 2204
rect 23815 2148 23819 2204
rect 23755 2144 23819 2148
rect 23835 2204 23899 2208
rect 23835 2148 23839 2204
rect 23839 2148 23895 2204
rect 23895 2148 23899 2204
rect 23835 2144 23899 2148
rect 23915 2204 23979 2208
rect 23915 2148 23919 2204
rect 23919 2148 23975 2204
rect 23975 2148 23979 2204
rect 23915 2144 23979 2148
rect 7972 1940 8036 2004
<< metal4 >>
rect 3784 22336 4104 22352
rect 3784 22272 3792 22336
rect 3856 22272 3872 22336
rect 3936 22272 3952 22336
rect 4016 22272 4032 22336
rect 4096 22272 4104 22336
rect 3784 21248 4104 22272
rect 3784 21184 3792 21248
rect 3856 21184 3872 21248
rect 3936 21184 3952 21248
rect 4016 21184 4032 21248
rect 4096 21184 4104 21248
rect 3784 20160 4104 21184
rect 6624 21792 6944 22352
rect 6624 21728 6632 21792
rect 6696 21728 6712 21792
rect 6776 21728 6792 21792
rect 6856 21728 6872 21792
rect 6936 21728 6944 21792
rect 4291 20772 4357 20773
rect 4291 20708 4292 20772
rect 4356 20708 4357 20772
rect 4291 20707 4357 20708
rect 3784 20096 3792 20160
rect 3856 20096 3872 20160
rect 3936 20096 3952 20160
rect 4016 20096 4032 20160
rect 4096 20096 4104 20160
rect 3555 19412 3621 19413
rect 3555 19348 3556 19412
rect 3620 19348 3621 19412
rect 3555 19347 3621 19348
rect 3371 16692 3437 16693
rect 3371 16628 3372 16692
rect 3436 16628 3437 16692
rect 3371 16627 3437 16628
rect 3374 7445 3434 16627
rect 3371 7444 3437 7445
rect 3371 7380 3372 7444
rect 3436 7380 3437 7444
rect 3371 7379 3437 7380
rect 3558 4045 3618 19347
rect 3784 19072 4104 20096
rect 3784 19008 3792 19072
rect 3856 19008 3872 19072
rect 3936 19008 3952 19072
rect 4016 19008 4032 19072
rect 4096 19008 4104 19072
rect 3784 17984 4104 19008
rect 3784 17920 3792 17984
rect 3856 17920 3872 17984
rect 3936 17920 3952 17984
rect 4016 17920 4032 17984
rect 4096 17920 4104 17984
rect 3784 16896 4104 17920
rect 3784 16832 3792 16896
rect 3856 16832 3872 16896
rect 3936 16832 3952 16896
rect 4016 16832 4032 16896
rect 4096 16832 4104 16896
rect 3784 15808 4104 16832
rect 3784 15744 3792 15808
rect 3856 15744 3872 15808
rect 3936 15744 3952 15808
rect 4016 15744 4032 15808
rect 4096 15744 4104 15808
rect 3784 14720 4104 15744
rect 3784 14656 3792 14720
rect 3856 14656 3872 14720
rect 3936 14656 3952 14720
rect 4016 14656 4032 14720
rect 4096 14656 4104 14720
rect 3784 13632 4104 14656
rect 3784 13568 3792 13632
rect 3856 13568 3872 13632
rect 3936 13568 3952 13632
rect 4016 13568 4032 13632
rect 4096 13568 4104 13632
rect 3784 12544 4104 13568
rect 3784 12480 3792 12544
rect 3856 12480 3872 12544
rect 3936 12480 3952 12544
rect 4016 12480 4032 12544
rect 4096 12480 4104 12544
rect 3784 11456 4104 12480
rect 4294 12341 4354 20707
rect 6624 20704 6944 21728
rect 9465 22336 9785 22352
rect 9465 22272 9473 22336
rect 9537 22272 9553 22336
rect 9617 22272 9633 22336
rect 9697 22272 9713 22336
rect 9777 22272 9785 22336
rect 9465 21248 9785 22272
rect 9465 21184 9473 21248
rect 9537 21184 9553 21248
rect 9617 21184 9633 21248
rect 9697 21184 9713 21248
rect 9777 21184 9785 21248
rect 7603 20772 7669 20773
rect 7603 20708 7604 20772
rect 7668 20708 7669 20772
rect 7603 20707 7669 20708
rect 6624 20640 6632 20704
rect 6696 20640 6712 20704
rect 6776 20640 6792 20704
rect 6856 20640 6872 20704
rect 6936 20640 6944 20704
rect 6624 19616 6944 20640
rect 6624 19552 6632 19616
rect 6696 19552 6712 19616
rect 6776 19552 6792 19616
rect 6856 19552 6872 19616
rect 6936 19552 6944 19616
rect 6315 19412 6381 19413
rect 6315 19348 6316 19412
rect 6380 19348 6381 19412
rect 6315 19347 6381 19348
rect 5027 12612 5093 12613
rect 5027 12548 5028 12612
rect 5092 12548 5093 12612
rect 5027 12547 5093 12548
rect 4291 12340 4357 12341
rect 4291 12276 4292 12340
rect 4356 12276 4357 12340
rect 4291 12275 4357 12276
rect 4294 11933 4354 12275
rect 4291 11932 4357 11933
rect 4291 11868 4292 11932
rect 4356 11868 4357 11932
rect 4291 11867 4357 11868
rect 3784 11392 3792 11456
rect 3856 11392 3872 11456
rect 3936 11392 3952 11456
rect 4016 11392 4032 11456
rect 4096 11392 4104 11456
rect 3784 10368 4104 11392
rect 3784 10304 3792 10368
rect 3856 10304 3872 10368
rect 3936 10304 3952 10368
rect 4016 10304 4032 10368
rect 4096 10304 4104 10368
rect 3784 9280 4104 10304
rect 3784 9216 3792 9280
rect 3856 9216 3872 9280
rect 3936 9216 3952 9280
rect 4016 9216 4032 9280
rect 4096 9216 4104 9280
rect 3784 8192 4104 9216
rect 3784 8128 3792 8192
rect 3856 8128 3872 8192
rect 3936 8128 3952 8192
rect 4016 8128 4032 8192
rect 4096 8128 4104 8192
rect 3784 7104 4104 8128
rect 3784 7040 3792 7104
rect 3856 7040 3872 7104
rect 3936 7040 3952 7104
rect 4016 7040 4032 7104
rect 4096 7040 4104 7104
rect 3784 6016 4104 7040
rect 3784 5952 3792 6016
rect 3856 5952 3872 6016
rect 3936 5952 3952 6016
rect 4016 5952 4032 6016
rect 4096 5952 4104 6016
rect 3784 4928 4104 5952
rect 3784 4864 3792 4928
rect 3856 4864 3872 4928
rect 3936 4864 3952 4928
rect 4016 4864 4032 4928
rect 4096 4864 4104 4928
rect 3555 4044 3621 4045
rect 3555 3980 3556 4044
rect 3620 3980 3621 4044
rect 3555 3979 3621 3980
rect 3784 3840 4104 4864
rect 3784 3776 3792 3840
rect 3856 3776 3872 3840
rect 3936 3776 3952 3840
rect 4016 3776 4032 3840
rect 4096 3776 4104 3840
rect 3784 2752 4104 3776
rect 4294 3501 4354 11867
rect 4291 3500 4357 3501
rect 4291 3436 4292 3500
rect 4356 3436 4357 3500
rect 4291 3435 4357 3436
rect 3784 2688 3792 2752
rect 3856 2688 3872 2752
rect 3936 2688 3952 2752
rect 4016 2688 4032 2752
rect 4096 2688 4104 2752
rect 3784 2128 4104 2688
rect 5030 2685 5090 12547
rect 6318 12205 6378 19347
rect 6624 18528 6944 19552
rect 6624 18464 6632 18528
rect 6696 18464 6712 18528
rect 6776 18464 6792 18528
rect 6856 18464 6872 18528
rect 6936 18464 6944 18528
rect 6624 17440 6944 18464
rect 7419 18052 7485 18053
rect 7419 17988 7420 18052
rect 7484 17988 7485 18052
rect 7419 17987 7485 17988
rect 6624 17376 6632 17440
rect 6696 17376 6712 17440
rect 6776 17376 6792 17440
rect 6856 17376 6872 17440
rect 6936 17376 6944 17440
rect 6624 16352 6944 17376
rect 6624 16288 6632 16352
rect 6696 16288 6712 16352
rect 6776 16288 6792 16352
rect 6856 16288 6872 16352
rect 6936 16288 6944 16352
rect 6624 15264 6944 16288
rect 6624 15200 6632 15264
rect 6696 15200 6712 15264
rect 6776 15200 6792 15264
rect 6856 15200 6872 15264
rect 6936 15200 6944 15264
rect 6624 14176 6944 15200
rect 6624 14112 6632 14176
rect 6696 14112 6712 14176
rect 6776 14112 6792 14176
rect 6856 14112 6872 14176
rect 6936 14112 6944 14176
rect 6624 13088 6944 14112
rect 6624 13024 6632 13088
rect 6696 13024 6712 13088
rect 6776 13024 6792 13088
rect 6856 13024 6872 13088
rect 6936 13024 6944 13088
rect 6315 12204 6381 12205
rect 6315 12140 6316 12204
rect 6380 12140 6381 12204
rect 6315 12139 6381 12140
rect 6624 12000 6944 13024
rect 6624 11936 6632 12000
rect 6696 11936 6712 12000
rect 6776 11936 6792 12000
rect 6856 11936 6872 12000
rect 6936 11936 6944 12000
rect 6624 10912 6944 11936
rect 6624 10848 6632 10912
rect 6696 10848 6712 10912
rect 6776 10848 6792 10912
rect 6856 10848 6872 10912
rect 6936 10848 6944 10912
rect 6624 9824 6944 10848
rect 6624 9760 6632 9824
rect 6696 9760 6712 9824
rect 6776 9760 6792 9824
rect 6856 9760 6872 9824
rect 6936 9760 6944 9824
rect 6624 8736 6944 9760
rect 7422 9485 7482 17987
rect 7606 11253 7666 20707
rect 9465 20160 9785 21184
rect 9465 20096 9473 20160
rect 9537 20096 9553 20160
rect 9617 20096 9633 20160
rect 9697 20096 9713 20160
rect 9777 20096 9785 20160
rect 9465 19072 9785 20096
rect 9465 19008 9473 19072
rect 9537 19008 9553 19072
rect 9617 19008 9633 19072
rect 9697 19008 9713 19072
rect 9777 19008 9785 19072
rect 9465 17984 9785 19008
rect 9465 17920 9473 17984
rect 9537 17920 9553 17984
rect 9617 17920 9633 17984
rect 9697 17920 9713 17984
rect 9777 17920 9785 17984
rect 9465 16896 9785 17920
rect 9465 16832 9473 16896
rect 9537 16832 9553 16896
rect 9617 16832 9633 16896
rect 9697 16832 9713 16896
rect 9777 16832 9785 16896
rect 9465 15808 9785 16832
rect 9465 15744 9473 15808
rect 9537 15744 9553 15808
rect 9617 15744 9633 15808
rect 9697 15744 9713 15808
rect 9777 15744 9785 15808
rect 9465 14720 9785 15744
rect 9465 14656 9473 14720
rect 9537 14656 9553 14720
rect 9617 14656 9633 14720
rect 9697 14656 9713 14720
rect 9777 14656 9785 14720
rect 9465 13632 9785 14656
rect 9465 13568 9473 13632
rect 9537 13568 9553 13632
rect 9617 13568 9633 13632
rect 9697 13568 9713 13632
rect 9777 13568 9785 13632
rect 9465 12544 9785 13568
rect 9465 12480 9473 12544
rect 9537 12480 9553 12544
rect 9617 12480 9633 12544
rect 9697 12480 9713 12544
rect 9777 12480 9785 12544
rect 8523 12068 8589 12069
rect 8523 12004 8524 12068
rect 8588 12004 8589 12068
rect 8523 12003 8589 12004
rect 8155 11932 8221 11933
rect 8155 11868 8156 11932
rect 8220 11868 8221 11932
rect 8155 11867 8221 11868
rect 7603 11252 7669 11253
rect 7603 11188 7604 11252
rect 7668 11188 7669 11252
rect 7603 11187 7669 11188
rect 7419 9484 7485 9485
rect 7419 9420 7420 9484
rect 7484 9420 7485 9484
rect 7419 9419 7485 9420
rect 7971 9348 8037 9349
rect 7971 9284 7972 9348
rect 8036 9284 8037 9348
rect 7971 9283 8037 9284
rect 6624 8672 6632 8736
rect 6696 8672 6712 8736
rect 6776 8672 6792 8736
rect 6856 8672 6872 8736
rect 6936 8672 6944 8736
rect 6624 7648 6944 8672
rect 7787 8396 7853 8397
rect 7787 8332 7788 8396
rect 7852 8332 7853 8396
rect 7787 8331 7853 8332
rect 6624 7584 6632 7648
rect 6696 7584 6712 7648
rect 6776 7584 6792 7648
rect 6856 7584 6872 7648
rect 6936 7584 6944 7648
rect 6624 6560 6944 7584
rect 6624 6496 6632 6560
rect 6696 6496 6712 6560
rect 6776 6496 6792 6560
rect 6856 6496 6872 6560
rect 6936 6496 6944 6560
rect 6624 5472 6944 6496
rect 6624 5408 6632 5472
rect 6696 5408 6712 5472
rect 6776 5408 6792 5472
rect 6856 5408 6872 5472
rect 6936 5408 6944 5472
rect 6624 4384 6944 5408
rect 6624 4320 6632 4384
rect 6696 4320 6712 4384
rect 6776 4320 6792 4384
rect 6856 4320 6872 4384
rect 6936 4320 6944 4384
rect 6624 3296 6944 4320
rect 6624 3232 6632 3296
rect 6696 3232 6712 3296
rect 6776 3232 6792 3296
rect 6856 3232 6872 3296
rect 6936 3232 6944 3296
rect 5027 2684 5093 2685
rect 5027 2620 5028 2684
rect 5092 2620 5093 2684
rect 5027 2619 5093 2620
rect 6624 2208 6944 3232
rect 7790 2685 7850 8331
rect 7974 3501 8034 9283
rect 7971 3500 8037 3501
rect 7971 3436 7972 3500
rect 8036 3436 8037 3500
rect 7971 3435 8037 3436
rect 7787 2684 7853 2685
rect 7787 2620 7788 2684
rect 7852 2620 7853 2684
rect 7787 2619 7853 2620
rect 6624 2144 6632 2208
rect 6696 2144 6712 2208
rect 6776 2144 6792 2208
rect 6856 2144 6872 2208
rect 6936 2144 6944 2208
rect 6624 2128 6944 2144
rect 7974 2005 8034 3435
rect 8158 2413 8218 11867
rect 8339 9756 8405 9757
rect 8339 9692 8340 9756
rect 8404 9692 8405 9756
rect 8339 9691 8405 9692
rect 8342 4725 8402 9691
rect 8339 4724 8405 4725
rect 8339 4660 8340 4724
rect 8404 4660 8405 4724
rect 8339 4659 8405 4660
rect 8526 4045 8586 12003
rect 9465 11456 9785 12480
rect 9465 11392 9473 11456
rect 9537 11392 9553 11456
rect 9617 11392 9633 11456
rect 9697 11392 9713 11456
rect 9777 11392 9785 11456
rect 9465 10368 9785 11392
rect 9465 10304 9473 10368
rect 9537 10304 9553 10368
rect 9617 10304 9633 10368
rect 9697 10304 9713 10368
rect 9777 10304 9785 10368
rect 9259 9756 9325 9757
rect 9259 9692 9260 9756
rect 9324 9692 9325 9756
rect 9259 9691 9325 9692
rect 9262 5813 9322 9691
rect 9465 9280 9785 10304
rect 12305 21792 12625 22352
rect 12305 21728 12313 21792
rect 12377 21728 12393 21792
rect 12457 21728 12473 21792
rect 12537 21728 12553 21792
rect 12617 21728 12625 21792
rect 12305 20704 12625 21728
rect 12305 20640 12313 20704
rect 12377 20640 12393 20704
rect 12457 20640 12473 20704
rect 12537 20640 12553 20704
rect 12617 20640 12625 20704
rect 12305 19616 12625 20640
rect 12305 19552 12313 19616
rect 12377 19552 12393 19616
rect 12457 19552 12473 19616
rect 12537 19552 12553 19616
rect 12617 19552 12625 19616
rect 12305 18528 12625 19552
rect 12305 18464 12313 18528
rect 12377 18464 12393 18528
rect 12457 18464 12473 18528
rect 12537 18464 12553 18528
rect 12617 18464 12625 18528
rect 12305 17440 12625 18464
rect 12305 17376 12313 17440
rect 12377 17376 12393 17440
rect 12457 17376 12473 17440
rect 12537 17376 12553 17440
rect 12617 17376 12625 17440
rect 12305 16352 12625 17376
rect 12305 16288 12313 16352
rect 12377 16288 12393 16352
rect 12457 16288 12473 16352
rect 12537 16288 12553 16352
rect 12617 16288 12625 16352
rect 12305 15264 12625 16288
rect 12305 15200 12313 15264
rect 12377 15200 12393 15264
rect 12457 15200 12473 15264
rect 12537 15200 12553 15264
rect 12617 15200 12625 15264
rect 12305 14176 12625 15200
rect 12305 14112 12313 14176
rect 12377 14112 12393 14176
rect 12457 14112 12473 14176
rect 12537 14112 12553 14176
rect 12617 14112 12625 14176
rect 12305 13088 12625 14112
rect 12305 13024 12313 13088
rect 12377 13024 12393 13088
rect 12457 13024 12473 13088
rect 12537 13024 12553 13088
rect 12617 13024 12625 13088
rect 12305 12000 12625 13024
rect 15146 22336 15466 22352
rect 15146 22272 15154 22336
rect 15218 22272 15234 22336
rect 15298 22272 15314 22336
rect 15378 22272 15394 22336
rect 15458 22272 15466 22336
rect 15146 21248 15466 22272
rect 15146 21184 15154 21248
rect 15218 21184 15234 21248
rect 15298 21184 15314 21248
rect 15378 21184 15394 21248
rect 15458 21184 15466 21248
rect 15146 20160 15466 21184
rect 15146 20096 15154 20160
rect 15218 20096 15234 20160
rect 15298 20096 15314 20160
rect 15378 20096 15394 20160
rect 15458 20096 15466 20160
rect 15146 19072 15466 20096
rect 15146 19008 15154 19072
rect 15218 19008 15234 19072
rect 15298 19008 15314 19072
rect 15378 19008 15394 19072
rect 15458 19008 15466 19072
rect 15146 17984 15466 19008
rect 15146 17920 15154 17984
rect 15218 17920 15234 17984
rect 15298 17920 15314 17984
rect 15378 17920 15394 17984
rect 15458 17920 15466 17984
rect 15146 16896 15466 17920
rect 15146 16832 15154 16896
rect 15218 16832 15234 16896
rect 15298 16832 15314 16896
rect 15378 16832 15394 16896
rect 15458 16832 15466 16896
rect 15146 15808 15466 16832
rect 15146 15744 15154 15808
rect 15218 15744 15234 15808
rect 15298 15744 15314 15808
rect 15378 15744 15394 15808
rect 15458 15744 15466 15808
rect 15146 14720 15466 15744
rect 17986 21792 18306 22352
rect 17986 21728 17994 21792
rect 18058 21728 18074 21792
rect 18138 21728 18154 21792
rect 18218 21728 18234 21792
rect 18298 21728 18306 21792
rect 17986 20704 18306 21728
rect 17986 20640 17994 20704
rect 18058 20640 18074 20704
rect 18138 20640 18154 20704
rect 18218 20640 18234 20704
rect 18298 20640 18306 20704
rect 17986 19616 18306 20640
rect 17986 19552 17994 19616
rect 18058 19552 18074 19616
rect 18138 19552 18154 19616
rect 18218 19552 18234 19616
rect 18298 19552 18306 19616
rect 17986 18528 18306 19552
rect 17986 18464 17994 18528
rect 18058 18464 18074 18528
rect 18138 18464 18154 18528
rect 18218 18464 18234 18528
rect 18298 18464 18306 18528
rect 17986 17440 18306 18464
rect 17986 17376 17994 17440
rect 18058 17376 18074 17440
rect 18138 17376 18154 17440
rect 18218 17376 18234 17440
rect 18298 17376 18306 17440
rect 17986 16352 18306 17376
rect 17986 16288 17994 16352
rect 18058 16288 18074 16352
rect 18138 16288 18154 16352
rect 18218 16288 18234 16352
rect 18298 16288 18306 16352
rect 17986 15264 18306 16288
rect 17986 15200 17994 15264
rect 18058 15200 18074 15264
rect 18138 15200 18154 15264
rect 18218 15200 18234 15264
rect 18298 15200 18306 15264
rect 16435 15060 16501 15061
rect 16435 14996 16436 15060
rect 16500 14996 16501 15060
rect 16435 14995 16501 14996
rect 15146 14656 15154 14720
rect 15218 14656 15234 14720
rect 15298 14656 15314 14720
rect 15378 14656 15394 14720
rect 15458 14656 15466 14720
rect 15146 13632 15466 14656
rect 15699 13836 15765 13837
rect 15699 13772 15700 13836
rect 15764 13772 15765 13836
rect 15699 13771 15765 13772
rect 15146 13568 15154 13632
rect 15218 13568 15234 13632
rect 15298 13568 15314 13632
rect 15378 13568 15394 13632
rect 15458 13568 15466 13632
rect 15146 12544 15466 13568
rect 15146 12480 15154 12544
rect 15218 12480 15234 12544
rect 15298 12480 15314 12544
rect 15378 12480 15394 12544
rect 15458 12480 15466 12544
rect 12939 12204 13005 12205
rect 12939 12140 12940 12204
rect 13004 12140 13005 12204
rect 12939 12139 13005 12140
rect 12305 11936 12313 12000
rect 12377 11936 12393 12000
rect 12457 11936 12473 12000
rect 12537 11936 12553 12000
rect 12617 11936 12625 12000
rect 12305 10912 12625 11936
rect 12305 10848 12313 10912
rect 12377 10848 12393 10912
rect 12457 10848 12473 10912
rect 12537 10848 12553 10912
rect 12617 10848 12625 10912
rect 12305 9824 12625 10848
rect 12942 9893 13002 12139
rect 15146 11456 15466 12480
rect 15146 11392 15154 11456
rect 15218 11392 15234 11456
rect 15298 11392 15314 11456
rect 15378 11392 15394 11456
rect 15458 11392 15466 11456
rect 15146 10368 15466 11392
rect 15146 10304 15154 10368
rect 15218 10304 15234 10368
rect 15298 10304 15314 10368
rect 15378 10304 15394 10368
rect 15458 10304 15466 10368
rect 12939 9892 13005 9893
rect 12939 9828 12940 9892
rect 13004 9828 13005 9892
rect 12939 9827 13005 9828
rect 12305 9760 12313 9824
rect 12377 9760 12393 9824
rect 12457 9760 12473 9824
rect 12537 9760 12553 9824
rect 12617 9760 12625 9824
rect 10915 9756 10981 9757
rect 10915 9692 10916 9756
rect 10980 9692 10981 9756
rect 10915 9691 10981 9692
rect 9465 9216 9473 9280
rect 9537 9216 9553 9280
rect 9617 9216 9633 9280
rect 9697 9216 9713 9280
rect 9777 9216 9785 9280
rect 9465 8192 9785 9216
rect 9465 8128 9473 8192
rect 9537 8128 9553 8192
rect 9617 8128 9633 8192
rect 9697 8128 9713 8192
rect 9777 8128 9785 8192
rect 9465 7104 9785 8128
rect 10918 7989 10978 9691
rect 12305 8736 12625 9760
rect 12305 8672 12313 8736
rect 12377 8672 12393 8736
rect 12457 8672 12473 8736
rect 12537 8672 12553 8736
rect 12617 8672 12625 8736
rect 10915 7988 10981 7989
rect 10915 7924 10916 7988
rect 10980 7924 10981 7988
rect 10915 7923 10981 7924
rect 9465 7040 9473 7104
rect 9537 7040 9553 7104
rect 9617 7040 9633 7104
rect 9697 7040 9713 7104
rect 9777 7040 9785 7104
rect 9465 6016 9785 7040
rect 9465 5952 9473 6016
rect 9537 5952 9553 6016
rect 9617 5952 9633 6016
rect 9697 5952 9713 6016
rect 9777 5952 9785 6016
rect 9259 5812 9325 5813
rect 9259 5748 9260 5812
rect 9324 5748 9325 5812
rect 9259 5747 9325 5748
rect 9465 4928 9785 5952
rect 9465 4864 9473 4928
rect 9537 4864 9553 4928
rect 9617 4864 9633 4928
rect 9697 4864 9713 4928
rect 9777 4864 9785 4928
rect 8523 4044 8589 4045
rect 8523 3980 8524 4044
rect 8588 3980 8589 4044
rect 8523 3979 8589 3980
rect 8526 2549 8586 3979
rect 9465 3840 9785 4864
rect 9465 3776 9473 3840
rect 9537 3776 9553 3840
rect 9617 3776 9633 3840
rect 9697 3776 9713 3840
rect 9777 3776 9785 3840
rect 9465 2752 9785 3776
rect 9465 2688 9473 2752
rect 9537 2688 9553 2752
rect 9617 2688 9633 2752
rect 9697 2688 9713 2752
rect 9777 2688 9785 2752
rect 8523 2548 8589 2549
rect 8523 2484 8524 2548
rect 8588 2484 8589 2548
rect 8523 2483 8589 2484
rect 8155 2412 8221 2413
rect 8155 2348 8156 2412
rect 8220 2348 8221 2412
rect 8155 2347 8221 2348
rect 9465 2128 9785 2688
rect 12305 7648 12625 8672
rect 12305 7584 12313 7648
rect 12377 7584 12393 7648
rect 12457 7584 12473 7648
rect 12537 7584 12553 7648
rect 12617 7584 12625 7648
rect 12305 6560 12625 7584
rect 12305 6496 12313 6560
rect 12377 6496 12393 6560
rect 12457 6496 12473 6560
rect 12537 6496 12553 6560
rect 12617 6496 12625 6560
rect 12305 5472 12625 6496
rect 12305 5408 12313 5472
rect 12377 5408 12393 5472
rect 12457 5408 12473 5472
rect 12537 5408 12553 5472
rect 12617 5408 12625 5472
rect 12305 4384 12625 5408
rect 12305 4320 12313 4384
rect 12377 4320 12393 4384
rect 12457 4320 12473 4384
rect 12537 4320 12553 4384
rect 12617 4320 12625 4384
rect 12305 3296 12625 4320
rect 12305 3232 12313 3296
rect 12377 3232 12393 3296
rect 12457 3232 12473 3296
rect 12537 3232 12553 3296
rect 12617 3232 12625 3296
rect 12305 2208 12625 3232
rect 12305 2144 12313 2208
rect 12377 2144 12393 2208
rect 12457 2144 12473 2208
rect 12537 2144 12553 2208
rect 12617 2144 12625 2208
rect 12305 2128 12625 2144
rect 15146 9280 15466 10304
rect 15146 9216 15154 9280
rect 15218 9216 15234 9280
rect 15298 9216 15314 9280
rect 15378 9216 15394 9280
rect 15458 9216 15466 9280
rect 15146 8192 15466 9216
rect 15146 8128 15154 8192
rect 15218 8128 15234 8192
rect 15298 8128 15314 8192
rect 15378 8128 15394 8192
rect 15458 8128 15466 8192
rect 15146 7104 15466 8128
rect 15146 7040 15154 7104
rect 15218 7040 15234 7104
rect 15298 7040 15314 7104
rect 15378 7040 15394 7104
rect 15458 7040 15466 7104
rect 15146 6016 15466 7040
rect 15702 6493 15762 13771
rect 16438 9213 16498 14995
rect 17986 14176 18306 15200
rect 17986 14112 17994 14176
rect 18058 14112 18074 14176
rect 18138 14112 18154 14176
rect 18218 14112 18234 14176
rect 18298 14112 18306 14176
rect 17986 13088 18306 14112
rect 20827 22336 21147 22352
rect 20827 22272 20835 22336
rect 20899 22272 20915 22336
rect 20979 22272 20995 22336
rect 21059 22272 21075 22336
rect 21139 22272 21147 22336
rect 20827 21248 21147 22272
rect 20827 21184 20835 21248
rect 20899 21184 20915 21248
rect 20979 21184 20995 21248
rect 21059 21184 21075 21248
rect 21139 21184 21147 21248
rect 20827 20160 21147 21184
rect 20827 20096 20835 20160
rect 20899 20096 20915 20160
rect 20979 20096 20995 20160
rect 21059 20096 21075 20160
rect 21139 20096 21147 20160
rect 20827 19072 21147 20096
rect 20827 19008 20835 19072
rect 20899 19008 20915 19072
rect 20979 19008 20995 19072
rect 21059 19008 21075 19072
rect 21139 19008 21147 19072
rect 20827 17984 21147 19008
rect 20827 17920 20835 17984
rect 20899 17920 20915 17984
rect 20979 17920 20995 17984
rect 21059 17920 21075 17984
rect 21139 17920 21147 17984
rect 20827 16896 21147 17920
rect 20827 16832 20835 16896
rect 20899 16832 20915 16896
rect 20979 16832 20995 16896
rect 21059 16832 21075 16896
rect 21139 16832 21147 16896
rect 20827 15808 21147 16832
rect 20827 15744 20835 15808
rect 20899 15744 20915 15808
rect 20979 15744 20995 15808
rect 21059 15744 21075 15808
rect 21139 15744 21147 15808
rect 20827 14720 21147 15744
rect 20827 14656 20835 14720
rect 20899 14656 20915 14720
rect 20979 14656 20995 14720
rect 21059 14656 21075 14720
rect 21139 14656 21147 14720
rect 20115 13836 20181 13837
rect 20115 13772 20116 13836
rect 20180 13772 20181 13836
rect 20115 13771 20181 13772
rect 17986 13024 17994 13088
rect 18058 13024 18074 13088
rect 18138 13024 18154 13088
rect 18218 13024 18234 13088
rect 18298 13024 18306 13088
rect 17986 12000 18306 13024
rect 17986 11936 17994 12000
rect 18058 11936 18074 12000
rect 18138 11936 18154 12000
rect 18218 11936 18234 12000
rect 18298 11936 18306 12000
rect 17986 10912 18306 11936
rect 17986 10848 17994 10912
rect 18058 10848 18074 10912
rect 18138 10848 18154 10912
rect 18218 10848 18234 10912
rect 18298 10848 18306 10912
rect 17986 9824 18306 10848
rect 17986 9760 17994 9824
rect 18058 9760 18074 9824
rect 18138 9760 18154 9824
rect 18218 9760 18234 9824
rect 18298 9760 18306 9824
rect 16435 9212 16501 9213
rect 16435 9148 16436 9212
rect 16500 9148 16501 9212
rect 16435 9147 16501 9148
rect 17986 8736 18306 9760
rect 17986 8672 17994 8736
rect 18058 8672 18074 8736
rect 18138 8672 18154 8736
rect 18218 8672 18234 8736
rect 18298 8672 18306 8736
rect 17986 7648 18306 8672
rect 20118 8125 20178 13771
rect 20827 13632 21147 14656
rect 20827 13568 20835 13632
rect 20899 13568 20915 13632
rect 20979 13568 20995 13632
rect 21059 13568 21075 13632
rect 21139 13568 21147 13632
rect 20827 12544 21147 13568
rect 20827 12480 20835 12544
rect 20899 12480 20915 12544
rect 20979 12480 20995 12544
rect 21059 12480 21075 12544
rect 21139 12480 21147 12544
rect 20827 11456 21147 12480
rect 20827 11392 20835 11456
rect 20899 11392 20915 11456
rect 20979 11392 20995 11456
rect 21059 11392 21075 11456
rect 21139 11392 21147 11456
rect 20827 10368 21147 11392
rect 20827 10304 20835 10368
rect 20899 10304 20915 10368
rect 20979 10304 20995 10368
rect 21059 10304 21075 10368
rect 21139 10304 21147 10368
rect 20299 9484 20365 9485
rect 20299 9420 20300 9484
rect 20364 9420 20365 9484
rect 20299 9419 20365 9420
rect 20115 8124 20181 8125
rect 20115 8060 20116 8124
rect 20180 8060 20181 8124
rect 20115 8059 20181 8060
rect 17986 7584 17994 7648
rect 18058 7584 18074 7648
rect 18138 7584 18154 7648
rect 18218 7584 18234 7648
rect 18298 7584 18306 7648
rect 17986 6560 18306 7584
rect 17986 6496 17994 6560
rect 18058 6496 18074 6560
rect 18138 6496 18154 6560
rect 18218 6496 18234 6560
rect 18298 6496 18306 6560
rect 15699 6492 15765 6493
rect 15699 6428 15700 6492
rect 15764 6428 15765 6492
rect 15699 6427 15765 6428
rect 15146 5952 15154 6016
rect 15218 5952 15234 6016
rect 15298 5952 15314 6016
rect 15378 5952 15394 6016
rect 15458 5952 15466 6016
rect 15146 4928 15466 5952
rect 15146 4864 15154 4928
rect 15218 4864 15234 4928
rect 15298 4864 15314 4928
rect 15378 4864 15394 4928
rect 15458 4864 15466 4928
rect 15146 3840 15466 4864
rect 15146 3776 15154 3840
rect 15218 3776 15234 3840
rect 15298 3776 15314 3840
rect 15378 3776 15394 3840
rect 15458 3776 15466 3840
rect 15146 2752 15466 3776
rect 15146 2688 15154 2752
rect 15218 2688 15234 2752
rect 15298 2688 15314 2752
rect 15378 2688 15394 2752
rect 15458 2688 15466 2752
rect 15146 2128 15466 2688
rect 17986 5472 18306 6496
rect 20302 5541 20362 9419
rect 20827 9280 21147 10304
rect 20827 9216 20835 9280
rect 20899 9216 20915 9280
rect 20979 9216 20995 9280
rect 21059 9216 21075 9280
rect 21139 9216 21147 9280
rect 20827 8192 21147 9216
rect 20827 8128 20835 8192
rect 20899 8128 20915 8192
rect 20979 8128 20995 8192
rect 21059 8128 21075 8192
rect 21139 8128 21147 8192
rect 20827 7104 21147 8128
rect 20827 7040 20835 7104
rect 20899 7040 20915 7104
rect 20979 7040 20995 7104
rect 21059 7040 21075 7104
rect 21139 7040 21147 7104
rect 20827 6016 21147 7040
rect 20827 5952 20835 6016
rect 20899 5952 20915 6016
rect 20979 5952 20995 6016
rect 21059 5952 21075 6016
rect 21139 5952 21147 6016
rect 20299 5540 20365 5541
rect 20299 5476 20300 5540
rect 20364 5476 20365 5540
rect 20299 5475 20365 5476
rect 17986 5408 17994 5472
rect 18058 5408 18074 5472
rect 18138 5408 18154 5472
rect 18218 5408 18234 5472
rect 18298 5408 18306 5472
rect 17986 4384 18306 5408
rect 17986 4320 17994 4384
rect 18058 4320 18074 4384
rect 18138 4320 18154 4384
rect 18218 4320 18234 4384
rect 18298 4320 18306 4384
rect 17986 3296 18306 4320
rect 17986 3232 17994 3296
rect 18058 3232 18074 3296
rect 18138 3232 18154 3296
rect 18218 3232 18234 3296
rect 18298 3232 18306 3296
rect 17986 2208 18306 3232
rect 17986 2144 17994 2208
rect 18058 2144 18074 2208
rect 18138 2144 18154 2208
rect 18218 2144 18234 2208
rect 18298 2144 18306 2208
rect 17986 2128 18306 2144
rect 20827 4928 21147 5952
rect 20827 4864 20835 4928
rect 20899 4864 20915 4928
rect 20979 4864 20995 4928
rect 21059 4864 21075 4928
rect 21139 4864 21147 4928
rect 20827 3840 21147 4864
rect 20827 3776 20835 3840
rect 20899 3776 20915 3840
rect 20979 3776 20995 3840
rect 21059 3776 21075 3840
rect 21139 3776 21147 3840
rect 20827 2752 21147 3776
rect 20827 2688 20835 2752
rect 20899 2688 20915 2752
rect 20979 2688 20995 2752
rect 21059 2688 21075 2752
rect 21139 2688 21147 2752
rect 20827 2128 21147 2688
rect 23667 21792 23987 22352
rect 23667 21728 23675 21792
rect 23739 21728 23755 21792
rect 23819 21728 23835 21792
rect 23899 21728 23915 21792
rect 23979 21728 23987 21792
rect 23667 20704 23987 21728
rect 23667 20640 23675 20704
rect 23739 20640 23755 20704
rect 23819 20640 23835 20704
rect 23899 20640 23915 20704
rect 23979 20640 23987 20704
rect 23667 19616 23987 20640
rect 23667 19552 23675 19616
rect 23739 19552 23755 19616
rect 23819 19552 23835 19616
rect 23899 19552 23915 19616
rect 23979 19552 23987 19616
rect 23667 18528 23987 19552
rect 23667 18464 23675 18528
rect 23739 18464 23755 18528
rect 23819 18464 23835 18528
rect 23899 18464 23915 18528
rect 23979 18464 23987 18528
rect 23667 17440 23987 18464
rect 23667 17376 23675 17440
rect 23739 17376 23755 17440
rect 23819 17376 23835 17440
rect 23899 17376 23915 17440
rect 23979 17376 23987 17440
rect 23667 16352 23987 17376
rect 23667 16288 23675 16352
rect 23739 16288 23755 16352
rect 23819 16288 23835 16352
rect 23899 16288 23915 16352
rect 23979 16288 23987 16352
rect 23667 15264 23987 16288
rect 23667 15200 23675 15264
rect 23739 15200 23755 15264
rect 23819 15200 23835 15264
rect 23899 15200 23915 15264
rect 23979 15200 23987 15264
rect 23667 14176 23987 15200
rect 23667 14112 23675 14176
rect 23739 14112 23755 14176
rect 23819 14112 23835 14176
rect 23899 14112 23915 14176
rect 23979 14112 23987 14176
rect 23667 13088 23987 14112
rect 23667 13024 23675 13088
rect 23739 13024 23755 13088
rect 23819 13024 23835 13088
rect 23899 13024 23915 13088
rect 23979 13024 23987 13088
rect 23667 12000 23987 13024
rect 23667 11936 23675 12000
rect 23739 11936 23755 12000
rect 23819 11936 23835 12000
rect 23899 11936 23915 12000
rect 23979 11936 23987 12000
rect 23667 10912 23987 11936
rect 23667 10848 23675 10912
rect 23739 10848 23755 10912
rect 23819 10848 23835 10912
rect 23899 10848 23915 10912
rect 23979 10848 23987 10912
rect 23667 9824 23987 10848
rect 23667 9760 23675 9824
rect 23739 9760 23755 9824
rect 23819 9760 23835 9824
rect 23899 9760 23915 9824
rect 23979 9760 23987 9824
rect 23667 8736 23987 9760
rect 23667 8672 23675 8736
rect 23739 8672 23755 8736
rect 23819 8672 23835 8736
rect 23899 8672 23915 8736
rect 23979 8672 23987 8736
rect 23667 7648 23987 8672
rect 23667 7584 23675 7648
rect 23739 7584 23755 7648
rect 23819 7584 23835 7648
rect 23899 7584 23915 7648
rect 23979 7584 23987 7648
rect 23667 6560 23987 7584
rect 23667 6496 23675 6560
rect 23739 6496 23755 6560
rect 23819 6496 23835 6560
rect 23899 6496 23915 6560
rect 23979 6496 23987 6560
rect 23667 5472 23987 6496
rect 23667 5408 23675 5472
rect 23739 5408 23755 5472
rect 23819 5408 23835 5472
rect 23899 5408 23915 5472
rect 23979 5408 23987 5472
rect 23667 4384 23987 5408
rect 23667 4320 23675 4384
rect 23739 4320 23755 4384
rect 23819 4320 23835 4384
rect 23899 4320 23915 4384
rect 23979 4320 23987 4384
rect 23667 3296 23987 4320
rect 23667 3232 23675 3296
rect 23739 3232 23755 3296
rect 23819 3232 23835 3296
rect 23899 3232 23915 3296
rect 23979 3232 23987 3296
rect 23667 2208 23987 3232
rect 23667 2144 23675 2208
rect 23739 2144 23755 2208
rect 23819 2144 23835 2208
rect 23899 2144 23915 2208
rect 23979 2144 23987 2208
rect 23667 2128 23987 2144
rect 7971 2004 8037 2005
rect 7971 1940 7972 2004
rect 8036 1940 8037 2004
rect 7971 1939 8037 1940
use sky130_fd_sc_hd__diode_2  ANTENNA__407__A2 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 1840 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__411__A
timestamp 1666464484
transform -1 0 1748 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__415__B
timestamp 1666464484
transform -1 0 9016 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__417__A
timestamp 1666464484
transform 1 0 3312 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__419__A
timestamp 1666464484
transform 1 0 10212 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__421__A
timestamp 1666464484
transform -1 0 1748 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__423__B_N
timestamp 1666464484
transform 1 0 1840 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__425__B
timestamp 1666464484
transform 1 0 2116 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__429__B
timestamp 1666464484
transform -1 0 1840 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__433__B
timestamp 1666464484
transform 1 0 2116 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__437__B
timestamp 1666464484
transform 1 0 4048 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__440__C
timestamp 1666464484
transform -1 0 4324 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__445__A
timestamp 1666464484
transform -1 0 1748 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__447__A_N
timestamp 1666464484
transform -1 0 1748 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__454__B1
timestamp 1666464484
transform 1 0 2024 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__457__B1
timestamp 1666464484
transform 1 0 1840 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__464__B1
timestamp 1666464484
transform -1 0 15088 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__466__B1
timestamp 1666464484
transform 1 0 7084 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__470__B1
timestamp 1666464484
transform -1 0 6716 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__473__A
timestamp 1666464484
transform 1 0 14352 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__474__A
timestamp 1666464484
transform -1 0 13984 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__475__A
timestamp 1666464484
transform 1 0 8464 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__481__A
timestamp 1666464484
transform 1 0 7820 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__486__A
timestamp 1666464484
transform 1 0 14260 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__487__A
timestamp 1666464484
transform 1 0 12880 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__493__A
timestamp 1666464484
transform -1 0 17020 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__494__A
timestamp 1666464484
transform 1 0 14904 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__495__A1
timestamp 1666464484
transform 1 0 14260 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__496__B1
timestamp 1666464484
transform 1 0 6624 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__499__B1
timestamp 1666464484
transform 1 0 13432 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__509__A1
timestamp 1666464484
transform 1 0 21344 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__519__A2
timestamp 1666464484
transform 1 0 14812 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__522__A
timestamp 1666464484
transform -1 0 16652 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__530__A
timestamp 1666464484
transform 1 0 13616 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__539__A2
timestamp 1666464484
transform 1 0 21344 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__546__B
timestamp 1666464484
transform -1 0 21528 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__557__A2
timestamp 1666464484
transform 1 0 21160 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__558__B
timestamp 1666464484
transform -1 0 22632 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__565__S
timestamp 1666464484
transform 1 0 17940 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__568__A
timestamp 1666464484
transform 1 0 12788 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__573__B1
timestamp 1666464484
transform 1 0 22356 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__578__A2
timestamp 1666464484
transform 1 0 18768 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__580__C1
timestamp 1666464484
transform 1 0 18584 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__585__A1
timestamp 1666464484
transform 1 0 22908 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__591__C1
timestamp 1666464484
transform -1 0 22172 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__594__A2
timestamp 1666464484
transform 1 0 16008 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__597__A1
timestamp 1666464484
transform 1 0 22172 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__597__C1
timestamp 1666464484
transform -1 0 22908 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__600__B
timestamp 1666464484
transform 1 0 16928 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__601__A2
timestamp 1666464484
transform 1 0 16376 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__602__C1
timestamp 1666464484
transform -1 0 18308 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__604__A1
timestamp 1666464484
transform 1 0 21252 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__605__A2
timestamp 1666464484
transform -1 0 19044 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__607__B
timestamp 1666464484
transform -1 0 16928 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__609__B
timestamp 1666464484
transform -1 0 17296 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__611__A1
timestamp 1666464484
transform -1 0 19596 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__616__A1
timestamp 1666464484
transform -1 0 18860 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__616__C1
timestamp 1666464484
transform -1 0 17756 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__618__A
timestamp 1666464484
transform 1 0 15824 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__621__A2
timestamp 1666464484
transform -1 0 17664 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__622__A1
timestamp 1666464484
transform 1 0 10120 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__624__A1
timestamp 1666464484
transform 1 0 14812 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__625__A1
timestamp 1666464484
transform 1 0 11684 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__626__B1
timestamp 1666464484
transform -1 0 23184 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__627__A1
timestamp 1666464484
transform -1 0 23184 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__627__C1
timestamp 1666464484
transform 1 0 21988 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__629__A
timestamp 1666464484
transform -1 0 22080 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__633__B1
timestamp 1666464484
transform 1 0 10212 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__637__A
timestamp 1666464484
transform 1 0 11224 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__641__A1
timestamp 1666464484
transform 1 0 16836 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__642__D1
timestamp 1666464484
transform 1 0 13892 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__643__A
timestamp 1666464484
transform 1 0 11040 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__644__A1
timestamp 1666464484
transform 1 0 11040 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__646__A1
timestamp 1666464484
transform -1 0 15640 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__648__C1
timestamp 1666464484
transform 1 0 14260 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__651__B1
timestamp 1666464484
transform 1 0 13432 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__653__A1
timestamp 1666464484
transform 1 0 21988 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__659__A1
timestamp 1666464484
transform 1 0 16192 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__664__A1
timestamp 1666464484
transform 1 0 14076 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__670__A1
timestamp 1666464484
transform -1 0 19596 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__674__A1
timestamp 1666464484
transform 1 0 19412 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__675__A1
timestamp 1666464484
transform 1 0 17848 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__678__A1
timestamp 1666464484
transform 1 0 17572 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__679__S
timestamp 1666464484
transform 1 0 16008 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__687__S
timestamp 1666464484
transform 1 0 10212 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__688__A
timestamp 1666464484
transform -1 0 1840 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__701__A
timestamp 1666464484
transform 1 0 8280 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__702__A1
timestamp 1666464484
transform 1 0 8188 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__718__A
timestamp 1666464484
transform 1 0 9568 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__719__B2
timestamp 1666464484
transform 1 0 4048 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__721__S
timestamp 1666464484
transform 1 0 10488 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__734__A1
timestamp 1666464484
transform 1 0 7728 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__736__S
timestamp 1666464484
transform 1 0 11040 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__748__B
timestamp 1666464484
transform 1 0 3312 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__752__B2
timestamp 1666464484
transform 1 0 8464 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__753__A
timestamp 1666464484
transform -1 0 9292 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__760__A1
timestamp 1666464484
transform -1 0 15640 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__769__B2
timestamp 1666464484
transform -1 0 4692 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__774__B1
timestamp 1666464484
transform 1 0 8648 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__781__A
timestamp 1666464484
transform 1 0 5888 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__798__A1
timestamp 1666464484
transform 1 0 4232 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__807__B2
timestamp 1666464484
transform 1 0 7728 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__816__D
timestamp 1666464484
transform 1 0 12236 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__818__D
timestamp 1666464484
transform -1 0 11868 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__819__D
timestamp 1666464484
transform 1 0 12144 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__821__D
timestamp 1666464484
transform 1 0 11684 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__822__D
timestamp 1666464484
transform 1 0 11684 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__827__D
timestamp 1666464484
transform -1 0 9384 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__868__A
timestamp 1666464484
transform -1 0 17480 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_clk_A
timestamp 1666464484
transform -1 0 7268 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1666464484
transform -1 0 15272 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1666464484
transform -1 0 18308 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1666464484
transform -1 0 23276 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1666464484
transform -1 0 7176 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output5_A
timestamp 1666464484
transform -1 0 18032 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output8_A
timestamp 1666464484
transform -1 0 18952 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output9_A
timestamp 1666464484
transform -1 0 17572 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output10_A
timestamp 1666464484
transform -1 0 17020 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output11_A
timestamp 1666464484
transform 1 0 16008 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output12_A
timestamp 1666464484
transform 1 0 16192 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 1380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 1932 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 2300 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18
timestamp 1666464484
transform 1 0 2760 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26
timestamp 1666464484
transform 1 0 3496 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29
timestamp 1666464484
transform 1 0 3772 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35
timestamp 1666464484
transform 1 0 4324 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43
timestamp 1666464484
transform 1 0 5060 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_51
timestamp 1666464484
transform 1 0 5796 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55
timestamp 1666464484
transform 1 0 6164 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57
timestamp 1666464484
transform 1 0 6348 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_63
timestamp 1666464484
transform 1 0 6900 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67
timestamp 1666464484
transform 1 0 7268 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_74
timestamp 1666464484
transform 1 0 7912 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_78
timestamp 1666464484
transform 1 0 8280 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_82
timestamp 1666464484
transform 1 0 8648 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_85
timestamp 1666464484
transform 1 0 8924 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_92 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 9568 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_103
timestamp 1666464484
transform 1 0 10580 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_110
timestamp 1666464484
transform 1 0 11224 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_113
timestamp 1666464484
transform 1 0 11500 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_118 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 11960 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_127
timestamp 1666464484
transform 1 0 12788 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_134
timestamp 1666464484
transform 1 0 13432 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_141
timestamp 1666464484
transform 1 0 14076 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_146
timestamp 1666464484
transform 1 0 14536 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_153
timestamp 1666464484
transform 1 0 15180 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_160
timestamp 1666464484
transform 1 0 15824 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_166
timestamp 1666464484
transform 1 0 16376 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_169
timestamp 1666464484
transform 1 0 16652 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_174
timestamp 1666464484
transform 1 0 17112 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_181
timestamp 1666464484
transform 1 0 17756 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_188
timestamp 1666464484
transform 1 0 18400 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_194
timestamp 1666464484
transform 1 0 18952 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_197
timestamp 1666464484
transform 1 0 19228 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_202
timestamp 1666464484
transform 1 0 19688 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_209
timestamp 1666464484
transform 1 0 20332 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_216
timestamp 1666464484
transform 1 0 20976 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_225
timestamp 1666464484
transform 1 0 21804 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_230
timestamp 1666464484
transform 1 0 22264 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_237
timestamp 1666464484
transform 1 0 22908 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_243
timestamp 1666464484
transform 1 0 23460 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_1_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 1380 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_8
timestamp 1666464484
transform 1 0 1840 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_16
timestamp 1666464484
transform 1 0 2576 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_27
timestamp 1666464484
transform 1 0 3588 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_34
timestamp 1666464484
transform 1 0 4232 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_41
timestamp 1666464484
transform 1 0 4876 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_51
timestamp 1666464484
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1666464484
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_57
timestamp 1666464484
transform 1 0 6348 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_61
timestamp 1666464484
transform 1 0 6716 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_73
timestamp 1666464484
transform 1 0 7820 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_83
timestamp 1666464484
transform 1 0 8740 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_92
timestamp 1666464484
transform 1 0 9568 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_103
timestamp 1666464484
transform 1 0 10580 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_110
timestamp 1666464484
transform 1 0 11224 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_113
timestamp 1666464484
transform 1 0 11500 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_120
timestamp 1666464484
transform 1 0 12144 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_127
timestamp 1666464484
transform 1 0 12788 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_134
timestamp 1666464484
transform 1 0 13432 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_140
timestamp 1666464484
transform 1 0 13984 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_146
timestamp 1666464484
transform 1 0 14536 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_152
timestamp 1666464484
transform 1 0 15088 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_158
timestamp 1666464484
transform 1 0 15640 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_162
timestamp 1666464484
transform 1 0 16008 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_1_169
timestamp 1666464484
transform 1 0 16652 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_173
timestamp 1666464484
transform 1 0 17020 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_179
timestamp 1666464484
transform 1 0 17572 0 -1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_1_190 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 18584 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_202
timestamp 1666464484
transform 1 0 19688 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_214
timestamp 1666464484
transform 1 0 20792 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_218
timestamp 1666464484
transform 1 0 21160 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_1_225
timestamp 1666464484
transform 1 0 21804 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_233
timestamp 1666464484
transform 1 0 22540 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_239
timestamp 1666464484
transform 1 0 23092 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_243
timestamp 1666464484
transform 1 0 23460 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_3
timestamp 1666464484
transform 1 0 1380 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_12
timestamp 1666464484
transform 1 0 2208 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_19
timestamp 1666464484
transform 1 0 2852 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_26
timestamp 1666464484
transform 1 0 3496 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_29
timestamp 1666464484
transform 1 0 3772 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_42
timestamp 1666464484
transform 1 0 4968 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_49
timestamp 1666464484
transform 1 0 5612 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_61
timestamp 1666464484
transform 1 0 6716 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_72
timestamp 1666464484
transform 1 0 7728 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_2_81
timestamp 1666464484
transform 1 0 8556 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_85
timestamp 1666464484
transform 1 0 8924 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_95
timestamp 1666464484
transform 1 0 9844 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_106
timestamp 1666464484
transform 1 0 10856 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_113
timestamp 1666464484
transform 1 0 11500 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_124
timestamp 1666464484
transform 1 0 12512 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_130
timestamp 1666464484
transform 1 0 13064 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_136
timestamp 1666464484
transform 1 0 13616 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_141
timestamp 1666464484
transform 1 0 14076 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_145
timestamp 1666464484
transform 1 0 14444 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_149
timestamp 1666464484
transform 1 0 14812 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_152
timestamp 1666464484
transform 1 0 15088 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_158
timestamp 1666464484
transform 1 0 15640 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_164
timestamp 1666464484
transform 1 0 16192 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_172
timestamp 1666464484
transform 1 0 16928 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_178
timestamp 1666464484
transform 1 0 17480 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_184
timestamp 1666464484
transform 1 0 18032 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_197
timestamp 1666464484
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_209
timestamp 1666464484
transform 1 0 20332 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_221
timestamp 1666464484
transform 1 0 21436 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_233
timestamp 1666464484
transform 1 0 22540 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_2_242
timestamp 1666464484
transform 1 0 23368 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_3
timestamp 1666464484
transform 1 0 1380 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_7
timestamp 1666464484
transform 1 0 1748 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_13
timestamp 1666464484
transform 1 0 2300 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_20
timestamp 1666464484
transform 1 0 2944 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_27
timestamp 1666464484
transform 1 0 3588 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_37
timestamp 1666464484
transform 1 0 4508 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_44
timestamp 1666464484
transform 1 0 5152 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_54
timestamp 1666464484
transform 1 0 6072 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_57
timestamp 1666464484
transform 1 0 6348 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_67
timestamp 1666464484
transform 1 0 7268 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_77
timestamp 1666464484
transform 1 0 8188 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_3_107
timestamp 1666464484
transform 1 0 10948 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1666464484
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_113
timestamp 1666464484
transform 1 0 11500 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_123
timestamp 1666464484
transform 1 0 12420 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_132
timestamp 1666464484
transform 1 0 13248 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_138
timestamp 1666464484
transform 1 0 13800 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_142
timestamp 1666464484
transform 1 0 14168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_145
timestamp 1666464484
transform 1 0 14444 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_151
timestamp 1666464484
transform 1 0 14996 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_155
timestamp 1666464484
transform 1 0 15364 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_159
timestamp 1666464484
transform 1 0 15732 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_162
timestamp 1666464484
transform 1 0 16008 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_169
timestamp 1666464484
transform 1 0 16652 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_173
timestamp 1666464484
transform 1 0 17020 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_176
timestamp 1666464484
transform 1 0 17296 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_188
timestamp 1666464484
transform 1 0 18400 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_192
timestamp 1666464484
transform 1 0 18768 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_195
timestamp 1666464484
transform 1 0 19044 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_207
timestamp 1666464484
transform 1 0 20148 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_219
timestamp 1666464484
transform 1 0 21252 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_223
timestamp 1666464484
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_225
timestamp 1666464484
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_237
timestamp 1666464484
transform 1 0 22908 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_243
timestamp 1666464484
transform 1 0 23460 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_3
timestamp 1666464484
transform 1 0 1380 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_7
timestamp 1666464484
transform 1 0 1748 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_18
timestamp 1666464484
transform 1 0 2760 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_22
timestamp 1666464484
transform 1 0 3128 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_26
timestamp 1666464484
transform 1 0 3496 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_29
timestamp 1666464484
transform 1 0 3772 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_40
timestamp 1666464484
transform 1 0 4784 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_52
timestamp 1666464484
transform 1 0 5888 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_60
timestamp 1666464484
transform 1 0 6624 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_69
timestamp 1666464484
transform 1 0 7452 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_73
timestamp 1666464484
transform 1 0 7820 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_80
timestamp 1666464484
transform 1 0 8464 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_85
timestamp 1666464484
transform 1 0 8924 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_93
timestamp 1666464484
transform 1 0 9660 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_101
timestamp 1666464484
transform 1 0 10396 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_105
timestamp 1666464484
transform 1 0 10764 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_114
timestamp 1666464484
transform 1 0 11592 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_127
timestamp 1666464484
transform 1 0 12788 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_136
timestamp 1666464484
transform 1 0 13616 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_141
timestamp 1666464484
transform 1 0 14076 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_152
timestamp 1666464484
transform 1 0 15088 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_161
timestamp 1666464484
transform 1 0 15916 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_165
timestamp 1666464484
transform 1 0 16284 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_168
timestamp 1666464484
transform 1 0 16560 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_174
timestamp 1666464484
transform 1 0 17112 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_178
timestamp 1666464484
transform 1 0 17480 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_181
timestamp 1666464484
transform 1 0 17756 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_187
timestamp 1666464484
transform 1 0 18308 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_4_193
timestamp 1666464484
transform 1 0 18860 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_197
timestamp 1666464484
transform 1 0 19228 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_201
timestamp 1666464484
transform 1 0 19596 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_213
timestamp 1666464484
transform 1 0 20700 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_225
timestamp 1666464484
transform 1 0 21804 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_237
timestamp 1666464484
transform 1 0 22908 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_243
timestamp 1666464484
transform 1 0 23460 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_3
timestamp 1666464484
transform 1 0 1380 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_17
timestamp 1666464484
transform 1 0 2668 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_28
timestamp 1666464484
transform 1 0 3680 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_34
timestamp 1666464484
transform 1 0 4232 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_45
timestamp 1666464484
transform 1 0 5244 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_52
timestamp 1666464484
transform 1 0 5888 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_5_57
timestamp 1666464484
transform 1 0 6348 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_62
timestamp 1666464484
transform 1 0 6808 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_73
timestamp 1666464484
transform 1 0 7820 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_79
timestamp 1666464484
transform 1 0 8372 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_89
timestamp 1666464484
transform 1 0 9292 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_98
timestamp 1666464484
transform 1 0 10120 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_5_109
timestamp 1666464484
transform 1 0 11132 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_113
timestamp 1666464484
transform 1 0 11500 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_122
timestamp 1666464484
transform 1 0 12328 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_131
timestamp 1666464484
transform 1 0 13156 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_143
timestamp 1666464484
transform 1 0 14260 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_152
timestamp 1666464484
transform 1 0 15088 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_158
timestamp 1666464484
transform 1 0 15640 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_164
timestamp 1666464484
transform 1 0 16192 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_169
timestamp 1666464484
transform 1 0 16652 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_174
timestamp 1666464484
transform 1 0 17112 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_180
timestamp 1666464484
transform 1 0 17664 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_186
timestamp 1666464484
transform 1 0 18216 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_193
timestamp 1666464484
transform 1 0 18860 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_205
timestamp 1666464484
transform 1 0 19964 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_212
timestamp 1666464484
transform 1 0 20608 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_225
timestamp 1666464484
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_237
timestamp 1666464484
transform 1 0 22908 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_243
timestamp 1666464484
transform 1 0 23460 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_3
timestamp 1666464484
transform 1 0 1380 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_6_17
timestamp 1666464484
transform 1 0 2668 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_24
timestamp 1666464484
transform 1 0 3312 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_29
timestamp 1666464484
transform 1 0 3772 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_34
timestamp 1666464484
transform 1 0 4232 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_38
timestamp 1666464484
transform 1 0 4600 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_60
timestamp 1666464484
transform 1 0 6624 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_66
timestamp 1666464484
transform 1 0 7176 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_74
timestamp 1666464484
transform 1 0 7912 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_6_82
timestamp 1666464484
transform 1 0 8648 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_85
timestamp 1666464484
transform 1 0 8924 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_93
timestamp 1666464484
transform 1 0 9660 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_103
timestamp 1666464484
transform 1 0 10580 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_115
timestamp 1666464484
transform 1 0 11684 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_125
timestamp 1666464484
transform 1 0 12604 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_138
timestamp 1666464484
transform 1 0 13800 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_141
timestamp 1666464484
transform 1 0 14076 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_6_149
timestamp 1666464484
transform 1 0 14812 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_155
timestamp 1666464484
transform 1 0 15364 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_163
timestamp 1666464484
transform 1 0 16100 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_170
timestamp 1666464484
transform 1 0 16744 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_6_180
timestamp 1666464484
transform 1 0 17664 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_6_194
timestamp 1666464484
transform 1 0 18952 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_197
timestamp 1666464484
transform 1 0 19228 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_205
timestamp 1666464484
transform 1 0 19964 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_214
timestamp 1666464484
transform 1 0 20792 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_6_220
timestamp 1666464484
transform 1 0 21344 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_232
timestamp 1666464484
transform 1 0 22448 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_3
timestamp 1666464484
transform 1 0 1380 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_12
timestamp 1666464484
transform 1 0 2208 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_24
timestamp 1666464484
transform 1 0 3312 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_38
timestamp 1666464484
transform 1 0 4600 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_50
timestamp 1666464484
transform 1 0 5704 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_7_57
timestamp 1666464484
transform 1 0 6348 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_7_67
timestamp 1666464484
transform 1 0 7268 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_7_75
timestamp 1666464484
transform 1 0 8004 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_87
timestamp 1666464484
transform 1 0 9108 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_97
timestamp 1666464484
transform 1 0 10028 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_7_110
timestamp 1666464484
transform 1 0 11224 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_113
timestamp 1666464484
transform 1 0 11500 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_117
timestamp 1666464484
transform 1 0 11868 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_127
timestamp 1666464484
transform 1 0 12788 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_140
timestamp 1666464484
transform 1 0 13984 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_144
timestamp 1666464484
transform 1 0 14352 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_151
timestamp 1666464484
transform 1 0 14996 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_159
timestamp 1666464484
transform 1 0 15732 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_166
timestamp 1666464484
transform 1 0 16376 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_169
timestamp 1666464484
transform 1 0 16652 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_7_174
timestamp 1666464484
transform 1 0 17112 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_182
timestamp 1666464484
transform 1 0 17848 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_190
timestamp 1666464484
transform 1 0 18584 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_199
timestamp 1666464484
transform 1 0 19412 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_211
timestamp 1666464484
transform 1 0 20516 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_220
timestamp 1666464484
transform 1 0 21344 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_225
timestamp 1666464484
transform 1 0 21804 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_229
timestamp 1666464484
transform 1 0 22172 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_7_241
timestamp 1666464484
transform 1 0 23276 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_8_3
timestamp 1666464484
transform 1 0 1380 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_9
timestamp 1666464484
transform 1 0 1932 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_16
timestamp 1666464484
transform 1 0 2576 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_24
timestamp 1666464484
transform 1 0 3312 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_29
timestamp 1666464484
transform 1 0 3772 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_38
timestamp 1666464484
transform 1 0 4600 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_49
timestamp 1666464484
transform 1 0 5612 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_61
timestamp 1666464484
transform 1 0 6716 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_67
timestamp 1666464484
transform 1 0 7268 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_78
timestamp 1666464484
transform 1 0 8280 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_8_85
timestamp 1666464484
transform 1 0 8924 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_8_94
timestamp 1666464484
transform 1 0 9752 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_8_110
timestamp 1666464484
transform 1 0 11224 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_118
timestamp 1666464484
transform 1 0 11960 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_125
timestamp 1666464484
transform 1 0 12604 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_129
timestamp 1666464484
transform 1 0 12972 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp 1666464484
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1666464484
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_141
timestamp 1666464484
transform 1 0 14076 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_145
timestamp 1666464484
transform 1 0 14444 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_151
timestamp 1666464484
transform 1 0 14996 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_160
timestamp 1666464484
transform 1 0 15824 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_172
timestamp 1666464484
transform 1 0 16928 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_184
timestamp 1666464484
transform 1 0 18032 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_194
timestamp 1666464484
transform 1 0 18952 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_197
timestamp 1666464484
transform 1 0 19228 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_201
timestamp 1666464484
transform 1 0 19596 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_210
timestamp 1666464484
transform 1 0 20424 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_222
timestamp 1666464484
transform 1 0 21528 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_8_230
timestamp 1666464484
transform 1 0 22264 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_8_242
timestamp 1666464484
transform 1 0 23368 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_3
timestamp 1666464484
transform 1 0 1380 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_11
timestamp 1666464484
transform 1 0 2116 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_21
timestamp 1666464484
transform 1 0 3036 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_30
timestamp 1666464484
transform 1 0 3864 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_9_43
timestamp 1666464484
transform 1 0 5060 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_49
timestamp 1666464484
transform 1 0 5612 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_54
timestamp 1666464484
transform 1 0 6072 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_9_57
timestamp 1666464484
transform 1 0 6348 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_63
timestamp 1666464484
transform 1 0 6900 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_80
timestamp 1666464484
transform 1 0 8464 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_90
timestamp 1666464484
transform 1 0 9384 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_100
timestamp 1666464484
transform 1 0 10304 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_110
timestamp 1666464484
transform 1 0 11224 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_113
timestamp 1666464484
transform 1 0 11500 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_122
timestamp 1666464484
transform 1 0 12328 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_133
timestamp 1666464484
transform 1 0 13340 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_141
timestamp 1666464484
transform 1 0 14076 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_150
timestamp 1666464484
transform 1 0 14904 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_161
timestamp 1666464484
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1666464484
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_169
timestamp 1666464484
transform 1 0 16652 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_178
timestamp 1666464484
transform 1 0 17480 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_188
timestamp 1666464484
transform 1 0 18400 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_195
timestamp 1666464484
transform 1 0 19044 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_201
timestamp 1666464484
transform 1 0 19596 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_208
timestamp 1666464484
transform 1 0 20240 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_217
timestamp 1666464484
transform 1 0 21068 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_223
timestamp 1666464484
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_225
timestamp 1666464484
transform 1 0 21804 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_234
timestamp 1666464484
transform 1 0 22632 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_240
timestamp 1666464484
transform 1 0 23184 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_10_3
timestamp 1666464484
transform 1 0 1380 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_8
timestamp 1666464484
transform 1 0 1840 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_18
timestamp 1666464484
transform 1 0 2760 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_26
timestamp 1666464484
transform 1 0 3496 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_29
timestamp 1666464484
transform 1 0 3772 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_35
timestamp 1666464484
transform 1 0 4324 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_46
timestamp 1666464484
transform 1 0 5336 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_10_60
timestamp 1666464484
transform 1 0 6624 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_10_73
timestamp 1666464484
transform 1 0 7820 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_80
timestamp 1666464484
transform 1 0 8464 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_85
timestamp 1666464484
transform 1 0 8924 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_94
timestamp 1666464484
transform 1 0 9752 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_100
timestamp 1666464484
transform 1 0 10304 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_108
timestamp 1666464484
transform 1 0 11040 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_10_121
timestamp 1666464484
transform 1 0 12236 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_127
timestamp 1666464484
transform 1 0 12788 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_135
timestamp 1666464484
transform 1 0 13524 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1666464484
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_141
timestamp 1666464484
transform 1 0 14076 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_10_155
timestamp 1666464484
transform 1 0 15364 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_166
timestamp 1666464484
transform 1 0 16376 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_174
timestamp 1666464484
transform 1 0 17112 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_180
timestamp 1666464484
transform 1 0 17664 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_188
timestamp 1666464484
transform 1 0 18400 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_194
timestamp 1666464484
transform 1 0 18952 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_197
timestamp 1666464484
transform 1 0 19228 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_204
timestamp 1666464484
transform 1 0 19872 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_215
timestamp 1666464484
transform 1 0 20884 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_225
timestamp 1666464484
transform 1 0 21804 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_231
timestamp 1666464484
transform 1 0 22356 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_237
timestamp 1666464484
transform 1 0 22908 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_243
timestamp 1666464484
transform 1 0 23460 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_3
timestamp 1666464484
transform 1 0 1380 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_11
timestamp 1666464484
transform 1 0 2116 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_21
timestamp 1666464484
transform 1 0 3036 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_27
timestamp 1666464484
transform 1 0 3588 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_35
timestamp 1666464484
transform 1 0 4324 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_11_49
timestamp 1666464484
transform 1 0 5612 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1666464484
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_57
timestamp 1666464484
transform 1 0 6348 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_63
timestamp 1666464484
transform 1 0 6900 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_67
timestamp 1666464484
transform 1 0 7268 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_76
timestamp 1666464484
transform 1 0 8096 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_83
timestamp 1666464484
transform 1 0 8740 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_96
timestamp 1666464484
transform 1 0 9936 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_105
timestamp 1666464484
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1666464484
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_113
timestamp 1666464484
transform 1 0 11500 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_117
timestamp 1666464484
transform 1 0 11868 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_129
timestamp 1666464484
transform 1 0 12972 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_138
timestamp 1666464484
transform 1 0 13800 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_145
timestamp 1666464484
transform 1 0 14444 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_156
timestamp 1666464484
transform 1 0 15456 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_160
timestamp 1666464484
transform 1 0 15824 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_166
timestamp 1666464484
transform 1 0 16376 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_169
timestamp 1666464484
transform 1 0 16652 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_179
timestamp 1666464484
transform 1 0 17572 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_190
timestamp 1666464484
transform 1 0 18584 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_198
timestamp 1666464484
transform 1 0 19320 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_207
timestamp 1666464484
transform 1 0 20148 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_218
timestamp 1666464484
transform 1 0 21160 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_11_225
timestamp 1666464484
transform 1 0 21804 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_233
timestamp 1666464484
transform 1 0 22540 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_11_241
timestamp 1666464484
transform 1 0 23276 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_3
timestamp 1666464484
transform 1 0 1380 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_7
timestamp 1666464484
transform 1 0 1748 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_13
timestamp 1666464484
transform 1 0 2300 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_26
timestamp 1666464484
transform 1 0 3496 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_12_29
timestamp 1666464484
transform 1 0 3772 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_35
timestamp 1666464484
transform 1 0 4324 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_41
timestamp 1666464484
transform 1 0 4876 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_51
timestamp 1666464484
transform 1 0 5796 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_60
timestamp 1666464484
transform 1 0 6624 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_68
timestamp 1666464484
transform 1 0 7360 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_12_82
timestamp 1666464484
transform 1 0 8648 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_85
timestamp 1666464484
transform 1 0 8924 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_95
timestamp 1666464484
transform 1 0 9844 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_104
timestamp 1666464484
transform 1 0 10672 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_12_117
timestamp 1666464484
transform 1 0 11868 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_127
timestamp 1666464484
transform 1 0 12788 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_138
timestamp 1666464484
transform 1 0 13800 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_141
timestamp 1666464484
transform 1 0 14076 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_12_150
timestamp 1666464484
transform 1 0 14904 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_12_162
timestamp 1666464484
transform 1 0 16008 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_173
timestamp 1666464484
transform 1 0 17020 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_185
timestamp 1666464484
transform 1 0 18124 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_194
timestamp 1666464484
transform 1 0 18952 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_197
timestamp 1666464484
transform 1 0 19228 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_201
timestamp 1666464484
transform 1 0 19596 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_206
timestamp 1666464484
transform 1 0 20056 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_217
timestamp 1666464484
transform 1 0 21068 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_227
timestamp 1666464484
transform 1 0 21988 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_237
timestamp 1666464484
transform 1 0 22908 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_243
timestamp 1666464484
transform 1 0 23460 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_3
timestamp 1666464484
transform 1 0 1380 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_7
timestamp 1666464484
transform 1 0 1748 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_10
timestamp 1666464484
transform 1 0 2024 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_19
timestamp 1666464484
transform 1 0 2852 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_29
timestamp 1666464484
transform 1 0 3772 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_13_39
timestamp 1666464484
transform 1 0 4692 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_45
timestamp 1666464484
transform 1 0 5244 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_54
timestamp 1666464484
transform 1 0 6072 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_57
timestamp 1666464484
transform 1 0 6348 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_68
timestamp 1666464484
transform 1 0 7360 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_74
timestamp 1666464484
transform 1 0 7912 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_80
timestamp 1666464484
transform 1 0 8464 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_86
timestamp 1666464484
transform 1 0 9016 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_13_94
timestamp 1666464484
transform 1 0 9752 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_103
timestamp 1666464484
transform 1 0 10580 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_107
timestamp 1666464484
transform 1 0 10948 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_110
timestamp 1666464484
transform 1 0 11224 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_113
timestamp 1666464484
transform 1 0 11500 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_120
timestamp 1666464484
transform 1 0 12144 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_132
timestamp 1666464484
transform 1 0 13248 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_136
timestamp 1666464484
transform 1 0 13616 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_140
timestamp 1666464484
transform 1 0 13984 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_152
timestamp 1666464484
transform 1 0 15088 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_164
timestamp 1666464484
transform 1 0 16192 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_169
timestamp 1666464484
transform 1 0 16652 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_173
timestamp 1666464484
transform 1 0 17020 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_177
timestamp 1666464484
transform 1 0 17388 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_186
timestamp 1666464484
transform 1 0 18216 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_192
timestamp 1666464484
transform 1 0 18768 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_13_203
timestamp 1666464484
transform 1 0 19780 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_215
timestamp 1666464484
transform 1 0 20884 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_13_221
timestamp 1666464484
transform 1 0 21436 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_225
timestamp 1666464484
transform 1 0 21804 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_231
timestamp 1666464484
transform 1 0 22356 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_239
timestamp 1666464484
transform 1 0 23092 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_243
timestamp 1666464484
transform 1 0 23460 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_14_3
timestamp 1666464484
transform 1 0 1380 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_8
timestamp 1666464484
transform 1 0 1840 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_19
timestamp 1666464484
transform 1 0 2852 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_23
timestamp 1666464484
transform 1 0 3220 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_26
timestamp 1666464484
transform 1 0 3496 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_29
timestamp 1666464484
transform 1 0 3772 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_14_37
timestamp 1666464484
transform 1 0 4508 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_14_47
timestamp 1666464484
transform 1 0 5428 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_56
timestamp 1666464484
transform 1 0 6256 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_60
timestamp 1666464484
transform 1 0 6624 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_65
timestamp 1666464484
transform 1 0 7084 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_71
timestamp 1666464484
transform 1 0 7636 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_80
timestamp 1666464484
transform 1 0 8464 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_85
timestamp 1666464484
transform 1 0 8924 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_94
timestamp 1666464484
transform 1 0 9752 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_98
timestamp 1666464484
transform 1 0 10120 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_101
timestamp 1666464484
transform 1 0 10396 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_108
timestamp 1666464484
transform 1 0 11040 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_119
timestamp 1666464484
transform 1 0 12052 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_130
timestamp 1666464484
transform 1 0 13064 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_138
timestamp 1666464484
transform 1 0 13800 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_141
timestamp 1666464484
transform 1 0 14076 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_14_148
timestamp 1666464484
transform 1 0 14720 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_154
timestamp 1666464484
transform 1 0 15272 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_163
timestamp 1666464484
transform 1 0 16100 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_169
timestamp 1666464484
transform 1 0 16652 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_173
timestamp 1666464484
transform 1 0 17020 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_181
timestamp 1666464484
transform 1 0 17756 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_14_193
timestamp 1666464484
transform 1 0 18860 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_197
timestamp 1666464484
transform 1 0 19228 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_202
timestamp 1666464484
transform 1 0 19688 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_210
timestamp 1666464484
transform 1 0 20424 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_216
timestamp 1666464484
transform 1 0 20976 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_222
timestamp 1666464484
transform 1 0 21528 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_228
timestamp 1666464484
transform 1 0 22080 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_234
timestamp 1666464484
transform 1 0 22632 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_240
timestamp 1666464484
transform 1 0 23184 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_15_3
timestamp 1666464484
transform 1 0 1380 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_12
timestamp 1666464484
transform 1 0 2208 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_24
timestamp 1666464484
transform 1 0 3312 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_28
timestamp 1666464484
transform 1 0 3680 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_35
timestamp 1666464484
transform 1 0 4324 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_43
timestamp 1666464484
transform 1 0 5060 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_50
timestamp 1666464484
transform 1 0 5704 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_15_57
timestamp 1666464484
transform 1 0 6348 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_64
timestamp 1666464484
transform 1 0 6992 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_72
timestamp 1666464484
transform 1 0 7728 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_76
timestamp 1666464484
transform 1 0 8096 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_88
timestamp 1666464484
transform 1 0 9200 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_99
timestamp 1666464484
transform 1 0 10212 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_105
timestamp 1666464484
transform 1 0 10764 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_110
timestamp 1666464484
transform 1 0 11224 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_113
timestamp 1666464484
transform 1 0 11500 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_122
timestamp 1666464484
transform 1 0 12328 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_135
timestamp 1666464484
transform 1 0 13524 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_141
timestamp 1666464484
transform 1 0 14076 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_149
timestamp 1666464484
transform 1 0 14812 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_153
timestamp 1666464484
transform 1 0 15180 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_159
timestamp 1666464484
transform 1 0 15732 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_166
timestamp 1666464484
transform 1 0 16376 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_169
timestamp 1666464484
transform 1 0 16652 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_15_173
timestamp 1666464484
transform 1 0 17020 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_15_182
timestamp 1666464484
transform 1 0 17848 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_186
timestamp 1666464484
transform 1 0 18216 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_194
timestamp 1666464484
transform 1 0 18952 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_205
timestamp 1666464484
transform 1 0 19964 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_216
timestamp 1666464484
transform 1 0 20976 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_222
timestamp 1666464484
transform 1 0 21528 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_225
timestamp 1666464484
transform 1 0 21804 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_229
timestamp 1666464484
transform 1 0 22172 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_15_241
timestamp 1666464484
transform 1 0 23276 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_3
timestamp 1666464484
transform 1 0 1380 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_7
timestamp 1666464484
transform 1 0 1748 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_17
timestamp 1666464484
transform 1 0 2668 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_26
timestamp 1666464484
transform 1 0 3496 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_29
timestamp 1666464484
transform 1 0 3772 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_34
timestamp 1666464484
transform 1 0 4232 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_16_47
timestamp 1666464484
transform 1 0 5428 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_57
timestamp 1666464484
transform 1 0 6348 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_16_71
timestamp 1666464484
transform 1 0 7636 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_16_82
timestamp 1666464484
transform 1 0 8648 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_85
timestamp 1666464484
transform 1 0 8924 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_94
timestamp 1666464484
transform 1 0 9752 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_101
timestamp 1666464484
transform 1 0 10396 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_127
timestamp 1666464484
transform 1 0 12788 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_135
timestamp 1666464484
transform 1 0 13524 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 1666464484
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_141
timestamp 1666464484
transform 1 0 14076 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_151
timestamp 1666464484
transform 1 0 14996 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_158
timestamp 1666464484
transform 1 0 15640 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_168
timestamp 1666464484
transform 1 0 16560 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_176
timestamp 1666464484
transform 1 0 17296 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_184
timestamp 1666464484
transform 1 0 18032 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_194
timestamp 1666464484
transform 1 0 18952 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_197
timestamp 1666464484
transform 1 0 19228 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_205
timestamp 1666464484
transform 1 0 19964 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_217
timestamp 1666464484
transform 1 0 21068 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_226
timestamp 1666464484
transform 1 0 21896 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_233
timestamp 1666464484
transform 1 0 22540 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_16_241
timestamp 1666464484
transform 1 0 23276 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_17_3
timestamp 1666464484
transform 1 0 1380 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_9
timestamp 1666464484
transform 1 0 1932 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_13
timestamp 1666464484
transform 1 0 2300 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_21
timestamp 1666464484
transform 1 0 3036 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_28
timestamp 1666464484
transform 1 0 3680 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_34
timestamp 1666464484
transform 1 0 4232 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_41
timestamp 1666464484
transform 1 0 4876 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_54
timestamp 1666464484
transform 1 0 6072 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_57
timestamp 1666464484
transform 1 0 6348 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_17_67
timestamp 1666464484
transform 1 0 7268 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_73
timestamp 1666464484
transform 1 0 7820 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_81
timestamp 1666464484
transform 1 0 8556 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_17_94
timestamp 1666464484
transform 1 0 9752 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_102
timestamp 1666464484
transform 1 0 10488 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_17_110
timestamp 1666464484
transform 1 0 11224 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_113
timestamp 1666464484
transform 1 0 11500 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_122
timestamp 1666464484
transform 1 0 12328 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_132
timestamp 1666464484
transform 1 0 13248 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_141
timestamp 1666464484
transform 1 0 14076 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_150
timestamp 1666464484
transform 1 0 14904 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_154
timestamp 1666464484
transform 1 0 15272 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_164
timestamp 1666464484
transform 1 0 16192 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_169
timestamp 1666464484
transform 1 0 16652 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_178
timestamp 1666464484
transform 1 0 17480 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_184
timestamp 1666464484
transform 1 0 18032 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_195
timestamp 1666464484
transform 1 0 19044 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_201
timestamp 1666464484
transform 1 0 19596 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_205
timestamp 1666464484
transform 1 0 19964 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_214
timestamp 1666464484
transform 1 0 20792 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_222
timestamp 1666464484
transform 1 0 21528 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_225
timestamp 1666464484
transform 1 0 21804 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_233
timestamp 1666464484
transform 1 0 22540 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_239
timestamp 1666464484
transform 1 0 23092 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_243
timestamp 1666464484
transform 1 0 23460 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_3
timestamp 1666464484
transform 1 0 1380 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_18_13
timestamp 1666464484
transform 1 0 2300 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_23
timestamp 1666464484
transform 1 0 3220 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1666464484
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_29
timestamp 1666464484
transform 1 0 3772 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_18_38
timestamp 1666464484
transform 1 0 4600 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_18_51
timestamp 1666464484
transform 1 0 5796 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_63
timestamp 1666464484
transform 1 0 6900 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_75
timestamp 1666464484
transform 1 0 8004 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_79
timestamp 1666464484
transform 1 0 8372 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_82
timestamp 1666464484
transform 1 0 8648 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_85
timestamp 1666464484
transform 1 0 8924 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_95
timestamp 1666464484
transform 1 0 9844 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_101
timestamp 1666464484
transform 1 0 10396 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_109
timestamp 1666464484
transform 1 0 11132 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_112
timestamp 1666464484
transform 1 0 11408 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_119
timestamp 1666464484
transform 1 0 12052 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_130
timestamp 1666464484
transform 1 0 13064 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_136
timestamp 1666464484
transform 1 0 13616 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_141
timestamp 1666464484
transform 1 0 14076 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_18_151
timestamp 1666464484
transform 1 0 14996 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_157
timestamp 1666464484
transform 1 0 15548 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_161
timestamp 1666464484
transform 1 0 15916 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_171
timestamp 1666464484
transform 1 0 16836 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_175
timestamp 1666464484
transform 1 0 17204 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_182
timestamp 1666464484
transform 1 0 17848 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_194
timestamp 1666464484
transform 1 0 18952 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_18_197
timestamp 1666464484
transform 1 0 19228 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_18_208
timestamp 1666464484
transform 1 0 20240 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_18_220
timestamp 1666464484
transform 1 0 21344 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_227
timestamp 1666464484
transform 1 0 21988 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_233
timestamp 1666464484
transform 1 0 22540 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_241
timestamp 1666464484
transform 1 0 23276 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_3
timestamp 1666464484
transform 1 0 1380 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_9
timestamp 1666464484
transform 1 0 1932 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_20
timestamp 1666464484
transform 1 0 2944 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_19_33
timestamp 1666464484
transform 1 0 4140 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_39
timestamp 1666464484
transform 1 0 4692 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_49
timestamp 1666464484
transform 1 0 5612 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1666464484
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_57
timestamp 1666464484
transform 1 0 6348 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_19_66
timestamp 1666464484
transform 1 0 7176 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_19_74
timestamp 1666464484
transform 1 0 7912 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_19_84
timestamp 1666464484
transform 1 0 8832 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_95
timestamp 1666464484
transform 1 0 9844 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_106
timestamp 1666464484
transform 1 0 10856 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_19_113
timestamp 1666464484
transform 1 0 11500 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_121
timestamp 1666464484
transform 1 0 12236 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_145
timestamp 1666464484
transform 1 0 14444 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_156
timestamp 1666464484
transform 1 0 15456 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_166
timestamp 1666464484
transform 1 0 16376 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_169
timestamp 1666464484
transform 1 0 16652 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_19_179
timestamp 1666464484
transform 1 0 17572 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_185
timestamp 1666464484
transform 1 0 18124 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_192
timestamp 1666464484
transform 1 0 18768 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_201
timestamp 1666464484
transform 1 0 19596 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_19_216
timestamp 1666464484
transform 1 0 20976 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_222
timestamp 1666464484
transform 1 0 21528 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_225
timestamp 1666464484
transform 1 0 21804 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_229
timestamp 1666464484
transform 1 0 22172 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_19_241
timestamp 1666464484
transform 1 0 23276 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_3
timestamp 1666464484
transform 1 0 1380 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_7
timestamp 1666464484
transform 1 0 1748 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_11
timestamp 1666464484
transform 1 0 2116 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_20
timestamp 1666464484
transform 1 0 2944 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_26
timestamp 1666464484
transform 1 0 3496 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_29
timestamp 1666464484
transform 1 0 3772 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_33
timestamp 1666464484
transform 1 0 4140 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_36
timestamp 1666464484
transform 1 0 4416 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_48
timestamp 1666464484
transform 1 0 5520 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_20_63
timestamp 1666464484
transform 1 0 6900 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_70
timestamp 1666464484
transform 1 0 7544 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_77
timestamp 1666464484
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1666464484
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_85
timestamp 1666464484
transform 1 0 8924 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_98
timestamp 1666464484
transform 1 0 10120 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_104
timestamp 1666464484
transform 1 0 10672 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_110
timestamp 1666464484
transform 1 0 11224 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_117
timestamp 1666464484
transform 1 0 11868 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_125
timestamp 1666464484
transform 1 0 12604 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_132
timestamp 1666464484
transform 1 0 13248 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_20_141
timestamp 1666464484
transform 1 0 14076 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_20_151
timestamp 1666464484
transform 1 0 14996 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_159
timestamp 1666464484
transform 1 0 15732 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_166
timestamp 1666464484
transform 1 0 16376 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_173
timestamp 1666464484
transform 1 0 17020 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_20_187
timestamp 1666464484
transform 1 0 18308 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_194
timestamp 1666464484
transform 1 0 18952 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_197
timestamp 1666464484
transform 1 0 19228 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_207
timestamp 1666464484
transform 1 0 20148 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_216
timestamp 1666464484
transform 1 0 20976 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_224
timestamp 1666464484
transform 1 0 21712 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_236
timestamp 1666464484
transform 1 0 22816 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_21_3
timestamp 1666464484
transform 1 0 1380 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_7
timestamp 1666464484
transform 1 0 1748 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_10
timestamp 1666464484
transform 1 0 2024 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_18
timestamp 1666464484
transform 1 0 2760 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_25
timestamp 1666464484
transform 1 0 3404 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_21_36
timestamp 1666464484
transform 1 0 4416 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_40
timestamp 1666464484
transform 1 0 4784 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_48
timestamp 1666464484
transform 1 0 5520 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_54
timestamp 1666464484
transform 1 0 6072 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_57
timestamp 1666464484
transform 1 0 6348 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_21_67
timestamp 1666464484
transform 1 0 7268 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_21_79
timestamp 1666464484
transform 1 0 8372 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_21_96
timestamp 1666464484
transform 1 0 9936 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_100
timestamp 1666464484
transform 1 0 10304 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_110
timestamp 1666464484
transform 1 0 11224 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_113
timestamp 1666464484
transform 1 0 11500 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_123
timestamp 1666464484
transform 1 0 12420 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_129
timestamp 1666464484
transform 1 0 12972 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_21_141
timestamp 1666464484
transform 1 0 14076 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_149
timestamp 1666464484
transform 1 0 14812 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_160
timestamp 1666464484
transform 1 0 15824 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_166
timestamp 1666464484
transform 1 0 16376 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_169
timestamp 1666464484
transform 1 0 16652 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_177
timestamp 1666464484
transform 1 0 17388 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_181
timestamp 1666464484
transform 1 0 17756 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_189
timestamp 1666464484
transform 1 0 18492 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_195
timestamp 1666464484
transform 1 0 19044 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_203
timestamp 1666464484
transform 1 0 19780 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_210
timestamp 1666464484
transform 1 0 20424 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_222
timestamp 1666464484
transform 1 0 21528 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_225
timestamp 1666464484
transform 1 0 21804 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_237
timestamp 1666464484
transform 1 0 22908 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_243
timestamp 1666464484
transform 1 0 23460 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_3
timestamp 1666464484
transform 1 0 1380 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_9
timestamp 1666464484
transform 1 0 1932 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_12
timestamp 1666464484
transform 1 0 2208 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_21
timestamp 1666464484
transform 1 0 3036 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1666464484
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_22_29
timestamp 1666464484
transform 1 0 3772 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_36
timestamp 1666464484
transform 1 0 4416 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_59
timestamp 1666464484
transform 1 0 6532 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_68
timestamp 1666464484
transform 1 0 7360 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_72
timestamp 1666464484
transform 1 0 7728 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_80
timestamp 1666464484
transform 1 0 8464 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_85
timestamp 1666464484
transform 1 0 8924 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_91
timestamp 1666464484
transform 1 0 9476 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_98
timestamp 1666464484
transform 1 0 10120 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_106
timestamp 1666464484
transform 1 0 10856 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_116
timestamp 1666464484
transform 1 0 11776 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_126
timestamp 1666464484
transform 1 0 12696 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_134
timestamp 1666464484
transform 1 0 13432 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_138
timestamp 1666464484
transform 1 0 13800 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_141
timestamp 1666464484
transform 1 0 14076 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_22_149
timestamp 1666464484
transform 1 0 14812 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_155
timestamp 1666464484
transform 1 0 15364 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_164
timestamp 1666464484
transform 1 0 16192 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_176
timestamp 1666464484
transform 1 0 17296 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_184
timestamp 1666464484
transform 1 0 18032 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_194
timestamp 1666464484
transform 1 0 18952 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_197
timestamp 1666464484
transform 1 0 19228 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_22_202
timestamp 1666464484
transform 1 0 19688 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_208
timestamp 1666464484
transform 1 0 20240 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_213
timestamp 1666464484
transform 1 0 20700 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_225
timestamp 1666464484
transform 1 0 21804 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_237
timestamp 1666464484
transform 1 0 22908 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_243
timestamp 1666464484
transform 1 0 23460 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_3
timestamp 1666464484
transform 1 0 1380 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_11
timestamp 1666464484
transform 1 0 2116 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_20
timestamp 1666464484
transform 1 0 2944 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_31
timestamp 1666464484
transform 1 0 3956 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_42
timestamp 1666464484
transform 1 0 4968 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_52
timestamp 1666464484
transform 1 0 5888 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_57
timestamp 1666464484
transform 1 0 6348 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_65
timestamp 1666464484
transform 1 0 7084 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_73
timestamp 1666464484
transform 1 0 7820 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_81
timestamp 1666464484
transform 1 0 8556 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_92
timestamp 1666464484
transform 1 0 9568 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_100
timestamp 1666464484
transform 1 0 10304 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_110
timestamp 1666464484
transform 1 0 11224 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_113
timestamp 1666464484
transform 1 0 11500 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_121
timestamp 1666464484
transform 1 0 12236 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_128
timestamp 1666464484
transform 1 0 12880 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_134
timestamp 1666464484
transform 1 0 13432 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_141
timestamp 1666464484
transform 1 0 14076 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_148
timestamp 1666464484
transform 1 0 14720 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_23_161
timestamp 1666464484
transform 1 0 15916 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_167
timestamp 1666464484
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_169
timestamp 1666464484
transform 1 0 16652 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_175
timestamp 1666464484
transform 1 0 17204 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_181
timestamp 1666464484
transform 1 0 17756 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_23_193
timestamp 1666464484
transform 1 0 18860 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_203
timestamp 1666464484
transform 1 0 19780 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_215
timestamp 1666464484
transform 1 0 20884 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_223
timestamp 1666464484
transform 1 0 21620 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_225
timestamp 1666464484
transform 1 0 21804 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_237
timestamp 1666464484
transform 1 0 22908 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_243
timestamp 1666464484
transform 1 0 23460 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_3
timestamp 1666464484
transform 1 0 1380 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_11
timestamp 1666464484
transform 1 0 2116 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_24
timestamp 1666464484
transform 1 0 3312 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_29
timestamp 1666464484
transform 1 0 3772 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_47
timestamp 1666464484
transform 1 0 5428 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_54
timestamp 1666464484
transform 1 0 6072 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_67
timestamp 1666464484
transform 1 0 7268 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_80
timestamp 1666464484
transform 1 0 8464 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_85
timestamp 1666464484
transform 1 0 8924 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_90
timestamp 1666464484
transform 1 0 9384 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_110
timestamp 1666464484
transform 1 0 11224 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_123
timestamp 1666464484
transform 1 0 12420 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_134
timestamp 1666464484
transform 1 0 13432 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_24_141
timestamp 1666464484
transform 1 0 14076 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_150
timestamp 1666464484
transform 1 0 14904 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_164
timestamp 1666464484
transform 1 0 16192 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_177
timestamp 1666464484
transform 1 0 17388 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_24_185
timestamp 1666464484
transform 1 0 18124 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_24_193
timestamp 1666464484
transform 1 0 18860 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_197
timestamp 1666464484
transform 1 0 19228 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_201
timestamp 1666464484
transform 1 0 19596 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_213
timestamp 1666464484
transform 1 0 20700 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_225
timestamp 1666464484
transform 1 0 21804 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_237
timestamp 1666464484
transform 1 0 22908 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_243
timestamp 1666464484
transform 1 0 23460 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_25_3
timestamp 1666464484
transform 1 0 1380 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_11
timestamp 1666464484
transform 1 0 2116 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_15
timestamp 1666464484
transform 1 0 2484 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_36
timestamp 1666464484
transform 1 0 4416 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_47
timestamp 1666464484
transform 1 0 5428 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_54
timestamp 1666464484
transform 1 0 6072 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_57
timestamp 1666464484
transform 1 0 6348 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_61
timestamp 1666464484
transform 1 0 6716 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_69
timestamp 1666464484
transform 1 0 7452 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_93
timestamp 1666464484
transform 1 0 9660 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_25_101
timestamp 1666464484
transform 1 0 10396 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_107
timestamp 1666464484
transform 1 0 10948 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_110
timestamp 1666464484
transform 1 0 11224 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_113
timestamp 1666464484
transform 1 0 11500 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_25_122
timestamp 1666464484
transform 1 0 12328 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_134
timestamp 1666464484
transform 1 0 13432 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_140
timestamp 1666464484
transform 1 0 13984 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_143
timestamp 1666464484
transform 1 0 14260 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_155
timestamp 1666464484
transform 1 0 15364 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_25_167
timestamp 1666464484
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_169
timestamp 1666464484
transform 1 0 16652 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_181
timestamp 1666464484
transform 1 0 17756 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_193
timestamp 1666464484
transform 1 0 18860 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_205
timestamp 1666464484
transform 1 0 19964 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_217
timestamp 1666464484
transform 1 0 21068 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_223
timestamp 1666464484
transform 1 0 21620 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_225
timestamp 1666464484
transform 1 0 21804 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_237
timestamp 1666464484
transform 1 0 22908 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_243
timestamp 1666464484
transform 1 0 23460 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_3
timestamp 1666464484
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_18
timestamp 1666464484
transform 1 0 2760 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_26
timestamp 1666464484
transform 1 0 3496 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_29
timestamp 1666464484
transform 1 0 3772 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_37
timestamp 1666464484
transform 1 0 4508 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_54
timestamp 1666464484
transform 1 0 6072 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_62
timestamp 1666464484
transform 1 0 6808 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_79
timestamp 1666464484
transform 1 0 8372 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1666464484
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_85
timestamp 1666464484
transform 1 0 8924 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_89
timestamp 1666464484
transform 1 0 9292 0 1 16320
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_26_113
timestamp 1666464484
transform 1 0 11500 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_125
timestamp 1666464484
transform 1 0 12604 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_26_137
timestamp 1666464484
transform 1 0 13708 0 1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_26_141
timestamp 1666464484
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_153
timestamp 1666464484
transform 1 0 15180 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_161
timestamp 1666464484
transform 1 0 15916 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_166
timestamp 1666464484
transform 1 0 16376 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_178
timestamp 1666464484
transform 1 0 17480 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_190
timestamp 1666464484
transform 1 0 18584 0 1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_26_197
timestamp 1666464484
transform 1 0 19228 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_209
timestamp 1666464484
transform 1 0 20332 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_221
timestamp 1666464484
transform 1 0 21436 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_233
timestamp 1666464484
transform 1 0 22540 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_26_241
timestamp 1666464484
transform 1 0 23276 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_27_3
timestamp 1666464484
transform 1 0 1380 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_27_27
timestamp 1666464484
transform 1 0 3588 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_48
timestamp 1666464484
transform 1 0 5520 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_27_57
timestamp 1666464484
transform 1 0 6348 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_63
timestamp 1666464484
transform 1 0 6900 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_81
timestamp 1666464484
transform 1 0 8556 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_93
timestamp 1666464484
transform 1 0 9660 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_110
timestamp 1666464484
transform 1 0 11224 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_113
timestamp 1666464484
transform 1 0 11500 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_117
timestamp 1666464484
transform 1 0 11868 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_129
timestamp 1666464484
transform 1 0 12972 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_141
timestamp 1666464484
transform 1 0 14076 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_153
timestamp 1666464484
transform 1 0 15180 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_165
timestamp 1666464484
transform 1 0 16284 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_27_169
timestamp 1666464484
transform 1 0 16652 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_181
timestamp 1666464484
transform 1 0 17756 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_193
timestamp 1666464484
transform 1 0 18860 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_205
timestamp 1666464484
transform 1 0 19964 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_217
timestamp 1666464484
transform 1 0 21068 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_223
timestamp 1666464484
transform 1 0 21620 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_225
timestamp 1666464484
transform 1 0 21804 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_237
timestamp 1666464484
transform 1 0 22908 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_243
timestamp 1666464484
transform 1 0 23460 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_28_3
timestamp 1666464484
transform 1 0 1380 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_9
timestamp 1666464484
transform 1 0 1932 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_26
timestamp 1666464484
transform 1 0 3496 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_29
timestamp 1666464484
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_41
timestamp 1666464484
transform 1 0 4876 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_65
timestamp 1666464484
transform 1 0 7084 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_73
timestamp 1666464484
transform 1 0 7820 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_79
timestamp 1666464484
transform 1 0 8372 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_83
timestamp 1666464484
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_85
timestamp 1666464484
transform 1 0 8924 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_93
timestamp 1666464484
transform 1 0 9660 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_111
timestamp 1666464484
transform 1 0 11316 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_132
timestamp 1666464484
transform 1 0 13248 0 1 17408
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_28_141
timestamp 1666464484
transform 1 0 14076 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_153
timestamp 1666464484
transform 1 0 15180 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_165
timestamp 1666464484
transform 1 0 16284 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_177
timestamp 1666464484
transform 1 0 17388 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_189
timestamp 1666464484
transform 1 0 18492 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_195
timestamp 1666464484
transform 1 0 19044 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_197
timestamp 1666464484
transform 1 0 19228 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_209
timestamp 1666464484
transform 1 0 20332 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_221
timestamp 1666464484
transform 1 0 21436 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_233
timestamp 1666464484
transform 1 0 22540 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_28_241
timestamp 1666464484
transform 1 0 23276 0 1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_29_3
timestamp 1666464484
transform 1 0 1380 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_15
timestamp 1666464484
transform 1 0 2484 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_23
timestamp 1666464484
transform 1 0 3220 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_42
timestamp 1666464484
transform 1 0 4968 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_54
timestamp 1666464484
transform 1 0 6072 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_57
timestamp 1666464484
transform 1 0 6348 0 -1 18496
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_29_81
timestamp 1666464484
transform 1 0 8556 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_29_93
timestamp 1666464484
transform 1 0 9660 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_110
timestamp 1666464484
transform 1 0 11224 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_113
timestamp 1666464484
transform 1 0 11500 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_117
timestamp 1666464484
transform 1 0 11868 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_29_123
timestamp 1666464484
transform 1 0 12420 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_135
timestamp 1666464484
transform 1 0 13524 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_147
timestamp 1666464484
transform 1 0 14628 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_159
timestamp 1666464484
transform 1 0 15732 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_167
timestamp 1666464484
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_169
timestamp 1666464484
transform 1 0 16652 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_181
timestamp 1666464484
transform 1 0 17756 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_193
timestamp 1666464484
transform 1 0 18860 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_205
timestamp 1666464484
transform 1 0 19964 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_217
timestamp 1666464484
transform 1 0 21068 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_223
timestamp 1666464484
transform 1 0 21620 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_225
timestamp 1666464484
transform 1 0 21804 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_237
timestamp 1666464484
transform 1 0 22908 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_243
timestamp 1666464484
transform 1 0 23460 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_3
timestamp 1666464484
transform 1 0 1380 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_11
timestamp 1666464484
transform 1 0 2116 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_16
timestamp 1666464484
transform 1 0 2576 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_29
timestamp 1666464484
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_41
timestamp 1666464484
transform 1 0 4876 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_58
timestamp 1666464484
transform 1 0 6440 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_79
timestamp 1666464484
transform 1 0 8372 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp 1666464484
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_85
timestamp 1666464484
transform 1 0 8924 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_30_90
timestamp 1666464484
transform 1 0 9384 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_96
timestamp 1666464484
transform 1 0 9936 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_116
timestamp 1666464484
transform 1 0 11776 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_30_122
timestamp 1666464484
transform 1 0 12328 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_134
timestamp 1666464484
transform 1 0 13432 0 1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_30_141
timestamp 1666464484
transform 1 0 14076 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_153
timestamp 1666464484
transform 1 0 15180 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_165
timestamp 1666464484
transform 1 0 16284 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_177
timestamp 1666464484
transform 1 0 17388 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_185
timestamp 1666464484
transform 1 0 18124 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_30_189
timestamp 1666464484
transform 1 0 18492 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_195
timestamp 1666464484
transform 1 0 19044 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_197
timestamp 1666464484
transform 1 0 19228 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_209
timestamp 1666464484
transform 1 0 20332 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_221
timestamp 1666464484
transform 1 0 21436 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_233
timestamp 1666464484
transform 1 0 22540 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_30_241
timestamp 1666464484
transform 1 0 23276 0 1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_31_3
timestamp 1666464484
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_15
timestamp 1666464484
transform 1 0 2484 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_31_27
timestamp 1666464484
transform 1 0 3588 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_44
timestamp 1666464484
transform 1 0 5152 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_57
timestamp 1666464484
transform 1 0 6348 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_31_67
timestamp 1666464484
transform 1 0 7268 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_31_91
timestamp 1666464484
transform 1 0 9476 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_103
timestamp 1666464484
transform 1 0 10580 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_111
timestamp 1666464484
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_113
timestamp 1666464484
transform 1 0 11500 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_125
timestamp 1666464484
transform 1 0 12604 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_137
timestamp 1666464484
transform 1 0 13708 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_149
timestamp 1666464484
transform 1 0 14812 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_161
timestamp 1666464484
transform 1 0 15916 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_167
timestamp 1666464484
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_169
timestamp 1666464484
transform 1 0 16652 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_181
timestamp 1666464484
transform 1 0 17756 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_193
timestamp 1666464484
transform 1 0 18860 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_205
timestamp 1666464484
transform 1 0 19964 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_217
timestamp 1666464484
transform 1 0 21068 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_223
timestamp 1666464484
transform 1 0 21620 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_225
timestamp 1666464484
transform 1 0 21804 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_237
timestamp 1666464484
transform 1 0 22908 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_243
timestamp 1666464484
transform 1 0 23460 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_3
timestamp 1666464484
transform 1 0 1380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_15
timestamp 1666464484
transform 1 0 2484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1666464484
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_29
timestamp 1666464484
transform 1 0 3772 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_48
timestamp 1666464484
transform 1 0 5520 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_60
timestamp 1666464484
transform 1 0 6624 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_32_78
timestamp 1666464484
transform 1 0 8280 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_32_85
timestamp 1666464484
transform 1 0 8924 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_93
timestamp 1666464484
transform 1 0 9660 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_110
timestamp 1666464484
transform 1 0 11224 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_130
timestamp 1666464484
transform 1 0 13064 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_138
timestamp 1666464484
transform 1 0 13800 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_141
timestamp 1666464484
transform 1 0 14076 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_153
timestamp 1666464484
transform 1 0 15180 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_165
timestamp 1666464484
transform 1 0 16284 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_177
timestamp 1666464484
transform 1 0 17388 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_189
timestamp 1666464484
transform 1 0 18492 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_195
timestamp 1666464484
transform 1 0 19044 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_197
timestamp 1666464484
transform 1 0 19228 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_209
timestamp 1666464484
transform 1 0 20332 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_221
timestamp 1666464484
transform 1 0 21436 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_233
timestamp 1666464484
transform 1 0 22540 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_32_241
timestamp 1666464484
transform 1 0 23276 0 1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_33_3
timestamp 1666464484
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_15
timestamp 1666464484
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_27
timestamp 1666464484
transform 1 0 3588 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_33
timestamp 1666464484
transform 1 0 4140 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_50
timestamp 1666464484
transform 1 0 5704 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_33_57
timestamp 1666464484
transform 1 0 6348 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_65
timestamp 1666464484
transform 1 0 7084 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_82
timestamp 1666464484
transform 1 0 8648 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_110
timestamp 1666464484
transform 1 0 11224 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_113
timestamp 1666464484
transform 1 0 11500 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_117
timestamp 1666464484
transform 1 0 11868 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_33_125
timestamp 1666464484
transform 1 0 12604 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_33_131
timestamp 1666464484
transform 1 0 13156 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_143
timestamp 1666464484
transform 1 0 14260 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_155
timestamp 1666464484
transform 1 0 15364 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_33_167
timestamp 1666464484
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_169
timestamp 1666464484
transform 1 0 16652 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_181
timestamp 1666464484
transform 1 0 17756 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_193
timestamp 1666464484
transform 1 0 18860 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_205
timestamp 1666464484
transform 1 0 19964 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_217
timestamp 1666464484
transform 1 0 21068 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_223
timestamp 1666464484
transform 1 0 21620 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_225
timestamp 1666464484
transform 1 0 21804 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_237
timestamp 1666464484
transform 1 0 22908 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_243
timestamp 1666464484
transform 1 0 23460 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_3
timestamp 1666464484
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_15
timestamp 1666464484
transform 1 0 2484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1666464484
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_29
timestamp 1666464484
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_57
timestamp 1666464484
transform 1 0 6348 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_77
timestamp 1666464484
transform 1 0 8188 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_83
timestamp 1666464484
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_85
timestamp 1666464484
transform 1 0 8924 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_97
timestamp 1666464484
transform 1 0 10028 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_121
timestamp 1666464484
transform 1 0 12236 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_34_136
timestamp 1666464484
transform 1 0 13616 0 1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_34_141
timestamp 1666464484
transform 1 0 14076 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_153
timestamp 1666464484
transform 1 0 15180 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_165
timestamp 1666464484
transform 1 0 16284 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_177
timestamp 1666464484
transform 1 0 17388 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_189
timestamp 1666464484
transform 1 0 18492 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_195
timestamp 1666464484
transform 1 0 19044 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_197
timestamp 1666464484
transform 1 0 19228 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_209
timestamp 1666464484
transform 1 0 20332 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_221
timestamp 1666464484
transform 1 0 21436 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_233
timestamp 1666464484
transform 1 0 22540 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_34_241
timestamp 1666464484
transform 1 0 23276 0 1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_35_3
timestamp 1666464484
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_15
timestamp 1666464484
transform 1 0 2484 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_27
timestamp 1666464484
transform 1 0 3588 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_39
timestamp 1666464484
transform 1 0 4692 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_51
timestamp 1666464484
transform 1 0 5796 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_55
timestamp 1666464484
transform 1 0 6164 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_35_57
timestamp 1666464484
transform 1 0 6348 0 -1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_35_76
timestamp 1666464484
transform 1 0 8096 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_88
timestamp 1666464484
transform 1 0 9200 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_35_110
timestamp 1666464484
transform 1 0 11224 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_113
timestamp 1666464484
transform 1 0 11500 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_131
timestamp 1666464484
transform 1 0 13156 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_143
timestamp 1666464484
transform 1 0 14260 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_35_150
timestamp 1666464484
transform 1 0 14904 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_162
timestamp 1666464484
transform 1 0 16008 0 -1 21760
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_35_169
timestamp 1666464484
transform 1 0 16652 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_181
timestamp 1666464484
transform 1 0 17756 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_193
timestamp 1666464484
transform 1 0 18860 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_205
timestamp 1666464484
transform 1 0 19964 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_217
timestamp 1666464484
transform 1 0 21068 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_223
timestamp 1666464484
transform 1 0 21620 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_225
timestamp 1666464484
transform 1 0 21804 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_237
timestamp 1666464484
transform 1 0 22908 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_243
timestamp 1666464484
transform 1 0 23460 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_3
timestamp 1666464484
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_15
timestamp 1666464484
transform 1 0 2484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 1666464484
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_29
timestamp 1666464484
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_41
timestamp 1666464484
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_36_53
timestamp 1666464484
transform 1 0 5980 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_36_57
timestamp 1666464484
transform 1 0 6348 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_63
timestamp 1666464484
transform 1 0 6900 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_66
timestamp 1666464484
transform 1 0 7176 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_74
timestamp 1666464484
transform 1 0 7912 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_82
timestamp 1666464484
transform 1 0 8648 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_36_85
timestamp 1666464484
transform 1 0 8924 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_36_90
timestamp 1666464484
transform 1 0 9384 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_110
timestamp 1666464484
transform 1 0 11224 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_113
timestamp 1666464484
transform 1 0 11500 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_131
timestamp 1666464484
transform 1 0 13156 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_138
timestamp 1666464484
transform 1 0 13800 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_141
timestamp 1666464484
transform 1 0 14076 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_148
timestamp 1666464484
transform 1 0 14720 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_36_154
timestamp 1666464484
transform 1 0 15272 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_36_166
timestamp 1666464484
transform 1 0 16376 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_36_169
timestamp 1666464484
transform 1 0 16652 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_177
timestamp 1666464484
transform 1 0 17388 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_181
timestamp 1666464484
transform 1 0 17756 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_187
timestamp 1666464484
transform 1 0 18308 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_195
timestamp 1666464484
transform 1 0 19044 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_197
timestamp 1666464484
transform 1 0 19228 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_209
timestamp 1666464484
transform 1 0 20332 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_36_221
timestamp 1666464484
transform 1 0 21436 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_36_225
timestamp 1666464484
transform 1 0 21804 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_231
timestamp 1666464484
transform 1 0 22356 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_235
timestamp 1666464484
transform 1 0 22724 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_36_241
timestamp 1666464484
transform 1 0 23276 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1666464484
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1666464484
transform -1 0 23828 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1666464484
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1666464484
transform -1 0 23828 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1666464484
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1666464484
transform -1 0 23828 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1666464484
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1666464484
transform -1 0 23828 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1666464484
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1666464484
transform -1 0 23828 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1666464484
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1666464484
transform -1 0 23828 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1666464484
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1666464484
transform -1 0 23828 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1666464484
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1666464484
transform -1 0 23828 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1666464484
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1666464484
transform -1 0 23828 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1666464484
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1666464484
transform -1 0 23828 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1666464484
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1666464484
transform -1 0 23828 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1666464484
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1666464484
transform -1 0 23828 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1666464484
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1666464484
transform -1 0 23828 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1666464484
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1666464484
transform -1 0 23828 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1666464484
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1666464484
transform -1 0 23828 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1666464484
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1666464484
transform -1 0 23828 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1666464484
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1666464484
transform -1 0 23828 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1666464484
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1666464484
transform -1 0 23828 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1666464484
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1666464484
transform -1 0 23828 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1666464484
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1666464484
transform -1 0 23828 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1666464484
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1666464484
transform -1 0 23828 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1666464484
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1666464484
transform -1 0 23828 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1666464484
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1666464484
transform -1 0 23828 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1666464484
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1666464484
transform -1 0 23828 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1666464484
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1666464484
transform -1 0 23828 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1666464484
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1666464484
transform -1 0 23828 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1666464484
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1666464484
transform -1 0 23828 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1666464484
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1666464484
transform -1 0 23828 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1666464484
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1666464484
transform -1 0 23828 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1666464484
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1666464484
transform -1 0 23828 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1666464484
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1666464484
transform -1 0 23828 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1666464484
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1666464484
transform -1 0 23828 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1666464484
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1666464484
transform -1 0 23828 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1666464484
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1666464484
transform -1 0 23828 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1666464484
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1666464484
transform -1 0 23828 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1666464484
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1666464484
transform -1 0 23828 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1666464484
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1666464484
transform -1 0 23828 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1666464484
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1666464484
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1666464484
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1666464484
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1666464484
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1666464484
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1666464484
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1666464484
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1666464484
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1666464484
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1666464484
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1666464484
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1666464484
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1666464484
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1666464484
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1666464484
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1666464484
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1666464484
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1666464484
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1666464484
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1666464484
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1666464484
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1666464484
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1666464484
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1666464484
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1666464484
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1666464484
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1666464484
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1666464484
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1666464484
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1666464484
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1666464484
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1666464484
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1666464484
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1666464484
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1666464484
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1666464484
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1666464484
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1666464484
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1666464484
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1666464484
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1666464484
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1666464484
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1666464484
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1666464484
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1666464484
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1666464484
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1666464484
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1666464484
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1666464484
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1666464484
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1666464484
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1666464484
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1666464484
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1666464484
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1666464484
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1666464484
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1666464484
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1666464484
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1666464484
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1666464484
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1666464484
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1666464484
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1666464484
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1666464484
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1666464484
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1666464484
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1666464484
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1666464484
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1666464484
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1666464484
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1666464484
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1666464484
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1666464484
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1666464484
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1666464484
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1666464484
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1666464484
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1666464484
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1666464484
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1666464484
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1666464484
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1666464484
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1666464484
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1666464484
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1666464484
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1666464484
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1666464484
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1666464484
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1666464484
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1666464484
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1666464484
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1666464484
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1666464484
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1666464484
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1666464484
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1666464484
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1666464484
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1666464484
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1666464484
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1666464484
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1666464484
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1666464484
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1666464484
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1666464484
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1666464484
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1666464484
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1666464484
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1666464484
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1666464484
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1666464484
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1666464484
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1666464484
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1666464484
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1666464484
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1666464484
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1666464484
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1666464484
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1666464484
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1666464484
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1666464484
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1666464484
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1666464484
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1666464484
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1666464484
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1666464484
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1666464484
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1666464484
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1666464484
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1666464484
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1666464484
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1666464484
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1666464484
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1666464484
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1666464484
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1666464484
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1666464484
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1666464484
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1666464484
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1666464484
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1666464484
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1666464484
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1666464484
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1666464484
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1666464484
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1666464484
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1666464484
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1666464484
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1666464484
transform 1 0 6256 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1666464484
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1666464484
transform 1 0 11408 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1666464484
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1666464484
transform 1 0 16560 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1666464484
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1666464484
transform 1 0 21712 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_4  _404_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 6440 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _405_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 7544 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _406_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 2300 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_1  _407_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 4324 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _408_
timestamp 1666464484
transform 1 0 2944 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _409_
timestamp 1666464484
transform 1 0 3956 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _410_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 7360 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _411_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 2668 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _412_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 5704 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _413_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 4692 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _414_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 5336 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _415_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 2392 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nor2b_4  _416_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 8924 0 -1 14144
box -38 -48 1050 592
use sky130_fd_sc_hd__nor2_1  _417_
timestamp 1666464484
transform -1 0 4416 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__nand4b_4  _418_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 6532 0 1 14144
box -38 -48 1786 592
use sky130_fd_sc_hd__nor3_1  _419_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 10120 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_2  _420_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 10120 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__or2b_1  _421_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 1656 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _422_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 2300 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _423_
timestamp 1666464484
transform 1 0 2116 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _424_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 3496 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_1  _425_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 2852 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _426_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 2576 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _427_
timestamp 1666464484
transform 1 0 1564 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__and3_2  _428_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 2024 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_2  _429_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 3680 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _430_
timestamp 1666464484
transform 1 0 8096 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__or2b_2  _431_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 9568 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _432_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 9292 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__and2_2  _433_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 2484 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _434_
timestamp 1666464484
transform 1 0 3220 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__a211oi_4  _435_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 8464 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__xor2_1  _436_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 9844 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _437_
timestamp 1666464484
transform 1 0 4600 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _438_
timestamp 1666464484
transform 1 0 6532 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _439_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 3128 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _440_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 4416 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__or4b_1  _441_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 7912 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _442_
timestamp 1666464484
transform -1 0 2116 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__or3_2  _443_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 5244 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _444_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 9844 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _445_
timestamp 1666464484
transform -1 0 5888 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and4_2  _446_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 4968 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__nand3b_1  _447_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 2208 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _448_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 2116 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _449_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 2668 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__or2_2  _450_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 3404 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__and4bb_1  _451_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 3680 0 -1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__nor2b_4  _452_
timestamp 1666464484
transform 1 0 9108 0 1 13056
box -38 -48 1050 592
use sky130_fd_sc_hd__buf_2  _453_
timestamp 1666464484
transform -1 0 3496 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_2  _454_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 2668 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _455_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 5244 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__o311ai_4  _456_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 4692 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__o311a_1  _457_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 2668 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__o31a_1  _458_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 2208 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_1  _459_
timestamp 1666464484
transform 1 0 2116 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _460_
timestamp 1666464484
transform 1 0 9108 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _461_
timestamp 1666464484
transform 1 0 2484 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _462_
timestamp 1666464484
transform 1 0 2576 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _463_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 8188 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__a41o_1  _464_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 9844 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _465_
timestamp 1666464484
transform -1 0 5612 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _466_
timestamp 1666464484
transform -1 0 9660 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _467_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 10672 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _468_
timestamp 1666464484
transform 1 0 12052 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _469_
timestamp 1666464484
transform 1 0 10212 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__a41oi_4  _470_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 10948 0 -1 4352
box -38 -48 2062 592
use sky130_fd_sc_hd__clkbuf_4  _471_
timestamp 1666464484
transform 1 0 6532 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _472_
timestamp 1666464484
transform 1 0 10948 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _473_
timestamp 1666464484
transform -1 0 11960 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _474_
timestamp 1666464484
transform 1 0 11224 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__or4b_1  _475_
timestamp 1666464484
transform 1 0 10488 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  _476_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 11224 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_4  _477_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 12420 0 -1 13056
box -38 -48 2062 592
use sky130_fd_sc_hd__nor2_2  _478_
timestamp 1666464484
transform 1 0 18952 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _479_
timestamp 1666464484
transform 1 0 22264 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _480_
timestamp 1666464484
transform -1 0 21344 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkinv_2  _481_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 11960 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _482_
timestamp 1666464484
transform 1 0 10672 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__o31a_2  _483_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 11684 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _484_
timestamp 1666464484
transform -1 0 10580 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _485_
timestamp 1666464484
transform -1 0 12420 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__or3_2  _486_
timestamp 1666464484
transform 1 0 14444 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _487_
timestamp 1666464484
transform -1 0 12604 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _488_
timestamp 1666464484
transform -1 0 11224 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_2  _489_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 12236 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_2  _490_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 20608 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _491_
timestamp 1666464484
transform 1 0 12788 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__or4_4  _492_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 11960 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__or2_2  _493_
timestamp 1666464484
transform 1 0 15272 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _494_
timestamp 1666464484
transform -1 0 15364 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _495_
timestamp 1666464484
transform -1 0 12512 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _496_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 10396 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_1  _497_
timestamp 1666464484
transform -1 0 10856 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _498_
timestamp 1666464484
transform 1 0 15456 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_1  _499_
timestamp 1666464484
transform -1 0 12328 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _500_
timestamp 1666464484
transform -1 0 11592 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_2  _501_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 14260 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _502_
timestamp 1666464484
transform -1 0 17112 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _503_
timestamp 1666464484
transform -1 0 12052 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__nor3_1  _504_
timestamp 1666464484
transform -1 0 10856 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _505_
timestamp 1666464484
transform -1 0 11868 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__nor3_2  _506_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 11684 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _507_
timestamp 1666464484
transform -1 0 21712 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _508_
timestamp 1666464484
transform -1 0 17296 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__o211ai_1  _509_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 17848 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__or3_2  _510_
timestamp 1666464484
transform 1 0 10028 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _511_
timestamp 1666464484
transform 1 0 11224 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _512_
timestamp 1666464484
transform 1 0 11684 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__and3_2  _513_
timestamp 1666464484
transform 1 0 12144 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _514_
timestamp 1666464484
transform -1 0 19688 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _515_
timestamp 1666464484
transform 1 0 19228 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_2  _516_
timestamp 1666464484
transform -1 0 13156 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _517_
timestamp 1666464484
transform -1 0 19044 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _518_
timestamp 1666464484
transform 1 0 19412 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _519_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 14812 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _520_
timestamp 1666464484
transform 1 0 14628 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _521_
timestamp 1666464484
transform 1 0 15364 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _522_
timestamp 1666464484
transform 1 0 14260 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _523_
timestamp 1666464484
transform -1 0 14812 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__or3_2  _524_
timestamp 1666464484
transform 1 0 14260 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _525_
timestamp 1666464484
transform 1 0 21712 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _526_
timestamp 1666464484
transform 1 0 19320 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _527_
timestamp 1666464484
transform -1 0 18860 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _528_
timestamp 1666464484
transform -1 0 19688 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_2  _529_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 14260 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__or4_4  _530_
timestamp 1666464484
transform 1 0 13156 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__and4_1  _531_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 20976 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _532_
timestamp 1666464484
transform -1 0 16376 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_4  _533_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 10764 0 1 10880
box -38 -48 2062 592
use sky130_fd_sc_hd__o311a_1  _534_
timestamp 1666464484
transform -1 0 16928 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _535_
timestamp 1666464484
transform -1 0 18032 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _536_
timestamp 1666464484
transform 1 0 22908 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_1  _537_
timestamp 1666464484
transform 1 0 21988 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__o311a_1  _538_
timestamp 1666464484
transform 1 0 20056 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _539_
timestamp 1666464484
transform 1 0 18400 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _540_
timestamp 1666464484
transform 1 0 21160 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _541_
timestamp 1666464484
transform -1 0 18952 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _542_
timestamp 1666464484
transform -1 0 20148 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _543_
timestamp 1666464484
transform 1 0 17848 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_2  _544_
timestamp 1666464484
transform -1 0 13800 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkinv_2  _545_
timestamp 1666464484
transform 1 0 17296 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__and4_1  _546_
timestamp 1666464484
transform 1 0 17112 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _547_
timestamp 1666464484
transform -1 0 18952 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _548_
timestamp 1666464484
transform -1 0 19596 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _549_
timestamp 1666464484
transform 1 0 13156 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _550_
timestamp 1666464484
transform 1 0 11684 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__a2111o_1  _551_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 12788 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _552_
timestamp 1666464484
transform -1 0 20608 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _553_
timestamp 1666464484
transform 1 0 20884 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _554_
timestamp 1666464484
transform -1 0 20424 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _555_
timestamp 1666464484
transform -1 0 20240 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _556_
timestamp 1666464484
transform 1 0 21252 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _557_
timestamp 1666464484
transform 1 0 20792 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _558_
timestamp 1666464484
transform 1 0 19504 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _559_
timestamp 1666464484
transform 1 0 20424 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _560_
timestamp 1666464484
transform 1 0 20240 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _561_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 19780 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _562_
timestamp 1666464484
transform -1 0 12880 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _563_
timestamp 1666464484
transform 1 0 12788 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_4  _564_
timestamp 1666464484
transform -1 0 12328 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _565_
timestamp 1666464484
transform 1 0 18124 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _566_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 18216 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _567_
timestamp 1666464484
transform -1 0 20700 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _568_
timestamp 1666464484
transform 1 0 12236 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _569_
timestamp 1666464484
transform -1 0 22264 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _570_
timestamp 1666464484
transform 1 0 20516 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _571_
timestamp 1666464484
transform 1 0 19780 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _572_
timestamp 1666464484
transform 1 0 21436 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _573_
timestamp 1666464484
transform -1 0 22540 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _574_
timestamp 1666464484
transform -1 0 23092 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _575_
timestamp 1666464484
transform -1 0 22540 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _576_
timestamp 1666464484
transform 1 0 21988 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _577_
timestamp 1666464484
transform -1 0 13800 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__o32a_1  _578_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 15456 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__a311o_1  _579_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 17480 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _580_
timestamp 1666464484
transform 1 0 14352 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _581_
timestamp 1666464484
transform 1 0 14260 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _582_
timestamp 1666464484
transform 1 0 13432 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _583_
timestamp 1666464484
transform -1 0 13800 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _584_
timestamp 1666464484
transform 1 0 12972 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _585_
timestamp 1666464484
transform 1 0 16836 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _586_
timestamp 1666464484
transform 1 0 15180 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__o211ai_1  _587_
timestamp 1666464484
transform -1 0 14812 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _588_
timestamp 1666464484
transform -1 0 15916 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _589_
timestamp 1666464484
transform 1 0 20516 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _590_
timestamp 1666464484
transform 1 0 20148 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _591_
timestamp 1666464484
transform 1 0 20332 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _592_
timestamp 1666464484
transform -1 0 20424 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a22oi_1  _593_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 14076 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _594_
timestamp 1666464484
transform -1 0 14904 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _595_
timestamp 1666464484
transform 1 0 15364 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__a211oi_1  _596_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 18952 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _597_
timestamp 1666464484
transform 1 0 16928 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _598_
timestamp 1666464484
transform -1 0 13340 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _599_
timestamp 1666464484
transform 1 0 15916 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _600_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 15456 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _601_
timestamp 1666464484
transform 1 0 15732 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _602_
timestamp 1666464484
transform -1 0 17480 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _603_
timestamp 1666464484
transform 1 0 17388 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _604_
timestamp 1666464484
transform 1 0 16376 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _605_
timestamp 1666464484
transform -1 0 18860 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _606_
timestamp 1666464484
transform 1 0 19412 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _607_
timestamp 1666464484
transform -1 0 16744 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nor4_1  _608_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 20792 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _609_
timestamp 1666464484
transform 1 0 16836 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _610_
timestamp 1666464484
transform -1 0 18584 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__o32a_1  _611_
timestamp 1666464484
transform 1 0 18216 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _612_
timestamp 1666464484
transform 1 0 19780 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _613_
timestamp 1666464484
transform -1 0 22908 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _614_
timestamp 1666464484
transform 1 0 19412 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _615_
timestamp 1666464484
transform 1 0 19412 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _616_
timestamp 1666464484
transform 1 0 17756 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _617_
timestamp 1666464484
transform 1 0 15456 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _618_
timestamp 1666464484
transform -1 0 15824 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _619_
timestamp 1666464484
transform 1 0 14812 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a21boi_1  _620_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 12788 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _621_
timestamp 1666464484
transform 1 0 15272 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _622_
timestamp 1666464484
transform 1 0 11684 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _623_
timestamp 1666464484
transform -1 0 13340 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _624_
timestamp 1666464484
transform 1 0 12880 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _625_
timestamp 1666464484
transform 1 0 11776 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _626_
timestamp 1666464484
transform -1 0 20056 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_1  _627_
timestamp 1666464484
transform 1 0 20516 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _628_
timestamp 1666464484
transform -1 0 18584 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _629_
timestamp 1666464484
transform -1 0 18952 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _630_
timestamp 1666464484
transform 1 0 15364 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _631_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 13524 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__a2111o_1  _632_
timestamp 1666464484
transform 1 0 18124 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__a31o_1  _633_
timestamp 1666464484
transform 1 0 12420 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _634_
timestamp 1666464484
transform 1 0 11224 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _635_
timestamp 1666464484
transform -1 0 17112 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _636_
timestamp 1666464484
transform -1 0 11040 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _637_
timestamp 1666464484
transform -1 0 12052 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _638_
timestamp 1666464484
transform -1 0 14904 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _639_
timestamp 1666464484
transform 1 0 12420 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _640_
timestamp 1666464484
transform 1 0 12236 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _641_
timestamp 1666464484
transform 1 0 12512 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__o2111a_1  _642_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 12696 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__nor3_1  _643_
timestamp 1666464484
transform -1 0 11224 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _644_
timestamp 1666464484
transform -1 0 12328 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _645_
timestamp 1666464484
transform 1 0 14168 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _646_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 14628 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _647_
timestamp 1666464484
transform -1 0 13984 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _648_
timestamp 1666464484
transform 1 0 13156 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _649_
timestamp 1666464484
transform -1 0 16376 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__o32a_1  _650_
timestamp 1666464484
transform 1 0 14260 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _651_
timestamp 1666464484
transform 1 0 12696 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _652_
timestamp 1666464484
transform -1 0 12328 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _653_
timestamp 1666464484
transform 1 0 20332 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _654_
timestamp 1666464484
transform 1 0 14812 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_1  _655_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 14260 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _656_
timestamp 1666464484
transform 1 0 14444 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _657_
timestamp 1666464484
transform -1 0 14076 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _658_
timestamp 1666464484
transform 1 0 16284 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__o311a_1  _659_
timestamp 1666464484
transform 1 0 15456 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__a2111o_1  _660_
timestamp 1666464484
transform -1 0 16192 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_1  _661_
timestamp 1666464484
transform -1 0 18308 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _662_
timestamp 1666464484
transform 1 0 15824 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _663_
timestamp 1666464484
transform -1 0 15916 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _664_
timestamp 1666464484
transform 1 0 14260 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _665_
timestamp 1666464484
transform 1 0 17572 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _666_
timestamp 1666464484
transform -1 0 21896 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _667_
timestamp 1666464484
transform 1 0 19412 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_1  _668_
timestamp 1666464484
transform 1 0 18216 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _669_
timestamp 1666464484
transform 1 0 18216 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _670_
timestamp 1666464484
transform 1 0 18308 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _671_
timestamp 1666464484
transform 1 0 17848 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _672_
timestamp 1666464484
transform -1 0 16376 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _673_
timestamp 1666464484
transform 1 0 16744 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _674_
timestamp 1666464484
transform -1 0 16560 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_1  _675_
timestamp 1666464484
transform 1 0 16836 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _676_
timestamp 1666464484
transform 1 0 16836 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _677_
timestamp 1666464484
transform 1 0 16560 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _678_
timestamp 1666464484
transform 1 0 16836 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _679_
timestamp 1666464484
transform 1 0 16560 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _680_
timestamp 1666464484
transform 1 0 16100 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _681_
timestamp 1666464484
transform 1 0 14260 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _682_
timestamp 1666464484
transform 1 0 12880 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _683_
timestamp 1666464484
transform -1 0 14904 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _684_
timestamp 1666464484
transform -1 0 13616 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _685_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 14260 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__nor3_2  _686_
timestamp 1666464484
transform 1 0 2576 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_2  _687_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 10396 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _688_
timestamp 1666464484
transform 1 0 4692 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _689_
timestamp 1666464484
transform -1 0 7728 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _690_
timestamp 1666464484
transform -1 0 5152 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _691_
timestamp 1666464484
transform -1 0 3588 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_2  _692_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 3956 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _693_
timestamp 1666464484
transform 1 0 2668 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _694_
timestamp 1666464484
transform 1 0 5520 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__a2bb2o_1  _695_
timestamp 1666464484
transform -1 0 6716 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__or2b_2  _696_
timestamp 1666464484
transform 1 0 10212 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _697_
timestamp 1666464484
transform 1 0 6532 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _698_
timestamp 1666464484
transform 1 0 6164 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _699_
timestamp 1666464484
transform 1 0 8188 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _700_
timestamp 1666464484
transform -1 0 8280 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _701_
timestamp 1666464484
transform 1 0 4324 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _702_
timestamp 1666464484
transform 1 0 6808 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _703_
timestamp 1666464484
transform -1 0 7360 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_1  _704_
timestamp 1666464484
transform 1 0 5704 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__a21bo_1  _705_
timestamp 1666464484
transform 1 0 5980 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _706_
timestamp 1666464484
transform 1 0 6072 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _707_
timestamp 1666464484
transform -1 0 7912 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _708_
timestamp 1666464484
transform -1 0 10120 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _709_
timestamp 1666464484
transform -1 0 8464 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _710_
timestamp 1666464484
transform 1 0 9108 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _711_
timestamp 1666464484
transform -1 0 6992 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _712_
timestamp 1666464484
transform 1 0 3956 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _713_
timestamp 1666464484
transform 1 0 3956 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _714_
timestamp 1666464484
transform 1 0 3772 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__nor3_1  _715_
timestamp 1666464484
transform 1 0 5060 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _716_
timestamp 1666464484
transform 1 0 4968 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _717_
timestamp 1666464484
transform -1 0 6072 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _718_
timestamp 1666464484
transform -1 0 10396 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _719_
timestamp 1666464484
transform 1 0 6164 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _720_
timestamp 1666464484
transform 1 0 8464 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _721_
timestamp 1666464484
transform 1 0 10396 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _722_
timestamp 1666464484
transform -1 0 5612 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _723_
timestamp 1666464484
transform 1 0 10304 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _724_
timestamp 1666464484
transform 1 0 9108 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__o2111a_1  _725_
timestamp 1666464484
transform 1 0 9108 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _726_
timestamp 1666464484
transform 1 0 7636 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_1  _727_
timestamp 1666464484
transform -1 0 7268 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _728_
timestamp 1666464484
transform -1 0 7452 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _729_
timestamp 1666464484
transform 1 0 9476 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _730_
timestamp 1666464484
transform -1 0 9384 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__or4b_1  _731_
timestamp 1666464484
transform 1 0 5336 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _732_
timestamp 1666464484
transform 1 0 5796 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _733_
timestamp 1666464484
transform -1 0 7268 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _734_
timestamp 1666464484
transform -1 0 8556 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _735_
timestamp 1666464484
transform -1 0 7084 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _736_
timestamp 1666464484
transform 1 0 11592 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _737_
timestamp 1666464484
transform -1 0 8096 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _738_
timestamp 1666464484
transform 1 0 9568 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _739_
timestamp 1666464484
transform -1 0 9752 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _740_
timestamp 1666464484
transform 1 0 3036 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__a21boi_1  _741_
timestamp 1666464484
transform 1 0 3956 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__a41o_1  _742_
timestamp 1666464484
transform -1 0 5888 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_1  _743_
timestamp 1666464484
transform 1 0 4048 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _744_
timestamp 1666464484
transform 1 0 7728 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _745_
timestamp 1666464484
transform 1 0 8464 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _746_
timestamp 1666464484
transform 1 0 8188 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nand3b_1  _747_
timestamp 1666464484
transform 1 0 5796 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _748_
timestamp 1666464484
transform -1 0 4876 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _749_
timestamp 1666464484
transform 1 0 3956 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _750_
timestamp 1666464484
transform -1 0 5796 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _751_
timestamp 1666464484
transform -1 0 6900 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _752_
timestamp 1666464484
transform 1 0 9108 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _753_
timestamp 1666464484
transform 1 0 9108 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _754_
timestamp 1666464484
transform 1 0 9844 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _755_
timestamp 1666464484
transform 1 0 9108 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _756_
timestamp 1666464484
transform 1 0 3220 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__o21bai_1  _757_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 5244 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _758_
timestamp 1666464484
transform -1 0 9568 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _759_
timestamp 1666464484
transform -1 0 2208 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__o41a_1  _760_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 4968 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__a21bo_1  _761_
timestamp 1666464484
transform 1 0 7084 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _762_
timestamp 1666464484
transform 1 0 7176 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _763_
timestamp 1666464484
transform 1 0 9752 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _764_
timestamp 1666464484
transform 1 0 9108 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _765_
timestamp 1666464484
transform -1 0 9108 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _766_
timestamp 1666464484
transform 1 0 9108 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__or2b_1  _767_
timestamp 1666464484
transform 1 0 5060 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _768_
timestamp 1666464484
transform -1 0 7176 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _769_
timestamp 1666464484
transform 1 0 7268 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _770_
timestamp 1666464484
transform 1 0 7452 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _771_
timestamp 1666464484
transform -1 0 3680 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _772_
timestamp 1666464484
transform -1 0 3036 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _773_
timestamp 1666464484
transform 1 0 6900 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _774_
timestamp 1666464484
transform 1 0 9108 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_1  _775_
timestamp 1666464484
transform 1 0 7820 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _776_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 7820 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _777_
timestamp 1666464484
transform -1 0 8464 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _778_
timestamp 1666464484
transform 1 0 9108 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _779_
timestamp 1666464484
transform -1 0 8556 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _780_
timestamp 1666464484
transform 1 0 5796 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _781_
timestamp 1666464484
transform 1 0 5796 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _782_
timestamp 1666464484
transform -1 0 5520 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _783_
timestamp 1666464484
transform 1 0 7912 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _784_
timestamp 1666464484
transform 1 0 6624 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a41o_1  _785_
timestamp 1666464484
transform 1 0 4784 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _786_
timestamp 1666464484
transform -1 0 4968 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a31oi_1  _787_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 2484 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _788_
timestamp 1666464484
transform 1 0 2668 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _789_
timestamp 1666464484
transform -1 0 4140 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _790_
timestamp 1666464484
transform 1 0 3128 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _791_
timestamp 1666464484
transform 1 0 2300 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _792_
timestamp 1666464484
transform 1 0 1840 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _793_
timestamp 1666464484
transform 1 0 3312 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _794_
timestamp 1666464484
transform 1 0 2392 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _795_
timestamp 1666464484
transform 1 0 1748 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _796_
timestamp 1666464484
transform -1 0 5428 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _797_
timestamp 1666464484
transform 1 0 2484 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _798_
timestamp 1666464484
transform 1 0 4048 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _799_
timestamp 1666464484
transform 1 0 1564 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _800_
timestamp 1666464484
transform 1 0 1656 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _801_
timestamp 1666464484
transform -1 0 2576 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _802_
timestamp 1666464484
transform 1 0 2484 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _803_
timestamp 1666464484
transform 1 0 2484 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _804_
timestamp 1666464484
transform -1 0 7912 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__o221ai_1  _805_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 7820 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _806_
timestamp 1666464484
transform 1 0 7360 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__a32o_1  _807_
timestamp 1666464484
transform 1 0 6900 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _808_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 6348 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _809_
timestamp 1666464484
transform -1 0 8372 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _810_
timestamp 1666464484
transform -1 0 8280 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _811_
timestamp 1666464484
transform -1 0 6440 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _812_
timestamp 1666464484
transform -1 0 8096 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _813_
timestamp 1666464484
transform -1 0 13156 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _814_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 6808 0 1 18496
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _815_
timestamp 1666464484
transform 1 0 6992 0 -1 17408
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _816_
timestamp 1666464484
transform 1 0 9752 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _817_
timestamp 1666464484
transform 1 0 11684 0 1 17408
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _818_
timestamp 1666464484
transform -1 0 11316 0 1 17408
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_4  _819_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 11776 0 1 18496
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_1  _820_
timestamp 1666464484
transform -1 0 11224 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _821_
timestamp 1666464484
transform 1 0 9752 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _822_
timestamp 1666464484
transform 1 0 9752 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _823_
timestamp 1666464484
transform -1 0 5152 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _824_
timestamp 1666464484
transform 1 0 4600 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _825_
timestamp 1666464484
transform -1 0 13064 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _826_
timestamp 1666464484
transform -1 0 13156 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _827_
timestamp 1666464484
transform 1 0 9752 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _828_
timestamp 1666464484
transform 1 0 7084 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _829_
timestamp 1666464484
transform -1 0 11224 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _830_
timestamp 1666464484
transform -1 0 11224 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _831_
timestamp 1666464484
transform 1 0 10028 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _832_
timestamp 1666464484
transform -1 0 5704 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _833_
timestamp 1666464484
transform 1 0 7176 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _834_
timestamp 1666464484
transform -1 0 4968 0 -1 18496
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _835_
timestamp 1666464484
transform -1 0 3588 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _836_
timestamp 1666464484
transform 1 0 3956 0 -1 17408
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _837_
timestamp 1666464484
transform -1 0 5428 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _838_
timestamp 1666464484
transform 1 0 3956 0 1 19584
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _839_
timestamp 1666464484
transform 1 0 2024 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _840_
timestamp 1666464484
transform 1 0 6716 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  _868_
timestamp 1666464484
transform 1 0 3220 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 7636 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_0__f_clk
timestamp 1666464484
transform -1 0 4416 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_1__f_clk
timestamp 1666464484
transform -1 0 7084 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_2__f_clk
timestamp 1666464484
transform -1 0 9660 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_3__f_clk
timestamp 1666464484
transform 1 0 10396 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1666464484
transform -1 0 13800 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1666464484
transform 1 0 17480 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1666464484
transform 1 0 22448 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input4
timestamp 1666464484
transform -1 0 7912 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output5
timestamp 1666464484
transform -1 0 1932 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output6
timestamp 1666464484
transform -1 0 2576 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output7
timestamp 1666464484
transform -1 0 2760 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output8
timestamp 1666464484
transform -1 0 3496 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output9
timestamp 1666464484
transform -1 0 4324 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output10
timestamp 1666464484
transform -1 0 5060 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output11
timestamp 1666464484
transform -1 0 5796 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output12
timestamp 1666464484
transform -1 0 6900 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  tt2_tholin_namebadge_13 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 3312 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt2_tholin_namebadge_14
timestamp 1666464484
transform 1 0 3956 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt2_tholin_namebadge_15
timestamp 1666464484
transform 1 0 4600 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt2_tholin_namebadge_16
timestamp 1666464484
transform 1 0 5336 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt2_tholin_namebadge_17
timestamp 1666464484
transform -1 0 13432 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt2_tholin_namebadge_18
timestamp 1666464484
transform -1 0 12788 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt2_tholin_namebadge_19
timestamp 1666464484
transform 1 0 8372 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt2_tholin_namebadge_20
timestamp 1666464484
transform 1 0 10304 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt2_tholin_namebadge_21
timestamp 1666464484
transform 1 0 10948 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt2_tholin_namebadge_22
timestamp 1666464484
transform -1 0 12788 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt2_tholin_namebadge_23
timestamp 1666464484
transform -1 0 13432 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt2_tholin_namebadge_24
timestamp 1666464484
transform -1 0 14536 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt2_tholin_namebadge_25
timestamp 1666464484
transform -1 0 15180 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt2_tholin_namebadge_26
timestamp 1666464484
transform -1 0 15824 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt2_tholin_namebadge_27
timestamp 1666464484
transform -1 0 16008 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt2_tholin_namebadge_28
timestamp 1666464484
transform -1 0 17112 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt2_tholin_namebadge_29
timestamp 1666464484
transform -1 0 17756 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt2_tholin_namebadge_30
timestamp 1666464484
transform -1 0 18400 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt2_tholin_namebadge_31
timestamp 1666464484
transform -1 0 18584 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt2_tholin_namebadge_32
timestamp 1666464484
transform -1 0 19688 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt2_tholin_namebadge_33
timestamp 1666464484
transform -1 0 20332 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt2_tholin_namebadge_34
timestamp 1666464484
transform -1 0 20976 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt2_tholin_namebadge_35
timestamp 1666464484
transform -1 0 21160 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt2_tholin_namebadge_36
timestamp 1666464484
transform -1 0 22264 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt2_tholin_namebadge_37
timestamp 1666464484
transform -1 0 22908 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt2_tholin_namebadge_38
timestamp 1666464484
transform -1 0 23092 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt2_tholin_namebadge_39
timestamp 1666464484
transform 1 0 23092 0 1 3264
box -38 -48 314 592
<< labels >>
flabel metal2 s 2502 24200 2558 25000 0 FreeSans 224 90 0 0 clk
port 0 nsew signal input
flabel metal2 s 12438 24200 12494 25000 0 FreeSans 224 90 0 0 io_in[0]
port 1 nsew signal input
flabel metal2 s 17406 24200 17462 25000 0 FreeSans 224 90 0 0 io_in[1]
port 2 nsew signal input
flabel metal2 s 22374 24200 22430 25000 0 FreeSans 224 90 0 0 io_in[2]
port 3 nsew signal input
flabel metal2 s 6642 0 6698 800 0 FreeSans 224 90 0 0 io_oeb[0]
port 4 nsew signal tristate
flabel metal2 s 13082 0 13138 800 0 FreeSans 224 90 0 0 io_oeb[10]
port 5 nsew signal tristate
flabel metal2 s 13726 0 13782 800 0 FreeSans 224 90 0 0 io_oeb[11]
port 6 nsew signal tristate
flabel metal2 s 14370 0 14426 800 0 FreeSans 224 90 0 0 io_oeb[12]
port 7 nsew signal tristate
flabel metal2 s 15014 0 15070 800 0 FreeSans 224 90 0 0 io_oeb[13]
port 8 nsew signal tristate
flabel metal2 s 15658 0 15714 800 0 FreeSans 224 90 0 0 io_oeb[14]
port 9 nsew signal tristate
flabel metal2 s 16302 0 16358 800 0 FreeSans 224 90 0 0 io_oeb[15]
port 10 nsew signal tristate
flabel metal2 s 16946 0 17002 800 0 FreeSans 224 90 0 0 io_oeb[16]
port 11 nsew signal tristate
flabel metal2 s 17590 0 17646 800 0 FreeSans 224 90 0 0 io_oeb[17]
port 12 nsew signal tristate
flabel metal2 s 18234 0 18290 800 0 FreeSans 224 90 0 0 io_oeb[18]
port 13 nsew signal tristate
flabel metal2 s 18878 0 18934 800 0 FreeSans 224 90 0 0 io_oeb[19]
port 14 nsew signal tristate
flabel metal2 s 7286 0 7342 800 0 FreeSans 224 90 0 0 io_oeb[1]
port 15 nsew signal tristate
flabel metal2 s 19522 0 19578 800 0 FreeSans 224 90 0 0 io_oeb[20]
port 16 nsew signal tristate
flabel metal2 s 20166 0 20222 800 0 FreeSans 224 90 0 0 io_oeb[21]
port 17 nsew signal tristate
flabel metal2 s 20810 0 20866 800 0 FreeSans 224 90 0 0 io_oeb[22]
port 18 nsew signal tristate
flabel metal2 s 21454 0 21510 800 0 FreeSans 224 90 0 0 io_oeb[23]
port 19 nsew signal tristate
flabel metal2 s 22098 0 22154 800 0 FreeSans 224 90 0 0 io_oeb[24]
port 20 nsew signal tristate
flabel metal2 s 22742 0 22798 800 0 FreeSans 224 90 0 0 io_oeb[25]
port 21 nsew signal tristate
flabel metal2 s 23386 0 23442 800 0 FreeSans 224 90 0 0 io_oeb[26]
port 22 nsew signal tristate
flabel metal2 s 7930 0 7986 800 0 FreeSans 224 90 0 0 io_oeb[2]
port 23 nsew signal tristate
flabel metal2 s 8574 0 8630 800 0 FreeSans 224 90 0 0 io_oeb[3]
port 24 nsew signal tristate
flabel metal2 s 9218 0 9274 800 0 FreeSans 224 90 0 0 io_oeb[4]
port 25 nsew signal tristate
flabel metal2 s 9862 0 9918 800 0 FreeSans 224 90 0 0 io_oeb[5]
port 26 nsew signal tristate
flabel metal2 s 10506 0 10562 800 0 FreeSans 224 90 0 0 io_oeb[6]
port 27 nsew signal tristate
flabel metal2 s 11150 0 11206 800 0 FreeSans 224 90 0 0 io_oeb[7]
port 28 nsew signal tristate
flabel metal2 s 11794 0 11850 800 0 FreeSans 224 90 0 0 io_oeb[8]
port 29 nsew signal tristate
flabel metal2 s 12438 0 12494 800 0 FreeSans 224 90 0 0 io_oeb[9]
port 30 nsew signal tristate
flabel metal2 s 1490 0 1546 800 0 FreeSans 224 90 0 0 io_out[0]
port 31 nsew signal tristate
flabel metal2 s 2134 0 2190 800 0 FreeSans 224 90 0 0 io_out[1]
port 32 nsew signal tristate
flabel metal2 s 2778 0 2834 800 0 FreeSans 224 90 0 0 io_out[2]
port 33 nsew signal tristate
flabel metal2 s 3422 0 3478 800 0 FreeSans 224 90 0 0 io_out[3]
port 34 nsew signal tristate
flabel metal2 s 4066 0 4122 800 0 FreeSans 224 90 0 0 io_out[4]
port 35 nsew signal tristate
flabel metal2 s 4710 0 4766 800 0 FreeSans 224 90 0 0 io_out[5]
port 36 nsew signal tristate
flabel metal2 s 5354 0 5410 800 0 FreeSans 224 90 0 0 io_out[6]
port 37 nsew signal tristate
flabel metal2 s 5998 0 6054 800 0 FreeSans 224 90 0 0 io_out[7]
port 38 nsew signal tristate
flabel metal2 s 7470 24200 7526 25000 0 FreeSans 224 90 0 0 rst
port 39 nsew signal input
flabel metal4 s 3784 2128 4104 22352 0 FreeSans 1920 90 0 0 vccd1
port 40 nsew power bidirectional
flabel metal4 s 9465 2128 9785 22352 0 FreeSans 1920 90 0 0 vccd1
port 40 nsew power bidirectional
flabel metal4 s 15146 2128 15466 22352 0 FreeSans 1920 90 0 0 vccd1
port 40 nsew power bidirectional
flabel metal4 s 20827 2128 21147 22352 0 FreeSans 1920 90 0 0 vccd1
port 40 nsew power bidirectional
flabel metal4 s 6624 2128 6944 22352 0 FreeSans 1920 90 0 0 vssd1
port 41 nsew ground bidirectional
flabel metal4 s 12305 2128 12625 22352 0 FreeSans 1920 90 0 0 vssd1
port 41 nsew ground bidirectional
flabel metal4 s 17986 2128 18306 22352 0 FreeSans 1920 90 0 0 vssd1
port 41 nsew ground bidirectional
flabel metal4 s 23667 2128 23987 22352 0 FreeSans 1920 90 0 0 vssd1
port 41 nsew ground bidirectional
rlabel metal1 12466 22304 12466 22304 0 vccd1
rlabel via1 12545 21760 12545 21760 0 vssd1
rlabel metal1 18308 18938 18308 18938 0 _000_
rlabel metal1 13800 14790 13800 14790 0 _001_
rlabel metal1 10115 21930 10115 21930 0 _002_
rlabel via3 7429 18020 7429 18020 0 _003_
rlabel metal1 10948 19686 10948 19686 0 _004_
rlabel metal1 14306 15368 14306 15368 0 _005_
rlabel metal1 14283 16422 14283 16422 0 _006_
rlabel metal1 7176 13906 7176 13906 0 _007_
rlabel metal1 13217 21590 13217 21590 0 _008_
rlabel metal2 9338 21284 9338 21284 0 _009_
rlabel metal1 6133 20842 6133 20842 0 _010_
rlabel metal2 7958 14178 7958 14178 0 _011_
rlabel metal1 8234 19720 8234 19720 0 _012_
rlabel via1 6122 18666 6122 18666 0 _013_
rlabel metal1 8137 18666 8137 18666 0 _014_
rlabel metal1 7866 15130 7866 15130 0 _015_
rlabel metal1 19826 11798 19826 11798 0 _016_
rlabel metal1 13064 13430 13064 13430 0 _017_
rlabel metal1 14168 13838 14168 13838 0 _018_
rlabel via1 22103 12614 22103 12614 0 _019_
rlabel metal1 11837 20502 11837 20502 0 _020_
rlabel metal1 20838 8262 20838 8262 0 _021_
rlabel via2 21022 10948 21022 10948 0 _022_
rlabel metal2 5934 17816 5934 17816 0 _023_
rlabel metal2 4922 17238 4922 17238 0 _024_
rlabel metal1 7268 14042 7268 14042 0 _025_
rlabel metal2 4370 16694 4370 16694 0 _026_
rlabel metal1 3404 12954 3404 12954 0 _027_
rlabel metal1 4094 15130 4094 15130 0 _028_
rlabel metal1 4972 15402 4972 15402 0 _029_
rlabel metal2 4278 19346 4278 19346 0 _030_
rlabel metal2 2530 17170 2530 17170 0 _031_
rlabel metal1 7355 20842 7355 20842 0 _032_
rlabel metal1 3312 15538 3312 15538 0 _033_
rlabel metal1 10258 7412 10258 7412 0 _034_
rlabel metal1 8832 12750 8832 12750 0 _035_
rlabel metal1 5290 7514 5290 7514 0 _036_
rlabel metal1 6302 7888 6302 7888 0 _037_
rlabel metal1 3450 8058 3450 8058 0 _038_
rlabel viali 6427 8908 6427 8908 0 _039_
rlabel metal1 9338 8976 9338 8976 0 _040_
rlabel metal2 2438 14144 2438 14144 0 _041_
rlabel metal2 7268 13260 7268 13260 0 _042_
rlabel metal2 9982 6460 9982 6460 0 _043_
rlabel metal1 5474 6426 5474 6426 0 _044_
rlabel metal1 4416 4114 4416 4114 0 _045_
rlabel metal2 2898 8500 2898 8500 0 _046_
rlabel metal2 2070 8772 2070 8772 0 _047_
rlabel metal1 5106 5712 5106 5712 0 _048_
rlabel metal1 6026 9486 6026 9486 0 _049_
rlabel metal1 5014 6086 5014 6086 0 _050_
rlabel metal1 6762 4658 6762 4658 0 _051_
rlabel metal1 2714 13396 2714 13396 0 _052_
rlabel metal1 4738 5236 4738 5236 0 _053_
rlabel metal2 6302 5508 6302 5508 0 _054_
rlabel metal1 9338 4114 9338 4114 0 _055_
rlabel metal1 2576 5542 2576 5542 0 _056_
rlabel metal1 2116 4590 2116 4590 0 _057_
rlabel metal1 4278 4454 4278 4454 0 _058_
rlabel metal1 8694 2992 8694 2992 0 _059_
rlabel metal1 2622 3536 2622 3536 0 _060_
rlabel metal2 2714 3145 2714 3145 0 _061_
rlabel metal2 9154 3332 9154 3332 0 _062_
rlabel metal2 10902 5644 10902 5644 0 _063_
rlabel metal1 7590 4658 7590 4658 0 _064_
rlabel metal1 11148 5270 11148 5270 0 _065_
rlabel metal1 12029 6154 12029 6154 0 _066_
rlabel metal1 13386 15504 13386 15504 0 _067_
rlabel metal1 10672 7854 10672 7854 0 _068_
rlabel metal1 10396 4046 10396 4046 0 _069_
rlabel metal1 6992 14790 6992 14790 0 _070_
rlabel metal1 11316 3162 11316 3162 0 _071_
rlabel metal1 11960 5202 11960 5202 0 _072_
rlabel metal1 11040 6222 11040 6222 0 _073_
rlabel metal2 11178 7174 11178 7174 0 _074_
rlabel metal1 11040 14382 11040 14382 0 _075_
rlabel metal1 18492 7174 18492 7174 0 _076_
rlabel metal1 21298 6698 21298 6698 0 _077_
rlabel metal1 21758 11084 21758 11084 0 _078_
rlabel metal1 7130 9588 7130 9588 0 _079_
rlabel metal2 12742 4930 12742 4930 0 _080_
rlabel metal2 14674 5542 14674 5542 0 _081_
rlabel metal1 12098 4182 12098 4182 0 _082_
rlabel metal2 13662 4522 13662 4522 0 _083_
rlabel metal1 17066 6256 17066 6256 0 _084_
rlabel metal2 13110 6256 13110 6256 0 _085_
rlabel metal1 11730 7854 11730 7854 0 _086_
rlabel metal1 14263 8466 14263 8466 0 _087_
rlabel metal1 21160 7446 21160 7446 0 _088_
rlabel metal2 13478 5032 13478 5032 0 _089_
rlabel via1 17434 6764 17434 6764 0 _090_
rlabel metal1 17641 13294 17641 13294 0 _091_
rlabel metal1 16008 4522 16008 4522 0 _092_
rlabel metal1 15318 4658 15318 4658 0 _093_
rlabel metal1 10488 4726 10488 4726 0 _094_
rlabel metal2 15042 4080 15042 4080 0 _095_
rlabel metal2 16882 4998 16882 4998 0 _096_
rlabel metal2 13938 5542 13938 5542 0 _097_
rlabel metal1 12834 5168 12834 5168 0 _098_
rlabel metal1 18032 14042 18032 14042 0 _099_
rlabel metal1 18078 9894 18078 9894 0 _100_
rlabel metal1 12880 10438 12880 10438 0 _101_
rlabel metal1 11316 14790 11316 14790 0 _102_
rlabel metal1 12006 13498 12006 13498 0 _103_
rlabel metal2 21666 13804 21666 13804 0 _104_
rlabel metal1 20102 13328 20102 13328 0 _105_
rlabel metal1 17250 12716 17250 12716 0 _106_
rlabel metal1 18124 11730 18124 11730 0 _107_
rlabel metal1 11730 7344 11730 7344 0 _108_
rlabel metal2 12834 14790 12834 14790 0 _109_
rlabel metal2 12374 14552 12374 14552 0 _110_
rlabel metal1 15962 13294 15962 13294 0 _111_
rlabel metal1 19596 14246 19596 14246 0 _112_
rlabel metal1 14168 12682 14168 12682 0 _113_
rlabel metal1 16514 6936 16514 6936 0 _114_
rlabel metal1 17135 10030 17135 10030 0 _115_
rlabel metal1 15272 5338 15272 5338 0 _116_
rlabel metal2 19872 7956 19872 7956 0 _117_
rlabel metal2 14674 10438 14674 10438 0 _118_
rlabel metal1 19642 10064 19642 10064 0 _119_
rlabel metal1 14996 8398 14996 8398 0 _120_
rlabel metal1 20148 10642 20148 10642 0 _121_
rlabel metal1 18676 10030 18676 10030 0 _122_
rlabel metal1 18722 10234 18722 10234 0 _123_
rlabel metal2 19642 10914 19642 10914 0 _124_
rlabel metal1 21114 6800 21114 6800 0 _125_
rlabel metal3 20194 12852 20194 12852 0 _126_
rlabel metal1 20424 10778 20424 10778 0 _127_
rlabel metal1 15594 7854 15594 7854 0 _128_
rlabel metal2 12650 8534 12650 8534 0 _129_
rlabel metal1 21988 7378 21988 7378 0 _130_
rlabel metal1 18446 6834 18446 6834 0 _131_
rlabel metal2 22586 7820 22586 7820 0 _132_
rlabel metal1 21988 7514 21988 7514 0 _133_
rlabel metal1 19504 11662 19504 11662 0 _134_
rlabel metal1 18492 11866 18492 11866 0 _135_
rlabel metal2 16284 9316 16284 9316 0 _136_
rlabel metal1 19826 13192 19826 13192 0 _137_
rlabel metal2 19458 13702 19458 13702 0 _138_
rlabel metal1 18584 8466 18584 8466 0 _139_
rlabel metal1 13248 5814 13248 5814 0 _140_
rlabel metal1 18078 10234 18078 10234 0 _141_
rlabel metal1 19136 10778 19136 10778 0 _142_
rlabel metal1 19274 12954 19274 12954 0 _143_
rlabel metal1 12190 4556 12190 4556 0 _144_
rlabel metal2 12098 3910 12098 3910 0 _145_
rlabel metal2 14582 5916 14582 5916 0 _146_
rlabel metal2 20700 7956 20700 7956 0 _147_
rlabel metal1 21298 12614 21298 12614 0 _148_
rlabel metal2 20378 7276 20378 7276 0 _149_
rlabel metal1 19918 7514 19918 7514 0 _150_
rlabel metal1 21022 7922 21022 7922 0 _151_
rlabel metal1 20792 6834 20792 6834 0 _152_
rlabel metal1 20056 9622 20056 9622 0 _153_
rlabel metal2 20562 8330 20562 8330 0 _154_
rlabel metal3 19849 13804 19849 13804 0 _155_
rlabel metal2 19182 14144 19182 14144 0 _156_
rlabel metal1 13018 15130 13018 15130 0 _157_
rlabel metal2 12834 15878 12834 15878 0 _158_
rlabel metal1 18308 14586 18308 14586 0 _159_
rlabel metal1 20102 13906 20102 13906 0 _160_
rlabel metal2 14398 14586 14398 14586 0 _161_
rlabel metal1 15134 12852 15134 12852 0 _162_
rlabel metal1 21620 9554 21620 9554 0 _163_
rlabel metal1 20378 12818 20378 12818 0 _164_
rlabel metal2 21666 8636 21666 8636 0 _165_
rlabel metal1 22172 9554 22172 9554 0 _166_
rlabel metal2 14674 9486 14674 9486 0 _167_
rlabel metal2 22494 9044 22494 9044 0 _168_
rlabel metal2 14582 8993 14582 8993 0 _169_
rlabel metal1 13938 8602 13938 8602 0 _170_
rlabel metal1 14766 9520 14766 9520 0 _171_
rlabel metal1 14858 9588 14858 9588 0 _172_
rlabel metal2 14766 9180 14766 9180 0 _173_
rlabel metal1 13938 14858 13938 14858 0 _174_
rlabel metal1 14168 14450 14168 14450 0 _175_
rlabel metal1 16008 13838 16008 13838 0 _176_
rlabel metal1 14858 14042 14858 14042 0 _177_
rlabel metal2 13846 14790 13846 14790 0 _178_
rlabel metal2 20562 12954 20562 12954 0 _179_
rlabel metal2 19734 11271 19734 11271 0 _180_
rlabel metal1 20792 9418 20792 9418 0 _181_
rlabel metal2 20378 12614 20378 12614 0 _182_
rlabel metal1 19780 14042 19780 14042 0 _183_
rlabel via1 15433 7786 15433 7786 0 _184_
rlabel metal2 16698 9588 16698 9588 0 _185_
rlabel metal2 18446 7582 18446 7582 0 _186_
rlabel metal1 16790 8602 16790 8602 0 _187_
rlabel metal1 16108 8602 16108 8602 0 _188_
rlabel metal1 16422 8602 16422 8602 0 _189_
rlabel metal1 16652 5814 16652 5814 0 _190_
rlabel metal2 15778 8262 15778 8262 0 _191_
rlabel metal1 17664 7514 17664 7514 0 _192_
rlabel metal1 17158 9010 17158 9010 0 _193_
rlabel metal1 16146 9010 16146 9010 0 _194_
rlabel metal1 18630 5338 18630 5338 0 _195_
rlabel metal1 19228 5338 19228 5338 0 _196_
rlabel metal1 16790 12070 16790 12070 0 _197_
rlabel metal1 19320 5678 19320 5678 0 _198_
rlabel metal1 17618 6426 17618 6426 0 _199_
rlabel metal2 18722 5916 18722 5916 0 _200_
rlabel metal1 18308 5882 18308 5882 0 _201_
rlabel metal1 19642 8466 19642 8466 0 _202_
rlabel metal1 19826 8500 19826 8500 0 _203_
rlabel metal1 19872 8058 19872 8058 0 _204_
rlabel metal1 18262 7888 18262 7888 0 _205_
rlabel metal2 17802 8432 17802 8432 0 _206_
rlabel metal1 15410 11084 15410 11084 0 _207_
rlabel metal1 14858 8568 14858 8568 0 _208_
rlabel metal2 11914 9214 11914 9214 0 _209_
rlabel metal1 14674 7514 14674 7514 0 _210_
rlabel metal1 12604 7514 12604 7514 0 _211_
rlabel metal1 13064 7446 13064 7446 0 _212_
rlabel metal1 13156 8058 13156 8058 0 _213_
rlabel metal1 11868 9146 11868 9146 0 _214_
rlabel metal2 21022 8772 21022 8772 0 _215_
rlabel metal1 20470 8602 20470 8602 0 _216_
rlabel metal1 18630 8602 18630 8602 0 _217_
rlabel metal2 18538 8857 18538 8857 0 _218_
rlabel metal1 16698 11254 16698 11254 0 _219_
rlabel metal1 12788 10098 12788 10098 0 _220_
rlabel via2 12650 10115 12650 10115 0 _221_
rlabel metal1 12604 10234 12604 10234 0 _222_
rlabel via2 16882 7973 16882 7973 0 _223_
rlabel metal1 12006 10540 12006 10540 0 _224_
rlabel metal1 14444 12750 14444 12750 0 _225_
rlabel metal1 14766 11594 14766 11594 0 _226_
rlabel metal2 12834 11356 12834 11356 0 _227_
rlabel metal1 12972 8602 12972 8602 0 _228_
rlabel metal2 11086 10064 11086 10064 0 _229_
rlabel metal1 11178 10676 11178 10676 0 _230_
rlabel metal1 11178 10540 11178 10540 0 _231_
rlabel metal1 12098 10778 12098 10778 0 _232_
rlabel metal2 14950 8092 14950 8092 0 _233_
rlabel metal2 14674 8432 14674 8432 0 _234_
rlabel metal1 13662 8976 13662 8976 0 _235_
rlabel metal1 13248 9078 13248 9078 0 _236_
rlabel metal1 15870 14518 15870 14518 0 _237_
rlabel metal1 13708 11322 13708 11322 0 _238_
rlabel metal1 12512 11730 12512 11730 0 _239_
rlabel metal1 19918 12614 19918 12614 0 _240_
rlabel metal1 14904 12274 14904 12274 0 _241_
rlabel metal1 14306 12138 14306 12138 0 _242_
rlabel metal2 14582 15300 14582 15300 0 _243_
rlabel metal1 14214 15470 14214 15470 0 _244_
rlabel metal1 16974 14348 16974 14348 0 _245_
rlabel metal1 15686 14586 15686 14586 0 _246_
rlabel metal1 16192 11866 16192 11866 0 _247_
rlabel metal1 16330 13328 16330 13328 0 _248_
rlabel metal1 15686 13498 15686 13498 0 _249_
rlabel metal2 15318 15300 15318 15300 0 _250_
rlabel metal1 18078 10778 18078 10778 0 _251_
rlabel metal1 21114 11322 21114 11322 0 _252_
rlabel metal2 19458 11662 19458 11662 0 _253_
rlabel metal1 18308 12410 18308 12410 0 _254_
rlabel metal1 18354 12954 18354 12954 0 _255_
rlabel metal1 18170 13940 18170 13940 0 _256_
rlabel metal1 17434 13974 17434 13974 0 _257_
rlabel metal1 16744 12886 16744 12886 0 _258_
rlabel metal2 17066 12988 17066 12988 0 _259_
rlabel metal1 16882 12954 16882 12954 0 _260_
rlabel metal1 17020 12750 17020 12750 0 _261_
rlabel metal1 16974 14042 16974 14042 0 _262_
rlabel metal2 16606 14790 16606 14790 0 _263_
rlabel metal1 16974 14858 16974 14858 0 _264_
rlabel metal2 16606 16116 16606 16116 0 _265_
rlabel metal1 14214 21522 14214 21522 0 _266_
rlabel metal2 14214 21012 14214 21012 0 _267_
rlabel metal2 13478 21148 13478 21148 0 _268_
rlabel metal1 6946 6392 6946 6392 0 _269_
rlabel metal2 10534 13605 10534 13605 0 _270_
rlabel metal1 6808 3502 6808 3502 0 _271_
rlabel metal1 6026 3604 6026 3604 0 _272_
rlabel metal1 4646 4182 4646 4182 0 _273_
rlabel metal1 4692 3910 4692 3910 0 _274_
rlabel metal1 4646 6698 4646 6698 0 _275_
rlabel metal1 3404 4046 3404 4046 0 _276_
rlabel metal2 6118 3774 6118 3774 0 _277_
rlabel metal1 6578 3706 6578 3706 0 _278_
rlabel metal1 8786 6222 8786 6222 0 _279_
rlabel metal2 7222 6562 7222 6562 0 _280_
rlabel metal1 6624 9078 6624 9078 0 _281_
rlabel metal1 8004 7718 8004 7718 0 _282_
rlabel metal1 7406 5712 7406 5712 0 _283_
rlabel metal1 2714 12886 2714 12886 0 _284_
rlabel metal1 6716 15878 6716 15878 0 _285_
rlabel metal2 6578 8636 6578 8636 0 _286_
rlabel metal1 6164 6834 6164 6834 0 _287_
rlabel metal1 6578 6970 6578 6970 0 _288_
rlabel metal2 7314 6698 7314 6698 0 _289_
rlabel metal1 8004 5882 8004 5882 0 _290_
rlabel metal1 8786 5270 8786 5270 0 _291_
rlabel metal2 8418 5814 8418 5814 0 _292_
rlabel metal1 8878 6630 8878 6630 0 _293_
rlabel metal2 6578 11458 6578 11458 0 _294_
rlabel metal1 4186 10438 4186 10438 0 _295_
rlabel metal1 3864 10234 3864 10234 0 _296_
rlabel metal2 5658 11254 5658 11254 0 _297_
rlabel metal1 5160 11050 5160 11050 0 _298_
rlabel metal2 5474 11866 5474 11866 0 _299_
rlabel metal2 6026 12002 6026 12002 0 _300_
rlabel metal2 9890 11696 9890 11696 0 _301_
rlabel metal1 9246 8398 9246 8398 0 _302_
rlabel metal1 10488 13702 10488 13702 0 _303_
rlabel metal1 7636 7854 7636 7854 0 _304_
rlabel metal1 9338 7888 9338 7888 0 _305_
rlabel metal1 9798 8058 9798 8058 0 _306_
rlabel metal2 9154 7718 9154 7718 0 _307_
rlabel metal1 7360 4114 7360 4114 0 _308_
rlabel metal2 7222 4386 7222 4386 0 _309_
rlabel metal1 7682 4794 7682 4794 0 _310_
rlabel metal1 9430 6426 9430 6426 0 _311_
rlabel metal1 8602 7514 8602 7514 0 _312_
rlabel metal1 5934 9690 5934 9690 0 _313_
rlabel metal2 6210 10948 6210 10948 0 _314_
rlabel metal1 8510 11696 8510 11696 0 _315_
rlabel metal2 9890 10268 9890 10268 0 _316_
rlabel metal1 11408 15334 11408 15334 0 _317_
rlabel metal1 9476 10098 9476 10098 0 _318_
rlabel metal1 9476 10778 9476 10778 0 _319_
rlabel metal2 8418 11424 8418 11424 0 _320_
rlabel metal2 4278 5100 4278 5100 0 _321_
rlabel metal1 4186 4250 4186 4250 0 _322_
rlabel metal1 5244 4658 5244 4658 0 _323_
rlabel metal2 4094 4743 4094 4743 0 _324_
rlabel metal1 8694 10234 8694 10234 0 _325_
rlabel metal2 8510 10914 8510 10914 0 _326_
rlabel metal2 8602 11730 8602 11730 0 _327_
rlabel metal1 6578 12818 6578 12818 0 _328_
rlabel metal1 4922 12818 4922 12818 0 _329_
rlabel metal1 5014 13260 5014 13260 0 _330_
rlabel metal1 6210 12750 6210 12750 0 _331_
rlabel metal1 9338 12240 9338 12240 0 _332_
rlabel metal2 9890 14892 9890 14892 0 _333_
rlabel metal1 9200 2414 9200 2414 0 _334_
rlabel metal2 9154 10676 9154 10676 0 _335_
rlabel metal2 4554 4114 4554 4114 0 _336_
rlabel metal1 7038 2958 7038 2958 0 _337_
rlabel metal1 8832 2618 8832 2618 0 _338_
rlabel metal1 3266 3638 3266 3638 0 _339_
rlabel metal1 6026 3162 6026 3162 0 _340_
rlabel metal1 7590 3162 7590 3162 0 _341_
rlabel metal1 8234 5338 8234 5338 0 _342_
rlabel metal1 9752 5678 9752 5678 0 _343_
rlabel metal1 8878 5882 8878 5882 0 _344_
rlabel metal2 9062 8738 9062 8738 0 _345_
rlabel metal1 8510 10982 8510 10982 0 _346_
rlabel metal1 7268 12818 7268 12818 0 _347_
rlabel metal1 7314 12614 7314 12614 0 _348_
rlabel metal2 2530 15198 2530 15198 0 _349_
rlabel metal1 2714 11696 2714 11696 0 _350_
rlabel metal1 1840 14994 1840 14994 0 _351_
rlabel metal1 8096 14994 8096 14994 0 _352_
rlabel metal1 8326 14416 8326 14416 0 _353_
rlabel metal2 8142 14008 8142 14008 0 _354_
rlabel metal2 8326 15232 8326 15232 0 _355_
rlabel metal2 8418 17204 8418 17204 0 _356_
rlabel metal1 5704 13906 5704 13906 0 _357_
rlabel metal2 6854 13736 6854 13736 0 _358_
rlabel metal1 4784 13498 4784 13498 0 _359_
rlabel metal2 2806 12376 2806 12376 0 _360_
rlabel metal1 3450 12886 3450 12886 0 _361_
rlabel metal1 2990 12818 2990 12818 0 _362_
rlabel metal1 2116 12954 2116 12954 0 _363_
rlabel metal2 3542 14246 3542 14246 0 _364_
rlabel metal1 2211 14042 2211 14042 0 _365_
rlabel metal1 3818 15096 3818 15096 0 _366_
rlabel metal2 2898 14586 2898 14586 0 _367_
rlabel metal1 3588 15402 3588 15402 0 _368_
rlabel metal2 1610 15878 1610 15878 0 _369_
rlabel metal1 2208 16218 2208 16218 0 _370_
rlabel metal2 2530 16116 2530 16116 0 _371_
rlabel via2 7866 2635 7866 2635 0 _372_
rlabel metal1 7682 8058 7682 8058 0 _373_
rlabel metal1 7268 8602 7268 8602 0 _374_
rlabel metal1 9430 12886 9430 12886 0 _375_
rlabel metal1 2116 11730 2116 11730 0 _376_
rlabel metal1 5244 8602 5244 8602 0 _377_
rlabel metal2 2714 6188 2714 6188 0 _378_
rlabel metal2 5198 6154 5198 6154 0 _379_
rlabel metal1 1978 5270 1978 5270 0 _380_
rlabel metal2 1932 10540 1932 10540 0 _381_
rlabel metal1 6394 6902 6394 6902 0 _382_
rlabel metal1 9706 11152 9706 11152 0 _383_
rlabel metal2 6486 14586 6486 14586 0 _384_
rlabel metal1 5980 14382 5980 14382 0 _385_
rlabel metal1 5428 13158 5428 13158 0 _386_
rlabel metal1 5428 13294 5428 13294 0 _387_
rlabel metal1 2070 13260 2070 13260 0 _388_
rlabel metal2 10350 11322 10350 11322 0 _389_
rlabel metal1 10672 6222 10672 6222 0 _390_
rlabel metal1 2990 10540 2990 10540 0 _391_
rlabel metal1 3450 11764 3450 11764 0 _392_
rlabel metal1 2898 10710 2898 10710 0 _393_
rlabel metal2 2806 10812 2806 10812 0 _394_
rlabel metal2 2254 10438 2254 10438 0 _395_
rlabel metal2 8878 7344 8878 7344 0 _396_
rlabel metal1 2116 6698 2116 6698 0 _397_
rlabel metal1 2530 12716 2530 12716 0 _398_
rlabel metal1 3404 4114 3404 4114 0 _399_
rlabel metal1 8648 3706 8648 3706 0 _400_
rlabel metal1 9016 14790 9016 14790 0 _401_
rlabel metal1 9384 3570 9384 3570 0 _402_
rlabel metal2 7406 7565 7406 7565 0 _403_
rlabel metal2 2530 22688 2530 22688 0 clk
rlabel metal2 7038 16898 7038 16898 0 clknet_0_clk
rlabel metal1 7084 17170 7084 17170 0 clknet_2_0__leaf_clk
rlabel metal1 5336 19346 5336 19346 0 clknet_2_1__leaf_clk
rlabel metal1 8280 19822 8280 19822 0 clknet_2_2__leaf_clk
rlabel metal1 13110 21386 13110 21386 0 clknet_2_3__leaf_clk
rlabel metal1 14352 21998 14352 21998 0 io_in[0]
rlabel metal1 17572 21998 17572 21998 0 io_in[1]
rlabel metal1 22540 21998 22540 21998 0 io_in[2]
rlabel metal2 1518 1520 1518 1520 0 io_out[0]
rlabel metal2 2162 1792 2162 1792 0 io_out[1]
rlabel metal2 2806 1520 2806 1520 0 io_out[2]
rlabel metal2 3450 1520 3450 1520 0 io_out[3]
rlabel metal2 4094 1520 4094 1520 0 io_out[4]
rlabel metal2 4738 1520 4738 1520 0 io_out[5]
rlabel metal2 5382 1520 5382 1520 0 io_out[6]
rlabel metal2 6026 1520 6026 1520 0 io_out[7]
rlabel metal1 7038 16048 7038 16048 0 lcd.num_state\[0\]
rlabel metal1 9200 16014 9200 16014 0 lcd.num_state\[1\]
rlabel metal1 11546 18122 11546 18122 0 lcd.rom_addr\[0\]
rlabel metal1 14582 17510 14582 17510 0 lcd.rom_addr\[1\]
rlabel metal1 12926 12852 12926 12852 0 lcd.rom_addr\[3\]
rlabel metal1 10580 14518 10580 14518 0 lcd.rom_addr\[4\]
rlabel metal1 11638 14994 11638 14994 0 lcd.rom_addr\[5\]
rlabel metal2 13110 16252 13110 16252 0 lcd.rom_addr\[6\]
rlabel metal1 7958 15538 7958 15538 0 lcd.round\[0\]
rlabel metal2 8510 15980 8510 15980 0 lcd.round\[1\]
rlabel metal1 11316 15130 11316 15130 0 lcd.s_ROM\[0\]
rlabel metal1 11730 21896 11730 21896 0 lcd.s_ROM\[1\]
rlabel metal1 11776 15538 11776 15538 0 lcd.s_ROM\[2\]
rlabel metal2 9154 16762 9154 16762 0 lcd.s_ROM\[3\]
rlabel metal2 10810 17374 10810 17374 0 lcd.s_ROM\[4\]
rlabel metal1 10810 13838 10810 13838 0 lcd.s_ROM\[5\]
rlabel metal2 12006 15946 12006 15946 0 lcd.s_ROM\[6\]
rlabel metal1 4370 20230 4370 20230 0 lcd.seq\[0\]
rlabel metal1 2346 11118 2346 11118 0 lcd.seq\[1\]
rlabel metal2 2254 6154 2254 6154 0 lcd.seq\[2\]
rlabel metal1 1932 5814 1932 5814 0 lcd.seq\[3\]
rlabel metal1 1932 11322 1932 11322 0 lcd.seq\[4\]
rlabel metal1 3174 6766 3174 6766 0 lcd.seq\[5\]
rlabel metal1 1748 11254 1748 11254 0 lcd.seq\[6\]
rlabel via3 3427 16660 3427 16660 0 lcd.seq\[7\]
rlabel metal1 6762 15436 6762 15436 0 lcd.toggle
rlabel metal2 13754 21148 13754 21148 0 net1
rlabel metal2 16882 2720 16882 2720 0 net10
rlabel metal1 12558 6800 12558 6800 0 net11
rlabel metal1 16238 2448 16238 2448 0 net12
rlabel metal2 6670 1095 6670 1095 0 net13
rlabel metal1 6900 3026 6900 3026 0 net14
rlabel metal1 6394 3094 6394 3094 0 net15
rlabel metal2 8602 2064 8602 2064 0 net16
rlabel metal2 9246 1928 9246 1928 0 net17
rlabel metal2 9890 1826 9890 1826 0 net18
rlabel metal2 10534 1554 10534 1554 0 net19
rlabel metal1 13846 21420 13846 21420 0 net2
rlabel metal2 11178 1656 11178 1656 0 net20
rlabel metal2 11822 1554 11822 1554 0 net21
rlabel metal2 12466 823 12466 823 0 net22
rlabel metal2 13110 1588 13110 1588 0 net23
rlabel metal2 13754 1588 13754 1588 0 net24
rlabel metal2 14398 1588 14398 1588 0 net25
rlabel metal2 15042 1588 15042 1588 0 net26
rlabel metal1 15732 2822 15732 2822 0 net27
rlabel metal2 16330 1588 16330 1588 0 net28
rlabel metal2 16974 1588 16974 1588 0 net29
rlabel metal1 22494 21896 22494 21896 0 net3
rlabel metal2 17618 1588 17618 1588 0 net30
rlabel metal2 18262 1095 18262 1095 0 net31
rlabel metal2 18906 1588 18906 1588 0 net32
rlabel metal2 19550 1588 19550 1588 0 net33
rlabel metal2 20194 1588 20194 1588 0 net34
rlabel metal2 20838 1095 20838 1095 0 net35
rlabel metal2 21482 1588 21482 1588 0 net36
rlabel metal2 22126 1588 22126 1588 0 net37
rlabel metal1 22816 2822 22816 2822 0 net38
rlabel metal1 23368 3502 23368 3502 0 net39
rlabel metal1 7314 15470 7314 15470 0 net4
rlabel metal2 1886 2193 1886 2193 0 net5
rlabel metal2 2530 3519 2530 3519 0 net6
rlabel metal1 2990 2414 2990 2414 0 net7
rlabel metal2 16422 2210 16422 2210 0 net8
rlabel metal2 17434 3587 17434 3587 0 net9
rlabel metal1 7452 21930 7452 21930 0 rst
<< properties >>
string FIXED_BBOX 0 0 25000 25000
<< end >>
