magic
tech sky130B
magscale 1 2
timestamp 1680615612
<< metal1 >>
rect 267642 700816 267648 700868
rect 267700 700856 267706 700868
rect 445110 700856 445116 700868
rect 267700 700828 445116 700856
rect 267700 700816 267706 700828
rect 445110 700816 445116 700828
rect 445168 700816 445174 700868
rect 235166 700748 235172 700800
rect 235224 700788 235230 700800
rect 449250 700788 449256 700800
rect 235224 700760 449256 700788
rect 235224 700748 235230 700760
rect 449250 700748 449256 700760
rect 449308 700748 449314 700800
rect 218974 700680 218980 700732
rect 219032 700720 219038 700732
rect 446490 700720 446496 700732
rect 219032 700692 446496 700720
rect 219032 700680 219038 700692
rect 446490 700680 446496 700692
rect 446548 700680 446554 700732
rect 154114 700612 154120 700664
rect 154172 700652 154178 700664
rect 418798 700652 418804 700664
rect 154172 700624 418804 700652
rect 154172 700612 154178 700624
rect 418798 700612 418804 700624
rect 418856 700612 418862 700664
rect 429838 700612 429844 700664
rect 429896 700652 429902 700664
rect 444098 700652 444104 700664
rect 429896 700624 444104 700652
rect 429896 700612 429902 700624
rect 444098 700612 444104 700624
rect 444156 700612 444162 700664
rect 170306 700544 170312 700596
rect 170364 700584 170370 700596
rect 446398 700584 446404 700596
rect 170364 700556 446404 700584
rect 170364 700544 170370 700556
rect 446398 700544 446404 700556
rect 446456 700544 446462 700596
rect 137830 700476 137836 700528
rect 137888 700516 137894 700528
rect 445202 700516 445208 700528
rect 137888 700488 445208 700516
rect 137888 700476 137894 700488
rect 445202 700476 445208 700488
rect 445260 700476 445266 700528
rect 105446 700408 105452 700460
rect 105504 700448 105510 700460
rect 444190 700448 444196 700460
rect 105504 700420 444196 700448
rect 105504 700408 105510 700420
rect 444190 700408 444196 700420
rect 444248 700408 444254 700460
rect 447870 700408 447876 700460
rect 447928 700448 447934 700460
rect 478506 700448 478512 700460
rect 447928 700420 478512 700448
rect 447928 700408 447934 700420
rect 478506 700408 478512 700420
rect 478564 700408 478570 700460
rect 40494 700340 40500 700392
rect 40552 700380 40558 700392
rect 449158 700380 449164 700392
rect 40552 700352 449164 700380
rect 40552 700340 40558 700352
rect 449158 700340 449164 700352
rect 449216 700340 449222 700392
rect 8110 700272 8116 700324
rect 8168 700312 8174 700324
rect 445018 700312 445024 700324
rect 8168 700284 445024 700312
rect 8168 700272 8174 700284
rect 445018 700272 445024 700284
rect 445076 700272 445082 700324
rect 447778 700272 447784 700324
rect 447836 700312 447842 700324
rect 494790 700312 494796 700324
rect 447836 700284 494796 700312
rect 447836 700272 447842 700284
rect 494790 700272 494796 700284
rect 494848 700272 494854 700324
rect 348786 686536 348792 686588
rect 348844 686576 348850 686588
rect 446582 686576 446588 686588
rect 348844 686548 446588 686576
rect 348844 686536 348850 686548
rect 446582 686536 446588 686548
rect 446640 686536 446646 686588
rect 283834 686468 283840 686520
rect 283892 686508 283898 686520
rect 446674 686508 446680 686520
rect 283892 686480 446680 686508
rect 283892 686468 283898 686480
rect 446674 686468 446680 686480
rect 446732 686468 446738 686520
rect 332502 685312 332508 685364
rect 332560 685352 332566 685364
rect 418890 685352 418896 685364
rect 332560 685324 418896 685352
rect 332560 685312 332566 685324
rect 418890 685312 418896 685324
rect 418948 685312 418954 685364
rect 202782 685244 202788 685296
rect 202840 685284 202846 685296
rect 445294 685284 445300 685296
rect 202840 685256 445300 685284
rect 202840 685244 202846 685256
rect 445294 685244 445300 685256
rect 445352 685244 445358 685296
rect 89162 685176 89168 685228
rect 89220 685216 89226 685228
rect 416038 685216 416044 685228
rect 89220 685188 416044 685216
rect 89220 685176 89226 685188
rect 416038 685176 416044 685188
rect 416096 685176 416102 685228
rect 72970 685108 72976 685160
rect 73028 685148 73034 685160
rect 449342 685148 449348 685160
rect 73028 685120 449348 685148
rect 73028 685108 73034 685120
rect 449342 685108 449348 685120
rect 449400 685108 449406 685160
rect 19978 684564 19984 684616
rect 20036 684604 20042 684616
rect 418982 684604 418988 684616
rect 20036 684576 418988 684604
rect 20036 684564 20042 684576
rect 418982 684564 418988 684576
rect 419040 684564 419046 684616
rect 3786 684496 3792 684548
rect 3844 684536 3850 684548
rect 420178 684536 420184 684548
rect 3844 684508 420184 684536
rect 3844 684496 3850 684508
rect 420178 684496 420184 684508
rect 420236 684496 420242 684548
rect 18322 683748 18328 683800
rect 18380 683788 18386 683800
rect 359458 683788 359464 683800
rect 18380 683760 359464 683788
rect 18380 683748 18386 683760
rect 359458 683748 359464 683760
rect 359516 683748 359522 683800
rect 21358 683680 21364 683732
rect 21416 683720 21422 683732
rect 420730 683720 420736 683732
rect 21416 683692 420736 683720
rect 21416 683680 21422 683692
rect 420730 683680 420736 683692
rect 420788 683680 420794 683732
rect 4062 683612 4068 683664
rect 4120 683652 4126 683664
rect 420270 683652 420276 683664
rect 4120 683624 420276 683652
rect 4120 683612 4126 683624
rect 420270 683612 420276 683624
rect 420328 683612 420334 683664
rect 3510 683544 3516 683596
rect 3568 683584 3574 683596
rect 420362 683584 420368 683596
rect 3568 683556 420368 683584
rect 3568 683544 3574 683556
rect 420362 683544 420368 683556
rect 420420 683544 420426 683596
rect 3694 683476 3700 683528
rect 3752 683516 3758 683528
rect 420638 683516 420644 683528
rect 3752 683488 420644 683516
rect 3752 683476 3758 683488
rect 420638 683476 420644 683488
rect 420696 683476 420702 683528
rect 3418 683408 3424 683460
rect 3476 683448 3482 683460
rect 420546 683448 420552 683460
rect 3476 683420 420552 683448
rect 3476 683408 3482 683420
rect 420546 683408 420552 683420
rect 420604 683408 420610 683460
rect 3878 683340 3884 683392
rect 3936 683380 3942 683392
rect 445478 683380 445484 683392
rect 3936 683352 445484 683380
rect 3936 683340 3942 683352
rect 445478 683340 445484 683352
rect 445536 683340 445542 683392
rect 3602 683272 3608 683324
rect 3660 683312 3666 683324
rect 445386 683312 445392 683324
rect 3660 683284 445392 683312
rect 3660 683272 3666 683284
rect 445386 683272 445392 683284
rect 445444 683272 445450 683324
rect 3970 683204 3976 683256
rect 4028 683244 4034 683256
rect 446858 683244 446864 683256
rect 4028 683216 446864 683244
rect 4028 683204 4034 683216
rect 446858 683204 446864 683216
rect 446916 683204 446922 683256
rect 3326 683136 3332 683188
rect 3384 683176 3390 683188
rect 446306 683176 446312 683188
rect 3384 683148 446312 683176
rect 3384 683136 3390 683148
rect 446306 683136 446312 683148
rect 446364 683136 446370 683188
rect 576118 683136 576124 683188
rect 576176 683176 576182 683188
rect 579614 683176 579620 683188
rect 576176 683148 579620 683176
rect 576176 683136 576182 683148
rect 579614 683136 579620 683148
rect 579672 683136 579678 683188
rect 3234 682660 3240 682712
rect 3292 682700 3298 682712
rect 447042 682700 447048 682712
rect 3292 682672 447048 682700
rect 3292 682660 3298 682672
rect 447042 682660 447048 682672
rect 447100 682660 447106 682712
rect 17218 680348 17224 680400
rect 17276 680388 17282 680400
rect 18322 680388 18328 680400
rect 17276 680360 18328 680388
rect 17276 680348 17282 680360
rect 18322 680348 18328 680360
rect 18380 680348 18386 680400
rect 359458 672052 359464 672104
rect 359516 672092 359522 672104
rect 360838 672092 360844 672104
rect 359516 672064 360844 672092
rect 359516 672052 359522 672064
rect 360838 672052 360844 672064
rect 360896 672052 360902 672104
rect 361758 667904 361764 667956
rect 361816 667944 361822 667956
rect 378870 667944 378876 667956
rect 361816 667916 378876 667944
rect 361816 667904 361822 667916
rect 378870 667904 378876 667916
rect 378928 667904 378934 667956
rect 17218 661076 17224 661088
rect 16546 661048 17224 661076
rect 14182 660968 14188 661020
rect 14240 661008 14246 661020
rect 16546 661008 16574 661048
rect 17218 661036 17224 661048
rect 17276 661036 17282 661088
rect 14240 660980 16574 661008
rect 14240 660968 14246 660980
rect 3142 658180 3148 658232
rect 3200 658220 3206 658232
rect 19978 658220 19984 658232
rect 3200 658192 19984 658220
rect 3200 658180 3206 658192
rect 19978 658180 19984 658192
rect 20036 658180 20042 658232
rect 361758 656888 361764 656940
rect 361816 656928 361822 656940
rect 376018 656928 376024 656940
rect 361816 656900 376024 656928
rect 361816 656888 361822 656900
rect 376018 656888 376024 656900
rect 376076 656888 376082 656940
rect 11698 656616 11704 656668
rect 11756 656656 11762 656668
rect 14182 656656 14188 656668
rect 11756 656628 14188 656656
rect 11756 656616 11762 656628
rect 14182 656616 14188 656628
rect 14240 656616 14246 656668
rect 361758 645872 361764 645924
rect 361816 645912 361822 645924
rect 374638 645912 374644 645924
rect 361816 645884 374644 645912
rect 361816 645872 361822 645884
rect 374638 645872 374644 645884
rect 374696 645872 374702 645924
rect 10594 645804 10600 645856
rect 10652 645844 10658 645856
rect 11698 645844 11704 645856
rect 10652 645816 11704 645844
rect 10652 645804 10658 645816
rect 11698 645804 11704 645816
rect 11756 645804 11762 645856
rect 5534 643696 5540 643748
rect 5592 643736 5598 643748
rect 10594 643736 10600 643748
rect 5592 643708 10600 643736
rect 5592 643696 5598 643708
rect 10594 643696 10600 643708
rect 10652 643696 10658 643748
rect 4798 640296 4804 640348
rect 4856 640336 4862 640348
rect 5534 640336 5540 640348
rect 4856 640308 5540 640336
rect 4856 640296 4862 640308
rect 5534 640296 5540 640308
rect 5592 640296 5598 640348
rect 361574 634788 361580 634840
rect 361632 634828 361638 634840
rect 400858 634828 400864 634840
rect 361632 634800 400864 634828
rect 361632 634788 361638 634800
rect 400858 634788 400864 634800
rect 400916 634788 400922 634840
rect 3602 631320 3608 631372
rect 3660 631360 3666 631372
rect 20898 631360 20904 631372
rect 3660 631332 20904 631360
rect 3660 631320 3666 631332
rect 20898 631320 20904 631332
rect 20956 631320 20962 631372
rect 361574 623772 361580 623824
rect 361632 623812 361638 623824
rect 371878 623812 371884 623824
rect 361632 623784 371884 623812
rect 361632 623772 361638 623784
rect 371878 623772 371884 623784
rect 371936 623772 371942 623824
rect 570598 616836 570604 616888
rect 570656 616876 570662 616888
rect 579614 616876 579620 616888
rect 570656 616848 579620 616876
rect 570656 616836 570662 616848
rect 579614 616836 579620 616848
rect 579672 616836 579678 616888
rect 361574 612824 361580 612876
rect 361632 612864 361638 612876
rect 363598 612864 363604 612876
rect 361632 612836 363604 612864
rect 361632 612824 361638 612836
rect 363598 612824 363604 612836
rect 363656 612824 363662 612876
rect 458818 604120 458824 604172
rect 458876 604120 458882 604172
rect 458836 603968 458864 604120
rect 458818 603916 458824 603968
rect 458876 603916 458882 603968
rect 459002 603712 459008 603764
rect 459060 603752 459066 603764
rect 459462 603752 459468 603764
rect 459060 603724 459468 603752
rect 459060 603712 459066 603724
rect 459462 603712 459468 603724
rect 459520 603712 459526 603764
rect 459830 602080 459836 602132
rect 459888 602120 459894 602132
rect 460106 602120 460112 602132
rect 459888 602092 460112 602120
rect 459888 602080 459894 602092
rect 460106 602080 460112 602092
rect 460164 602080 460170 602132
rect 361758 601672 361764 601724
rect 361816 601712 361822 601724
rect 370498 601712 370504 601724
rect 361816 601684 370504 601712
rect 361816 601672 361822 601684
rect 370498 601672 370504 601684
rect 370556 601672 370562 601724
rect 460106 600244 460112 600296
rect 460164 600284 460170 600296
rect 462314 600284 462320 600296
rect 460164 600256 462320 600284
rect 460164 600244 460170 600256
rect 462314 600244 462320 600256
rect 462372 600244 462378 600296
rect 457346 600176 457352 600228
rect 457404 600216 457410 600228
rect 462958 600216 462964 600228
rect 457404 600188 462964 600216
rect 457404 600176 457410 600188
rect 462958 600176 462964 600188
rect 463016 600176 463022 600228
rect 457530 599768 457536 599820
rect 457588 599808 457594 599820
rect 464338 599808 464344 599820
rect 457588 599780 464344 599808
rect 457588 599768 457594 599780
rect 464338 599768 464344 599780
rect 464396 599768 464402 599820
rect 459002 599700 459008 599752
rect 459060 599740 459066 599752
rect 466454 599740 466460 599752
rect 459060 599712 466460 599740
rect 459060 599700 459066 599712
rect 466454 599700 466460 599712
rect 466512 599700 466518 599752
rect 458726 599632 458732 599684
rect 458784 599672 458790 599684
rect 469214 599672 469220 599684
rect 458784 599644 469220 599672
rect 458784 599632 458790 599644
rect 469214 599632 469220 599644
rect 469272 599632 469278 599684
rect 457438 599564 457444 599616
rect 457496 599604 457502 599616
rect 468478 599604 468484 599616
rect 457496 599576 468484 599604
rect 457496 599564 457502 599576
rect 468478 599564 468484 599576
rect 468536 599564 468542 599616
rect 515398 599564 515404 599616
rect 515456 599604 515462 599616
rect 580534 599604 580540 599616
rect 515456 599576 580540 599604
rect 515456 599564 515462 599576
rect 580534 599564 580540 599576
rect 580592 599564 580598 599616
rect 457254 598680 457260 598732
rect 457312 598720 457318 598732
rect 461578 598720 461584 598732
rect 457312 598692 461584 598720
rect 457312 598680 457318 598692
rect 461578 598680 461584 598692
rect 461636 598680 461642 598732
rect 459462 598408 459468 598460
rect 459520 598448 459526 598460
rect 463694 598448 463700 598460
rect 459520 598420 463700 598448
rect 459520 598408 459526 598420
rect 463694 598408 463700 598420
rect 463752 598408 463758 598460
rect 458634 598272 458640 598324
rect 458692 598312 458698 598324
rect 465074 598312 465080 598324
rect 458692 598284 465080 598312
rect 458692 598272 458698 598284
rect 465074 598272 465080 598284
rect 465132 598272 465138 598324
rect 488626 598272 488632 598324
rect 488684 598312 488690 598324
rect 494330 598312 494336 598324
rect 488684 598284 494336 598312
rect 488684 598272 488690 598284
rect 494330 598272 494336 598284
rect 494388 598272 494394 598324
rect 360838 598204 360844 598256
rect 360896 598244 360902 598256
rect 367738 598244 367744 598256
rect 360896 598216 367744 598244
rect 360896 598204 360902 598216
rect 367738 598204 367744 598216
rect 367796 598204 367802 598256
rect 457714 598204 457720 598256
rect 457772 598244 457778 598256
rect 465718 598244 465724 598256
rect 457772 598216 465724 598244
rect 457772 598204 457778 598216
rect 465718 598204 465724 598216
rect 465776 598204 465782 598256
rect 493318 598204 493324 598256
rect 493376 598244 493382 598256
rect 526714 598244 526720 598256
rect 493376 598216 526720 598244
rect 493376 598204 493382 598216
rect 526714 598204 526720 598216
rect 526772 598204 526778 598256
rect 459830 596844 459836 596896
rect 459888 596884 459894 596896
rect 466546 596884 466552 596896
rect 459888 596856 466552 596884
rect 459888 596844 459894 596856
rect 466546 596844 466552 596856
rect 466604 596844 466610 596896
rect 450538 596776 450544 596828
rect 450596 596816 450602 596828
rect 494974 596816 494980 596828
rect 450596 596788 494980 596816
rect 450596 596776 450602 596788
rect 494974 596776 494980 596788
rect 495032 596776 495038 596828
rect 457898 595892 457904 595944
rect 457956 595932 457962 595944
rect 461670 595932 461676 595944
rect 457956 595904 461676 595932
rect 457956 595892 457962 595904
rect 461670 595892 461676 595904
rect 461728 595892 461734 595944
rect 460198 595484 460204 595536
rect 460256 595524 460262 595536
rect 467926 595524 467932 595536
rect 460256 595496 467932 595524
rect 460256 595484 460262 595496
rect 467926 595484 467932 595496
rect 467984 595484 467990 595536
rect 457622 595416 457628 595468
rect 457680 595456 457686 595468
rect 468570 595456 468576 595468
rect 457680 595428 468576 595456
rect 457680 595416 457686 595428
rect 468570 595416 468576 595428
rect 468628 595416 468634 595468
rect 460014 594124 460020 594176
rect 460072 594164 460078 594176
rect 465166 594164 465172 594176
rect 460072 594136 465172 594164
rect 460072 594124 460078 594136
rect 465166 594124 465172 594136
rect 465224 594124 465230 594176
rect 457806 594056 457812 594108
rect 457864 594096 457870 594108
rect 467098 594096 467104 594108
rect 457864 594068 467104 594096
rect 457864 594056 457870 594068
rect 467098 594056 467104 594068
rect 467156 594056 467162 594108
rect 361574 590792 361580 590844
rect 361632 590832 361638 590844
rect 363690 590832 363696 590844
rect 361632 590804 363696 590832
rect 361632 590792 361638 590804
rect 363690 590792 363696 590804
rect 363748 590792 363754 590844
rect 511258 590656 511264 590708
rect 511316 590696 511322 590708
rect 580166 590696 580172 590708
rect 511316 590668 580172 590696
rect 511316 590656 511322 590668
rect 580166 590656 580172 590668
rect 580224 590656 580230 590708
rect 367738 587800 367744 587852
rect 367796 587840 367802 587852
rect 370590 587840 370596 587852
rect 367796 587812 370596 587840
rect 367796 587800 367802 587812
rect 370590 587800 370596 587812
rect 370648 587800 370654 587852
rect 361758 579640 361764 579692
rect 361816 579680 361822 579692
rect 368014 579680 368020 579692
rect 361816 579652 368020 579680
rect 361816 579640 361822 579652
rect 368014 579640 368020 579652
rect 368072 579640 368078 579692
rect 370590 579572 370596 579624
rect 370648 579612 370654 579624
rect 371970 579612 371976 579624
rect 370648 579584 371976 579612
rect 370648 579572 370654 579584
rect 371970 579572 371976 579584
rect 372028 579572 372034 579624
rect 511350 576852 511356 576904
rect 511408 576892 511414 576904
rect 579982 576892 579988 576904
rect 511408 576864 579988 576892
rect 511408 576852 511414 576864
rect 579982 576852 579988 576864
rect 580040 576852 580046 576904
rect 371970 571276 371976 571328
rect 372028 571316 372034 571328
rect 373258 571316 373264 571328
rect 372028 571288 373264 571316
rect 372028 571276 372034 571288
rect 373258 571276 373264 571288
rect 373316 571276 373322 571328
rect 361574 568760 361580 568812
rect 361632 568800 361638 568812
rect 363782 568800 363788 568812
rect 361632 568772 363788 568800
rect 361632 568760 361638 568772
rect 363782 568760 363788 568772
rect 363840 568760 363846 568812
rect 373258 564340 373264 564392
rect 373316 564380 373322 564392
rect 375282 564380 375288 564392
rect 373316 564352 375288 564380
rect 373316 564340 373322 564352
rect 375282 564340 375288 564352
rect 375340 564340 375346 564392
rect 515490 563048 515496 563100
rect 515548 563088 515554 563100
rect 580166 563088 580172 563100
rect 515548 563060 580172 563088
rect 515548 563048 515554 563060
rect 580166 563048 580172 563060
rect 580224 563048 580230 563100
rect 361666 557540 361672 557592
rect 361724 557580 361730 557592
rect 403618 557580 403624 557592
rect 361724 557552 403624 557580
rect 361724 557540 361730 557552
rect 403618 557540 403624 557552
rect 403676 557540 403682 557592
rect 375374 557132 375380 557184
rect 375432 557172 375438 557184
rect 377766 557172 377772 557184
rect 375432 557144 377772 557172
rect 375432 557132 375438 557144
rect 377766 557132 377772 557144
rect 377824 557132 377830 557184
rect 377766 550604 377772 550656
rect 377824 550644 377830 550656
rect 377824 550616 378180 550644
rect 377824 550604 377830 550616
rect 378152 550576 378180 550616
rect 380158 550576 380164 550588
rect 378152 550548 380164 550576
rect 380158 550536 380164 550548
rect 380216 550536 380222 550588
rect 361758 546456 361764 546508
rect 361816 546496 361822 546508
rect 419074 546496 419080 546508
rect 361816 546468 419080 546496
rect 361816 546456 361822 546468
rect 419074 546456 419080 546468
rect 419132 546456 419138 546508
rect 459922 542988 459928 543040
rect 459980 543028 459986 543040
rect 463786 543028 463792 543040
rect 459980 543000 463792 543028
rect 459980 542988 459986 543000
rect 463786 542988 463792 543000
rect 463844 542988 463850 543040
rect 380158 540880 380164 540932
rect 380216 540920 380222 540932
rect 382274 540920 382280 540932
rect 380216 540892 382280 540920
rect 380216 540880 380222 540892
rect 382274 540880 382280 540892
rect 382332 540880 382338 540932
rect 519538 536800 519544 536852
rect 519596 536840 519602 536852
rect 580166 536840 580172 536852
rect 519596 536812 580172 536840
rect 519596 536800 519602 536812
rect 580166 536800 580172 536812
rect 580224 536800 580230 536852
rect 361758 535440 361764 535492
rect 361816 535480 361822 535492
rect 406378 535480 406384 535492
rect 361816 535452 406384 535480
rect 361816 535440 361822 535452
rect 406378 535440 406384 535452
rect 406436 535440 406442 535492
rect 382274 532652 382280 532704
rect 382332 532692 382338 532704
rect 384298 532692 384304 532704
rect 382332 532664 384304 532692
rect 382332 532652 382338 532664
rect 384298 532652 384304 532664
rect 384356 532652 384362 532704
rect 361758 524424 361764 524476
rect 361816 524464 361822 524476
rect 407758 524464 407764 524476
rect 361816 524436 407764 524464
rect 361816 524424 361822 524436
rect 407758 524424 407764 524436
rect 407816 524424 407822 524476
rect 518158 524424 518164 524476
rect 518216 524464 518222 524476
rect 580166 524464 580172 524476
rect 518216 524436 580172 524464
rect 518216 524424 518222 524436
rect 580166 524424 580172 524436
rect 580224 524424 580230 524476
rect 384298 524084 384304 524136
rect 384356 524124 384362 524136
rect 385678 524124 385684 524136
rect 384356 524096 385684 524124
rect 384356 524084 384362 524096
rect 385678 524084 385684 524096
rect 385736 524084 385742 524136
rect 457990 522316 457996 522368
rect 458048 522356 458054 522368
rect 464430 522356 464436 522368
rect 458048 522328 464436 522356
rect 458048 522316 458054 522328
rect 464430 522316 464436 522328
rect 464488 522316 464494 522368
rect 459186 522248 459192 522300
rect 459244 522288 459250 522300
rect 469398 522288 469404 522300
rect 459244 522260 469404 522288
rect 459244 522248 459250 522260
rect 469398 522248 469404 522260
rect 469456 522248 469462 522300
rect 459278 520888 459284 520940
rect 459336 520928 459342 520940
rect 470594 520928 470600 520940
rect 459336 520900 470600 520928
rect 459336 520888 459342 520900
rect 470594 520888 470600 520900
rect 470652 520888 470658 520940
rect 482922 520888 482928 520940
rect 482980 520928 482986 520940
rect 520274 520928 520280 520940
rect 482980 520900 520280 520928
rect 482980 520888 482986 520900
rect 520274 520888 520280 520900
rect 520332 520888 520338 520940
rect 458082 519596 458088 519648
rect 458140 519636 458146 519648
rect 468662 519636 468668 519648
rect 458140 519608 468668 519636
rect 458140 519596 458146 519608
rect 468662 519596 468668 519608
rect 468720 519596 468726 519648
rect 459370 519528 459376 519580
rect 459428 519568 459434 519580
rect 470870 519568 470876 519580
rect 459428 519540 470876 519568
rect 459428 519528 459434 519540
rect 470870 519528 470876 519540
rect 470928 519528 470934 519580
rect 449710 518168 449716 518220
rect 449768 518208 449774 518220
rect 469858 518208 469864 518220
rect 449768 518180 469864 518208
rect 449768 518168 449774 518180
rect 469858 518168 469864 518180
rect 469916 518208 469922 518220
rect 494238 518208 494244 518220
rect 469916 518180 494244 518208
rect 469916 518168 469922 518180
rect 494238 518168 494244 518180
rect 494296 518168 494302 518220
rect 476022 517624 476028 517676
rect 476080 517664 476086 517676
rect 494146 517664 494152 517676
rect 476080 517636 494152 517664
rect 476080 517624 476086 517636
rect 494146 517624 494152 517636
rect 494204 517624 494210 517676
rect 449802 517556 449808 517608
rect 449860 517596 449866 517608
rect 488626 517596 488632 517608
rect 449860 517568 488632 517596
rect 449860 517556 449866 517568
rect 488626 517556 488632 517568
rect 488684 517556 488690 517608
rect 450354 517488 450360 517540
rect 450412 517528 450418 517540
rect 494330 517528 494336 517540
rect 450412 517500 494336 517528
rect 450412 517488 450418 517500
rect 494330 517488 494336 517500
rect 494388 517488 494394 517540
rect 482278 517420 482284 517472
rect 482336 517420 482342 517472
rect 450630 516808 450636 516860
rect 450688 516848 450694 516860
rect 476022 516848 476028 516860
rect 450688 516820 476028 516848
rect 450688 516808 450694 516820
rect 476022 516808 476028 516820
rect 476080 516808 476086 516860
rect 449986 516740 449992 516792
rect 450044 516780 450050 516792
rect 482296 516780 482324 517420
rect 492122 516780 492128 516792
rect 450044 516752 492128 516780
rect 450044 516740 450050 516752
rect 492122 516740 492128 516752
rect 492180 516740 492186 516792
rect 385678 516128 385684 516180
rect 385736 516168 385742 516180
rect 385736 516140 386460 516168
rect 385736 516128 385742 516140
rect 386432 516100 386460 516140
rect 389174 516100 389180 516112
rect 386432 516072 389180 516100
rect 389174 516060 389180 516072
rect 389232 516060 389238 516112
rect 3970 514768 3976 514820
rect 4028 514808 4034 514820
rect 4798 514808 4804 514820
rect 4028 514780 4804 514808
rect 4028 514768 4034 514780
rect 4798 514768 4804 514780
rect 4856 514768 4862 514820
rect 502242 514020 502248 514072
rect 502300 514060 502306 514072
rect 545114 514060 545120 514072
rect 502300 514032 545120 514060
rect 502300 514020 502306 514032
rect 545114 514020 545120 514032
rect 545172 514020 545178 514072
rect 361758 513340 361764 513392
rect 361816 513380 361822 513392
rect 410518 513380 410524 513392
rect 361816 513352 410524 513380
rect 361816 513340 361822 513352
rect 410518 513340 410524 513352
rect 410576 513340 410582 513392
rect 492122 512592 492128 512644
rect 492180 512632 492186 512644
rect 535454 512632 535460 512644
rect 492180 512604 535460 512632
rect 492180 512592 492186 512604
rect 535454 512592 535460 512604
rect 535512 512592 535518 512644
rect 389174 511912 389180 511964
rect 389232 511952 389238 511964
rect 391198 511952 391204 511964
rect 389232 511924 391204 511952
rect 389232 511912 389238 511924
rect 391198 511912 391204 511924
rect 391256 511912 391262 511964
rect 516778 510620 516784 510672
rect 516836 510660 516842 510672
rect 580166 510660 580172 510672
rect 516836 510632 580172 510660
rect 516836 510620 516842 510632
rect 580166 510620 580172 510632
rect 580224 510620 580230 510672
rect 494330 509872 494336 509924
rect 494388 509912 494394 509924
rect 538214 509912 538220 509924
rect 494388 509884 538220 509912
rect 494388 509872 494394 509884
rect 538214 509872 538220 509884
rect 538272 509872 538278 509924
rect 494146 508512 494152 508564
rect 494204 508552 494210 508564
rect 532694 508552 532700 508564
rect 494204 508524 532700 508552
rect 494204 508512 494210 508524
rect 532694 508512 532700 508524
rect 532752 508512 532758 508564
rect 391198 505792 391204 505844
rect 391256 505832 391262 505844
rect 392578 505832 392584 505844
rect 391256 505804 392584 505832
rect 391256 505792 391262 505804
rect 392578 505792 392584 505804
rect 392636 505792 392642 505844
rect 495066 505724 495072 505776
rect 495124 505764 495130 505776
rect 529934 505764 529940 505776
rect 495124 505736 529940 505764
rect 495124 505724 495130 505736
rect 529934 505724 529940 505736
rect 529992 505724 529998 505776
rect 361758 502324 361764 502376
rect 361816 502364 361822 502376
rect 411898 502364 411904 502376
rect 361816 502336 411904 502364
rect 361816 502324 361822 502336
rect 411898 502324 411904 502336
rect 411956 502324 411962 502376
rect 463142 497700 463148 497752
rect 463200 497740 463206 497752
rect 480254 497740 480260 497752
rect 463200 497712 480260 497740
rect 463200 497700 463206 497712
rect 480254 497700 480260 497712
rect 480312 497700 480318 497752
rect 458818 497632 458824 497684
rect 458876 497672 458882 497684
rect 481634 497672 481640 497684
rect 458876 497644 481640 497672
rect 458876 497632 458882 497644
rect 481634 497632 481640 497644
rect 481692 497632 481698 497684
rect 457530 497564 457536 497616
rect 457588 497604 457594 497616
rect 482646 497604 482652 497616
rect 457588 497576 482652 497604
rect 457588 497564 457594 497576
rect 482646 497564 482652 497576
rect 482704 497564 482710 497616
rect 457438 497496 457444 497548
rect 457496 497536 457502 497548
rect 483842 497536 483848 497548
rect 457496 497508 483848 497536
rect 457496 497496 457502 497508
rect 483842 497496 483848 497508
rect 483900 497496 483906 497548
rect 454678 497428 454684 497480
rect 454736 497468 454742 497480
rect 486234 497468 486240 497480
rect 454736 497440 486240 497468
rect 454736 497428 454742 497440
rect 486234 497428 486240 497440
rect 486292 497428 486298 497480
rect 455322 497020 455328 497072
rect 455380 497060 455386 497072
rect 459554 497060 459560 497072
rect 455380 497032 459560 497060
rect 455380 497020 455386 497032
rect 459554 497020 459560 497032
rect 459612 497020 459618 497072
rect 456518 496952 456524 497004
rect 456576 496992 456582 497004
rect 461026 496992 461032 497004
rect 456576 496964 461032 496992
rect 456576 496952 456582 496964
rect 461026 496952 461032 496964
rect 461084 496952 461090 497004
rect 453942 496884 453948 496936
rect 454000 496924 454006 496936
rect 456610 496924 456616 496936
rect 454000 496896 456616 496924
rect 454000 496884 454006 496896
rect 456610 496884 456616 496896
rect 456668 496884 456674 496936
rect 452562 496816 452568 496868
rect 452620 496856 452626 496868
rect 453666 496856 453672 496868
rect 452620 496828 453672 496856
rect 452620 496816 452626 496828
rect 453666 496816 453672 496828
rect 453724 496816 453730 496868
rect 455138 496816 455144 496868
rect 455196 496856 455202 496868
rect 458082 496856 458088 496868
rect 455196 496828 458088 496856
rect 455196 496816 455202 496828
rect 458082 496816 458088 496828
rect 458140 496816 458146 496868
rect 483658 496816 483664 496868
rect 483716 496856 483722 496868
rect 485038 496856 485044 496868
rect 483716 496828 485044 496856
rect 483716 496816 483722 496828
rect 485038 496816 485044 496828
rect 485096 496816 485102 496868
rect 361758 491308 361764 491360
rect 361816 491348 361822 491360
rect 381630 491348 381636 491360
rect 361816 491320 381636 491348
rect 361816 491308 361822 491320
rect 381630 491308 381636 491320
rect 381688 491308 381694 491360
rect 518250 484372 518256 484424
rect 518308 484412 518314 484424
rect 580166 484412 580172 484424
rect 518308 484384 580172 484412
rect 518308 484372 518314 484384
rect 580166 484372 580172 484384
rect 580224 484372 580230 484424
rect 361758 480224 361764 480276
rect 361816 480264 361822 480276
rect 419166 480264 419172 480276
rect 361816 480236 419172 480264
rect 361816 480224 361822 480236
rect 419166 480224 419172 480236
rect 419224 480224 419230 480276
rect 361758 469208 361764 469260
rect 361816 469248 361822 469260
rect 396718 469248 396724 469260
rect 361816 469220 396724 469248
rect 361816 469208 361822 469220
rect 396718 469208 396724 469220
rect 396776 469208 396782 469260
rect 494698 462476 494704 462528
rect 494756 462516 494762 462528
rect 527634 462516 527640 462528
rect 494756 462488 527640 462516
rect 494756 462476 494762 462488
rect 527634 462476 527640 462488
rect 527692 462476 527698 462528
rect 453298 462408 453304 462460
rect 453356 462448 453362 462460
rect 524690 462448 524696 462460
rect 453356 462420 524696 462448
rect 453356 462408 453362 462420
rect 524690 462408 524696 462420
rect 524748 462408 524754 462460
rect 450538 462340 450544 462392
rect 450596 462380 450602 462392
rect 542354 462380 542360 462392
rect 450596 462352 542360 462380
rect 450596 462340 450602 462352
rect 542354 462340 542360 462352
rect 542412 462340 542418 462392
rect 467190 460980 467196 461032
rect 467248 461020 467254 461032
rect 553854 461020 553860 461032
rect 467248 460992 553860 461020
rect 467248 460980 467254 460992
rect 553854 460980 553860 460992
rect 553912 460980 553918 461032
rect 458910 460912 458916 460964
rect 458968 460952 458974 460964
rect 550910 460952 550916 460964
rect 458968 460924 550916 460952
rect 458968 460912 458974 460924
rect 550910 460912 550916 460924
rect 550968 460912 550974 460964
rect 447502 458804 447508 458856
rect 447560 458844 447566 458856
rect 483658 458844 483664 458856
rect 447560 458816 483664 458844
rect 447560 458804 447566 458816
rect 483658 458804 483664 458816
rect 483716 458804 483722 458856
rect 361758 458192 361764 458244
rect 361816 458232 361822 458244
rect 414658 458232 414664 458244
rect 361816 458204 414664 458232
rect 361816 458192 361822 458204
rect 414658 458192 414664 458204
rect 414716 458192 414722 458244
rect 569218 456764 569224 456816
rect 569276 456804 569282 456816
rect 580166 456804 580172 456816
rect 569276 456776 580172 456804
rect 569276 456764 569282 456776
rect 580166 456764 580172 456776
rect 580224 456764 580230 456816
rect 392578 456696 392584 456748
rect 392636 456736 392642 456748
rect 395338 456736 395344 456748
rect 392636 456708 395344 456736
rect 392636 456696 392642 456708
rect 395338 456696 395344 456708
rect 395396 456696 395402 456748
rect 488258 456016 488264 456068
rect 488316 456056 488322 456068
rect 494698 456056 494704 456068
rect 488316 456028 494704 456056
rect 488316 456016 488322 456028
rect 494698 456016 494704 456028
rect 494756 456016 494762 456068
rect 461762 455472 461768 455524
rect 461820 455512 461826 455524
rect 488258 455512 488264 455524
rect 461820 455484 488264 455512
rect 461820 455472 461826 455484
rect 488258 455472 488264 455484
rect 488316 455472 488322 455524
rect 452010 455404 452016 455456
rect 452068 455444 452074 455456
rect 480990 455444 480996 455456
rect 452068 455416 480996 455444
rect 452068 455404 452074 455416
rect 480990 455404 480996 455416
rect 481048 455404 481054 455456
rect 449710 454724 449716 454776
rect 449768 454764 449774 454776
rect 487154 454764 487160 454776
rect 449768 454736 487160 454764
rect 449768 454724 449774 454736
rect 487154 454724 487160 454736
rect 487212 454724 487218 454776
rect 449618 454656 449624 454708
rect 449676 454696 449682 454708
rect 489914 454696 489920 454708
rect 449676 454668 489920 454696
rect 449676 454656 449682 454668
rect 489914 454656 489920 454668
rect 489972 454656 489978 454708
rect 459002 454044 459008 454096
rect 459060 454084 459066 454096
rect 473722 454084 473728 454096
rect 459060 454056 473728 454084
rect 459060 454044 459066 454056
rect 473722 454044 473728 454056
rect 473780 454044 473786 454096
rect 447410 448468 447416 448520
rect 447468 448508 447474 448520
rect 458910 448508 458916 448520
rect 447468 448480 458916 448508
rect 447468 448468 447474 448480
rect 458910 448468 458916 448480
rect 458968 448468 458974 448520
rect 447226 447856 447232 447908
rect 447284 447896 447290 447908
rect 448330 447896 448336 447908
rect 447284 447868 448336 447896
rect 447284 447856 447290 447868
rect 448330 447856 448336 447868
rect 448388 447896 448394 447908
rect 459002 447896 459008 447908
rect 448388 447868 459008 447896
rect 448388 447856 448394 447868
rect 459002 447856 459008 447868
rect 459060 447856 459066 447908
rect 447134 447788 447140 447840
rect 447192 447828 447198 447840
rect 447962 447828 447968 447840
rect 447192 447800 447968 447828
rect 447192 447788 447198 447800
rect 447962 447788 447968 447800
rect 448020 447828 448026 447840
rect 467190 447828 467196 447840
rect 448020 447800 467196 447828
rect 448020 447788 448026 447800
rect 467190 447788 467196 447800
rect 467248 447788 467254 447840
rect 422478 447380 422484 447432
rect 422536 447420 422542 447432
rect 447226 447420 447232 447432
rect 422536 447392 447232 447420
rect 422536 447380 422542 447392
rect 447226 447380 447232 447392
rect 447284 447380 447290 447432
rect 437382 447312 437388 447364
rect 437440 447352 437446 447364
rect 447134 447352 447140 447364
rect 437440 447324 447140 447352
rect 437440 447312 437446 447324
rect 447134 447312 447140 447324
rect 447192 447312 447198 447364
rect 432414 447244 432420 447296
rect 432472 447284 432478 447296
rect 447410 447284 447416 447296
rect 432472 447256 447416 447284
rect 432472 447244 432478 447256
rect 447410 447244 447416 447256
rect 447468 447244 447474 447296
rect 427446 447176 427452 447228
rect 427504 447216 427510 447228
rect 445662 447216 445668 447228
rect 427504 447188 445668 447216
rect 427504 447176 427510 447188
rect 445662 447176 445668 447188
rect 445720 447176 445726 447228
rect 361758 447108 361764 447160
rect 361816 447148 361822 447160
rect 399478 447148 399484 447160
rect 361816 447120 399484 447148
rect 361816 447108 361822 447120
rect 399478 447108 399484 447120
rect 399536 447108 399542 447160
rect 442626 444320 442632 444372
rect 442684 444360 442690 444372
rect 446214 444360 446220 444372
rect 442684 444332 446220 444360
rect 442684 444320 442690 444332
rect 446214 444320 446220 444332
rect 446272 444320 446278 444372
rect 361758 436092 361764 436144
rect 361816 436132 361822 436144
rect 416130 436132 416136 436144
rect 361816 436104 416136 436132
rect 361816 436092 361822 436104
rect 416130 436092 416136 436104
rect 416188 436092 416194 436144
rect 395338 433236 395344 433288
rect 395396 433276 395402 433288
rect 398098 433276 398104 433288
rect 395396 433248 398104 433276
rect 395396 433236 395402 433248
rect 398098 433236 398104 433248
rect 398156 433236 398162 433288
rect 458082 429972 458088 430024
rect 458140 430012 458146 430024
rect 474274 430012 474280 430024
rect 458140 429984 474280 430012
rect 458140 429972 458146 429984
rect 474274 429972 474280 429984
rect 474332 429972 474338 430024
rect 459462 429904 459468 429956
rect 459520 429944 459526 429956
rect 476942 429944 476948 429956
rect 459520 429916 476948 429944
rect 459520 429904 459526 429916
rect 476942 429904 476948 429916
rect 477000 429904 477006 429956
rect 459370 429836 459376 429888
rect 459428 429876 459434 429888
rect 479610 429876 479616 429888
rect 459428 429848 479616 429876
rect 459428 429836 459434 429848
rect 479610 429836 479616 429848
rect 479668 429836 479674 429888
rect 480898 429156 480904 429208
rect 480956 429196 480962 429208
rect 482278 429196 482284 429208
rect 480956 429168 482284 429196
rect 480956 429156 480962 429168
rect 482278 429156 482284 429168
rect 482336 429156 482342 429208
rect 483658 429156 483664 429208
rect 483716 429196 483722 429208
rect 484946 429196 484952 429208
rect 483716 429168 484952 429196
rect 483716 429156 483722 429168
rect 484946 429156 484952 429168
rect 485004 429156 485010 429208
rect 457622 428408 457628 428460
rect 457680 428448 457686 428460
rect 471606 428448 471612 428460
rect 457680 428420 471612 428448
rect 457680 428408 457686 428420
rect 471606 428408 471612 428420
rect 471664 428408 471670 428460
rect 361758 425076 361764 425128
rect 361816 425116 361822 425128
rect 417418 425116 417424 425128
rect 361816 425088 417424 425116
rect 361816 425076 361822 425088
rect 417418 425076 417424 425088
rect 417476 425076 417482 425128
rect 503622 424328 503628 424380
rect 503680 424368 503686 424380
rect 557534 424368 557540 424380
rect 503680 424340 557540 424368
rect 503680 424328 503686 424340
rect 557534 424328 557540 424340
rect 557592 424328 557598 424380
rect 398098 423580 398104 423632
rect 398156 423620 398162 423632
rect 398834 423620 398840 423632
rect 398156 423592 398840 423620
rect 398156 423580 398162 423592
rect 398834 423580 398840 423592
rect 398892 423580 398898 423632
rect 529198 423580 529204 423632
rect 529256 423620 529262 423632
rect 530210 423620 530216 423632
rect 529256 423592 530216 423620
rect 529256 423580 529262 423592
rect 530210 423580 530216 423592
rect 530268 423580 530274 423632
rect 530578 423580 530584 423632
rect 530636 423620 530642 423632
rect 532786 423620 532792 423632
rect 530636 423592 532792 423620
rect 530636 423580 530642 423592
rect 532786 423580 532792 423592
rect 532844 423580 532850 423632
rect 511534 423512 511540 423564
rect 511592 423552 511598 423564
rect 523770 423552 523776 423564
rect 511592 423524 523776 423552
rect 511592 423512 511598 423524
rect 523770 423512 523776 423524
rect 523828 423512 523834 423564
rect 522298 423444 522304 423496
rect 522356 423484 522362 423496
rect 549530 423484 549536 423496
rect 522356 423456 549536 423484
rect 522356 423444 522362 423456
rect 549530 423444 549536 423456
rect 549588 423444 549594 423496
rect 502978 423376 502984 423428
rect 503036 423416 503042 423428
rect 522482 423416 522488 423428
rect 503036 423388 522488 423416
rect 503036 423376 503042 423388
rect 522482 423376 522488 423388
rect 522540 423376 522546 423428
rect 523678 423376 523684 423428
rect 523736 423416 523742 423428
rect 552106 423416 552112 423428
rect 523736 423388 552112 423416
rect 523736 423376 523742 423388
rect 552106 423376 552112 423388
rect 552164 423376 552170 423428
rect 487062 423308 487068 423360
rect 487120 423348 487126 423360
rect 526346 423348 526352 423360
rect 487120 423320 526352 423348
rect 487120 423308 487126 423320
rect 526346 423308 526352 423320
rect 526404 423308 526410 423360
rect 526438 423308 526444 423360
rect 526496 423348 526502 423360
rect 554682 423348 554688 423360
rect 526496 423320 554688 423348
rect 526496 423308 526502 423320
rect 554682 423308 554688 423320
rect 554740 423308 554746 423360
rect 488258 423240 488264 423292
rect 488316 423280 488322 423292
rect 528922 423280 528928 423292
rect 488316 423252 528928 423280
rect 488316 423240 488322 423252
rect 528922 423240 528928 423252
rect 528980 423240 528986 423292
rect 489638 423172 489644 423224
rect 489696 423212 489702 423224
rect 531498 423212 531504 423224
rect 489696 423184 531504 423212
rect 489696 423172 489702 423184
rect 531498 423172 531504 423184
rect 531556 423172 531562 423224
rect 498102 423104 498108 423156
rect 498160 423144 498166 423156
rect 545666 423144 545672 423156
rect 498160 423116 545672 423144
rect 498160 423104 498166 423116
rect 545666 423104 545672 423116
rect 545724 423104 545730 423156
rect 499298 423036 499304 423088
rect 499356 423076 499362 423088
rect 548242 423076 548248 423088
rect 499356 423048 548248 423076
rect 499356 423036 499362 423048
rect 548242 423036 548248 423048
rect 548300 423036 548306 423088
rect 444282 422968 444288 423020
rect 444340 423008 444346 423020
rect 447870 423008 447876 423020
rect 444340 422980 447876 423008
rect 444340 422968 444346 422980
rect 447870 422968 447876 422980
rect 447928 422968 447934 423020
rect 500678 422968 500684 423020
rect 500736 423008 500742 423020
rect 550818 423008 550824 423020
rect 500736 422980 550824 423008
rect 500736 422968 500742 422980
rect 550818 422968 550824 422980
rect 550876 422968 550882 423020
rect 502242 422900 502248 422952
rect 502300 422940 502306 422952
rect 553394 422940 553400 422952
rect 502300 422912 553400 422940
rect 502300 422900 502306 422912
rect 553394 422900 553400 422912
rect 553452 422900 553458 422952
rect 484302 421540 484308 421592
rect 484360 421580 484366 421592
rect 521194 421580 521200 421592
rect 484360 421552 521200 421580
rect 484360 421540 484366 421552
rect 521194 421540 521200 421552
rect 521252 421540 521258 421592
rect 495342 420180 495348 420232
rect 495400 420220 495406 420232
rect 541802 420220 541808 420232
rect 495400 420192 541808 420220
rect 495400 420180 495406 420192
rect 541802 420180 541808 420192
rect 541860 420180 541866 420232
rect 398834 418820 398840 418872
rect 398892 418860 398898 418872
rect 400674 418860 400680 418872
rect 398892 418832 400680 418860
rect 398892 418820 398898 418832
rect 400674 418820 400680 418832
rect 400732 418820 400738 418872
rect 425974 417732 425980 417784
rect 426032 417772 426038 417784
rect 507946 417772 507952 417784
rect 426032 417744 507952 417772
rect 426032 417732 426038 417744
rect 507946 417732 507952 417744
rect 508004 417732 508010 417784
rect 425330 417664 425336 417716
rect 425388 417704 425394 417716
rect 507854 417704 507860 417716
rect 425388 417676 507860 417704
rect 425388 417664 425394 417676
rect 507854 417664 507860 417676
rect 507912 417664 507918 417716
rect 422110 417596 422116 417648
rect 422168 417636 422174 417648
rect 503990 417636 503996 417648
rect 422168 417608 503996 417636
rect 422168 417596 422174 417608
rect 503990 417596 503996 417608
rect 504048 417596 504054 417648
rect 421466 417528 421472 417580
rect 421524 417568 421530 417580
rect 503714 417568 503720 417580
rect 421524 417540 503720 417568
rect 421524 417528 421530 417540
rect 503714 417528 503720 417540
rect 503772 417528 503778 417580
rect 424686 417460 424692 417512
rect 424744 417500 424750 417512
rect 506474 417500 506480 417512
rect 424744 417472 506480 417500
rect 424744 417460 424750 417472
rect 506474 417460 506480 417472
rect 506532 417460 506538 417512
rect 424042 417392 424048 417444
rect 424100 417432 424106 417444
rect 506566 417432 506572 417444
rect 424100 417404 506572 417432
rect 424100 417392 424106 417404
rect 506566 417392 506572 417404
rect 506624 417392 506630 417444
rect 423122 416304 423128 416356
rect 423180 416344 423186 416356
rect 423582 416344 423588 416356
rect 423180 416316 423588 416344
rect 423180 416304 423186 416316
rect 423582 416304 423588 416316
rect 423640 416304 423646 416356
rect 486970 416032 486976 416084
rect 487028 416072 487034 416084
rect 527634 416072 527640 416084
rect 487028 416044 527640 416072
rect 487028 416032 487034 416044
rect 527634 416032 527640 416044
rect 527692 416032 527698 416084
rect 361574 413992 361580 414044
rect 361632 414032 361638 414044
rect 443638 414032 443644 414044
rect 361632 414004 443644 414032
rect 361632 413992 361638 414004
rect 443638 413992 443644 414004
rect 443696 413992 443702 414044
rect 400674 413924 400680 413976
rect 400732 413964 400738 413976
rect 402330 413964 402336 413976
rect 400732 413936 402336 413964
rect 400732 413924 400738 413936
rect 402330 413924 402336 413936
rect 402388 413924 402394 413976
rect 402330 410524 402336 410576
rect 402388 410564 402394 410576
rect 409138 410564 409144 410576
rect 402388 410536 409144 410564
rect 402388 410524 402394 410536
rect 409138 410524 409144 410536
rect 409196 410524 409202 410576
rect 511442 404336 511448 404388
rect 511500 404376 511506 404388
rect 580166 404376 580172 404388
rect 511500 404348 580172 404376
rect 511500 404336 511506 404348
rect 580166 404336 580172 404348
rect 580224 404336 580230 404388
rect 361574 402976 361580 403028
rect 361632 403016 361638 403028
rect 439498 403016 439504 403028
rect 361632 402988 439504 403016
rect 361632 402976 361638 402988
rect 439498 402976 439504 402988
rect 439556 402976 439562 403028
rect 497918 400868 497924 400920
rect 497976 400908 497982 400920
rect 546494 400908 546500 400920
rect 497976 400880 546500 400908
rect 497976 400868 497982 400880
rect 546494 400868 546500 400880
rect 546552 400868 546558 400920
rect 494606 399440 494612 399492
rect 494664 399480 494670 399492
rect 539594 399480 539600 399492
rect 494664 399452 539600 399480
rect 494664 399440 494670 399452
rect 539594 399440 539600 399452
rect 539652 399440 539658 399492
rect 493962 398080 493968 398132
rect 494020 398120 494026 398132
rect 538214 398120 538220 398132
rect 494020 398092 538220 398120
rect 494020 398080 494026 398092
rect 538214 398080 538220 398092
rect 538272 398080 538278 398132
rect 493410 396720 493416 396772
rect 493468 396760 493474 396772
rect 536834 396760 536840 396772
rect 493468 396732 536840 396760
rect 493468 396720 493474 396732
rect 536834 396720 536840 396732
rect 536892 396720 536898 396772
rect 409138 396040 409144 396092
rect 409196 396080 409202 396092
rect 409196 396052 409920 396080
rect 409196 396040 409202 396052
rect 409892 396012 409920 396052
rect 411622 396012 411628 396024
rect 409892 395984 411628 396012
rect 411622 395972 411628 395984
rect 411680 395972 411686 396024
rect 460750 395292 460756 395344
rect 460808 395332 460814 395344
rect 483658 395332 483664 395344
rect 460808 395304 483664 395332
rect 460808 395292 460814 395304
rect 483658 395292 483664 395304
rect 483716 395292 483722 395344
rect 492398 395292 492404 395344
rect 492456 395332 492462 395344
rect 535454 395332 535460 395344
rect 492456 395304 535460 395332
rect 492456 395292 492462 395304
rect 535454 395292 535460 395304
rect 535512 395292 535518 395344
rect 496722 394000 496728 394052
rect 496780 394040 496786 394052
rect 543734 394040 543740 394052
rect 496780 394012 543740 394040
rect 496780 394000 496786 394012
rect 543734 394000 543740 394012
rect 543792 394000 543798 394052
rect 423490 393932 423496 393984
rect 423548 393972 423554 393984
rect 505554 393972 505560 393984
rect 423548 393944 505560 393972
rect 423548 393932 423554 393944
rect 505554 393932 505560 393944
rect 505612 393932 505618 393984
rect 463602 392572 463608 392624
rect 463660 392612 463666 392624
rect 487154 392612 487160 392624
rect 463660 392584 487160 392612
rect 463660 392572 463666 392584
rect 487154 392572 487160 392584
rect 487212 392572 487218 392624
rect 491570 392572 491576 392624
rect 491628 392612 491634 392624
rect 534166 392612 534172 392624
rect 491628 392584 534172 392612
rect 491628 392572 491634 392584
rect 534166 392572 534172 392584
rect 534224 392572 534230 392624
rect 361574 391960 361580 392012
rect 361632 392000 361638 392012
rect 443730 392000 443736 392012
rect 361632 391972 443736 392000
rect 361632 391960 361638 391972
rect 443730 391960 443736 391972
rect 443788 391960 443794 392012
rect 495710 391280 495716 391332
rect 495768 391320 495774 391332
rect 542354 391320 542360 391332
rect 495768 391292 542360 391320
rect 495768 391280 495774 391292
rect 542354 391280 542360 391292
rect 542412 391280 542418 391332
rect 411622 391212 411628 391264
rect 411680 391252 411686 391264
rect 415394 391252 415400 391264
rect 411680 391224 415400 391252
rect 411680 391212 411686 391224
rect 415394 391212 415400 391224
rect 415452 391212 415458 391264
rect 423582 391212 423588 391264
rect 423640 391252 423646 391264
rect 505278 391252 505284 391264
rect 423640 391224 505284 391252
rect 423640 391212 423646 391224
rect 505278 391212 505284 391224
rect 505336 391212 505342 391264
rect 459646 389852 459652 389904
rect 459704 389892 459710 389904
rect 480898 389892 480904 389904
rect 459704 389864 480904 389892
rect 459704 389852 459710 389864
rect 480898 389852 480904 389864
rect 480956 389852 480962 389904
rect 448054 389784 448060 389836
rect 448112 389824 448118 389836
rect 463142 389824 463148 389836
rect 448112 389796 463148 389824
rect 448112 389784 448118 389796
rect 463142 389784 463148 389796
rect 463200 389784 463206 389836
rect 464890 389784 464896 389836
rect 464948 389824 464954 389836
rect 489914 389824 489920 389836
rect 464948 389796 489920 389824
rect 464948 389784 464954 389796
rect 489914 389784 489920 389796
rect 489972 389784 489978 389836
rect 490558 389784 490564 389836
rect 490616 389824 490622 389836
rect 534074 389824 534080 389836
rect 490616 389796 534080 389824
rect 490616 389784 490622 389796
rect 534074 389784 534080 389796
rect 534132 389784 534138 389836
rect 458450 389240 458456 389292
rect 458508 389280 458514 389292
rect 459462 389280 459468 389292
rect 458508 389252 459468 389280
rect 458508 389240 458514 389252
rect 459462 389240 459468 389252
rect 459520 389240 459526 389292
rect 465074 389240 465080 389292
rect 465132 389280 465138 389292
rect 465902 389280 465908 389292
rect 465132 389252 465908 389280
rect 465132 389240 465138 389252
rect 465902 389240 465908 389252
rect 465960 389240 465966 389292
rect 466454 389240 466460 389292
rect 466512 389280 466518 389292
rect 467374 389280 467380 389292
rect 466512 389252 467380 389280
rect 466512 389240 466518 389252
rect 467374 389240 467380 389252
rect 467432 389240 467438 389292
rect 486418 389240 486424 389292
rect 486476 389280 486482 389292
rect 487062 389280 487068 389292
rect 486476 389252 487068 389280
rect 486476 389240 486482 389252
rect 487062 389240 487068 389252
rect 487120 389240 487126 389292
rect 497458 389240 497464 389292
rect 497516 389280 497522 389292
rect 498102 389280 498108 389292
rect 497516 389252 498108 389280
rect 497516 389240 497522 389252
rect 498102 389240 498108 389252
rect 498160 389240 498166 389292
rect 506474 389240 506480 389292
rect 506532 389280 506538 389292
rect 507118 389280 507124 389292
rect 506532 389252 507124 389280
rect 506532 389240 506538 389252
rect 507118 389240 507124 389252
rect 507176 389240 507182 389292
rect 415394 389104 415400 389156
rect 415452 389144 415458 389156
rect 417510 389144 417516 389156
rect 415452 389116 417516 389144
rect 415452 389104 415458 389116
rect 417510 389104 417516 389116
rect 417568 389104 417574 389156
rect 453022 389104 453028 389156
rect 453080 389144 453086 389156
rect 454034 389144 454040 389156
rect 453080 389116 454040 389144
rect 453080 389104 453086 389116
rect 454034 389104 454040 389116
rect 454092 389104 454098 389156
rect 456702 389104 456708 389156
rect 456760 389144 456766 389156
rect 457622 389144 457628 389156
rect 456760 389116 457628 389144
rect 456760 389104 456766 389116
rect 457622 389104 457628 389116
rect 457680 389104 457686 389156
rect 468478 389036 468484 389088
rect 468536 389076 468542 389088
rect 475838 389076 475844 389088
rect 468536 389048 475844 389076
rect 468536 389036 468542 389048
rect 475838 389036 475844 389048
rect 475896 389036 475902 389088
rect 468570 388968 468576 389020
rect 468628 389008 468634 389020
rect 478046 389008 478052 389020
rect 468628 388980 478052 389008
rect 468628 388968 468634 388980
rect 478046 388968 478052 388980
rect 478104 388968 478110 389020
rect 502334 388968 502340 389020
rect 502392 389008 502398 389020
rect 502392 388980 509234 389008
rect 502392 388968 502398 388980
rect 467098 388900 467104 388952
rect 467156 388940 467162 388952
rect 478782 388940 478788 388952
rect 467156 388912 478788 388940
rect 467156 388900 467162 388912
rect 478782 388900 478788 388912
rect 478840 388900 478846 388952
rect 461578 388832 461584 388884
rect 461636 388872 461642 388884
rect 473630 388872 473636 388884
rect 461636 388844 473636 388872
rect 461636 388832 461642 388844
rect 473630 388832 473636 388844
rect 473688 388832 473694 388884
rect 483934 388832 483940 388884
rect 483992 388872 483998 388884
rect 502978 388872 502984 388884
rect 483992 388844 502984 388872
rect 483992 388832 483998 388844
rect 502978 388832 502984 388844
rect 503036 388832 503042 388884
rect 509206 388872 509234 388980
rect 526438 388872 526444 388884
rect 509206 388844 526444 388872
rect 526438 388832 526444 388844
rect 526496 388832 526502 388884
rect 461118 388764 461124 388816
rect 461176 388804 461182 388816
rect 463602 388804 463608 388816
rect 461176 388776 463608 388804
rect 461176 388764 461182 388776
rect 463602 388764 463608 388776
rect 463660 388764 463666 388816
rect 464338 388764 464344 388816
rect 464396 388804 464402 388816
rect 476574 388804 476580 388816
rect 464396 388776 476580 388804
rect 464396 388764 464402 388776
rect 476574 388764 476580 388776
rect 476632 388764 476638 388816
rect 500862 388764 500868 388816
rect 500920 388804 500926 388816
rect 523678 388804 523684 388816
rect 500920 388776 523684 388804
rect 500920 388764 500926 388776
rect 523678 388764 523684 388776
rect 523736 388764 523742 388816
rect 462958 388696 462964 388748
rect 463016 388736 463022 388748
rect 475102 388736 475108 388748
rect 463016 388708 475108 388736
rect 463016 388696 463022 388708
rect 475102 388696 475108 388708
rect 475160 388696 475166 388748
rect 499390 388696 499396 388748
rect 499448 388736 499454 388748
rect 522298 388736 522304 388748
rect 499448 388708 522304 388736
rect 499448 388696 499454 388708
rect 522298 388696 522304 388708
rect 522356 388696 522362 388748
rect 468662 388628 468668 388680
rect 468720 388668 468726 388680
rect 481726 388668 481732 388680
rect 468720 388640 481732 388668
rect 468720 388628 468726 388640
rect 481726 388628 481732 388640
rect 481784 388628 481790 388680
rect 484670 388628 484676 388680
rect 484728 388668 484734 388680
rect 511534 388668 511540 388680
rect 484728 388640 511540 388668
rect 484728 388628 484734 388640
rect 511534 388628 511540 388640
rect 511592 388628 511598 388680
rect 447778 388560 447784 388612
rect 447836 388600 447842 388612
rect 457438 388600 457444 388612
rect 447836 388572 457444 388600
rect 447836 388560 447842 388572
rect 457438 388560 457444 388572
rect 457496 388560 457502 388612
rect 465718 388560 465724 388612
rect 465776 388600 465782 388612
rect 480254 388600 480260 388612
rect 465776 388572 480260 388600
rect 465776 388560 465782 388572
rect 480254 388560 480260 388572
rect 480312 388560 480318 388612
rect 485406 388560 485412 388612
rect 485464 388600 485470 388612
rect 524414 388600 524420 388612
rect 485464 388572 524420 388600
rect 485464 388560 485470 388572
rect 524414 388560 524420 388572
rect 524472 388560 524478 388612
rect 447686 388492 447692 388544
rect 447744 388532 447750 388544
rect 457530 388532 457536 388544
rect 447744 388504 457536 388532
rect 447744 388492 447750 388504
rect 457530 388492 457536 388504
rect 457588 388492 457594 388544
rect 464522 388492 464528 388544
rect 464580 388532 464586 388544
rect 480990 388532 480996 388544
rect 464580 388504 480996 388532
rect 464580 388492 464586 388504
rect 480990 388492 480996 388504
rect 481048 388492 481054 388544
rect 488350 388492 488356 388544
rect 488408 388532 488414 388544
rect 529198 388532 529204 388544
rect 488408 388504 529204 388532
rect 488408 388492 488414 388504
rect 529198 388492 529204 388504
rect 529256 388492 529262 388544
rect 450722 388424 450728 388476
rect 450780 388464 450786 388476
rect 461762 388464 461768 388476
rect 450780 388436 461768 388464
rect 450780 388424 450786 388436
rect 461762 388424 461768 388436
rect 461820 388424 461826 388476
rect 463050 388424 463056 388476
rect 463108 388464 463114 388476
rect 482462 388464 482468 388476
rect 463108 388436 482468 388464
rect 463108 388424 463114 388436
rect 482462 388424 482468 388436
rect 482520 388424 482526 388476
rect 489822 388424 489828 388476
rect 489880 388464 489886 388476
rect 530578 388464 530584 388476
rect 489880 388436 530584 388464
rect 489880 388424 489886 388436
rect 530578 388424 530584 388436
rect 530636 388424 530642 388476
rect 461670 387880 461676 387932
rect 461728 387920 461734 387932
rect 462590 387920 462596 387932
rect 461728 387892 462596 387920
rect 461728 387880 461734 387892
rect 462590 387880 462596 387892
rect 462648 387880 462654 387932
rect 461854 387812 461860 387864
rect 461912 387852 461918 387864
rect 464890 387852 464896 387864
rect 461912 387824 464896 387852
rect 461912 387812 461918 387824
rect 464890 387812 464896 387824
rect 464948 387812 464954 387864
rect 447870 387200 447876 387252
rect 447928 387240 447934 387252
rect 458818 387240 458824 387252
rect 447928 387212 458824 387240
rect 447928 387200 447934 387212
rect 458818 387200 458824 387212
rect 458876 387200 458882 387252
rect 448974 387132 448980 387184
rect 449032 387172 449038 387184
rect 491294 387172 491300 387184
rect 449032 387144 491300 387172
rect 449032 387132 449038 387144
rect 491294 387132 491300 387144
rect 491352 387132 491358 387184
rect 449526 387064 449532 387116
rect 449584 387104 449590 387116
rect 513374 387104 513380 387116
rect 449584 387076 513380 387104
rect 449584 387064 449590 387076
rect 513374 387064 513380 387076
rect 513432 387064 513438 387116
rect 448330 386656 448336 386708
rect 448388 386696 448394 386708
rect 553946 386696 553952 386708
rect 448388 386668 553952 386696
rect 448388 386656 448394 386668
rect 553946 386656 553952 386668
rect 554004 386656 554010 386708
rect 381538 386588 381544 386640
rect 381596 386628 381602 386640
rect 512086 386628 512092 386640
rect 381596 386600 512092 386628
rect 381596 386588 381602 386600
rect 512086 386588 512092 386600
rect 512144 386588 512150 386640
rect 378778 386520 378784 386572
rect 378836 386560 378842 386572
rect 512546 386560 512552 386572
rect 378836 386532 512552 386560
rect 378836 386520 378842 386532
rect 512546 386520 512552 386532
rect 512604 386520 512610 386572
rect 367738 386452 367744 386504
rect 367796 386492 367802 386504
rect 511994 386492 512000 386504
rect 367796 386464 512000 386492
rect 367796 386452 367802 386464
rect 511994 386452 512000 386464
rect 512052 386452 512058 386504
rect 367830 386384 367836 386436
rect 367888 386424 367894 386436
rect 512270 386424 512276 386436
rect 367888 386396 512276 386424
rect 367888 386384 367894 386396
rect 512270 386384 512276 386396
rect 512328 386384 512334 386436
rect 448238 385976 448244 386028
rect 448296 386016 448302 386028
rect 453298 386016 453304 386028
rect 448296 385988 453304 386016
rect 448296 385976 448302 385988
rect 453298 385976 453304 385988
rect 453356 385976 453362 386028
rect 448422 385636 448428 385688
rect 448480 385676 448486 385688
rect 454402 385676 454408 385688
rect 448480 385648 454408 385676
rect 448480 385636 448486 385648
rect 454402 385636 454408 385648
rect 454460 385636 454466 385688
rect 448146 385364 448152 385416
rect 448204 385404 448210 385416
rect 452010 385404 452016 385416
rect 448204 385376 452016 385404
rect 448204 385364 448210 385376
rect 452010 385364 452016 385376
rect 452068 385364 452074 385416
rect 449434 385092 449440 385144
rect 449492 385132 449498 385144
rect 563422 385132 563428 385144
rect 449492 385104 563428 385132
rect 449492 385092 449498 385104
rect 563422 385092 563428 385104
rect 563480 385092 563486 385144
rect 367922 385024 367928 385076
rect 367980 385064 367986 385076
rect 512362 385064 512368 385076
rect 367980 385036 512368 385064
rect 367980 385024 367986 385036
rect 512362 385024 512368 385036
rect 512420 385024 512426 385076
rect 513190 383732 513196 383784
rect 513248 383772 513254 383784
rect 534718 383772 534724 383784
rect 513248 383744 534724 383772
rect 513248 383732 513254 383744
rect 534718 383732 534724 383744
rect 534776 383732 534782 383784
rect 513282 383664 513288 383716
rect 513340 383704 513346 383716
rect 548518 383704 548524 383716
rect 513340 383676 548524 383704
rect 513340 383664 513346 383676
rect 548518 383664 548524 383676
rect 548576 383664 548582 383716
rect 362218 383596 362224 383648
rect 362276 383636 362282 383648
rect 447134 383636 447140 383648
rect 362276 383608 447140 383636
rect 362276 383596 362282 383608
rect 447134 383596 447140 383608
rect 447192 383596 447198 383648
rect 378870 383528 378876 383580
rect 378928 383568 378934 383580
rect 447226 383568 447232 383580
rect 378928 383540 447232 383568
rect 378928 383528 378934 383540
rect 447226 383528 447232 383540
rect 447284 383528 447290 383580
rect 512638 382916 512644 382968
rect 512696 382956 512702 382968
rect 519722 382956 519728 382968
rect 512696 382928 519728 382956
rect 512696 382916 512702 382928
rect 519722 382916 519728 382928
rect 519780 382916 519786 382968
rect 513006 382712 513012 382764
rect 513064 382752 513070 382764
rect 518342 382752 518348 382764
rect 513064 382724 518348 382752
rect 513064 382712 513070 382724
rect 518342 382712 518348 382724
rect 518400 382712 518406 382764
rect 512454 382440 512460 382492
rect 512512 382480 512518 382492
rect 515582 382480 515588 382492
rect 512512 382452 515588 382480
rect 512512 382440 512518 382452
rect 515582 382440 515588 382452
rect 515640 382440 515646 382492
rect 374638 382168 374644 382220
rect 374696 382208 374702 382220
rect 447226 382208 447232 382220
rect 374696 382180 447232 382208
rect 374696 382168 374702 382180
rect 447226 382168 447232 382180
rect 447284 382168 447290 382220
rect 376018 382100 376024 382152
rect 376076 382140 376082 382152
rect 447134 382140 447140 382152
rect 376076 382112 447140 382140
rect 376076 382100 376082 382112
rect 447134 382100 447140 382112
rect 447192 382100 447198 382152
rect 361574 380876 361580 380928
rect 361632 380916 361638 380928
rect 443822 380916 443828 380928
rect 361632 380888 443828 380916
rect 361632 380876 361638 380888
rect 443822 380876 443828 380888
rect 443880 380876 443886 380928
rect 512454 380876 512460 380928
rect 512512 380916 512518 380928
rect 547138 380916 547144 380928
rect 512512 380888 547144 380916
rect 512512 380876 512518 380888
rect 547138 380876 547144 380888
rect 547196 380876 547202 380928
rect 363598 380808 363604 380860
rect 363656 380848 363662 380860
rect 447410 380848 447416 380860
rect 363656 380820 447416 380848
rect 363656 380808 363662 380820
rect 447410 380808 447416 380820
rect 447468 380808 447474 380860
rect 371878 380740 371884 380792
rect 371936 380780 371942 380792
rect 447134 380780 447140 380792
rect 371936 380752 447140 380780
rect 371936 380740 371942 380752
rect 447134 380740 447140 380752
rect 447192 380740 447198 380792
rect 400858 380672 400864 380724
rect 400916 380712 400922 380724
rect 447226 380712 447232 380724
rect 400916 380684 447232 380712
rect 400916 380672 400922 380684
rect 447226 380672 447232 380684
rect 447284 380672 447290 380724
rect 512546 379720 512552 379772
rect 512604 379760 512610 379772
rect 515674 379760 515680 379772
rect 512604 379732 515680 379760
rect 512604 379720 512610 379732
rect 515674 379720 515680 379732
rect 515732 379720 515738 379772
rect 513282 379516 513288 379568
rect 513340 379556 513346 379568
rect 549898 379556 549904 379568
rect 513340 379528 549904 379556
rect 513340 379516 513346 379528
rect 549898 379516 549904 379528
rect 549956 379516 549962 379568
rect 363690 379448 363696 379500
rect 363748 379488 363754 379500
rect 447318 379488 447324 379500
rect 363748 379460 447324 379488
rect 363748 379448 363754 379460
rect 447318 379448 447324 379460
rect 447376 379448 447382 379500
rect 370498 379380 370504 379432
rect 370556 379420 370562 379432
rect 447134 379420 447140 379432
rect 370556 379392 447140 379420
rect 370556 379380 370562 379392
rect 447134 379380 447140 379392
rect 447192 379380 447198 379432
rect 417510 378904 417516 378956
rect 417568 378944 417574 378956
rect 419258 378944 419264 378956
rect 417568 378916 419264 378944
rect 417568 378904 417574 378916
rect 419258 378904 419264 378916
rect 419316 378904 419322 378956
rect 513282 378292 513288 378344
rect 513340 378332 513346 378344
rect 522298 378332 522304 378344
rect 513340 378304 522304 378332
rect 513340 378292 513346 378304
rect 522298 378292 522304 378304
rect 522356 378292 522362 378344
rect 512822 378224 512828 378276
rect 512880 378264 512886 378276
rect 547230 378264 547236 378276
rect 512880 378236 547236 378264
rect 512880 378224 512886 378236
rect 547230 378224 547236 378236
rect 547288 378224 547294 378276
rect 514018 378156 514024 378208
rect 514076 378196 514082 378208
rect 580166 378196 580172 378208
rect 514076 378168 580172 378196
rect 514076 378156 514082 378168
rect 580166 378156 580172 378168
rect 580224 378156 580230 378208
rect 363782 378088 363788 378140
rect 363840 378128 363846 378140
rect 447226 378128 447232 378140
rect 363840 378100 447232 378128
rect 363840 378088 363846 378100
rect 447226 378088 447232 378100
rect 447284 378088 447290 378140
rect 368014 378020 368020 378072
rect 368072 378060 368078 378072
rect 447134 378060 447140 378072
rect 368072 378032 447140 378060
rect 368072 378020 368078 378032
rect 447134 378020 447140 378032
rect 447192 378020 447198 378072
rect 513190 377408 513196 377460
rect 513248 377448 513254 377460
rect 548610 377448 548616 377460
rect 513248 377420 548616 377448
rect 513248 377408 513254 377420
rect 548610 377408 548616 377420
rect 548668 377408 548674 377460
rect 513190 376728 513196 376780
rect 513248 376768 513254 376780
rect 516962 376768 516968 376780
rect 513248 376740 516968 376768
rect 513248 376728 513254 376740
rect 516962 376728 516968 376740
rect 517020 376728 517026 376780
rect 403618 376660 403624 376712
rect 403676 376700 403682 376712
rect 447134 376700 447140 376712
rect 403676 376672 447140 376700
rect 403676 376660 403682 376672
rect 447134 376660 447140 376672
rect 447192 376660 447198 376712
rect 419074 376592 419080 376644
rect 419132 376632 419138 376644
rect 447226 376632 447232 376644
rect 419132 376604 447232 376632
rect 419132 376592 419138 376604
rect 447226 376592 447232 376604
rect 447284 376592 447290 376644
rect 513006 375980 513012 376032
rect 513064 376020 513070 376032
rect 544378 376020 544384 376032
rect 513064 375992 544384 376020
rect 513064 375980 513070 375992
rect 544378 375980 544384 375992
rect 544436 375980 544442 376032
rect 406378 375300 406384 375352
rect 406436 375340 406442 375352
rect 447134 375340 447140 375352
rect 406436 375312 447140 375340
rect 406436 375300 406442 375312
rect 447134 375300 447140 375312
rect 447192 375300 447198 375352
rect 407758 375232 407764 375284
rect 407816 375272 407822 375284
rect 447226 375272 447232 375284
rect 407816 375244 447232 375272
rect 407816 375232 407822 375244
rect 447226 375232 447232 375244
rect 447284 375232 447290 375284
rect 513282 374144 513288 374196
rect 513340 374184 513346 374196
rect 517514 374184 517520 374196
rect 513340 374156 517520 374184
rect 513340 374144 513346 374156
rect 517514 374144 517520 374156
rect 517572 374144 517578 374196
rect 410518 373940 410524 373992
rect 410576 373980 410582 373992
rect 447134 373980 447140 373992
rect 410576 373952 447140 373980
rect 410576 373940 410582 373952
rect 447134 373940 447140 373952
rect 447192 373940 447198 373992
rect 411898 373872 411904 373924
rect 411956 373912 411962 373924
rect 447226 373912 447232 373924
rect 411956 373884 447232 373912
rect 411956 373872 411962 373884
rect 447226 373872 447232 373884
rect 447284 373872 447290 373924
rect 513282 372648 513288 372700
rect 513340 372688 513346 372700
rect 518894 372688 518900 372700
rect 513340 372660 518900 372688
rect 513340 372648 513346 372660
rect 518894 372648 518900 372660
rect 518952 372648 518958 372700
rect 512638 372580 512644 372632
rect 512696 372620 512702 372632
rect 521654 372620 521660 372632
rect 512696 372592 521660 372620
rect 512696 372580 512702 372592
rect 521654 372580 521660 372592
rect 521712 372580 521718 372632
rect 381630 372512 381636 372564
rect 381688 372552 381694 372564
rect 447134 372552 447140 372564
rect 381688 372524 447140 372552
rect 381688 372512 381694 372524
rect 447134 372512 447140 372524
rect 447192 372512 447198 372564
rect 419166 372444 419172 372496
rect 419224 372484 419230 372496
rect 447226 372484 447232 372496
rect 419224 372456 447232 372484
rect 419224 372444 419230 372456
rect 447226 372444 447232 372456
rect 447284 372444 447290 372496
rect 511994 371696 512000 371748
rect 512052 371736 512058 371748
rect 513834 371736 513840 371748
rect 512052 371708 513840 371736
rect 512052 371696 512058 371708
rect 513834 371696 513840 371708
rect 513892 371696 513898 371748
rect 396718 371152 396724 371204
rect 396776 371192 396782 371204
rect 447134 371192 447140 371204
rect 396776 371164 447140 371192
rect 396776 371152 396782 371164
rect 447134 371152 447140 371164
rect 447192 371152 447198 371204
rect 414658 371084 414664 371136
rect 414716 371124 414722 371136
rect 447226 371124 447232 371136
rect 414716 371096 447232 371124
rect 414716 371084 414722 371096
rect 447226 371084 447232 371096
rect 447284 371084 447290 371136
rect 512086 370200 512092 370252
rect 512144 370240 512150 370252
rect 514754 370240 514760 370252
rect 512144 370212 514760 370240
rect 512144 370200 512150 370212
rect 514754 370200 514760 370212
rect 514812 370200 514818 370252
rect 513282 370064 513288 370116
rect 513340 370104 513346 370116
rect 517606 370104 517612 370116
rect 513340 370076 517612 370104
rect 513340 370064 513346 370076
rect 517606 370064 517612 370076
rect 517664 370064 517670 370116
rect 361574 369860 361580 369912
rect 361632 369900 361638 369912
rect 409874 369900 409880 369912
rect 361632 369872 409880 369900
rect 361632 369860 361638 369872
rect 409874 369860 409880 369872
rect 409932 369860 409938 369912
rect 513282 369860 513288 369912
rect 513340 369900 513346 369912
rect 523034 369900 523040 369912
rect 513340 369872 523040 369900
rect 513340 369860 513346 369872
rect 523034 369860 523040 369872
rect 523092 369860 523098 369912
rect 399478 369792 399484 369844
rect 399536 369832 399542 369844
rect 447134 369832 447140 369844
rect 399536 369804 447140 369832
rect 399536 369792 399542 369804
rect 447134 369792 447140 369804
rect 447192 369792 447198 369844
rect 416130 369724 416136 369776
rect 416188 369764 416194 369776
rect 447226 369764 447232 369776
rect 416188 369736 447232 369764
rect 416188 369724 416194 369736
rect 447226 369724 447232 369736
rect 447284 369724 447290 369776
rect 419258 369316 419264 369368
rect 419316 369356 419322 369368
rect 421558 369356 421564 369368
rect 419316 369328 421564 369356
rect 419316 369316 419322 369328
rect 421558 369316 421564 369328
rect 421616 369316 421622 369368
rect 512086 369112 512092 369164
rect 512144 369152 512150 369164
rect 520274 369152 520280 369164
rect 512144 369124 520280 369152
rect 512144 369112 512150 369124
rect 520274 369112 520280 369124
rect 520332 369112 520338 369164
rect 512270 368568 512276 368620
rect 512328 368608 512334 368620
rect 515122 368608 515128 368620
rect 512328 368580 515128 368608
rect 512328 368568 512334 368580
rect 515122 368568 515128 368580
rect 515180 368568 515186 368620
rect 417418 368432 417424 368484
rect 417476 368472 417482 368484
rect 447134 368472 447140 368484
rect 417476 368444 447140 368472
rect 417476 368432 417482 368444
rect 447134 368432 447140 368444
rect 447192 368432 447198 368484
rect 443638 368364 443644 368416
rect 443696 368404 443702 368416
rect 447226 368404 447232 368416
rect 443696 368376 447232 368404
rect 443696 368364 443702 368376
rect 447226 368364 447232 368376
rect 447284 368364 447290 368416
rect 513282 367344 513288 367396
rect 513340 367384 513346 367396
rect 520366 367384 520372 367396
rect 513340 367356 520372 367384
rect 513340 367344 513346 367356
rect 520366 367344 520372 367356
rect 520424 367344 520430 367396
rect 439498 367004 439504 367056
rect 439556 367044 439562 367056
rect 447134 367044 447140 367056
rect 439556 367016 447140 367044
rect 439556 367004 439562 367016
rect 447134 367004 447140 367016
rect 447192 367004 447198 367056
rect 443730 366936 443736 366988
rect 443788 366976 443794 366988
rect 447226 366976 447232 366988
rect 443788 366948 447232 366976
rect 443788 366936 443794 366948
rect 447226 366936 447232 366948
rect 447284 366936 447290 366988
rect 513282 365712 513288 365764
rect 513340 365752 513346 365764
rect 521746 365752 521752 365764
rect 513340 365724 521752 365752
rect 513340 365712 513346 365724
rect 521746 365712 521752 365724
rect 521804 365712 521810 365764
rect 409874 365644 409880 365696
rect 409932 365684 409938 365696
rect 447134 365684 447140 365696
rect 409932 365656 447140 365684
rect 409932 365644 409938 365656
rect 447134 365644 447140 365656
rect 447192 365644 447198 365696
rect 443822 365576 443828 365628
rect 443880 365616 443886 365628
rect 447226 365616 447232 365628
rect 443880 365588 447232 365616
rect 443880 365576 443886 365588
rect 447226 365576 447232 365588
rect 447284 365576 447290 365628
rect 511994 365576 512000 365628
rect 512052 365616 512058 365628
rect 514202 365616 514208 365628
rect 512052 365588 514208 365616
rect 512052 365576 512058 365588
rect 514202 365576 514208 365588
rect 514260 365576 514266 365628
rect 513282 365032 513288 365084
rect 513340 365072 513346 365084
rect 519078 365072 519084 365084
rect 513340 365044 519084 365072
rect 513340 365032 513346 365044
rect 519078 365032 519084 365044
rect 519136 365032 519142 365084
rect 512822 364352 512828 364404
rect 512880 364392 512886 364404
rect 518986 364392 518992 364404
rect 512880 364364 518992 364392
rect 512880 364352 512886 364364
rect 518986 364352 518992 364364
rect 519044 364352 519050 364404
rect 573358 364352 573364 364404
rect 573416 364392 573422 364404
rect 580166 364392 580172 364404
rect 573416 364364 580172 364392
rect 573416 364352 573422 364364
rect 580166 364352 580172 364364
rect 580224 364352 580230 364404
rect 511994 363196 512000 363248
rect 512052 363236 512058 363248
rect 514846 363236 514852 363248
rect 512052 363208 514852 363236
rect 512052 363196 512058 363208
rect 514846 363196 514852 363208
rect 514904 363196 514910 363248
rect 432874 362992 432880 363044
rect 432932 363032 432938 363044
rect 447226 363032 447232 363044
rect 432932 363004 447232 363032
rect 432932 362992 432938 363004
rect 447226 362992 447232 363004
rect 447284 362992 447290 363044
rect 432782 362924 432788 362976
rect 432840 362964 432846 362976
rect 447134 362964 447140 362976
rect 432840 362936 447140 362964
rect 432840 362924 432846 362936
rect 447134 362924 447140 362936
rect 447192 362924 447198 362976
rect 421558 362448 421564 362500
rect 421616 362488 421622 362500
rect 423582 362488 423588 362500
rect 421616 362460 423588 362488
rect 421616 362448 421622 362460
rect 423582 362448 423588 362460
rect 423640 362448 423646 362500
rect 511994 362312 512000 362364
rect 512052 362352 512058 362364
rect 513650 362352 513656 362364
rect 512052 362324 513656 362352
rect 512052 362312 512058 362324
rect 513650 362312 513656 362324
rect 513708 362312 513714 362364
rect 442258 361632 442264 361684
rect 442316 361672 442322 361684
rect 447226 361672 447232 361684
rect 442316 361644 447232 361672
rect 442316 361632 442322 361644
rect 447226 361632 447232 361644
rect 447284 361632 447290 361684
rect 513006 361632 513012 361684
rect 513064 361672 513070 361684
rect 519170 361672 519176 361684
rect 513064 361644 519176 361672
rect 513064 361632 513070 361644
rect 519170 361632 519176 361644
rect 519228 361632 519234 361684
rect 432690 361564 432696 361616
rect 432748 361604 432754 361616
rect 447134 361604 447140 361616
rect 432748 361576 447140 361604
rect 432748 361564 432754 361576
rect 447134 361564 447140 361576
rect 447192 361564 447198 361616
rect 513282 361564 513288 361616
rect 513340 361604 513346 361616
rect 523126 361604 523132 361616
rect 513340 361576 523132 361604
rect 513340 361564 513346 361576
rect 523126 361564 523132 361576
rect 523184 361564 523190 361616
rect 512638 360680 512644 360732
rect 512696 360720 512702 360732
rect 520550 360720 520556 360732
rect 512696 360692 520556 360720
rect 512696 360680 512702 360692
rect 520550 360680 520556 360692
rect 520608 360680 520614 360732
rect 511994 360408 512000 360460
rect 512052 360448 512058 360460
rect 514938 360448 514944 360460
rect 512052 360420 514944 360448
rect 512052 360408 512058 360420
rect 514938 360408 514944 360420
rect 514996 360408 515002 360460
rect 439682 360272 439688 360324
rect 439740 360312 439746 360324
rect 447226 360312 447232 360324
rect 439740 360284 447232 360312
rect 439740 360272 439746 360284
rect 447226 360272 447232 360284
rect 447284 360272 447290 360324
rect 436922 360204 436928 360256
rect 436980 360244 436986 360256
rect 447134 360244 447140 360256
rect 436980 360216 447140 360244
rect 436980 360204 436986 360216
rect 447134 360204 447140 360216
rect 447192 360204 447198 360256
rect 547230 360136 547236 360188
rect 547288 360176 547294 360188
rect 552014 360176 552020 360188
rect 547288 360148 552020 360176
rect 547288 360136 547294 360148
rect 552014 360136 552020 360148
rect 552072 360136 552078 360188
rect 534718 360068 534724 360120
rect 534776 360108 534782 360120
rect 566734 360108 566740 360120
rect 534776 360080 566740 360108
rect 534776 360068 534782 360080
rect 566734 360068 566740 360080
rect 566792 360068 566798 360120
rect 549898 360000 549904 360052
rect 549956 360040 549962 360052
rect 554958 360040 554964 360052
rect 549956 360012 554964 360040
rect 549956 360000 549962 360012
rect 554958 360000 554964 360012
rect 555016 360000 555022 360052
rect 548518 359932 548524 359984
rect 548576 359972 548582 359984
rect 565262 359972 565268 359984
rect 548576 359944 565268 359972
rect 548576 359932 548582 359944
rect 565262 359932 565268 359944
rect 565320 359932 565326 359984
rect 547138 359864 547144 359916
rect 547196 359904 547202 359916
rect 558178 359904 558184 359916
rect 547196 359876 558184 359904
rect 547196 359864 547202 359876
rect 558178 359864 558184 359876
rect 558236 359864 558242 359916
rect 515674 359796 515680 359848
rect 515732 359836 515738 359848
rect 553762 359836 553768 359848
rect 515732 359808 553768 359836
rect 515732 359796 515738 359808
rect 553762 359796 553768 359808
rect 553820 359796 553826 359848
rect 522298 359728 522304 359780
rect 522356 359768 522362 359780
rect 550818 359768 550824 359780
rect 522356 359740 550824 359768
rect 522356 359728 522362 359740
rect 550818 359728 550824 359740
rect 550876 359728 550882 359780
rect 443822 358844 443828 358896
rect 443880 358884 443886 358896
rect 447226 358884 447232 358896
rect 443880 358856 447232 358884
rect 443880 358844 443886 358856
rect 447226 358844 447232 358856
rect 447284 358844 447290 358896
rect 435450 358776 435456 358828
rect 435508 358816 435514 358828
rect 447134 358816 447140 358828
rect 435508 358788 447140 358816
rect 435508 358776 435514 358788
rect 447134 358776 447140 358788
rect 447192 358776 447198 358828
rect 513006 358776 513012 358828
rect 513064 358816 513070 358828
rect 519262 358816 519268 358828
rect 513064 358788 519268 358816
rect 513064 358776 513070 358788
rect 519262 358776 519268 358788
rect 519320 358776 519326 358828
rect 548610 358708 548616 358760
rect 548668 358748 548674 358760
rect 556706 358748 556712 358760
rect 548668 358720 556712 358748
rect 548668 358708 548674 358720
rect 556706 358708 556712 358720
rect 556764 358708 556770 358760
rect 519722 358640 519728 358692
rect 519780 358680 519786 358692
rect 564066 358680 564072 358692
rect 519780 358652 564072 358680
rect 519780 358640 519786 358652
rect 564066 358640 564072 358652
rect 564124 358640 564130 358692
rect 518342 358572 518348 358624
rect 518400 358612 518406 358624
rect 562594 358612 562600 358624
rect 518400 358584 562600 358612
rect 518400 358572 518406 358584
rect 562594 358572 562600 358584
rect 562652 358572 562658 358624
rect 544378 358504 544384 358556
rect 544436 358544 544442 358556
rect 559650 358544 559656 358556
rect 544436 358516 559656 358544
rect 544436 358504 544442 358516
rect 559650 358504 559656 358516
rect 559708 358504 559714 358556
rect 515582 358436 515588 358488
rect 515640 358476 515646 358488
rect 561122 358476 561128 358488
rect 515640 358448 561128 358476
rect 515640 358436 515646 358448
rect 561122 358436 561128 358448
rect 561180 358436 561186 358488
rect 423582 357416 423588 357468
rect 423640 357456 423646 357468
rect 423640 357428 423720 357456
rect 423640 357416 423646 357428
rect 423692 357388 423720 357428
rect 426342 357388 426348 357400
rect 423692 357360 426348 357388
rect 426342 357348 426348 357360
rect 426400 357348 426406 357400
rect 512822 356328 512828 356380
rect 512880 356368 512886 356380
rect 516226 356368 516232 356380
rect 512880 356340 516232 356368
rect 512880 356328 512886 356340
rect 516226 356328 516232 356340
rect 516284 356328 516290 356380
rect 513282 356192 513288 356244
rect 513340 356232 513346 356244
rect 520458 356232 520464 356244
rect 513340 356204 520464 356232
rect 513340 356192 513346 356204
rect 520458 356192 520464 356204
rect 520516 356192 520522 356244
rect 513282 354968 513288 355020
rect 513340 355008 513346 355020
rect 517698 355008 517704 355020
rect 513340 354980 517704 355008
rect 513340 354968 513346 354980
rect 517698 354968 517704 354980
rect 517756 354968 517762 355020
rect 513282 354696 513288 354748
rect 513340 354736 513346 354748
rect 517882 354736 517888 354748
rect 513340 354708 517888 354736
rect 513340 354696 513346 354708
rect 517882 354696 517888 354708
rect 517940 354696 517946 354748
rect 512086 354152 512092 354204
rect 512144 354192 512150 354204
rect 513742 354192 513748 354204
rect 512144 354164 513748 354192
rect 512144 354152 512150 354164
rect 513742 354152 513748 354164
rect 513800 354152 513806 354204
rect 445662 353948 445668 354000
rect 445720 353988 445726 354000
rect 448422 353988 448428 354000
rect 445720 353960 448428 353988
rect 445720 353948 445726 353960
rect 448422 353948 448428 353960
rect 448480 353948 448486 354000
rect 513282 353472 513288 353524
rect 513340 353512 513346 353524
rect 517790 353512 517796 353524
rect 513340 353484 517796 353512
rect 513340 353472 513346 353484
rect 517790 353472 517796 353484
rect 517848 353472 517854 353524
rect 446214 352520 446220 352572
rect 446272 352560 446278 352572
rect 447778 352560 447784 352572
rect 446272 352532 447784 352560
rect 446272 352520 446278 352532
rect 447778 352520 447784 352532
rect 447836 352520 447842 352572
rect 512454 352248 512460 352300
rect 512512 352288 512518 352300
rect 515214 352288 515220 352300
rect 512512 352260 515220 352288
rect 512512 352248 512518 352260
rect 515214 352248 515220 352260
rect 515272 352248 515278 352300
rect 426434 351908 426440 351960
rect 426492 351948 426498 351960
rect 426492 351920 427860 351948
rect 426492 351908 426498 351920
rect 427832 351880 427860 351920
rect 432966 351880 432972 351892
rect 427832 351852 432972 351880
rect 432966 351840 432972 351852
rect 433024 351840 433030 351892
rect 512454 350820 512460 350872
rect 512512 350860 512518 350872
rect 515582 350860 515588 350872
rect 512512 350832 515588 350860
rect 512512 350820 512518 350832
rect 515582 350820 515588 350832
rect 515640 350820 515646 350872
rect 512914 350616 512920 350668
rect 512972 350656 512978 350668
rect 516318 350656 516324 350668
rect 512972 350628 516324 350656
rect 512972 350616 512978 350628
rect 516318 350616 516324 350628
rect 516376 350616 516382 350668
rect 407022 350548 407028 350600
rect 407080 350588 407086 350600
rect 447134 350588 447140 350600
rect 407080 350560 447140 350588
rect 407080 350548 407086 350560
rect 447134 350548 447140 350560
rect 447192 350548 447198 350600
rect 364978 349800 364984 349852
rect 365036 349840 365042 349852
rect 442350 349840 442356 349852
rect 365036 349812 442356 349840
rect 365036 349800 365042 349812
rect 442350 349800 442356 349812
rect 442408 349800 442414 349852
rect 512822 349664 512828 349716
rect 512880 349704 512886 349716
rect 517974 349704 517980 349716
rect 512880 349676 517980 349704
rect 512880 349664 512886 349676
rect 517974 349664 517980 349676
rect 518032 349664 518038 349716
rect 432966 349528 432972 349580
rect 433024 349568 433030 349580
rect 433978 349568 433984 349580
rect 433024 349540 433984 349568
rect 433024 349528 433030 349540
rect 433978 349528 433984 349540
rect 434036 349528 434042 349580
rect 513282 349392 513288 349444
rect 513340 349432 513346 349444
rect 519354 349432 519360 349444
rect 513340 349404 519360 349432
rect 513340 349392 513346 349404
rect 519354 349392 519360 349404
rect 519412 349392 519418 349444
rect 512086 349256 512092 349308
rect 512144 349296 512150 349308
rect 513926 349296 513932 349308
rect 512144 349268 513932 349296
rect 512144 349256 512150 349268
rect 513926 349256 513932 349268
rect 513984 349256 513990 349308
rect 513282 348440 513288 348492
rect 513340 348480 513346 348492
rect 520642 348480 520648 348492
rect 513340 348452 520648 348480
rect 513340 348440 513346 348452
rect 520642 348440 520648 348452
rect 520700 348440 520706 348492
rect 513282 348168 513288 348220
rect 513340 348208 513346 348220
rect 518066 348208 518072 348220
rect 513340 348180 518072 348208
rect 513340 348168 513346 348180
rect 518066 348168 518072 348180
rect 518124 348168 518130 348220
rect 361758 347760 361764 347812
rect 361816 347800 361822 347812
rect 402238 347800 402244 347812
rect 361816 347772 402244 347800
rect 361816 347760 361822 347772
rect 402238 347760 402244 347772
rect 402296 347760 402302 347812
rect 362218 347692 362224 347744
rect 362276 347732 362282 347744
rect 447134 347732 447140 347744
rect 362276 347704 447140 347732
rect 362276 347692 362282 347704
rect 447134 347692 447140 347704
rect 447192 347692 447198 347744
rect 512086 346740 512092 346792
rect 512144 346780 512150 346792
rect 515030 346780 515036 346792
rect 512144 346752 515036 346780
rect 512144 346740 512150 346752
rect 515030 346740 515036 346752
rect 515088 346740 515094 346792
rect 512638 346536 512644 346588
rect 512696 346576 512702 346588
rect 516502 346576 516508 346588
rect 512696 346548 516508 346576
rect 512696 346536 512702 346548
rect 516502 346536 516508 346548
rect 516560 346536 516566 346588
rect 512914 343680 512920 343732
rect 512972 343720 512978 343732
rect 516410 343720 516416 343732
rect 512972 343692 516416 343720
rect 512972 343680 512978 343692
rect 516410 343680 516416 343692
rect 516468 343680 516474 343732
rect 513190 342592 513196 342644
rect 513248 342632 513254 342644
rect 518342 342632 518348 342644
rect 513248 342604 518348 342632
rect 513248 342592 513254 342604
rect 518342 342592 518348 342604
rect 518400 342592 518406 342644
rect 513282 342252 513288 342304
rect 513340 342292 513346 342304
rect 521838 342292 521844 342304
rect 513340 342264 521844 342292
rect 513340 342252 513346 342264
rect 521838 342252 521844 342264
rect 521896 342252 521902 342304
rect 512638 341232 512644 341284
rect 512696 341272 512702 341284
rect 515306 341272 515312 341284
rect 512696 341244 515312 341272
rect 512696 341232 512702 341244
rect 515306 341232 515312 341244
rect 515364 341232 515370 341284
rect 444190 340960 444196 341012
rect 444248 341000 444254 341012
rect 447226 341000 447232 341012
rect 444248 340972 447232 341000
rect 444248 340960 444254 340972
rect 447226 340960 447232 340972
rect 447284 340960 447290 341012
rect 512822 340960 512828 341012
rect 512880 341000 512886 341012
rect 516594 341000 516600 341012
rect 512880 340972 516600 341000
rect 512880 340960 512886 340972
rect 516594 340960 516600 340972
rect 516652 340960 516658 341012
rect 361758 340892 361764 340944
rect 361816 340932 361822 340944
rect 447134 340932 447140 340944
rect 361816 340904 447140 340932
rect 361816 340892 361822 340904
rect 447134 340892 447140 340904
rect 447192 340892 447198 340944
rect 513282 340008 513288 340060
rect 513340 340048 513346 340060
rect 519446 340048 519452 340060
rect 513340 340020 519452 340048
rect 513340 340008 513346 340020
rect 519446 340008 519452 340020
rect 519504 340008 519510 340060
rect 431218 339532 431224 339584
rect 431276 339572 431282 339584
rect 447134 339572 447140 339584
rect 431276 339544 447140 339572
rect 431276 339532 431282 339544
rect 447134 339532 447140 339544
rect 447192 339532 447198 339584
rect 371878 339464 371884 339516
rect 371936 339504 371942 339516
rect 447226 339504 447232 339516
rect 371936 339476 447232 339504
rect 371936 339464 371942 339476
rect 447226 339464 447232 339476
rect 447284 339464 447290 339516
rect 513190 339464 513196 339516
rect 513248 339504 513254 339516
rect 521930 339504 521936 339516
rect 513248 339476 521936 339504
rect 513248 339464 513254 339476
rect 521930 339464 521936 339476
rect 521988 339464 521994 339516
rect 513282 338512 513288 338564
rect 513340 338552 513346 338564
rect 520734 338552 520740 338564
rect 513340 338524 520740 338552
rect 513340 338512 513346 338524
rect 520734 338512 520740 338524
rect 520792 338512 520798 338564
rect 436830 338172 436836 338224
rect 436888 338212 436894 338224
rect 447134 338212 447140 338224
rect 436888 338184 447140 338212
rect 436888 338172 436894 338184
rect 447134 338172 447140 338184
rect 447192 338172 447198 338224
rect 435358 338104 435364 338156
rect 435416 338144 435422 338156
rect 447226 338144 447232 338156
rect 435416 338116 447232 338144
rect 435416 338104 435422 338116
rect 447226 338104 447232 338116
rect 447284 338104 447290 338156
rect 402238 338036 402244 338088
rect 402296 338076 402302 338088
rect 448422 338076 448428 338088
rect 402296 338048 448428 338076
rect 402296 338036 402302 338048
rect 448422 338036 448428 338048
rect 448480 338076 448486 338088
rect 449434 338076 449440 338088
rect 448480 338048 449440 338076
rect 448480 338036 448486 338048
rect 449434 338036 449440 338048
rect 449492 338036 449498 338088
rect 433978 337968 433984 338020
rect 434036 338008 434042 338020
rect 436370 338008 436376 338020
rect 434036 337980 436376 338008
rect 434036 337968 434042 337980
rect 436370 337968 436376 337980
rect 436428 337968 436434 338020
rect 450078 337424 450084 337476
rect 450136 337464 450142 337476
rect 450354 337464 450360 337476
rect 450136 337436 450360 337464
rect 450136 337424 450142 337436
rect 450354 337424 450360 337436
rect 450412 337424 450418 337476
rect 513282 337288 513288 337340
rect 513340 337328 513346 337340
rect 519722 337328 519728 337340
rect 513340 337300 519728 337328
rect 513340 337288 513346 337300
rect 519722 337288 519728 337300
rect 519780 337288 519786 337340
rect 513098 337152 513104 337204
rect 513156 337192 513162 337204
rect 516870 337192 516876 337204
rect 513156 337164 516876 337192
rect 513156 337152 513162 337164
rect 516870 337152 516876 337164
rect 516928 337152 516934 337204
rect 416774 336880 416780 336932
rect 416832 336920 416838 336932
rect 450354 336920 450360 336932
rect 416832 336892 450360 336920
rect 416832 336880 416838 336892
rect 450354 336880 450360 336892
rect 450412 336880 450418 336932
rect 413094 336812 413100 336864
rect 413152 336852 413158 336864
rect 450170 336852 450176 336864
rect 413152 336824 450176 336852
rect 413152 336812 413158 336824
rect 450170 336812 450176 336824
rect 450228 336812 450234 336864
rect 409414 336744 409420 336796
rect 409472 336784 409478 336796
rect 450722 336784 450728 336796
rect 409472 336756 450728 336784
rect 409472 336744 409478 336756
rect 450722 336744 450728 336756
rect 450780 336744 450786 336796
rect 513190 336744 513196 336796
rect 513248 336784 513254 336796
rect 522022 336784 522028 336796
rect 513248 336756 522028 336784
rect 513248 336744 513254 336756
rect 522022 336744 522028 336756
rect 522080 336744 522086 336796
rect 448422 336676 448428 336728
rect 448480 336716 448486 336728
rect 449710 336716 449716 336728
rect 448480 336688 449716 336716
rect 448480 336676 448486 336688
rect 449710 336676 449716 336688
rect 449768 336676 449774 336728
rect 418798 336404 418804 336456
rect 418856 336444 418862 336456
rect 439866 336444 439872 336456
rect 418856 336416 439872 336444
rect 418856 336404 418862 336416
rect 439866 336404 439872 336416
rect 439924 336404 439930 336456
rect 418890 336336 418896 336388
rect 418948 336376 418954 336388
rect 442534 336376 442540 336388
rect 418948 336348 442540 336376
rect 418948 336336 418954 336348
rect 442534 336336 442540 336348
rect 442592 336336 442598 336388
rect 416038 336268 416044 336320
rect 416096 336308 416102 336320
rect 439774 336308 439780 336320
rect 416096 336280 439780 336308
rect 416096 336268 416102 336280
rect 439774 336268 439780 336280
rect 439832 336268 439838 336320
rect 440878 336268 440884 336320
rect 440936 336308 440942 336320
rect 447134 336308 447140 336320
rect 440936 336280 447140 336308
rect 440936 336268 440942 336280
rect 447134 336268 447140 336280
rect 447192 336268 447198 336320
rect 418982 336200 418988 336252
rect 419040 336240 419046 336252
rect 449526 336240 449532 336252
rect 419040 336212 449532 336240
rect 419040 336200 419046 336212
rect 449526 336200 449532 336212
rect 449584 336200 449590 336252
rect 413646 336132 413652 336184
rect 413704 336172 413710 336184
rect 449618 336172 449624 336184
rect 413704 336144 449624 336172
rect 413704 336132 413710 336144
rect 449618 336132 449624 336144
rect 449676 336132 449682 336184
rect 397454 336064 397460 336116
rect 397512 336104 397518 336116
rect 447686 336104 447692 336116
rect 397512 336076 447692 336104
rect 397512 336064 397518 336076
rect 447686 336064 447692 336076
rect 447744 336064 447750 336116
rect 362218 335996 362224 336048
rect 362276 336036 362282 336048
rect 444190 336036 444196 336048
rect 362276 336008 444196 336036
rect 362276 335996 362282 336008
rect 444190 335996 444196 336008
rect 444248 335996 444254 336048
rect 443730 335656 443736 335708
rect 443788 335696 443794 335708
rect 447134 335696 447140 335708
rect 443788 335668 447140 335696
rect 443788 335656 443794 335668
rect 447134 335656 447140 335668
rect 447192 335656 447198 335708
rect 399478 335316 399484 335368
rect 399536 335356 399542 335368
rect 447410 335356 447416 335368
rect 399536 335328 447416 335356
rect 399536 335316 399542 335328
rect 447410 335316 447416 335328
rect 447468 335316 447474 335368
rect 513282 335316 513288 335368
rect 513340 335356 513346 335368
rect 522114 335356 522120 335368
rect 513340 335328 522120 335356
rect 513340 335316 513346 335328
rect 522114 335316 522120 335328
rect 522172 335316 522178 335368
rect 432598 334908 432604 334960
rect 432656 334948 432662 334960
rect 447502 334948 447508 334960
rect 432656 334920 447508 334948
rect 432656 334908 432662 334920
rect 447502 334908 447508 334920
rect 447560 334908 447566 334960
rect 420546 334840 420552 334892
rect 420604 334880 420610 334892
rect 442442 334880 442448 334892
rect 420604 334852 442448 334880
rect 420604 334840 420610 334852
rect 442442 334840 442448 334852
rect 442500 334840 442506 334892
rect 420730 334772 420736 334824
rect 420788 334812 420794 334824
rect 442626 334812 442632 334824
rect 420788 334784 442632 334812
rect 420788 334772 420794 334784
rect 442626 334772 442632 334784
rect 442684 334772 442690 334824
rect 420178 334704 420184 334756
rect 420236 334744 420242 334756
rect 444926 334744 444932 334756
rect 420236 334716 444932 334744
rect 420236 334704 420242 334716
rect 444926 334704 444932 334716
rect 444984 334704 444990 334756
rect 420270 334636 420276 334688
rect 420328 334676 420334 334688
rect 445662 334676 445668 334688
rect 420328 334648 445668 334676
rect 420328 334636 420334 334648
rect 445662 334636 445668 334648
rect 445720 334636 445726 334688
rect 420638 334568 420644 334620
rect 420696 334608 420702 334620
rect 449710 334608 449716 334620
rect 420696 334580 449716 334608
rect 420696 334568 420702 334580
rect 449710 334568 449716 334580
rect 449768 334568 449774 334620
rect 513282 334568 513288 334620
rect 513340 334608 513346 334620
rect 520826 334608 520832 334620
rect 513340 334580 520832 334608
rect 513340 334568 513346 334580
rect 520826 334568 520832 334580
rect 520884 334568 520890 334620
rect 443638 334024 443644 334076
rect 443696 334064 443702 334076
rect 447226 334064 447232 334076
rect 443696 334036 447232 334064
rect 443696 334024 443702 334036
rect 447226 334024 447232 334036
rect 447284 334024 447290 334076
rect 363782 333956 363788 334008
rect 363840 333996 363846 334008
rect 447134 333996 447140 334008
rect 363840 333968 447140 333996
rect 363840 333956 363846 333968
rect 447134 333956 447140 333968
rect 447192 333956 447198 334008
rect 513282 333956 513288 334008
rect 513340 333996 513346 334008
rect 522206 333996 522212 334008
rect 513340 333968 522212 333996
rect 513340 333956 513346 333968
rect 522206 333956 522212 333968
rect 522264 333956 522270 334008
rect 513006 333072 513012 333124
rect 513064 333112 513070 333124
rect 516686 333112 516692 333124
rect 513064 333084 516692 333112
rect 513064 333072 513070 333084
rect 516686 333072 516692 333084
rect 516744 333072 516750 333124
rect 512638 332868 512644 332920
rect 512696 332908 512702 332920
rect 514110 332908 514116 332920
rect 512696 332880 514116 332908
rect 512696 332868 512702 332880
rect 514110 332868 514116 332880
rect 514168 332868 514174 332920
rect 439590 332664 439596 332716
rect 439648 332704 439654 332716
rect 447226 332704 447232 332716
rect 439648 332676 447232 332704
rect 439648 332664 439654 332676
rect 447226 332664 447232 332676
rect 447284 332664 447290 332716
rect 436738 332596 436744 332648
rect 436796 332636 436802 332648
rect 447134 332636 447140 332648
rect 436796 332608 447140 332636
rect 436796 332596 436802 332608
rect 447134 332596 447140 332608
rect 447192 332596 447198 332648
rect 512638 331440 512644 331492
rect 512696 331480 512702 331492
rect 516134 331480 516140 331492
rect 512696 331452 516140 331480
rect 512696 331440 512702 331452
rect 516134 331440 516140 331452
rect 516192 331440 516198 331492
rect 442902 330488 442908 330540
rect 442960 330528 442966 330540
rect 447962 330528 447968 330540
rect 442960 330500 447968 330528
rect 442960 330488 442966 330500
rect 447962 330488 447968 330500
rect 448020 330488 448026 330540
rect 450078 330488 450084 330540
rect 450136 330528 450142 330540
rect 450722 330528 450728 330540
rect 450136 330500 450728 330528
rect 450136 330488 450142 330500
rect 450722 330488 450728 330500
rect 450780 330488 450786 330540
rect 580718 330488 580724 330540
rect 580776 330528 580782 330540
rect 580902 330528 580908 330540
rect 580776 330500 580908 330528
rect 580776 330488 580782 330500
rect 580902 330488 580908 330500
rect 580960 330488 580966 330540
rect 432874 330148 432880 330200
rect 432932 330188 432938 330200
rect 439682 330188 439688 330200
rect 432932 330160 439688 330188
rect 432932 330148 432938 330160
rect 439682 330148 439688 330160
rect 439740 330148 439746 330200
rect 439498 329808 439504 329860
rect 439556 329848 439562 329860
rect 447134 329848 447140 329860
rect 439556 329820 447140 329848
rect 439556 329808 439562 329820
rect 447134 329808 447140 329820
rect 447192 329808 447198 329860
rect 436370 329740 436376 329792
rect 436428 329780 436434 329792
rect 438118 329780 438124 329792
rect 436428 329752 438124 329780
rect 436428 329740 436434 329752
rect 438118 329740 438124 329752
rect 438176 329740 438182 329792
rect 436002 328516 436008 328568
rect 436060 328556 436066 328568
rect 449894 328556 449900 328568
rect 436060 328528 449900 328556
rect 436060 328516 436066 328528
rect 449894 328516 449900 328528
rect 449952 328516 449958 328568
rect 431862 328448 431868 328500
rect 431920 328488 431926 328500
rect 450446 328488 450452 328500
rect 431920 328460 450452 328488
rect 431920 328448 431926 328460
rect 450446 328448 450452 328460
rect 450504 328448 450510 328500
rect 509510 326340 509516 326392
rect 509568 326380 509574 326392
rect 510154 326380 510160 326392
rect 509568 326352 510160 326380
rect 509568 326340 509574 326352
rect 510154 326340 510160 326352
rect 510212 326340 510218 326392
rect 509326 326204 509332 326256
rect 509384 326244 509390 326256
rect 509510 326244 509516 326256
rect 509384 326216 509516 326244
rect 509384 326204 509390 326216
rect 509510 326204 509516 326216
rect 509568 326204 509574 326256
rect 432874 324912 432880 324964
rect 432932 324952 432938 324964
rect 442258 324952 442264 324964
rect 432932 324924 442264 324952
rect 432932 324912 432938 324924
rect 442258 324912 442264 324924
rect 442316 324912 442322 324964
rect 438118 323960 438124 324012
rect 438176 324000 438182 324012
rect 439958 324000 439964 324012
rect 438176 323972 439964 324000
rect 438176 323960 438182 323972
rect 439958 323960 439964 323972
rect 440016 323960 440022 324012
rect 463804 323088 469720 323116
rect 432690 322940 432696 322992
rect 432748 322980 432754 322992
rect 436922 322980 436928 322992
rect 432748 322952 436928 322980
rect 432748 322940 432754 322952
rect 436922 322940 436928 322952
rect 436980 322940 436986 322992
rect 463804 322980 463832 323088
rect 463712 322952 463832 322980
rect 463712 322912 463740 322952
rect 458836 322884 463740 322912
rect 469692 322912 469720 323088
rect 570598 322912 570604 322924
rect 469692 322884 570604 322912
rect 444098 322804 444104 322856
rect 444156 322844 444162 322856
rect 444156 322816 451274 322844
rect 444156 322804 444162 322816
rect 451246 322708 451274 322816
rect 458836 322720 458864 322884
rect 570598 322872 570604 322884
rect 570656 322872 570662 322924
rect 580534 322844 580540 322856
rect 469600 322816 580540 322844
rect 459020 322748 469076 322776
rect 458266 322708 458272 322720
rect 451246 322680 458272 322708
rect 458266 322668 458272 322680
rect 458324 322668 458330 322720
rect 458818 322668 458824 322720
rect 458876 322668 458882 322720
rect 458542 322600 458548 322652
rect 458600 322640 458606 322652
rect 459020 322640 459048 322748
rect 469048 322720 469076 322748
rect 469600 322720 469628 322816
rect 580534 322804 580540 322816
rect 580592 322804 580598 322856
rect 569218 322776 569224 322788
rect 470980 322748 569224 322776
rect 459094 322668 459100 322720
rect 459152 322708 459158 322720
rect 468202 322708 468208 322720
rect 459152 322680 468208 322708
rect 459152 322668 459158 322680
rect 468202 322668 468208 322680
rect 468260 322668 468266 322720
rect 469030 322668 469036 322720
rect 469088 322668 469094 322720
rect 469582 322668 469588 322720
rect 469640 322668 469646 322720
rect 458600 322612 459048 322640
rect 458600 322600 458606 322612
rect 459370 322600 459376 322652
rect 459428 322640 459434 322652
rect 468478 322640 468484 322652
rect 459428 322612 468484 322640
rect 459428 322600 459434 322612
rect 468478 322600 468484 322612
rect 468536 322600 468542 322652
rect 470980 322584 471008 322748
rect 569218 322736 569224 322748
rect 569276 322736 569282 322788
rect 471238 322668 471244 322720
rect 471296 322708 471302 322720
rect 516778 322708 516784 322720
rect 471296 322680 516784 322708
rect 471296 322668 471302 322680
rect 516778 322668 516784 322680
rect 516836 322668 516842 322720
rect 471514 322600 471520 322652
rect 471572 322640 471578 322652
rect 515490 322640 515496 322652
rect 471572 322612 515496 322640
rect 471572 322600 471578 322612
rect 515490 322600 515496 322612
rect 515548 322600 515554 322652
rect 444926 322532 444932 322584
rect 444984 322572 444990 322584
rect 468754 322572 468760 322584
rect 444984 322544 468760 322572
rect 444984 322532 444990 322544
rect 468754 322532 468760 322544
rect 468812 322532 468818 322584
rect 470962 322532 470968 322584
rect 471020 322532 471026 322584
rect 484210 322572 484216 322584
rect 473326 322544 484216 322572
rect 458818 322464 458824 322516
rect 458876 322504 458882 322516
rect 459370 322504 459376 322516
rect 458876 322476 459376 322504
rect 458876 322464 458882 322476
rect 459370 322464 459376 322476
rect 459428 322464 459434 322516
rect 470134 322464 470140 322516
rect 470192 322504 470198 322516
rect 473326 322504 473354 322544
rect 484210 322532 484216 322544
rect 484268 322532 484274 322584
rect 470192 322476 473354 322504
rect 470192 322464 470198 322476
rect 479794 322464 479800 322516
rect 479852 322504 479858 322516
rect 518250 322504 518256 322516
rect 479852 322476 518256 322504
rect 479852 322464 479858 322476
rect 518250 322464 518256 322476
rect 518308 322464 518314 322516
rect 445662 322396 445668 322448
rect 445720 322436 445726 322448
rect 483934 322436 483940 322448
rect 445720 322408 483940 322436
rect 445720 322396 445726 322408
rect 483934 322396 483940 322408
rect 483992 322396 483998 322448
rect 449710 322328 449716 322380
rect 449768 322368 449774 322380
rect 455782 322368 455788 322380
rect 449768 322340 455788 322368
rect 449768 322328 449774 322340
rect 455782 322328 455788 322340
rect 455840 322328 455846 322380
rect 458266 322328 458272 322380
rect 458324 322368 458330 322380
rect 460474 322368 460480 322380
rect 458324 322340 460480 322368
rect 458324 322328 458330 322340
rect 460474 322328 460480 322340
rect 460532 322328 460538 322380
rect 468478 322328 468484 322380
rect 468536 322368 468542 322380
rect 471514 322368 471520 322380
rect 468536 322340 471520 322368
rect 468536 322328 468542 322340
rect 471514 322328 471520 322340
rect 471572 322328 471578 322380
rect 439866 322260 439872 322312
rect 439924 322300 439930 322312
rect 472066 322300 472072 322312
rect 439924 322272 472072 322300
rect 439924 322260 439930 322272
rect 472066 322260 472072 322272
rect 472124 322260 472130 322312
rect 507854 322260 507860 322312
rect 507912 322300 507918 322312
rect 580258 322300 580264 322312
rect 507912 322272 580264 322300
rect 507912 322260 507918 322272
rect 580258 322260 580264 322272
rect 580316 322260 580322 322312
rect 439958 322192 439964 322244
rect 440016 322232 440022 322244
rect 466546 322232 466552 322244
rect 440016 322204 466552 322232
rect 440016 322192 440022 322204
rect 466546 322192 466552 322204
rect 466604 322192 466610 322244
rect 468202 322192 468208 322244
rect 468260 322232 468266 322244
rect 471238 322232 471244 322244
rect 468260 322204 471244 322232
rect 468260 322192 468266 322204
rect 471238 322192 471244 322204
rect 471296 322192 471302 322244
rect 500218 322192 500224 322244
rect 500276 322232 500282 322244
rect 580166 322232 580172 322244
rect 500276 322204 580172 322232
rect 500276 322192 500282 322204
rect 580166 322192 580172 322204
rect 580224 322192 580230 322244
rect 447686 322124 447692 322176
rect 447744 322164 447750 322176
rect 481450 322164 481456 322176
rect 447744 322136 481456 322164
rect 447744 322124 447750 322136
rect 481450 322124 481456 322136
rect 481508 322124 481514 322176
rect 469306 322056 469312 322108
rect 469364 322096 469370 322108
rect 469582 322096 469588 322108
rect 469364 322068 469588 322096
rect 469364 322056 469370 322068
rect 469582 322056 469588 322068
rect 469640 322056 469646 322108
rect 455782 321988 455788 322040
rect 455840 322028 455846 322040
rect 463510 322028 463516 322040
rect 455840 322000 463516 322028
rect 455840 321988 455846 322000
rect 463510 321988 463516 322000
rect 463568 321988 463574 322040
rect 469030 321988 469036 322040
rect 469088 322028 469094 322040
rect 470962 322028 470968 322040
rect 469088 322000 470968 322028
rect 469088 321988 469094 322000
rect 470962 321988 470968 322000
rect 471020 321988 471026 322040
rect 507302 321648 507308 321700
rect 507360 321688 507366 321700
rect 509786 321688 509792 321700
rect 507360 321660 509792 321688
rect 507360 321648 507366 321660
rect 509786 321648 509792 321660
rect 509844 321648 509850 321700
rect 447042 321512 447048 321564
rect 447100 321552 447106 321564
rect 463050 321552 463056 321564
rect 447100 321524 463056 321552
rect 447100 321512 447106 321524
rect 463050 321512 463056 321524
rect 463108 321512 463114 321564
rect 468570 321512 468576 321564
rect 468628 321552 468634 321564
rect 573358 321552 573364 321564
rect 468628 321524 573364 321552
rect 468628 321512 468634 321524
rect 573358 321512 573364 321524
rect 573416 321512 573422 321564
rect 458358 321444 458364 321496
rect 458416 321484 458422 321496
rect 511442 321484 511448 321496
rect 458416 321456 511448 321484
rect 458416 321444 458422 321456
rect 511442 321444 511448 321456
rect 511500 321444 511506 321496
rect 449250 321376 449256 321428
rect 449308 321416 449314 321428
rect 461394 321416 461400 321428
rect 449308 321388 461400 321416
rect 449308 321376 449314 321388
rect 461394 321376 461400 321388
rect 461452 321376 461458 321428
rect 469398 321376 469404 321428
rect 469456 321416 469462 321428
rect 518158 321416 518164 321428
rect 469456 321388 518164 321416
rect 469456 321376 469462 321388
rect 518158 321376 518164 321388
rect 518216 321376 518222 321428
rect 446398 321308 446404 321360
rect 446456 321348 446462 321360
rect 461670 321348 461676 321360
rect 446456 321320 461676 321348
rect 446456 321308 446462 321320
rect 461670 321308 461676 321320
rect 461728 321308 461734 321360
rect 479058 321308 479064 321360
rect 479116 321348 479122 321360
rect 514018 321348 514024 321360
rect 479116 321320 514024 321348
rect 479116 321308 479122 321320
rect 514018 321308 514024 321320
rect 514076 321308 514082 321360
rect 445018 321240 445024 321292
rect 445076 321280 445082 321292
rect 483198 321280 483204 321292
rect 445076 321252 483204 321280
rect 445076 321240 445082 321252
rect 483198 321240 483204 321252
rect 483256 321240 483262 321292
rect 445478 321172 445484 321224
rect 445536 321212 445542 321224
rect 473814 321212 473820 321224
rect 445536 321184 473820 321212
rect 445536 321172 445542 321184
rect 473814 321172 473820 321184
rect 473872 321172 473878 321224
rect 507394 321172 507400 321224
rect 507452 321212 507458 321224
rect 513466 321212 513472 321224
rect 507452 321184 513472 321212
rect 507452 321172 507458 321184
rect 513466 321172 513472 321184
rect 513524 321172 513530 321224
rect 446490 321104 446496 321156
rect 446548 321144 446554 321156
rect 471882 321144 471888 321156
rect 446548 321116 471888 321144
rect 446548 321104 446554 321116
rect 471882 321104 471888 321116
rect 471940 321104 471946 321156
rect 507210 321104 507216 321156
rect 507268 321144 507274 321156
rect 516134 321144 516140 321156
rect 507268 321116 516140 321144
rect 507268 321104 507274 321116
rect 516134 321104 516140 321116
rect 516192 321104 516198 321156
rect 460198 321036 460204 321088
rect 460256 321076 460262 321088
rect 513834 321076 513840 321088
rect 460256 321048 513840 321076
rect 460256 321036 460262 321048
rect 513834 321036 513840 321048
rect 513892 321036 513898 321088
rect 445110 320968 445116 321020
rect 445168 321008 445174 321020
rect 482094 321008 482100 321020
rect 445168 320980 482100 321008
rect 445168 320968 445174 320980
rect 482094 320968 482100 320980
rect 482152 320968 482158 321020
rect 496814 320968 496820 321020
rect 496872 321008 496878 321020
rect 580626 321008 580632 321020
rect 496872 320980 580632 321008
rect 496872 320968 496878 320980
rect 580626 320968 580632 320980
rect 580684 320968 580690 321020
rect 459922 320900 459928 320952
rect 459980 320940 459986 320952
rect 580350 320940 580356 320952
rect 459980 320912 580356 320940
rect 459980 320900 459986 320912
rect 580350 320900 580356 320912
rect 580408 320900 580414 320952
rect 461854 320832 461860 320884
rect 461912 320872 461918 320884
rect 580810 320872 580816 320884
rect 461912 320844 580816 320872
rect 461912 320832 461918 320844
rect 580810 320832 580816 320844
rect 580868 320832 580874 320884
rect 446950 320764 446956 320816
rect 447008 320804 447014 320816
rect 473262 320804 473268 320816
rect 447008 320776 473268 320804
rect 447008 320764 447014 320776
rect 473262 320764 473268 320776
rect 473320 320764 473326 320816
rect 439774 320696 439780 320748
rect 439832 320736 439838 320748
rect 472434 320736 472440 320748
rect 439832 320708 472440 320736
rect 439832 320696 439838 320708
rect 472434 320696 472440 320708
rect 472492 320696 472498 320748
rect 442534 320628 442540 320680
rect 442592 320668 442598 320680
rect 481818 320668 481824 320680
rect 442592 320640 481824 320668
rect 442592 320628 442598 320640
rect 481818 320628 481824 320640
rect 481876 320628 481882 320680
rect 442350 320084 442356 320136
rect 442408 320124 442414 320136
rect 442408 320096 456104 320124
rect 442408 320084 442414 320096
rect 446858 320016 446864 320068
rect 446916 320056 446922 320068
rect 456076 320056 456104 320096
rect 458082 320084 458088 320136
rect 458140 320124 458146 320136
rect 461854 320124 461860 320136
rect 458140 320096 461860 320124
rect 458140 320084 458146 320096
rect 461854 320084 461860 320096
rect 461912 320084 461918 320136
rect 480714 320084 480720 320136
rect 480772 320124 480778 320136
rect 507854 320124 507860 320136
rect 480772 320096 507860 320124
rect 480772 320084 480778 320096
rect 507854 320084 507860 320096
rect 507912 320084 507918 320136
rect 460842 320056 460848 320068
rect 446916 320028 451274 320056
rect 456076 320028 460848 320056
rect 446916 320016 446922 320028
rect 451246 319988 451274 320028
rect 460842 320016 460848 320028
rect 460900 320016 460906 320068
rect 466546 320016 466552 320068
rect 466604 320056 466610 320068
rect 474366 320056 474372 320068
rect 466604 320028 474372 320056
rect 466604 320016 466610 320028
rect 474366 320016 474372 320028
rect 474424 320016 474430 320068
rect 479334 320016 479340 320068
rect 479392 320056 479398 320068
rect 496814 320056 496820 320068
rect 479392 320028 496820 320056
rect 479392 320016 479398 320028
rect 496814 320016 496820 320028
rect 496872 320016 496878 320068
rect 463326 319988 463332 320000
rect 451246 319960 463332 319988
rect 463326 319948 463332 319960
rect 463384 319948 463390 320000
rect 470226 319948 470232 320000
rect 470284 319988 470290 320000
rect 576118 319988 576124 320000
rect 470284 319960 576124 319988
rect 470284 319948 470290 319960
rect 576118 319948 576124 319960
rect 576176 319948 576182 320000
rect 479886 319880 479892 319932
rect 479944 319920 479950 319932
rect 519538 319920 519544 319932
rect 479944 319892 519544 319920
rect 479944 319880 479950 319892
rect 519538 319880 519544 319892
rect 519596 319880 519602 319932
rect 442626 319812 442632 319864
rect 442684 319852 442690 319864
rect 463878 319852 463884 319864
rect 442684 319824 463884 319852
rect 442684 319812 442690 319824
rect 463878 319812 463884 319824
rect 463936 319812 463942 319864
rect 469674 319812 469680 319864
rect 469732 319852 469738 319864
rect 511350 319852 511356 319864
rect 469732 319824 511356 319852
rect 469732 319812 469738 319824
rect 511350 319812 511356 319824
rect 511408 319812 511414 319864
rect 449618 319744 449624 319796
rect 449676 319784 449682 319796
rect 471054 319784 471060 319796
rect 449676 319756 471060 319784
rect 449676 319744 449682 319756
rect 471054 319744 471060 319756
rect 471112 319744 471118 319796
rect 480990 319744 480996 319796
rect 481048 319784 481054 319796
rect 519630 319784 519636 319796
rect 481048 319756 519636 319784
rect 481048 319744 481054 319756
rect 519630 319744 519636 319756
rect 519688 319744 519694 319796
rect 445386 319676 445392 319728
rect 445444 319716 445450 319728
rect 462774 319716 462780 319728
rect 445444 319688 462780 319716
rect 445444 319676 445450 319688
rect 462774 319676 462780 319688
rect 462832 319676 462838 319728
rect 480438 319676 480444 319728
rect 480496 319716 480502 319728
rect 515398 319716 515404 319728
rect 480496 319688 515404 319716
rect 480496 319676 480502 319688
rect 515398 319676 515404 319688
rect 515456 319676 515462 319728
rect 460382 319608 460388 319660
rect 460440 319648 460446 319660
rect 465810 319648 465816 319660
rect 460440 319620 465816 319648
rect 460440 319608 460446 319620
rect 465810 319608 465816 319620
rect 465868 319608 465874 319660
rect 480162 319608 480168 319660
rect 480220 319648 480226 319660
rect 511258 319648 511264 319660
rect 480220 319620 511264 319648
rect 480220 319608 480226 319620
rect 511258 319608 511264 319620
rect 511316 319608 511322 319660
rect 459002 319540 459008 319592
rect 459060 319580 459066 319592
rect 465534 319580 465540 319592
rect 459060 319552 465540 319580
rect 459060 319540 459066 319552
rect 465534 319540 465540 319552
rect 465592 319540 465598 319592
rect 498654 319540 498660 319592
rect 498712 319580 498718 319592
rect 534718 319580 534724 319592
rect 498712 319552 534724 319580
rect 498712 319540 498718 319552
rect 534718 319540 534724 319552
rect 534776 319540 534782 319592
rect 460290 319472 460296 319524
rect 460348 319512 460354 319524
rect 476298 319512 476304 319524
rect 460348 319484 476304 319512
rect 460348 319472 460354 319484
rect 476298 319472 476304 319484
rect 476356 319472 476362 319524
rect 498102 319472 498108 319524
rect 498160 319512 498166 319524
rect 533338 319512 533344 319524
rect 498160 319484 533344 319512
rect 498160 319472 498166 319484
rect 533338 319472 533344 319484
rect 533396 319472 533402 319524
rect 458818 319404 458824 319456
rect 458876 319444 458882 319456
rect 476022 319444 476028 319456
rect 458876 319416 476028 319444
rect 458876 319404 458882 319416
rect 476022 319404 476028 319416
rect 476080 319404 476086 319456
rect 478782 319404 478788 319456
rect 478840 319444 478846 319456
rect 500218 319444 500224 319456
rect 478840 319416 500224 319444
rect 478840 319404 478846 319416
rect 500218 319404 500224 319416
rect 500276 319404 500282 319456
rect 501690 319404 501696 319456
rect 501748 319444 501754 319456
rect 538858 319444 538864 319456
rect 501748 319416 538864 319444
rect 501748 319404 501754 319416
rect 538858 319404 538864 319416
rect 538916 319404 538922 319456
rect 446582 319336 446588 319388
rect 446640 319376 446646 319388
rect 471330 319376 471336 319388
rect 446640 319348 471336 319376
rect 446640 319336 446646 319348
rect 471330 319336 471336 319348
rect 471388 319336 471394 319388
rect 481266 319336 481272 319388
rect 481324 319376 481330 319388
rect 510614 319376 510620 319388
rect 481324 319348 510620 319376
rect 481324 319336 481330 319348
rect 510614 319336 510620 319348
rect 510672 319336 510678 319388
rect 445294 319268 445300 319320
rect 445352 319308 445358 319320
rect 482370 319308 482376 319320
rect 445352 319280 482376 319308
rect 445352 319268 445358 319280
rect 482370 319268 482376 319280
rect 482428 319268 482434 319320
rect 502794 319268 502800 319320
rect 502852 319308 502858 319320
rect 530578 319308 530584 319320
rect 502852 319280 530584 319308
rect 502852 319268 502858 319280
rect 530578 319268 530584 319280
rect 530636 319268 530642 319320
rect 468846 319200 468852 319252
rect 468904 319240 468910 319252
rect 580902 319240 580908 319252
rect 468904 319212 580908 319240
rect 468904 319200 468910 319212
rect 580902 319200 580908 319212
rect 580960 319200 580966 319252
rect 455782 319132 455788 319184
rect 455840 319172 455846 319184
rect 456058 319172 456064 319184
rect 455840 319144 456064 319172
rect 455840 319132 455846 319144
rect 456058 319132 456064 319144
rect 456116 319132 456122 319184
rect 457162 319132 457168 319184
rect 457220 319172 457226 319184
rect 457990 319172 457996 319184
rect 457220 319144 457996 319172
rect 457220 319132 457226 319144
rect 457990 319132 457996 319144
rect 458048 319132 458054 319184
rect 466822 319132 466828 319184
rect 466880 319172 466886 319184
rect 467374 319172 467380 319184
rect 466880 319144 467380 319172
rect 466880 319132 466886 319144
rect 467374 319132 467380 319144
rect 467432 319132 467438 319184
rect 469950 319132 469956 319184
rect 470008 319172 470014 319184
rect 580442 319172 580448 319184
rect 470008 319144 580448 319172
rect 470008 319132 470014 319144
rect 580442 319132 580448 319144
rect 580500 319132 580506 319184
rect 442442 319064 442448 319116
rect 442500 319104 442506 319116
rect 484302 319104 484308 319116
rect 442500 319076 484308 319104
rect 442500 319064 442506 319076
rect 484302 319064 484308 319076
rect 484360 319064 484366 319116
rect 497458 319064 497464 319116
rect 497516 319104 497522 319116
rect 498010 319104 498016 319116
rect 497516 319076 498016 319104
rect 497516 319064 497522 319076
rect 498010 319064 498016 319076
rect 498068 319064 498074 319116
rect 501598 319064 501604 319116
rect 501656 319104 501662 319116
rect 502150 319104 502156 319116
rect 501656 319076 502156 319104
rect 501656 319064 501662 319076
rect 502150 319064 502156 319076
rect 502208 319064 502214 319116
rect 446674 318996 446680 319048
rect 446732 319036 446738 319048
rect 446732 319008 470594 319036
rect 446732 318996 446738 319008
rect 466638 318928 466644 318980
rect 466696 318968 466702 318980
rect 467374 318968 467380 318980
rect 466696 318940 467380 318968
rect 466696 318928 466702 318940
rect 467374 318928 467380 318940
rect 467432 318928 467438 318980
rect 470566 318968 470594 319008
rect 471238 318996 471244 319048
rect 471296 319036 471302 319048
rect 474642 319036 474648 319048
rect 471296 319008 474648 319036
rect 471296 318996 471302 319008
rect 474642 318996 474648 319008
rect 474700 318996 474706 319048
rect 471606 318968 471612 318980
rect 470566 318940 471612 318968
rect 471606 318928 471612 318940
rect 471664 318928 471670 318980
rect 449526 318724 449532 318776
rect 449584 318764 449590 318776
rect 483474 318764 483480 318776
rect 449584 318736 483480 318764
rect 449584 318724 449590 318736
rect 483474 318724 483480 318736
rect 483532 318724 483538 318776
rect 444282 318656 444288 318708
rect 444340 318696 444346 318708
rect 470778 318696 470784 318708
rect 444340 318668 470784 318696
rect 444340 318656 444346 318668
rect 470778 318656 470784 318668
rect 470836 318656 470842 318708
rect 432046 318248 432052 318300
rect 432104 318288 432110 318300
rect 435450 318288 435456 318300
rect 432104 318260 435456 318288
rect 432104 318248 432110 318260
rect 435450 318248 435456 318260
rect 435508 318248 435514 318300
rect 454770 318180 454776 318232
rect 454828 318220 454834 318232
rect 491478 318220 491484 318232
rect 454828 318192 491484 318220
rect 454828 318180 454834 318192
rect 491478 318180 491484 318192
rect 491536 318180 491542 318232
rect 496170 318180 496176 318232
rect 496228 318220 496234 318232
rect 539594 318220 539600 318232
rect 496228 318192 539600 318220
rect 496228 318180 496234 318192
rect 539594 318180 539600 318192
rect 539652 318180 539658 318232
rect 456058 318112 456064 318164
rect 456116 318152 456122 318164
rect 512086 318152 512092 318164
rect 456116 318124 512092 318152
rect 456116 318112 456122 318124
rect 512086 318112 512092 318124
rect 512144 318112 512150 318164
rect 476850 318044 476856 318096
rect 476908 318084 476914 318096
rect 569218 318084 569224 318096
rect 476908 318056 569224 318084
rect 476908 318044 476914 318056
rect 569218 318044 569224 318056
rect 569276 318044 569282 318096
rect 478506 317704 478512 317756
rect 478564 317744 478570 317756
rect 479518 317744 479524 317756
rect 478564 317716 479524 317744
rect 478564 317704 478570 317716
rect 479518 317704 479524 317716
rect 479576 317704 479582 317756
rect 453390 317364 453396 317416
rect 453448 317404 453454 317416
rect 464982 317404 464988 317416
rect 453448 317376 464988 317404
rect 453448 317364 453454 317376
rect 464982 317364 464988 317376
rect 465040 317364 465046 317416
rect 456334 317296 456340 317348
rect 456392 317336 456398 317348
rect 475746 317336 475752 317348
rect 456392 317308 475752 317336
rect 456392 317296 456398 317308
rect 475746 317296 475752 317308
rect 475804 317296 475810 317348
rect 456426 317228 456432 317280
rect 456484 317268 456490 317280
rect 475470 317268 475476 317280
rect 456484 317240 475476 317268
rect 456484 317228 456490 317240
rect 475470 317228 475476 317240
rect 475528 317228 475534 317280
rect 453298 317160 453304 317212
rect 453356 317200 453362 317212
rect 475194 317200 475200 317212
rect 453356 317172 475200 317200
rect 453356 317160 453362 317172
rect 475194 317160 475200 317172
rect 475252 317160 475258 317212
rect 459186 317092 459192 317144
rect 459244 317132 459250 317144
rect 486510 317132 486516 317144
rect 459244 317104 486516 317132
rect 459244 317092 459250 317104
rect 486510 317092 486516 317104
rect 486568 317092 486574 317144
rect 458910 317024 458916 317076
rect 458968 317064 458974 317076
rect 485958 317064 485964 317076
rect 458968 317036 485964 317064
rect 458968 317024 458974 317036
rect 485958 317024 485964 317036
rect 486016 317024 486022 317076
rect 453482 316956 453488 317008
rect 453540 316996 453546 317008
rect 485682 316996 485688 317008
rect 453540 316968 485688 316996
rect 453540 316956 453546 316968
rect 485682 316956 485688 316968
rect 485740 316956 485746 317008
rect 491662 316996 491668 317008
rect 487172 316968 491668 316996
rect 450630 316888 450636 316940
rect 450688 316928 450694 316940
rect 457714 316928 457720 316940
rect 450688 316900 457720 316928
rect 450688 316888 450694 316900
rect 457714 316888 457720 316900
rect 457772 316888 457778 316940
rect 459094 316888 459100 316940
rect 459152 316928 459158 316940
rect 487172 316928 487200 316968
rect 491662 316956 491668 316968
rect 491720 316956 491726 317008
rect 459152 316900 487200 316928
rect 459152 316888 459158 316900
rect 487246 316888 487252 316940
rect 487304 316928 487310 316940
rect 488350 316928 488356 316940
rect 487304 316900 488356 316928
rect 487304 316888 487310 316900
rect 488350 316888 488356 316900
rect 488408 316888 488414 316940
rect 500310 316888 500316 316940
rect 500368 316928 500374 316940
rect 539778 316928 539784 316940
rect 500368 316900 539784 316928
rect 500368 316888 500374 316900
rect 539778 316888 539784 316900
rect 539836 316888 539842 316940
rect 451918 316820 451924 316872
rect 451976 316860 451982 316872
rect 495894 316860 495900 316872
rect 451976 316832 495900 316860
rect 451976 316820 451982 316832
rect 495894 316820 495900 316832
rect 495952 316820 495958 316872
rect 502518 316820 502524 316872
rect 502576 316860 502582 316872
rect 542630 316860 542636 316872
rect 502576 316832 542636 316860
rect 502576 316820 502582 316832
rect 542630 316820 542636 316832
rect 542688 316820 542694 316872
rect 450630 316752 450636 316804
rect 450688 316792 450694 316804
rect 509510 316792 509516 316804
rect 450688 316764 509516 316792
rect 450688 316752 450694 316764
rect 509510 316752 509516 316764
rect 509568 316752 509574 316804
rect 450814 316684 450820 316736
rect 450872 316724 450878 316736
rect 474918 316724 474924 316736
rect 450872 316696 474924 316724
rect 450872 316684 450878 316696
rect 474918 316684 474924 316696
rect 474976 316684 474982 316736
rect 477954 316684 477960 316736
rect 478012 316724 478018 316736
rect 547138 316724 547144 316736
rect 478012 316696 547144 316724
rect 478012 316684 478018 316696
rect 547138 316684 547144 316696
rect 547196 316684 547202 316736
rect 453574 316616 453580 316668
rect 453632 316656 453638 316668
rect 464706 316656 464712 316668
rect 453632 316628 464712 316656
rect 453632 316616 453638 316628
rect 464706 316616 464712 316628
rect 464764 316616 464770 316668
rect 481726 316616 481732 316668
rect 481784 316656 481790 316668
rect 484394 316656 484400 316668
rect 481784 316628 484400 316656
rect 481784 316616 481790 316628
rect 484394 316616 484400 316628
rect 484452 316616 484458 316668
rect 485866 316616 485872 316668
rect 485924 316656 485930 316668
rect 486970 316656 486976 316668
rect 485924 316628 486976 316656
rect 485924 316616 485930 316628
rect 486970 316616 486976 316628
rect 487028 316616 487034 316668
rect 487522 316616 487528 316668
rect 487580 316656 487586 316668
rect 487798 316656 487804 316668
rect 487580 316628 487804 316656
rect 487580 316616 487586 316628
rect 487798 316616 487804 316628
rect 487856 316616 487862 316668
rect 487890 316616 487896 316668
rect 487948 316656 487954 316668
rect 488350 316656 488356 316668
rect 487948 316628 488356 316656
rect 487948 316616 487954 316628
rect 488350 316616 488356 316628
rect 488408 316616 488414 316668
rect 488626 316616 488632 316668
rect 488684 316656 488690 316668
rect 489178 316656 489184 316668
rect 488684 316628 489184 316656
rect 488684 316616 488690 316628
rect 489178 316616 489184 316628
rect 489236 316616 489242 316668
rect 490282 316616 490288 316668
rect 490340 316656 490346 316668
rect 490834 316656 490840 316668
rect 490340 316628 490840 316656
rect 490340 316616 490346 316628
rect 490834 316616 490840 316628
rect 490892 316616 490898 316668
rect 493318 316616 493324 316668
rect 493376 316656 493382 316668
rect 493870 316656 493876 316668
rect 493376 316628 493876 316656
rect 493376 316616 493382 316628
rect 493870 316616 493876 316628
rect 493928 316616 493934 316668
rect 494146 316616 494152 316668
rect 494204 316656 494210 316668
rect 495250 316656 495256 316668
rect 494204 316628 495256 316656
rect 494204 316616 494210 316628
rect 495250 316616 495256 316628
rect 495308 316616 495314 316668
rect 456242 316548 456248 316600
rect 456300 316588 456306 316600
rect 465258 316588 465264 316600
rect 456300 316560 465264 316588
rect 456300 316548 456306 316560
rect 465258 316548 465264 316560
rect 465316 316548 465322 316600
rect 490006 316548 490012 316600
rect 490064 316588 490070 316600
rect 491110 316588 491116 316600
rect 490064 316560 491116 316588
rect 490064 316548 490070 316560
rect 491110 316548 491116 316560
rect 491168 316548 491174 316600
rect 491386 316480 491392 316532
rect 491444 316520 491450 316532
rect 492214 316520 492220 316532
rect 491444 316492 492220 316520
rect 491444 316480 491450 316492
rect 492214 316480 492220 316492
rect 492272 316480 492278 316532
rect 457806 316004 457812 316056
rect 457864 316044 457870 316056
rect 461578 316044 461584 316056
rect 457864 316016 461584 316044
rect 457864 316004 457870 316016
rect 461578 316004 461584 316016
rect 461636 316004 461642 316056
rect 361758 315936 361764 315988
rect 361816 315976 361822 315988
rect 371878 315976 371884 315988
rect 361816 315948 371884 315976
rect 361816 315936 361822 315948
rect 371878 315936 371884 315948
rect 371936 315936 371942 315988
rect 457438 315392 457444 315444
rect 457496 315432 457502 315444
rect 489730 315432 489736 315444
rect 457496 315404 489736 315432
rect 457496 315392 457502 315404
rect 489730 315392 489736 315404
rect 489788 315392 489794 315444
rect 501598 315392 501604 315444
rect 501656 315432 501662 315444
rect 539870 315432 539876 315444
rect 501656 315404 539876 315432
rect 501656 315392 501662 315404
rect 539870 315392 539876 315404
rect 539928 315392 539934 315444
rect 459278 315324 459284 315376
rect 459336 315364 459342 315376
rect 492490 315364 492496 315376
rect 459336 315336 492496 315364
rect 459336 315324 459342 315336
rect 492490 315324 492496 315336
rect 492548 315324 492554 315376
rect 496630 315324 496636 315376
rect 496688 315364 496694 315376
rect 539686 315364 539692 315376
rect 496688 315336 539692 315364
rect 496688 315324 496694 315336
rect 539686 315324 539692 315336
rect 539744 315324 539750 315376
rect 478138 315256 478144 315308
rect 478196 315296 478202 315308
rect 551278 315296 551284 315308
rect 478196 315268 551284 315296
rect 478196 315256 478202 315268
rect 551278 315256 551284 315268
rect 551336 315256 551342 315308
rect 450998 314032 451004 314084
rect 451056 314072 451062 314084
rect 484762 314072 484768 314084
rect 451056 314044 484768 314072
rect 451056 314032 451062 314044
rect 484762 314032 484768 314044
rect 484820 314032 484826 314084
rect 503162 314032 503168 314084
rect 503220 314072 503226 314084
rect 543182 314072 543188 314084
rect 503220 314044 543188 314072
rect 503220 314032 503226 314044
rect 543182 314032 543188 314044
rect 543240 314032 543246 314084
rect 459370 313964 459376 314016
rect 459428 314004 459434 314016
rect 493594 314004 493600 314016
rect 459428 313976 493600 314004
rect 459428 313964 459434 313976
rect 493594 313964 493600 313976
rect 493652 313964 493658 314016
rect 496722 313964 496728 314016
rect 496780 314004 496786 314016
rect 540974 314004 540980 314016
rect 496780 313976 540980 314004
rect 496780 313964 496786 313976
rect 540974 313964 540980 313976
rect 541032 313964 541038 314016
rect 433150 313896 433156 313948
rect 433208 313936 433214 313948
rect 443822 313936 443828 313948
rect 433208 313908 443828 313936
rect 433208 313896 433214 313908
rect 443822 313896 443828 313908
rect 443880 313896 443886 313948
rect 455782 313896 455788 313948
rect 455840 313936 455846 313948
rect 566458 313936 566464 313948
rect 455840 313908 566464 313936
rect 455840 313896 455846 313908
rect 566458 313896 566464 313908
rect 566516 313896 566522 313948
rect 482094 313556 482100 313608
rect 482152 313596 482158 313608
rect 484486 313596 484492 313608
rect 482152 313568 484492 313596
rect 482152 313556 482158 313568
rect 484486 313556 484492 313568
rect 484544 313556 484550 313608
rect 461670 313284 461676 313336
rect 461728 313324 461734 313336
rect 463786 313324 463792 313336
rect 461728 313296 463792 313324
rect 461728 313284 461734 313296
rect 463786 313284 463792 313296
rect 463844 313284 463850 313336
rect 469030 313216 469036 313268
rect 469088 313256 469094 313268
rect 580166 313256 580172 313268
rect 469088 313228 580172 313256
rect 469088 313216 469094 313228
rect 580166 313216 580172 313228
rect 580224 313216 580230 313268
rect 439682 312536 439688 312588
rect 439740 312576 439746 312588
rect 471238 312576 471244 312588
rect 439740 312548 471244 312576
rect 439740 312536 439746 312548
rect 471238 312536 471244 312548
rect 471296 312536 471302 312588
rect 478874 312536 478880 312588
rect 478932 312576 478938 312588
rect 481726 312576 481732 312588
rect 478932 312548 481732 312576
rect 478932 312536 478938 312548
rect 481726 312536 481732 312548
rect 481784 312536 481790 312588
rect 502058 312536 502064 312588
rect 502116 312576 502122 312588
rect 542538 312576 542544 312588
rect 502116 312548 542544 312576
rect 502116 312536 502122 312548
rect 542538 312536 542544 312548
rect 542596 312536 542602 312588
rect 494606 311856 494612 311908
rect 494664 311896 494670 311908
rect 494790 311896 494796 311908
rect 494664 311868 494796 311896
rect 494664 311856 494670 311868
rect 494790 311856 494796 311868
rect 494848 311856 494854 311908
rect 469858 311244 469864 311296
rect 469916 311284 469922 311296
rect 482094 311284 482100 311296
rect 469916 311256 482100 311284
rect 469916 311244 469922 311256
rect 482094 311244 482100 311256
rect 482152 311244 482158 311296
rect 454862 311176 454868 311228
rect 454920 311216 454926 311228
rect 494422 311216 494428 311228
rect 454920 311188 494428 311216
rect 454920 311176 454926 311188
rect 494422 311176 494428 311188
rect 494480 311176 494486 311228
rect 467374 311108 467380 311160
rect 467432 311148 467438 311160
rect 548518 311148 548524 311160
rect 467432 311120 548524 311148
rect 467432 311108 467438 311120
rect 548518 311108 548524 311120
rect 548576 311108 548582 311160
rect 456518 309884 456524 309936
rect 456576 309924 456582 309936
rect 495618 309924 495624 309936
rect 456576 309896 495624 309924
rect 456576 309884 456582 309896
rect 495618 309884 495624 309896
rect 495676 309884 495682 309936
rect 503530 309884 503536 309936
rect 503588 309924 503594 309936
rect 538950 309924 538956 309936
rect 503588 309896 538956 309924
rect 503588 309884 503594 309896
rect 538950 309884 538956 309896
rect 539008 309884 539014 309936
rect 487706 309816 487712 309868
rect 487764 309856 487770 309868
rect 530026 309856 530032 309868
rect 487764 309828 530032 309856
rect 487764 309816 487770 309828
rect 530026 309816 530032 309828
rect 530084 309816 530090 309868
rect 452010 309748 452016 309800
rect 452068 309788 452074 309800
rect 494790 309788 494796 309800
rect 452068 309760 494796 309788
rect 452068 309748 452074 309760
rect 494790 309748 494796 309760
rect 494848 309748 494854 309800
rect 502150 309748 502156 309800
rect 502208 309788 502214 309800
rect 541066 309788 541072 309800
rect 502208 309760 541072 309788
rect 502208 309748 502214 309760
rect 541066 309748 541072 309760
rect 541124 309748 541130 309800
rect 453666 308456 453672 308508
rect 453724 308496 453730 308508
rect 489178 308496 489184 308508
rect 453724 308468 489184 308496
rect 453724 308456 453730 308468
rect 489178 308456 489184 308468
rect 489236 308456 489242 308508
rect 503254 308456 503260 308508
rect 503312 308496 503318 308508
rect 539042 308496 539048 308508
rect 503312 308468 539048 308496
rect 503312 308456 503318 308468
rect 539042 308456 539048 308468
rect 539100 308456 539106 308508
rect 487798 308388 487804 308440
rect 487856 308428 487862 308440
rect 529934 308428 529940 308440
rect 487856 308400 529940 308428
rect 487856 308388 487862 308400
rect 529934 308388 529940 308400
rect 529992 308388 529998 308440
rect 476758 308320 476764 308372
rect 476816 308360 476822 308372
rect 478874 308360 478880 308372
rect 476816 308332 478880 308360
rect 476816 308320 476822 308332
rect 478874 308320 478880 308332
rect 478932 308320 478938 308372
rect 3510 307708 3516 307760
rect 3568 307748 3574 307760
rect 4798 307748 4804 307760
rect 3568 307720 4804 307748
rect 3568 307708 3574 307720
rect 4798 307708 4804 307720
rect 4856 307708 4862 307760
rect 453758 307096 453764 307148
rect 453816 307136 453822 307148
rect 490282 307136 490288 307148
rect 453816 307108 490288 307136
rect 453816 307096 453822 307108
rect 490282 307096 490288 307108
rect 490340 307096 490346 307148
rect 457346 307028 457352 307080
rect 457404 307068 457410 307080
rect 576118 307068 576124 307080
rect 457404 307040 576124 307068
rect 457404 307028 457410 307040
rect 576118 307028 576124 307040
rect 576176 307028 576182 307080
rect 446122 306280 446128 306332
rect 446180 306320 446186 306332
rect 469858 306320 469864 306332
rect 446180 306292 469864 306320
rect 446180 306280 446186 306292
rect 469858 306280 469864 306292
rect 469916 306280 469922 306332
rect 457530 306212 457536 306264
rect 457588 306252 457594 306264
rect 491386 306252 491392 306264
rect 457588 306224 491392 306252
rect 457588 306212 457594 306224
rect 491386 306212 491392 306224
rect 491444 306212 491450 306264
rect 400858 306144 400864 306196
rect 400916 306184 400922 306196
rect 465442 306184 465448 306196
rect 400916 306156 465448 306184
rect 400916 306144 400922 306156
rect 465442 306144 465448 306156
rect 465500 306144 465506 306196
rect 477310 306144 477316 306196
rect 477368 306184 477374 306196
rect 544378 306184 544384 306196
rect 477368 306156 544384 306184
rect 477368 306144 477374 306156
rect 544378 306144 544384 306156
rect 544436 306144 544442 306196
rect 406654 306076 406660 306128
rect 406712 306116 406718 306128
rect 509970 306116 509976 306128
rect 406712 306088 509976 306116
rect 406712 306076 406718 306088
rect 509970 306076 509976 306088
rect 510028 306076 510034 306128
rect 406470 306008 406476 306060
rect 406528 306048 406534 306060
rect 509602 306048 509608 306060
rect 406528 306020 509608 306048
rect 406528 306008 406534 306020
rect 509602 306008 509608 306020
rect 509660 306008 509666 306060
rect 403802 305940 403808 305992
rect 403860 305980 403866 305992
rect 511166 305980 511172 305992
rect 403860 305952 511172 305980
rect 403860 305940 403866 305952
rect 511166 305940 511172 305952
rect 511224 305940 511230 305992
rect 403618 305872 403624 305924
rect 403676 305912 403682 305924
rect 511074 305912 511080 305924
rect 403676 305884 511080 305912
rect 403676 305872 403682 305884
rect 511074 305872 511080 305884
rect 511132 305872 511138 305924
rect 403894 305804 403900 305856
rect 403952 305844 403958 305856
rect 513926 305844 513932 305856
rect 403952 305816 513932 305844
rect 403952 305804 403958 305816
rect 513926 305804 513932 305816
rect 513984 305804 513990 305856
rect 403710 305736 403716 305788
rect 403768 305776 403774 305788
rect 515582 305776 515588 305788
rect 403768 305748 515588 305776
rect 403768 305736 403774 305748
rect 515582 305736 515588 305748
rect 515640 305736 515646 305788
rect 363598 305668 363604 305720
rect 363656 305708 363662 305720
rect 512730 305708 512736 305720
rect 363656 305680 512736 305708
rect 363656 305668 363662 305680
rect 512730 305668 512736 305680
rect 512788 305668 512794 305720
rect 360838 305600 360844 305652
rect 360896 305640 360902 305652
rect 512638 305640 512644 305652
rect 360896 305612 512644 305640
rect 360896 305600 360902 305612
rect 512638 305600 512644 305612
rect 512696 305600 512702 305652
rect 361758 304920 361764 304972
rect 361816 304960 361822 304972
rect 431218 304960 431224 304972
rect 361816 304932 431224 304960
rect 361816 304920 361822 304932
rect 431218 304920 431224 304932
rect 431276 304920 431282 304972
rect 450446 304580 450452 304632
rect 450504 304620 450510 304632
rect 455966 304620 455972 304632
rect 450504 304592 455972 304620
rect 450504 304580 450510 304592
rect 455966 304580 455972 304592
rect 456024 304580 456030 304632
rect 444742 304512 444748 304564
rect 444800 304552 444806 304564
rect 461670 304552 461676 304564
rect 444800 304524 461676 304552
rect 444800 304512 444806 304524
rect 461670 304512 461676 304524
rect 461728 304512 461734 304564
rect 455874 304444 455880 304496
rect 455932 304484 455938 304496
rect 562318 304484 562324 304496
rect 455932 304456 562324 304484
rect 455932 304444 455938 304456
rect 562318 304444 562324 304456
rect 562376 304444 562382 304496
rect 363690 304376 363696 304428
rect 363748 304416 363754 304428
rect 512362 304416 512368 304428
rect 363748 304388 512368 304416
rect 363748 304376 363754 304388
rect 512362 304376 512368 304388
rect 512420 304376 512426 304428
rect 360930 304308 360936 304360
rect 360988 304348 360994 304360
rect 511994 304348 512000 304360
rect 360988 304320 512000 304348
rect 360988 304308 360994 304320
rect 511994 304308 512000 304320
rect 512052 304308 512058 304360
rect 361022 304240 361028 304292
rect 361080 304280 361086 304292
rect 512178 304280 512184 304292
rect 361080 304252 512184 304280
rect 361080 304240 361086 304252
rect 512178 304240 512184 304252
rect 512236 304240 512242 304292
rect 401042 303560 401048 303612
rect 401100 303600 401106 303612
rect 510982 303600 510988 303612
rect 401100 303572 510988 303600
rect 401100 303560 401106 303572
rect 510982 303560 510988 303572
rect 511040 303560 511046 303612
rect 403986 303492 403992 303544
rect 404044 303532 404050 303544
rect 515214 303532 515220 303544
rect 404044 303504 515220 303532
rect 404044 303492 404050 303504
rect 515214 303492 515220 303504
rect 515272 303492 515278 303544
rect 401134 303424 401140 303476
rect 401192 303464 401198 303476
rect 513742 303464 513748 303476
rect 401192 303436 513748 303464
rect 401192 303424 401198 303436
rect 513742 303424 513748 303436
rect 513800 303424 513806 303476
rect 395614 303356 395620 303408
rect 395672 303396 395678 303408
rect 510706 303396 510712 303408
rect 395672 303368 510712 303396
rect 395672 303356 395678 303368
rect 510706 303356 510712 303368
rect 510764 303356 510770 303408
rect 398282 303288 398288 303340
rect 398340 303328 398346 303340
rect 514202 303328 514208 303340
rect 398340 303300 514208 303328
rect 398340 303288 398346 303300
rect 514202 303288 514208 303300
rect 514260 303288 514266 303340
rect 456610 303220 456616 303272
rect 456668 303260 456674 303272
rect 571978 303260 571984 303272
rect 456668 303232 571984 303260
rect 456668 303220 456674 303232
rect 571978 303220 571984 303232
rect 572036 303220 572042 303272
rect 398098 303152 398104 303204
rect 398156 303192 398162 303204
rect 513650 303192 513656 303204
rect 398156 303164 513656 303192
rect 398156 303152 398162 303164
rect 513650 303152 513656 303164
rect 513708 303152 513714 303204
rect 398374 303084 398380 303136
rect 398432 303124 398438 303136
rect 514938 303124 514944 303136
rect 398432 303096 514944 303124
rect 398432 303084 398438 303096
rect 514938 303084 514944 303096
rect 514996 303084 515002 303136
rect 398190 303016 398196 303068
rect 398248 303056 398254 303068
rect 514846 303056 514852 303068
rect 398248 303028 514852 303056
rect 398248 303016 398254 303028
rect 514846 303016 514852 303028
rect 514904 303016 514910 303068
rect 395798 302948 395804 303000
rect 395856 302988 395862 303000
rect 517606 302988 517612 303000
rect 395856 302960 517612 302988
rect 395856 302948 395862 302960
rect 517606 302948 517612 302960
rect 517664 302948 517670 303000
rect 361114 302880 361120 302932
rect 361172 302920 361178 302932
rect 512454 302920 512460 302932
rect 361172 302892 512460 302920
rect 361172 302880 361178 302892
rect 512454 302880 512460 302892
rect 512512 302880 512518 302932
rect 401318 302812 401324 302864
rect 401376 302852 401382 302864
rect 510798 302852 510804 302864
rect 401376 302824 510804 302852
rect 401376 302812 401382 302824
rect 510798 302812 510804 302824
rect 510856 302812 510862 302864
rect 400950 302744 400956 302796
rect 401008 302784 401014 302796
rect 509418 302784 509424 302796
rect 401008 302756 509424 302784
rect 401008 302744 401014 302756
rect 509418 302744 509424 302756
rect 509476 302744 509482 302796
rect 395430 302676 395436 302728
rect 395488 302716 395494 302728
rect 485866 302716 485872 302728
rect 395488 302688 485872 302716
rect 395488 302676 395494 302688
rect 485866 302676 485872 302688
rect 485924 302676 485930 302728
rect 456702 301520 456708 301572
rect 456760 301560 456766 301572
rect 573358 301560 573364 301572
rect 456760 301532 573364 301560
rect 456760 301520 456766 301532
rect 573358 301520 573364 301532
rect 573416 301520 573422 301572
rect 362218 301452 362224 301504
rect 362276 301492 362282 301504
rect 512270 301492 512276 301504
rect 362276 301464 512276 301492
rect 362276 301452 362282 301464
rect 512270 301452 512276 301464
rect 512328 301452 512334 301504
rect 440970 300636 440976 300688
rect 441028 300676 441034 300688
rect 446122 300676 446128 300688
rect 441028 300648 446128 300676
rect 441028 300636 441034 300648
rect 446122 300636 446128 300648
rect 446180 300636 446186 300688
rect 457990 300636 457996 300688
rect 458048 300676 458054 300688
rect 533430 300676 533436 300688
rect 458048 300648 533436 300676
rect 458048 300636 458054 300648
rect 533430 300636 533436 300648
rect 533488 300636 533494 300688
rect 395706 300568 395712 300620
rect 395764 300608 395770 300620
rect 516962 300608 516968 300620
rect 395764 300580 516968 300608
rect 395764 300568 395770 300580
rect 516962 300568 516968 300580
rect 517020 300568 517026 300620
rect 393038 300500 393044 300552
rect 393096 300540 393102 300552
rect 516594 300540 516600 300552
rect 393096 300512 516600 300540
rect 393096 300500 393102 300512
rect 516594 300500 516600 300512
rect 516652 300500 516658 300552
rect 392670 300432 392676 300484
rect 392728 300472 392734 300484
rect 516870 300472 516876 300484
rect 392728 300444 516876 300472
rect 392728 300432 392734 300444
rect 516870 300432 516876 300444
rect 516928 300432 516934 300484
rect 392854 300364 392860 300416
rect 392912 300404 392918 300416
rect 518342 300404 518348 300416
rect 392912 300376 518348 300404
rect 392912 300364 392918 300376
rect 518342 300364 518348 300376
rect 518400 300364 518406 300416
rect 390186 300296 390192 300348
rect 390244 300336 390250 300348
rect 516502 300336 516508 300348
rect 390244 300308 516508 300336
rect 390244 300296 390250 300308
rect 516502 300296 516508 300308
rect 516560 300296 516566 300348
rect 389910 300228 389916 300280
rect 389968 300268 389974 300280
rect 516318 300268 516324 300280
rect 389968 300240 516324 300268
rect 389968 300228 389974 300240
rect 516318 300228 516324 300240
rect 516376 300228 516382 300280
rect 390278 300160 390284 300212
rect 390336 300200 390342 300212
rect 518066 300200 518072 300212
rect 390336 300172 518072 300200
rect 390336 300160 390342 300172
rect 518066 300160 518072 300172
rect 518124 300160 518130 300212
rect 389818 300092 389824 300144
rect 389876 300132 389882 300144
rect 517974 300132 517980 300144
rect 389876 300104 517980 300132
rect 389876 300092 389882 300104
rect 517974 300092 517980 300104
rect 518032 300092 518038 300144
rect 436922 299548 436928 299600
rect 436980 299588 436986 299600
rect 439682 299588 439688 299600
rect 436980 299560 439688 299588
rect 436980 299548 436986 299560
rect 439682 299548 439688 299560
rect 439740 299548 439746 299600
rect 461578 299412 461584 299464
rect 461636 299452 461642 299464
rect 580166 299452 580172 299464
rect 461636 299424 580172 299452
rect 461636 299412 461642 299424
rect 580166 299412 580172 299424
rect 580224 299412 580230 299464
rect 387426 298052 387432 298104
rect 387484 298092 387490 298104
rect 513558 298092 513564 298104
rect 387484 298064 513564 298092
rect 387484 298052 387490 298064
rect 513558 298052 513564 298064
rect 513616 298052 513622 298104
rect 390002 297984 390008 298036
rect 390060 298024 390066 298036
rect 517882 298024 517888 298036
rect 390060 297996 517888 298024
rect 390060 297984 390066 297996
rect 517882 297984 517888 297996
rect 517940 297984 517946 298036
rect 387334 297916 387340 297968
rect 387392 297956 387398 297968
rect 516226 297956 516232 297968
rect 387392 297928 516232 297956
rect 387392 297916 387398 297928
rect 516226 297916 516232 297928
rect 516284 297916 516290 297968
rect 384390 297848 384396 297900
rect 384448 297888 384454 297900
rect 513374 297888 513380 297900
rect 384448 297860 513380 297888
rect 384448 297848 384454 297860
rect 513374 297848 513380 297860
rect 513432 297848 513438 297900
rect 387518 297780 387524 297832
rect 387576 297820 387582 297832
rect 519262 297820 519268 297832
rect 387576 297792 519268 297820
rect 387576 297780 387582 297792
rect 519262 297780 519268 297792
rect 519320 297780 519326 297832
rect 387150 297712 387156 297764
rect 387208 297752 387214 297764
rect 519170 297752 519176 297764
rect 387208 297724 519176 297752
rect 387208 297712 387214 297724
rect 519170 297712 519176 297724
rect 519228 297712 519234 297764
rect 381722 297644 381728 297696
rect 381780 297684 381786 297696
rect 514754 297684 514760 297696
rect 381780 297656 514760 297684
rect 381780 297644 381786 297656
rect 514754 297644 514760 297656
rect 514812 297644 514818 297696
rect 387242 297576 387248 297628
rect 387300 297616 387306 297628
rect 520550 297616 520556 297628
rect 387300 297588 520556 297616
rect 387300 297576 387306 297588
rect 520550 297576 520556 297588
rect 520608 297576 520614 297628
rect 384298 297508 384304 297560
rect 384356 297548 384362 297560
rect 519078 297548 519084 297560
rect 384356 297520 519084 297548
rect 384356 297508 384362 297520
rect 519078 297508 519084 297520
rect 519136 297508 519142 297560
rect 384482 297440 384488 297492
rect 384540 297480 384546 297492
rect 520274 297480 520280 297492
rect 384540 297452 520280 297480
rect 384540 297440 384546 297452
rect 520274 297440 520280 297452
rect 520332 297440 520338 297492
rect 384574 297372 384580 297424
rect 384632 297412 384638 297424
rect 520366 297412 520372 297424
rect 384632 297384 520372 297412
rect 384632 297372 384638 297384
rect 520366 297372 520372 297384
rect 520424 297372 520430 297424
rect 387058 297304 387064 297356
rect 387116 297344 387122 297356
rect 509694 297344 509700 297356
rect 387116 297316 509700 297344
rect 387116 297304 387122 297316
rect 509694 297304 509700 297316
rect 509752 297304 509758 297356
rect 390094 297236 390100 297288
rect 390152 297276 390158 297288
rect 510890 297276 510896 297288
rect 390152 297248 510896 297276
rect 390152 297236 390158 297248
rect 510890 297236 510896 297248
rect 510948 297236 510954 297288
rect 439682 297168 439688 297220
rect 439740 297208 439746 297220
rect 444742 297208 444748 297220
rect 439740 297180 444748 297208
rect 439740 297168 439746 297180
rect 444742 297168 444748 297180
rect 444800 297168 444806 297220
rect 457622 297168 457628 297220
rect 457680 297208 457686 297220
rect 574830 297208 574836 297220
rect 457680 297180 574836 297208
rect 457680 297168 457686 297180
rect 574830 297168 574836 297180
rect 574888 297168 574894 297220
rect 477402 295944 477408 295996
rect 477460 295984 477466 295996
rect 570598 295984 570604 295996
rect 477460 295956 570604 295984
rect 477460 295944 477466 295956
rect 570598 295944 570604 295956
rect 570656 295944 570662 295996
rect 381906 295264 381912 295316
rect 381964 295304 381970 295316
rect 510062 295304 510068 295316
rect 381964 295276 510068 295304
rect 381964 295264 381970 295276
rect 510062 295264 510068 295276
rect 510120 295264 510126 295316
rect 376018 295196 376024 295248
rect 376076 295236 376082 295248
rect 507486 295236 507492 295248
rect 376076 295208 507492 295236
rect 376076 295196 376082 295208
rect 507486 295196 507492 295208
rect 507544 295196 507550 295248
rect 381814 295128 381820 295180
rect 381872 295168 381878 295180
rect 517514 295168 517520 295180
rect 381872 295140 517520 295168
rect 381872 295128 381878 295140
rect 517514 295128 517520 295140
rect 517572 295128 517578 295180
rect 381998 295060 382004 295112
rect 382056 295100 382062 295112
rect 518894 295100 518900 295112
rect 382056 295072 518900 295100
rect 382056 295060 382062 295072
rect 518894 295060 518900 295072
rect 518952 295060 518958 295112
rect 378870 294992 378876 295044
rect 378928 295032 378934 295044
rect 516686 295032 516692 295044
rect 378928 295004 516692 295032
rect 378928 294992 378934 295004
rect 516686 294992 516692 295004
rect 516744 294992 516750 295044
rect 376202 294924 376208 294976
rect 376260 294964 376266 294976
rect 515306 294964 515312 294976
rect 376260 294936 515312 294964
rect 376260 294924 376266 294936
rect 515306 294924 515312 294936
rect 515364 294924 515370 294976
rect 376110 294856 376116 294908
rect 376168 294896 376174 294908
rect 516410 294896 516416 294908
rect 376168 294868 516416 294896
rect 376168 294856 376174 294868
rect 516410 294856 516416 294868
rect 516468 294856 516474 294908
rect 379054 294788 379060 294840
rect 379112 294828 379118 294840
rect 519722 294828 519728 294840
rect 379112 294800 519728 294828
rect 379112 294788 379118 294800
rect 519722 294788 519728 294800
rect 519780 294788 519786 294840
rect 379238 294720 379244 294772
rect 379296 294760 379302 294772
rect 520734 294760 520740 294772
rect 379296 294732 520740 294760
rect 379296 294720 379302 294732
rect 520734 294720 520740 294732
rect 520792 294720 520798 294772
rect 379146 294652 379152 294704
rect 379204 294692 379210 294704
rect 520826 294692 520832 294704
rect 379204 294664 520832 294692
rect 379204 294652 379210 294664
rect 520826 294652 520832 294664
rect 520884 294652 520890 294704
rect 376294 294584 376300 294636
rect 376352 294624 376358 294636
rect 519446 294624 519452 294636
rect 376352 294596 519452 294624
rect 376352 294584 376358 294596
rect 519446 294584 519452 294596
rect 519504 294584 519510 294636
rect 396718 294516 396724 294568
rect 396776 294556 396782 294568
rect 486418 294556 486424 294568
rect 396776 294528 486424 294556
rect 396776 294516 396782 294528
rect 486418 294516 486424 294528
rect 486476 294516 486482 294568
rect 447870 294448 447876 294500
rect 447928 294488 447934 294500
rect 536098 294488 536104 294500
rect 447928 294460 536104 294488
rect 447928 294448 447934 294460
rect 536098 294448 536104 294460
rect 536156 294448 536162 294500
rect 361758 293904 361764 293956
rect 361816 293944 361822 293956
rect 435358 293944 435364 293956
rect 361816 293916 435364 293944
rect 361816 293904 361822 293916
rect 435358 293904 435364 293916
rect 435416 293904 435422 293956
rect 467282 293224 467288 293276
rect 467340 293264 467346 293276
rect 555418 293264 555424 293276
rect 467340 293236 555424 293264
rect 467340 293224 467346 293236
rect 555418 293224 555424 293236
rect 555476 293224 555482 293276
rect 3418 292544 3424 292596
rect 3476 292584 3482 292596
rect 4890 292584 4896 292596
rect 3476 292556 4896 292584
rect 3476 292544 3482 292556
rect 4890 292544 4896 292556
rect 4948 292544 4954 292596
rect 437474 292544 437480 292596
rect 437532 292584 437538 292596
rect 440970 292584 440976 292596
rect 437532 292556 440976 292584
rect 437532 292544 437538 292556
rect 440970 292544 440976 292556
rect 441028 292544 441034 292596
rect 376386 292476 376392 292528
rect 376444 292516 376450 292528
rect 515030 292516 515036 292528
rect 376444 292488 515036 292516
rect 376444 292476 376450 292488
rect 515030 292476 515036 292488
rect 515088 292476 515094 292528
rect 376478 292408 376484 292460
rect 376536 292448 376542 292460
rect 520642 292448 520648 292460
rect 376536 292420 520648 292448
rect 376536 292408 376542 292420
rect 520642 292408 520648 292420
rect 520700 292408 520706 292460
rect 373534 292340 373540 292392
rect 373592 292380 373598 292392
rect 517790 292380 517796 292392
rect 373592 292352 517796 292380
rect 373592 292340 373598 292352
rect 517790 292340 517796 292352
rect 517848 292340 517854 292392
rect 373258 292272 373264 292324
rect 373316 292312 373322 292324
rect 517698 292312 517704 292324
rect 373316 292284 517704 292312
rect 373316 292272 373322 292284
rect 517698 292272 517704 292284
rect 517756 292272 517762 292324
rect 373442 292204 373448 292256
rect 373500 292244 373506 292256
rect 519354 292244 519360 292256
rect 373500 292216 519360 292244
rect 373500 292204 373506 292216
rect 519354 292204 519360 292216
rect 519412 292204 519418 292256
rect 370866 292136 370872 292188
rect 370924 292176 370930 292188
rect 518986 292176 518992 292188
rect 370924 292148 518992 292176
rect 370924 292136 370930 292148
rect 518986 292136 518992 292148
rect 519044 292136 519050 292188
rect 370590 292068 370596 292120
rect 370648 292108 370654 292120
rect 520458 292108 520464 292120
rect 370648 292080 520464 292108
rect 370648 292068 370654 292080
rect 520458 292068 520464 292080
rect 520516 292068 520522 292120
rect 370774 292000 370780 292052
rect 370832 292040 370838 292052
rect 521746 292040 521752 292052
rect 370832 292012 521752 292040
rect 370832 292000 370838 292012
rect 521746 292000 521752 292012
rect 521804 292000 521810 292052
rect 370958 291932 370964 291984
rect 371016 291972 371022 291984
rect 523034 291972 523040 291984
rect 371016 291944 523040 291972
rect 371016 291932 371022 291944
rect 523034 291932 523040 291944
rect 523092 291932 523098 291984
rect 370498 291864 370504 291916
rect 370556 291904 370562 291916
rect 523126 291904 523132 291916
rect 370556 291876 523132 291904
rect 370556 291864 370562 291876
rect 523126 291864 523132 291876
rect 523184 291864 523190 291916
rect 368014 291796 368020 291848
rect 368072 291836 368078 291848
rect 521654 291836 521660 291848
rect 368072 291808 521660 291836
rect 368072 291796 368078 291808
rect 521654 291796 521660 291808
rect 521712 291796 521718 291848
rect 370682 291728 370688 291780
rect 370740 291768 370746 291780
rect 507394 291768 507400 291780
rect 370740 291740 507400 291768
rect 370740 291728 370746 291740
rect 507394 291728 507400 291740
rect 507452 291728 507458 291780
rect 373350 291660 373356 291712
rect 373408 291700 373414 291712
rect 507302 291700 507308 291712
rect 373408 291672 507308 291700
rect 373408 291660 373414 291672
rect 507302 291660 507308 291672
rect 507360 291660 507366 291712
rect 478414 291592 478420 291644
rect 478472 291632 478478 291644
rect 559650 291632 559656 291644
rect 478472 291604 559656 291632
rect 478472 291592 478478 291604
rect 559650 291592 559656 291604
rect 559708 291592 559714 291644
rect 467006 290436 467012 290488
rect 467064 290476 467070 290488
rect 558178 290476 558184 290488
rect 467064 290448 558184 290476
rect 467064 290436 467070 290448
rect 558178 290436 558184 290448
rect 558236 290436 558242 290488
rect 427078 289552 427084 289604
rect 427136 289592 427142 289604
rect 437474 289592 437480 289604
rect 427136 289564 437480 289592
rect 427136 289552 427142 289564
rect 437474 289552 437480 289564
rect 437532 289552 437538 289604
rect 447778 289552 447784 289604
rect 447836 289592 447842 289604
rect 464062 289592 464068 289604
rect 447836 289564 464068 289592
rect 447836 289552 447842 289564
rect 464062 289552 464068 289564
rect 464120 289552 464126 289604
rect 407758 289484 407764 289536
rect 407816 289524 407822 289536
rect 507210 289524 507216 289536
rect 407816 289496 507216 289524
rect 407816 289484 407822 289496
rect 507210 289484 507216 289496
rect 507268 289484 507274 289536
rect 365346 289416 365352 289468
rect 365404 289456 365410 289468
rect 507118 289456 507124 289468
rect 365404 289428 507124 289456
rect 365404 289416 365410 289428
rect 507118 289416 507124 289428
rect 507176 289416 507182 289468
rect 368198 289348 368204 289400
rect 368256 289388 368262 289400
rect 522206 289388 522212 289400
rect 368256 289360 522212 289388
rect 368256 289348 368262 289360
rect 522206 289348 522212 289360
rect 522264 289348 522270 289400
rect 365254 289280 365260 289332
rect 365312 289320 365318 289332
rect 521838 289320 521844 289332
rect 365312 289292 521844 289320
rect 365312 289280 365318 289292
rect 521838 289280 521844 289292
rect 521896 289280 521902 289332
rect 365070 289212 365076 289264
rect 365128 289252 365134 289264
rect 521930 289252 521936 289264
rect 365128 289224 521936 289252
rect 365128 289212 365134 289224
rect 521930 289212 521936 289224
rect 521988 289212 521994 289264
rect 365162 289144 365168 289196
rect 365220 289184 365226 289196
rect 522114 289184 522120 289196
rect 365220 289156 522120 289184
rect 365220 289144 365226 289156
rect 522114 289144 522120 289156
rect 522172 289144 522178 289196
rect 364978 289076 364984 289128
rect 365036 289116 365042 289128
rect 522022 289116 522028 289128
rect 365036 289088 522028 289116
rect 365036 289076 365042 289088
rect 522022 289076 522028 289088
rect 522080 289076 522086 289128
rect 488350 287648 488356 287700
rect 488408 287688 488414 287700
rect 531314 287688 531320 287700
rect 488408 287660 531320 287688
rect 488408 287648 488414 287660
rect 531314 287648 531320 287660
rect 531372 287648 531378 287700
rect 381630 286356 381636 286408
rect 381688 286396 381694 286408
rect 476482 286396 476488 286408
rect 381688 286368 476488 286396
rect 381688 286356 381694 286368
rect 476482 286356 476488 286368
rect 476540 286356 476546 286408
rect 500126 286356 500132 286408
rect 500184 286396 500190 286408
rect 541158 286396 541164 286408
rect 500184 286368 541164 286396
rect 500184 286356 500190 286368
rect 541158 286356 541164 286368
rect 541216 286356 541222 286408
rect 410518 286288 410524 286340
rect 410576 286328 410582 286340
rect 436922 286328 436928 286340
rect 410576 286300 436928 286328
rect 410576 286288 410582 286300
rect 436922 286288 436928 286300
rect 436980 286288 436986 286340
rect 467650 286288 467656 286340
rect 467708 286328 467714 286340
rect 580258 286328 580264 286340
rect 467708 286300 580264 286328
rect 467708 286288 467714 286300
rect 580258 286288 580264 286300
rect 580316 286288 580322 286340
rect 469214 284996 469220 285048
rect 469272 285036 469278 285048
rect 476758 285036 476764 285048
rect 469272 285008 476764 285036
rect 469272 284996 469278 285008
rect 476758 284996 476764 285008
rect 476816 284996 476822 285048
rect 498838 284996 498844 285048
rect 498896 285036 498902 285048
rect 539962 285036 539968 285048
rect 498896 285008 539968 285036
rect 498896 284996 498902 285008
rect 539962 284996 539968 285008
rect 540020 284996 540026 285048
rect 466822 284928 466828 284980
rect 466880 284968 466886 284980
rect 559558 284968 559564 284980
rect 466880 284940 559564 284968
rect 466880 284928 466886 284940
rect 559558 284928 559564 284940
rect 559616 284928 559622 284980
rect 452286 283568 452292 283620
rect 452344 283608 452350 283620
rect 494698 283608 494704 283620
rect 452344 283580 494704 283608
rect 452344 283568 452350 283580
rect 494698 283568 494704 283580
rect 494756 283568 494762 283620
rect 361758 282820 361764 282872
rect 361816 282860 361822 282872
rect 436830 282860 436836 282872
rect 361816 282832 436836 282860
rect 361816 282820 361822 282832
rect 436830 282820 436836 282832
rect 436888 282820 436894 282872
rect 459462 282140 459468 282192
rect 459520 282180 459526 282192
rect 488994 282180 489000 282192
rect 459520 282152 489000 282180
rect 459520 282140 459526 282152
rect 488994 282140 489000 282152
rect 489052 282140 489058 282192
rect 462958 281868 462964 281920
rect 463016 281908 463022 281920
rect 469214 281908 469220 281920
rect 463016 281880 469220 281908
rect 463016 281868 463022 281880
rect 469214 281868 469220 281880
rect 469272 281868 469278 281920
rect 455046 280780 455052 280832
rect 455104 280820 455110 280832
rect 493410 280820 493416 280832
rect 455104 280792 493416 280820
rect 455104 280780 455110 280792
rect 493410 280780 493416 280792
rect 493468 280780 493474 280832
rect 497642 280780 497648 280832
rect 497700 280820 497706 280832
rect 542446 280820 542452 280832
rect 497700 280792 542452 280820
rect 497700 280780 497706 280792
rect 542446 280780 542452 280792
rect 542504 280780 542510 280832
rect 447870 279488 447876 279540
rect 447928 279528 447934 279540
rect 462958 279528 462964 279540
rect 447928 279500 462964 279528
rect 447928 279488 447934 279500
rect 462958 279488 462964 279500
rect 463016 279488 463022 279540
rect 453942 279420 453948 279472
rect 454000 279460 454006 279472
rect 490558 279460 490564 279472
rect 454000 279432 490564 279460
rect 454000 279420 454006 279432
rect 490558 279420 490564 279432
rect 490616 279420 490622 279472
rect 498010 279420 498016 279472
rect 498068 279460 498074 279472
rect 543274 279460 543280 279472
rect 498068 279432 543280 279460
rect 498068 279420 498074 279432
rect 543274 279420 543280 279432
rect 543332 279420 543338 279472
rect 452378 277992 452384 278044
rect 452436 278032 452442 278044
rect 494146 278032 494152 278044
rect 452436 278004 494152 278032
rect 452436 277992 452442 278004
rect 494146 277992 494152 278004
rect 494204 277992 494210 278044
rect 455230 276632 455236 276684
rect 455288 276672 455294 276684
rect 494514 276672 494520 276684
rect 455288 276644 494520 276672
rect 455288 276632 455294 276644
rect 494514 276632 494520 276644
rect 494572 276632 494578 276684
rect 499942 276632 499948 276684
rect 500000 276672 500006 276684
rect 540054 276672 540060 276684
rect 500000 276644 540060 276672
rect 500000 276632 500006 276644
rect 540054 276632 540060 276644
rect 540112 276632 540118 276684
rect 488074 275340 488080 275392
rect 488132 275380 488138 275392
rect 530118 275380 530124 275392
rect 488132 275352 530124 275380
rect 488132 275340 488138 275352
rect 530118 275340 530124 275352
rect 530176 275340 530182 275392
rect 458634 275272 458640 275324
rect 458692 275312 458698 275324
rect 493318 275312 493324 275324
rect 458692 275284 493324 275312
rect 458692 275272 458698 275284
rect 493318 275272 493324 275284
rect 493376 275272 493382 275324
rect 499022 275272 499028 275324
rect 499080 275312 499086 275324
rect 541250 275312 541256 275324
rect 499080 275284 541256 275312
rect 499080 275272 499086 275284
rect 541250 275272 541256 275284
rect 541308 275272 541314 275324
rect 453850 273980 453856 274032
rect 453908 274020 453914 274032
rect 488626 274020 488632 274032
rect 453908 273992 488632 274020
rect 453908 273980 453914 273992
rect 488626 273980 488632 273992
rect 488684 273980 488690 274032
rect 431218 273912 431224 273964
rect 431276 273952 431282 273964
rect 439682 273952 439688 273964
rect 431276 273924 439688 273952
rect 431276 273912 431282 273924
rect 439682 273912 439688 273924
rect 439740 273912 439746 273964
rect 454954 273912 454960 273964
rect 455012 273952 455018 273964
rect 491662 273952 491668 273964
rect 455012 273924 491668 273952
rect 455012 273912 455018 273924
rect 491662 273912 491668 273924
rect 491720 273912 491726 273964
rect 499390 273912 499396 273964
rect 499448 273952 499454 273964
rect 541342 273952 541348 273964
rect 499448 273924 541348 273952
rect 499448 273912 499454 273924
rect 541342 273912 541348 273924
rect 541400 273912 541406 273964
rect 479518 273164 479524 273216
rect 479576 273204 479582 273216
rect 579890 273204 579896 273216
rect 479576 273176 579896 273204
rect 479576 273164 479582 273176
rect 579890 273164 579896 273176
rect 579948 273164 579954 273216
rect 455138 272552 455144 272604
rect 455196 272592 455202 272604
rect 492766 272592 492772 272604
rect 455196 272564 492772 272592
rect 455196 272552 455202 272564
rect 492766 272552 492772 272564
rect 492824 272552 492830 272604
rect 452102 272484 452108 272536
rect 452160 272524 452166 272536
rect 490098 272524 490104 272536
rect 452160 272496 490104 272524
rect 452160 272484 452166 272496
rect 490098 272484 490104 272496
rect 490156 272484 490162 272536
rect 500770 272484 500776 272536
rect 500828 272524 500834 272536
rect 541434 272524 541440 272536
rect 500828 272496 541440 272524
rect 500828 272484 500834 272496
rect 541434 272484 541440 272496
rect 541492 272484 541498 272536
rect 361758 271804 361764 271856
rect 361816 271844 361822 271856
rect 432598 271844 432604 271856
rect 361816 271816 432604 271844
rect 361816 271804 361822 271816
rect 432598 271804 432604 271816
rect 432656 271804 432662 271856
rect 458726 271260 458732 271312
rect 458784 271300 458790 271312
rect 488902 271300 488908 271312
rect 458784 271272 488908 271300
rect 458784 271260 458790 271272
rect 488902 271260 488908 271272
rect 488960 271260 488966 271312
rect 456610 271192 456616 271244
rect 456668 271232 456674 271244
rect 490006 271232 490012 271244
rect 456668 271204 490012 271232
rect 456668 271192 456674 271204
rect 490006 271192 490012 271204
rect 490064 271192 490070 271244
rect 500494 271192 500500 271244
rect 500552 271232 500558 271244
rect 540238 271232 540244 271244
rect 500552 271204 540244 271232
rect 500552 271192 500558 271204
rect 540238 271192 540244 271204
rect 540296 271192 540302 271244
rect 457622 271124 457628 271176
rect 457680 271164 457686 271176
rect 493134 271164 493140 271176
rect 457680 271136 493140 271164
rect 457680 271124 457686 271136
rect 493134 271124 493140 271136
rect 493192 271124 493198 271176
rect 499114 271124 499120 271176
rect 499172 271164 499178 271176
rect 540146 271164 540152 271176
rect 499172 271136 540152 271164
rect 499172 271124 499178 271136
rect 540146 271124 540152 271136
rect 540204 271124 540210 271176
rect 456702 269900 456708 269952
rect 456760 269940 456766 269952
rect 487246 269940 487252 269952
rect 456760 269912 487252 269940
rect 456760 269900 456766 269912
rect 487246 269900 487252 269912
rect 487304 269900 487310 269952
rect 505002 269900 505008 269952
rect 505060 269940 505066 269952
rect 543734 269940 543740 269952
rect 505060 269912 543740 269940
rect 505060 269900 505066 269912
rect 543734 269900 543740 269912
rect 543792 269900 543798 269952
rect 400122 269832 400128 269884
rect 400180 269872 400186 269884
rect 410518 269872 410524 269884
rect 400180 269844 410524 269872
rect 400180 269832 400186 269844
rect 410518 269832 410524 269844
rect 410576 269832 410582 269884
rect 468754 269832 468760 269884
rect 468812 269872 468818 269884
rect 580350 269872 580356 269884
rect 468812 269844 580356 269872
rect 468812 269832 468818 269844
rect 580350 269832 580356 269844
rect 580408 269832 580414 269884
rect 359458 269764 359464 269816
rect 359516 269804 359522 269816
rect 512822 269804 512828 269816
rect 359516 269776 512828 269804
rect 359516 269764 359522 269776
rect 512822 269764 512828 269776
rect 512880 269764 512886 269816
rect 452194 268404 452200 268456
rect 452252 268444 452258 268456
rect 490374 268444 490380 268456
rect 452252 268416 490380 268444
rect 452252 268404 452258 268416
rect 490374 268404 490380 268416
rect 490432 268404 490438 268456
rect 497734 268404 497740 268456
rect 497792 268444 497798 268456
rect 542814 268444 542820 268456
rect 497792 268416 542820 268444
rect 497792 268404 497798 268416
rect 542814 268404 542820 268416
rect 542872 268404 542878 268456
rect 466362 268336 466368 268388
rect 466420 268376 466426 268388
rect 574738 268376 574744 268388
rect 466420 268348 574744 268376
rect 466420 268336 466426 268348
rect 574738 268336 574744 268348
rect 574796 268336 574802 268388
rect 445018 264936 445024 264988
rect 445076 264976 445082 264988
rect 447870 264976 447876 264988
rect 445076 264948 447876 264976
rect 445076 264936 445082 264948
rect 447870 264936 447876 264948
rect 447928 264936 447934 264988
rect 396810 263576 396816 263628
rect 396868 263616 396874 263628
rect 400122 263616 400128 263628
rect 396868 263588 400128 263616
rect 396868 263576 396874 263588
rect 400122 263576 400128 263588
rect 400180 263576 400186 263628
rect 449802 263508 449808 263560
rect 449860 263548 449866 263560
rect 456794 263548 456800 263560
rect 449860 263520 456800 263548
rect 449860 263508 449866 263520
rect 456794 263508 456800 263520
rect 456852 263508 456858 263560
rect 417418 262828 417424 262880
rect 417476 262868 417482 262880
rect 427078 262868 427084 262880
rect 417476 262840 427084 262868
rect 417476 262828 417482 262840
rect 427078 262828 427084 262840
rect 427136 262828 427142 262880
rect 444650 262216 444656 262268
rect 444708 262256 444714 262268
rect 447778 262256 447784 262268
rect 444708 262228 447784 262256
rect 444708 262216 444714 262228
rect 447778 262216 447784 262228
rect 447836 262216 447842 262268
rect 361758 260788 361764 260840
rect 361816 260828 361822 260840
rect 440878 260828 440884 260840
rect 361816 260800 440884 260828
rect 361816 260788 361822 260800
rect 440878 260788 440884 260800
rect 440936 260788 440942 260840
rect 406838 260108 406844 260160
rect 406896 260148 406902 260160
rect 417418 260148 417424 260160
rect 406896 260120 417424 260148
rect 406896 260108 406902 260120
rect 417418 260108 417424 260120
rect 417476 260108 417482 260160
rect 439682 258680 439688 258732
rect 439740 258720 439746 258732
rect 444650 258720 444656 258732
rect 439740 258692 444656 258720
rect 439740 258680 439746 258692
rect 444650 258680 444656 258692
rect 444708 258680 444714 258732
rect 3970 253920 3976 253972
rect 4028 253960 4034 253972
rect 5074 253960 5080 253972
rect 4028 253932 5080 253960
rect 4028 253920 4034 253932
rect 5074 253920 5080 253932
rect 5132 253920 5138 253972
rect 422938 253920 422944 253972
rect 422996 253960 423002 253972
rect 431218 253960 431224 253972
rect 422996 253932 431224 253960
rect 422996 253920 423002 253932
rect 431218 253920 431224 253932
rect 431276 253920 431282 253972
rect 361758 249704 361764 249756
rect 361816 249744 361822 249756
rect 399478 249744 399484 249756
rect 361816 249716 399484 249744
rect 361816 249704 361822 249716
rect 399478 249704 399484 249716
rect 399536 249704 399542 249756
rect 449434 249024 449440 249076
rect 449492 249064 449498 249076
rect 457806 249064 457812 249076
rect 449492 249036 457812 249064
rect 449492 249024 449498 249036
rect 457806 249024 457812 249036
rect 457864 249024 457870 249076
rect 435634 245624 435640 245676
rect 435692 245664 435698 245676
rect 439682 245664 439688 245676
rect 435692 245636 439688 245664
rect 435692 245624 435698 245636
rect 439682 245624 439688 245636
rect 439740 245624 439746 245676
rect 574830 245556 574836 245608
rect 574888 245596 574894 245608
rect 580166 245596 580172 245608
rect 574888 245568 580172 245596
rect 574888 245556 574894 245568
rect 580166 245556 580172 245568
rect 580224 245556 580230 245608
rect 420178 245284 420184 245336
rect 420236 245324 420242 245336
rect 422938 245324 422944 245336
rect 420236 245296 422944 245324
rect 420236 245284 420242 245296
rect 422938 245284 422944 245296
rect 422996 245284 423002 245336
rect 400214 244876 400220 244928
rect 400272 244916 400278 244928
rect 406838 244916 406844 244928
rect 400272 244888 406844 244916
rect 400272 244876 400278 244888
rect 406838 244876 406844 244888
rect 406896 244876 406902 244928
rect 3786 243924 3792 243976
rect 3844 243964 3850 243976
rect 4982 243964 4988 243976
rect 3844 243936 4988 243964
rect 3844 243924 3850 243936
rect 4982 243924 4988 243936
rect 5040 243924 5046 243976
rect 388438 242156 388444 242208
rect 388496 242196 388502 242208
rect 400214 242196 400220 242208
rect 388496 242168 400220 242196
rect 388496 242156 388502 242168
rect 400214 242156 400220 242168
rect 400272 242156 400278 242208
rect 382918 239436 382924 239488
rect 382976 239476 382982 239488
rect 388438 239476 388444 239488
rect 382976 239448 388444 239476
rect 382976 239436 382982 239448
rect 388438 239436 388444 239448
rect 388496 239436 388502 239488
rect 369118 239368 369124 239420
rect 369176 239408 369182 239420
rect 396810 239408 396816 239420
rect 369176 239380 396816 239408
rect 369176 239368 369182 239380
rect 396810 239368 396816 239380
rect 396868 239368 396874 239420
rect 427078 239368 427084 239420
rect 427136 239408 427142 239420
rect 435634 239408 435640 239420
rect 427136 239380 435640 239408
rect 427136 239368 427142 239380
rect 435634 239368 435640 239380
rect 435692 239368 435698 239420
rect 361758 238688 361764 238740
rect 361816 238728 361822 238740
rect 443730 238728 443736 238740
rect 361816 238700 443736 238728
rect 361816 238688 361822 238700
rect 443730 238688 443736 238700
rect 443788 238688 443794 238740
rect 411898 235220 411904 235272
rect 411956 235260 411962 235272
rect 420178 235260 420184 235272
rect 411956 235232 420184 235260
rect 411956 235220 411962 235232
rect 420178 235220 420184 235232
rect 420236 235220 420242 235272
rect 455966 234948 455972 235000
rect 456024 234988 456030 235000
rect 457990 234988 457996 235000
rect 456024 234960 457996 234988
rect 456024 234948 456030 234960
rect 457990 234948 457996 234960
rect 458048 234948 458054 235000
rect 559650 233180 559656 233232
rect 559708 233220 559714 233232
rect 580166 233220 580172 233232
rect 559708 233192 580172 233220
rect 559708 233180 559714 233192
rect 580166 233180 580172 233192
rect 580224 233180 580230 233232
rect 442258 232908 442264 232960
rect 442316 232948 442322 232960
rect 445018 232948 445024 232960
rect 442316 232920 445024 232948
rect 442316 232908 442322 232920
rect 445018 232908 445024 232920
rect 445076 232908 445082 232960
rect 362310 229712 362316 229764
rect 362368 229752 362374 229764
rect 369118 229752 369124 229764
rect 362368 229724 369124 229752
rect 362368 229712 362374 229724
rect 369118 229712 369124 229724
rect 369176 229712 369182 229764
rect 361758 227672 361764 227724
rect 361816 227712 361822 227724
rect 443638 227712 443644 227724
rect 361816 227684 443644 227712
rect 361816 227672 361822 227684
rect 443638 227672 443644 227684
rect 443696 227672 443702 227724
rect 399478 225564 399484 225616
rect 399536 225604 399542 225616
rect 411898 225604 411904 225616
rect 399536 225576 411904 225604
rect 399536 225564 399542 225576
rect 411898 225564 411904 225576
rect 411956 225564 411962 225616
rect 439682 223524 439688 223576
rect 439740 223564 439746 223576
rect 442258 223564 442264 223576
rect 439740 223536 442264 223564
rect 439740 223524 439746 223536
rect 442258 223524 442264 223536
rect 442316 223524 442322 223576
rect 3878 222096 3884 222148
rect 3936 222136 3942 222148
rect 5166 222136 5172 222148
rect 3936 222108 5172 222136
rect 3936 222096 3942 222108
rect 5166 222096 5172 222108
rect 5224 222096 5230 222148
rect 450354 221416 450360 221468
rect 450412 221456 450418 221468
rect 457990 221456 457996 221468
rect 450412 221428 457996 221456
rect 450412 221416 450418 221428
rect 457990 221416 457996 221428
rect 458048 221416 458054 221468
rect 361206 220056 361212 220108
rect 361264 220096 361270 220108
rect 382918 220096 382924 220108
rect 361264 220068 382924 220096
rect 361264 220056 361270 220068
rect 382918 220056 382924 220068
rect 382976 220056 382982 220108
rect 436094 218016 436100 218068
rect 436152 218056 436158 218068
rect 439682 218056 439688 218068
rect 436152 218028 439688 218056
rect 436152 218016 436158 218028
rect 439682 218016 439688 218028
rect 439740 218016 439746 218068
rect 361574 216316 361580 216368
rect 361632 216356 361638 216368
rect 363782 216356 363788 216368
rect 361632 216328 363788 216356
rect 361632 216316 361638 216328
rect 363782 216316 363788 216328
rect 363840 216316 363846 216368
rect 413094 214548 413100 214600
rect 413152 214588 413158 214600
rect 436094 214588 436100 214600
rect 413152 214560 436100 214588
rect 413152 214548 413158 214560
rect 436094 214548 436100 214560
rect 436152 214548 436158 214600
rect 396258 213936 396264 213988
rect 396316 213976 396322 213988
rect 399478 213976 399484 213988
rect 396316 213948 399484 213976
rect 396316 213936 396322 213948
rect 399478 213936 399484 213948
rect 399536 213936 399542 213988
rect 377398 211760 377404 211812
rect 377456 211800 377462 211812
rect 396258 211800 396264 211812
rect 377456 211772 396264 211800
rect 377456 211760 377462 211772
rect 396258 211760 396264 211772
rect 396316 211760 396322 211812
rect 407850 210128 407856 210180
rect 407908 210168 407914 210180
rect 413094 210168 413100 210180
rect 407908 210140 413100 210168
rect 407908 210128 407914 210140
rect 413094 210128 413100 210140
rect 413152 210128 413158 210180
rect 411898 209040 411904 209092
rect 411956 209080 411962 209092
rect 427078 209080 427084 209092
rect 411956 209052 427084 209080
rect 411956 209040 411962 209052
rect 427078 209040 427084 209052
rect 427136 209040 427142 209092
rect 399478 207612 399484 207664
rect 399536 207652 399542 207664
rect 407850 207652 407856 207664
rect 399536 207624 407856 207652
rect 399536 207612 399542 207624
rect 407850 207612 407856 207624
rect 407908 207612 407914 207664
rect 576118 206932 576124 206984
rect 576176 206972 576182 206984
rect 579798 206972 579804 206984
rect 576176 206944 579804 206972
rect 576176 206932 576182 206944
rect 579798 206932 579804 206944
rect 579856 206932 579862 206984
rect 361758 205572 361764 205624
rect 361816 205612 361822 205624
rect 439590 205612 439596 205624
rect 361816 205584 439596 205612
rect 361816 205572 361822 205584
rect 439590 205572 439596 205584
rect 439648 205572 439654 205624
rect 408494 198704 408500 198756
rect 408552 198744 408558 198756
rect 411898 198744 411904 198756
rect 408552 198716 411904 198744
rect 408552 198704 408558 198716
rect 411898 198704 411904 198716
rect 411956 198704 411962 198756
rect 447318 197956 447324 198008
rect 447376 197996 447382 198008
rect 475378 197996 475384 198008
rect 447376 197968 475384 197996
rect 447376 197956 447382 197968
rect 475378 197956 475384 197968
rect 475436 197956 475442 198008
rect 374638 195100 374644 195152
rect 374696 195140 374702 195152
rect 377398 195140 377404 195152
rect 374696 195112 377404 195140
rect 374696 195100 374702 195112
rect 377398 195100 377404 195112
rect 377456 195100 377462 195152
rect 361666 194488 361672 194540
rect 361724 194528 361730 194540
rect 436738 194528 436744 194540
rect 361724 194500 436744 194528
rect 361724 194488 361730 194500
rect 436738 194488 436744 194500
rect 436796 194488 436802 194540
rect 393958 194420 393964 194472
rect 394016 194460 394022 194472
rect 399478 194460 399484 194472
rect 394016 194432 399484 194460
rect 394016 194420 394022 194432
rect 399478 194420 399484 194432
rect 399536 194420 399542 194472
rect 547138 193128 547144 193180
rect 547196 193168 547202 193180
rect 580166 193168 580172 193180
rect 547196 193140 580172 193168
rect 547196 193128 547202 193140
rect 580166 193128 580172 193140
rect 580224 193128 580230 193180
rect 401594 191088 401600 191140
rect 401652 191128 401658 191140
rect 408494 191128 408500 191140
rect 401652 191100 408500 191128
rect 401652 191088 401658 191100
rect 408494 191088 408500 191100
rect 408552 191088 408558 191140
rect 398466 186328 398472 186380
rect 398524 186368 398530 186380
rect 401594 186368 401600 186380
rect 398524 186340 401600 186368
rect 398524 186328 398530 186340
rect 401594 186328 401600 186340
rect 401652 186328 401658 186380
rect 390646 186260 390652 186312
rect 390704 186300 390710 186312
rect 393958 186300 393964 186312
rect 390704 186272 393964 186300
rect 390704 186260 390710 186272
rect 393958 186260 393964 186272
rect 394016 186260 394022 186312
rect 361666 183472 361672 183524
rect 361724 183512 361730 183524
rect 447594 183512 447600 183524
rect 361724 183484 447600 183512
rect 361724 183472 361730 183484
rect 447594 183472 447600 183484
rect 447652 183512 447658 183524
rect 448054 183512 448060 183524
rect 447652 183484 448060 183512
rect 447652 183472 447658 183484
rect 448054 183472 448060 183484
rect 448112 183472 448118 183524
rect 447594 182792 447600 182844
rect 447652 182832 447658 182844
rect 528554 182832 528560 182844
rect 447652 182804 528560 182832
rect 447652 182792 447658 182804
rect 528554 182792 528560 182804
rect 528612 182792 528618 182844
rect 388438 181568 388444 181620
rect 388496 181608 388502 181620
rect 390646 181608 390652 181620
rect 388496 181580 390652 181608
rect 388496 181568 388502 181580
rect 390646 181568 390652 181580
rect 390704 181568 390710 181620
rect 362954 180072 362960 180124
rect 363012 180112 363018 180124
rect 374638 180112 374644 180124
rect 363012 180084 374644 180112
rect 363012 180072 363018 180084
rect 374638 180072 374644 180084
rect 374696 180072 374702 180124
rect 559558 179324 559564 179376
rect 559616 179364 559622 179376
rect 580166 179364 580172 179376
rect 559616 179336 580172 179364
rect 559616 179324 559622 179336
rect 580166 179324 580172 179336
rect 580224 179324 580230 179376
rect 361298 174632 361304 174684
rect 361356 174672 361362 174684
rect 362954 174672 362960 174684
rect 361356 174644 362960 174672
rect 361356 174632 361362 174644
rect 362954 174632 362960 174644
rect 363012 174632 363018 174684
rect 361666 172456 361672 172508
rect 361724 172496 361730 172508
rect 447594 172496 447600 172508
rect 361724 172468 447600 172496
rect 361724 172456 361730 172468
rect 447594 172456 447600 172468
rect 447652 172496 447658 172508
rect 448238 172496 448244 172508
rect 447652 172468 448244 172496
rect 447652 172456 447658 172468
rect 448238 172456 448244 172468
rect 448296 172456 448302 172508
rect 447594 171776 447600 171828
rect 447652 171816 447658 171828
rect 524414 171816 524420 171828
rect 447652 171788 524420 171816
rect 447652 171776 447658 171788
rect 524414 171776 524420 171788
rect 524472 171776 524478 171828
rect 386046 168376 386052 168428
rect 386104 168416 386110 168428
rect 388438 168416 388444 168428
rect 386104 168388 388444 168416
rect 386104 168376 386110 168388
rect 388438 168376 388444 168388
rect 388496 168376 388502 168428
rect 533430 166948 533436 167000
rect 533488 166988 533494 167000
rect 580166 166988 580172 167000
rect 533488 166960 580172 166988
rect 533488 166948 533494 166960
rect 580166 166948 580172 166960
rect 580224 166948 580230 167000
rect 438578 163616 438584 163668
rect 438636 163656 438642 163668
rect 439498 163656 439504 163668
rect 438636 163628 439504 163656
rect 438636 163616 438642 163628
rect 439498 163616 439504 163628
rect 439556 163616 439562 163668
rect 378686 162868 378692 162920
rect 378744 162908 378750 162920
rect 386046 162908 386052 162920
rect 378744 162880 386052 162908
rect 378744 162868 378750 162880
rect 386046 162868 386052 162880
rect 386104 162868 386110 162920
rect 418706 162324 418712 162376
rect 418764 162364 418770 162376
rect 457898 162364 457904 162376
rect 418764 162336 457904 162364
rect 418764 162324 418770 162336
rect 457898 162324 457904 162336
rect 457956 162364 457962 162376
rect 489914 162364 489920 162376
rect 457956 162336 489920 162364
rect 457956 162324 457962 162336
rect 489914 162324 489920 162336
rect 489972 162324 489978 162376
rect 414750 162256 414756 162308
rect 414808 162296 414814 162308
rect 457990 162296 457996 162308
rect 414808 162268 457996 162296
rect 414808 162256 414814 162268
rect 457990 162256 457996 162268
rect 458048 162296 458054 162308
rect 485774 162296 485780 162308
rect 458048 162268 485780 162296
rect 458048 162256 458054 162268
rect 485774 162256 485780 162268
rect 485832 162256 485838 162308
rect 411622 162188 411628 162240
rect 411680 162228 411686 162240
rect 458082 162228 458088 162240
rect 411680 162200 458088 162228
rect 411680 162188 411686 162200
rect 458082 162188 458088 162200
rect 458140 162228 458146 162240
rect 481634 162228 481640 162240
rect 458140 162200 481640 162228
rect 458140 162188 458146 162200
rect 481634 162188 481640 162200
rect 481692 162188 481698 162240
rect 445202 162120 445208 162172
rect 445260 162160 445266 162172
rect 457806 162160 457812 162172
rect 445260 162132 457812 162160
rect 445260 162120 445266 162132
rect 457806 162120 457812 162132
rect 457864 162160 457870 162172
rect 533430 162160 533436 162172
rect 457864 162132 533436 162160
rect 457864 162120 457870 162132
rect 533430 162120 533436 162132
rect 533488 162120 533494 162172
rect 406838 161440 406844 161492
rect 406896 161480 406902 161492
rect 414750 161480 414756 161492
rect 406896 161452 414756 161480
rect 406896 161440 406902 161452
rect 414750 161440 414756 161452
rect 414808 161440 414814 161492
rect 361758 161372 361764 161424
rect 361816 161412 361822 161424
rect 448330 161412 448336 161424
rect 361816 161384 448336 161412
rect 361816 161372 361822 161384
rect 448330 161372 448336 161384
rect 448388 161372 448394 161424
rect 448330 160692 448336 160744
rect 448388 160732 448394 160744
rect 521654 160732 521660 160744
rect 448388 160704 521660 160732
rect 448388 160692 448394 160704
rect 521654 160692 521660 160704
rect 521712 160692 521718 160744
rect 425330 160488 425336 160540
rect 425388 160528 425394 160540
rect 426342 160528 426348 160540
rect 425388 160500 426348 160528
rect 425388 160488 425394 160500
rect 426342 160488 426348 160500
rect 426400 160528 426406 160540
rect 496814 160528 496820 160540
rect 426400 160500 496820 160528
rect 426400 160488 426406 160500
rect 496814 160488 496820 160500
rect 496872 160488 496878 160540
rect 428642 160420 428648 160472
rect 428700 160460 428706 160472
rect 500954 160460 500960 160472
rect 428700 160432 500960 160460
rect 428700 160420 428706 160432
rect 500954 160420 500960 160432
rect 501012 160420 501018 160472
rect 422018 160352 422024 160404
rect 422076 160392 422082 160404
rect 494054 160392 494060 160404
rect 422076 160364 494060 160392
rect 422076 160352 422082 160364
rect 494054 160352 494060 160364
rect 494112 160352 494118 160404
rect 431770 160284 431776 160336
rect 431828 160324 431834 160336
rect 505094 160324 505100 160336
rect 431828 160296 505100 160324
rect 431828 160284 431834 160296
rect 505094 160284 505100 160296
rect 505152 160284 505158 160336
rect 404078 160216 404084 160268
rect 404136 160256 404142 160268
rect 418154 160256 418160 160268
rect 404136 160228 418160 160256
rect 404136 160216 404142 160228
rect 418154 160216 418160 160228
rect 418212 160216 418218 160268
rect 435266 160216 435272 160268
rect 435324 160256 435330 160268
rect 436002 160256 436008 160268
rect 435324 160228 436008 160256
rect 435324 160216 435330 160228
rect 436002 160216 436008 160228
rect 436060 160256 436066 160268
rect 509234 160256 509240 160268
rect 436060 160228 509240 160256
rect 436060 160216 436066 160228
rect 509234 160216 509240 160228
rect 509292 160216 509298 160268
rect 407850 160148 407856 160200
rect 407908 160188 407914 160200
rect 411438 160188 411444 160200
rect 407908 160160 411444 160188
rect 407908 160148 407914 160160
rect 411438 160148 411444 160160
rect 411496 160148 411502 160200
rect 438578 160148 438584 160200
rect 438636 160188 438642 160200
rect 513374 160188 513380 160200
rect 438636 160160 513380 160188
rect 438636 160148 438642 160160
rect 513374 160148 513380 160160
rect 513432 160148 513438 160200
rect 409690 160080 409696 160132
rect 409748 160120 409754 160132
rect 441568 160120 441574 160132
rect 409748 160092 441574 160120
rect 409748 160080 409754 160092
rect 441568 160080 441574 160092
rect 441626 160120 441632 160132
rect 442902 160120 442908 160132
rect 441626 160092 442908 160120
rect 441626 160080 441632 160092
rect 442902 160080 442908 160092
rect 442960 160120 442966 160132
rect 517514 160120 517520 160132
rect 442960 160092 517520 160120
rect 442960 160080 442966 160092
rect 517514 160080 517520 160092
rect 517572 160080 517578 160132
rect 409138 159672 409144 159724
rect 409196 159712 409202 159724
rect 421374 159712 421380 159724
rect 409196 159684 421380 159712
rect 409196 159672 409202 159684
rect 421374 159672 421380 159684
rect 421432 159672 421438 159724
rect 409230 159604 409236 159656
rect 409288 159644 409294 159656
rect 425146 159644 425152 159656
rect 409288 159616 425152 159644
rect 409288 159604 409294 159616
rect 425146 159604 425152 159616
rect 425204 159604 425210 159656
rect 409322 159536 409328 159588
rect 409380 159576 409386 159588
rect 427998 159576 428004 159588
rect 409380 159548 428004 159576
rect 409380 159536 409386 159548
rect 427998 159536 428004 159548
rect 428056 159536 428062 159588
rect 409414 159468 409420 159520
rect 409472 159508 409478 159520
rect 431310 159508 431316 159520
rect 409472 159480 431316 159508
rect 409472 159468 409478 159480
rect 431310 159468 431316 159480
rect 431368 159468 431374 159520
rect 409506 159400 409512 159452
rect 409564 159440 409570 159452
rect 434806 159440 434812 159452
rect 409564 159412 434812 159440
rect 409564 159400 409570 159412
rect 434806 159400 434812 159412
rect 434864 159400 434870 159452
rect 409598 159332 409604 159384
rect 409656 159372 409662 159384
rect 437934 159372 437940 159384
rect 409656 159344 437940 159372
rect 409656 159332 409662 159344
rect 437934 159332 437940 159344
rect 437992 159332 437998 159384
rect 452562 158244 452568 158296
rect 452620 158284 452626 158296
rect 456702 158284 456708 158296
rect 452620 158256 456708 158284
rect 452620 158244 452626 158256
rect 456702 158244 456708 158256
rect 456760 158244 456766 158296
rect 373626 156612 373632 156664
rect 373684 156652 373690 156664
rect 378686 156652 378692 156664
rect 373684 156624 378692 156652
rect 373684 156612 373690 156624
rect 378686 156612 378692 156624
rect 378744 156612 378750 156664
rect 452562 155660 452568 155712
rect 452620 155700 452626 155712
rect 456518 155700 456524 155712
rect 452620 155672 456524 155700
rect 452620 155660 452626 155672
rect 456518 155660 456524 155672
rect 456576 155660 456582 155712
rect 551278 153144 551284 153196
rect 551336 153184 551342 153196
rect 580166 153184 580172 153196
rect 551336 153156 580172 153184
rect 551336 153144 551342 153156
rect 580166 153144 580172 153156
rect 580224 153144 580230 153196
rect 361758 150356 361764 150408
rect 361816 150396 361822 150408
rect 409690 150396 409696 150408
rect 361816 150368 409696 150396
rect 361816 150356 361822 150368
rect 409690 150356 409696 150368
rect 409748 150356 409754 150408
rect 451550 150220 451556 150272
rect 451608 150260 451614 150272
rect 455230 150260 455236 150272
rect 451608 150232 455236 150260
rect 451608 150220 451614 150232
rect 455230 150220 455236 150232
rect 455288 150220 455294 150272
rect 371234 149676 371240 149728
rect 371292 149716 371298 149728
rect 398466 149716 398472 149728
rect 371292 149688 398472 149716
rect 371292 149676 371298 149688
rect 398466 149676 398472 149688
rect 398524 149676 398530 149728
rect 451734 148996 451740 149048
rect 451792 149036 451798 149048
rect 454862 149036 454868 149048
rect 451792 149008 454868 149036
rect 451792 148996 451798 149008
rect 454862 148996 454868 149008
rect 454920 148996 454926 149048
rect 451734 147364 451740 147416
rect 451792 147404 451798 147416
rect 458634 147404 458640 147416
rect 451792 147376 458640 147404
rect 451792 147364 451798 147376
rect 458634 147364 458640 147376
rect 458692 147364 458698 147416
rect 452562 146140 452568 146192
rect 452620 146180 452626 146192
rect 459370 146180 459376 146192
rect 452620 146152 459376 146180
rect 452620 146140 452626 146152
rect 459370 146140 459376 146152
rect 459428 146140 459434 146192
rect 452562 144644 452568 144696
rect 452620 144684 452626 144696
rect 455046 144684 455052 144696
rect 452620 144656 455052 144684
rect 452620 144644 452626 144656
rect 455046 144644 455052 144656
rect 455104 144644 455110 144696
rect 364242 144168 364248 144220
rect 364300 144208 364306 144220
rect 371234 144208 371240 144220
rect 364300 144180 371240 144208
rect 364300 144168 364306 144180
rect 371234 144168 371240 144180
rect 371292 144168 371298 144220
rect 368382 143828 368388 143880
rect 368440 143868 368446 143880
rect 373626 143868 373632 143880
rect 368440 143840 373632 143868
rect 368440 143828 368446 143840
rect 373626 143828 373632 143840
rect 373684 143828 373690 143880
rect 533430 143488 533436 143540
rect 533488 143528 533494 143540
rect 533982 143528 533988 143540
rect 533488 143500 533988 143528
rect 533488 143488 533494 143500
rect 533982 143488 533988 143500
rect 534040 143488 534046 143540
rect 536098 143488 536104 143540
rect 536156 143528 536162 143540
rect 537294 143528 537300 143540
rect 536156 143500 537300 143528
rect 536156 143488 536162 143500
rect 537294 143488 537300 143500
rect 537352 143488 537358 143540
rect 452562 143284 452568 143336
rect 452620 143324 452626 143336
rect 457622 143324 457628 143336
rect 452620 143296 457628 143324
rect 452620 143284 452626 143296
rect 457622 143284 457628 143296
rect 457680 143284 457686 143336
rect 533982 142196 533988 142248
rect 534040 142236 534046 142248
rect 540330 142236 540336 142248
rect 534040 142208 540336 142236
rect 534040 142196 534046 142208
rect 540330 142196 540336 142208
rect 540388 142196 540394 142248
rect 452562 141924 452568 141976
rect 452620 141964 452626 141976
rect 455138 141964 455144 141976
rect 452620 141936 455144 141964
rect 452620 141924 452626 141936
rect 455138 141924 455144 141936
rect 455196 141924 455202 141976
rect 365438 140768 365444 140820
rect 365496 140808 365502 140820
rect 368382 140808 368388 140820
rect 365496 140780 368388 140808
rect 365496 140768 365502 140780
rect 368382 140768 368388 140780
rect 368440 140768 368446 140820
rect 452562 140632 452568 140684
rect 452620 140672 452626 140684
rect 459278 140672 459284 140684
rect 452620 140644 459284 140672
rect 452620 140632 452626 140644
rect 459278 140632 459284 140644
rect 459336 140632 459342 140684
rect 534718 140156 534724 140208
rect 534776 140196 534782 140208
rect 542906 140196 542912 140208
rect 534776 140168 542912 140196
rect 534776 140156 534782 140168
rect 542906 140156 542912 140168
rect 542964 140156 542970 140208
rect 533338 140088 533344 140140
rect 533396 140128 533402 140140
rect 542722 140128 542728 140140
rect 533396 140100 542728 140128
rect 533396 140088 533402 140100
rect 542722 140088 542728 140100
rect 542780 140088 542786 140140
rect 530578 140020 530584 140072
rect 530636 140060 530642 140072
rect 543090 140060 543096 140072
rect 530636 140032 543096 140060
rect 530636 140020 530642 140032
rect 543090 140020 543096 140032
rect 543148 140020 543154 140072
rect 361758 139340 361764 139392
rect 361816 139380 361822 139392
rect 409598 139380 409604 139392
rect 361816 139352 409604 139380
rect 361816 139340 361822 139352
rect 409598 139340 409604 139352
rect 409656 139340 409662 139392
rect 451550 139340 451556 139392
rect 451608 139380 451614 139392
rect 457530 139380 457536 139392
rect 451608 139352 457536 139380
rect 451608 139340 451614 139352
rect 457530 139340 457536 139352
rect 457588 139340 457594 139392
rect 555418 139340 555424 139392
rect 555476 139380 555482 139392
rect 580166 139380 580172 139392
rect 555476 139352 580172 139380
rect 555476 139340 555482 139352
rect 580166 139340 580172 139352
rect 580224 139340 580230 139392
rect 538858 138524 538864 138576
rect 538916 138564 538922 138576
rect 542998 138564 543004 138576
rect 538916 138536 543004 138564
rect 538916 138524 538922 138536
rect 542998 138524 543004 138536
rect 543056 138524 543062 138576
rect 361390 137980 361396 138032
rect 361448 138020 361454 138032
rect 364242 138020 364248 138032
rect 361448 137992 364248 138020
rect 361448 137980 361454 137992
rect 364242 137980 364248 137992
rect 364300 137980 364306 138032
rect 452562 137844 452568 137896
rect 452620 137884 452626 137896
rect 454954 137884 454960 137896
rect 452620 137856 454960 137884
rect 452620 137844 452626 137856
rect 454954 137844 454960 137856
rect 455012 137844 455018 137896
rect 452562 136484 452568 136536
rect 452620 136524 452626 136536
rect 459094 136524 459100 136536
rect 452620 136496 459100 136524
rect 452620 136484 452626 136496
rect 459094 136484 459100 136496
rect 459152 136484 459158 136536
rect 452562 135124 452568 135176
rect 452620 135164 452626 135176
rect 454770 135164 454776 135176
rect 452620 135136 454776 135164
rect 452620 135124 452626 135136
rect 454770 135124 454776 135136
rect 454828 135124 454834 135176
rect 452562 133764 452568 133816
rect 452620 133804 452626 133816
rect 456610 133804 456616 133816
rect 452620 133776 456616 133804
rect 452620 133764 452626 133776
rect 456610 133764 456616 133776
rect 456668 133764 456674 133816
rect 452470 132404 452476 132456
rect 452528 132444 452534 132456
rect 453758 132444 453764 132456
rect 452528 132416 453764 132444
rect 452528 132404 452534 132416
rect 453758 132404 453764 132416
rect 453816 132404 453822 132456
rect 452562 131044 452568 131096
rect 452620 131084 452626 131096
rect 453942 131084 453948 131096
rect 452620 131056 453948 131084
rect 452620 131044 452626 131056
rect 453942 131044 453948 131056
rect 454000 131044 454006 131096
rect 361482 130160 361488 130212
rect 361540 130200 361546 130212
rect 365438 130200 365444 130212
rect 361540 130172 365444 130200
rect 361540 130160 361546 130172
rect 365438 130160 365444 130172
rect 365496 130160 365502 130212
rect 361574 128256 361580 128308
rect 361632 128296 361638 128308
rect 409506 128296 409512 128308
rect 361632 128268 409512 128296
rect 361632 128256 361638 128268
rect 409506 128256 409512 128268
rect 409564 128256 409570 128308
rect 452562 126896 452568 126948
rect 452620 126936 452626 126948
rect 457438 126936 457444 126948
rect 452620 126908 457444 126936
rect 452620 126896 452626 126908
rect 457438 126896 457444 126908
rect 457496 126896 457502 126948
rect 573358 126896 573364 126948
rect 573416 126936 573422 126948
rect 580166 126936 580172 126948
rect 573416 126908 580172 126936
rect 573416 126896 573422 126908
rect 580166 126896 580172 126908
rect 580224 126896 580230 126948
rect 451918 126012 451924 126064
rect 451976 126052 451982 126064
rect 453666 126052 453672 126064
rect 451976 126024 453672 126052
rect 451976 126012 451982 126024
rect 453666 126012 453672 126024
rect 453724 126012 453730 126064
rect 451918 124720 451924 124772
rect 451976 124760 451982 124772
rect 453850 124760 453856 124772
rect 451976 124732 453856 124760
rect 451976 124720 451982 124732
rect 453850 124720 453856 124732
rect 453908 124720 453914 124772
rect 451918 123224 451924 123276
rect 451976 123264 451982 123276
rect 459462 123264 459468 123276
rect 451976 123236 459468 123264
rect 451976 123224 451982 123236
rect 459462 123224 459468 123236
rect 459520 123224 459526 123276
rect 451734 122204 451740 122256
rect 451792 122244 451798 122256
rect 458726 122244 458732 122256
rect 451792 122216 458732 122244
rect 451792 122204 451798 122216
rect 458726 122204 458732 122216
rect 458784 122204 458790 122256
rect 361574 117240 361580 117292
rect 361632 117280 361638 117292
rect 409414 117280 409420 117292
rect 361632 117252 409420 117280
rect 361632 117240 361638 117252
rect 409414 117240 409420 117252
rect 409472 117240 409478 117292
rect 570598 113092 570604 113144
rect 570656 113132 570662 113144
rect 579798 113132 579804 113144
rect 570656 113104 579804 113132
rect 570656 113092 570662 113104
rect 579798 113092 579804 113104
rect 579856 113092 579862 113144
rect 361574 106224 361580 106276
rect 361632 106264 361638 106276
rect 409322 106264 409328 106276
rect 361632 106236 409328 106264
rect 361632 106224 361638 106236
rect 409322 106224 409328 106236
rect 409380 106224 409386 106276
rect 558178 100648 558184 100700
rect 558236 100688 558242 100700
rect 580166 100688 580172 100700
rect 558236 100660 580172 100688
rect 558236 100648 558242 100660
rect 580166 100648 580172 100660
rect 580224 100648 580230 100700
rect 3694 98608 3700 98660
rect 3752 98648 3758 98660
rect 20898 98648 20904 98660
rect 3752 98620 20904 98648
rect 3752 98608 3758 98620
rect 20898 98608 20904 98620
rect 20956 98608 20962 98660
rect 361758 95140 361764 95192
rect 361816 95180 361822 95192
rect 409230 95180 409236 95192
rect 361816 95152 409236 95180
rect 361816 95140 361822 95152
rect 409230 95140 409236 95152
rect 409288 95140 409294 95192
rect 571978 86912 571984 86964
rect 572036 86952 572042 86964
rect 580166 86952 580172 86964
rect 572036 86924 580172 86952
rect 572036 86912 572042 86924
rect 580166 86912 580172 86924
rect 580224 86912 580230 86964
rect 3602 86232 3608 86284
rect 3660 86272 3666 86284
rect 20898 86272 20904 86284
rect 3660 86244 20904 86272
rect 3660 86232 3666 86244
rect 20898 86232 20904 86244
rect 20956 86232 20962 86284
rect 361758 84124 361764 84176
rect 361816 84164 361822 84176
rect 409138 84164 409144 84176
rect 361816 84136 409144 84164
rect 361816 84124 361822 84136
rect 409138 84124 409144 84136
rect 409196 84124 409202 84176
rect 361758 73108 361764 73160
rect 361816 73148 361822 73160
rect 404078 73148 404084 73160
rect 361816 73120 404084 73148
rect 361816 73108 361822 73120
rect 404078 73108 404084 73120
rect 404136 73108 404142 73160
rect 544378 73108 544384 73160
rect 544436 73148 544442 73160
rect 580166 73148 580172 73160
rect 544436 73120 580172 73148
rect 544436 73108 544442 73120
rect 580166 73108 580172 73120
rect 580224 73108 580230 73160
rect 5074 70388 5080 70440
rect 5132 70428 5138 70440
rect 5132 70400 6914 70428
rect 5132 70388 5138 70400
rect 6886 70360 6914 70400
rect 7558 70360 7564 70372
rect 6886 70332 7564 70360
rect 7558 70320 7564 70332
rect 7616 70320 7622 70372
rect 361758 62024 361764 62076
rect 361816 62064 361822 62076
rect 406838 62064 406844 62076
rect 361816 62036 406844 62064
rect 361816 62024 361822 62036
rect 406838 62024 406844 62036
rect 406896 62024 406902 62076
rect 7558 60732 7564 60784
rect 7616 60772 7622 60784
rect 7616 60744 8340 60772
rect 7616 60732 7622 60744
rect 8312 60704 8340 60744
rect 10042 60704 10048 60716
rect 8312 60676 10048 60704
rect 10042 60664 10048 60676
rect 10100 60664 10106 60716
rect 548518 60664 548524 60716
rect 548576 60704 548582 60716
rect 580166 60704 580172 60716
rect 548576 60676 580172 60704
rect 548576 60664 548582 60676
rect 580166 60664 580172 60676
rect 580224 60664 580230 60716
rect 3510 59984 3516 60036
rect 3568 60024 3574 60036
rect 20898 60024 20904 60036
rect 3568 59996 20904 60024
rect 3568 59984 3574 59996
rect 20898 59984 20904 59996
rect 20956 59984 20962 60036
rect 4798 59304 4804 59356
rect 4856 59344 4862 59356
rect 5810 59344 5816 59356
rect 4856 59316 5816 59344
rect 4856 59304 4862 59316
rect 5810 59304 5816 59316
rect 5868 59304 5874 59356
rect 5810 57196 5816 57248
rect 5868 57236 5874 57248
rect 9766 57236 9772 57248
rect 5868 57208 9772 57236
rect 5868 57196 5874 57208
rect 9766 57196 9772 57208
rect 9824 57196 9830 57248
rect 4890 56516 4896 56568
rect 4948 56556 4954 56568
rect 7282 56556 7288 56568
rect 4948 56528 7288 56556
rect 4948 56516 4954 56528
rect 7282 56516 7288 56528
rect 7340 56516 7346 56568
rect 10042 56516 10048 56568
rect 10100 56556 10106 56568
rect 12342 56556 12348 56568
rect 10100 56528 12348 56556
rect 10100 56516 10106 56528
rect 12342 56516 12348 56528
rect 12400 56516 12406 56568
rect 9766 56176 9772 56228
rect 9824 56216 9830 56228
rect 12618 56216 12624 56228
rect 9824 56188 12624 56216
rect 9824 56176 9830 56188
rect 12618 56176 12624 56188
rect 12676 56176 12682 56228
rect 7282 54612 7288 54664
rect 7340 54652 7346 54664
rect 11974 54652 11980 54664
rect 7340 54624 11980 54652
rect 7340 54612 7346 54624
rect 11974 54612 11980 54624
rect 12032 54612 12038 54664
rect 5534 54476 5540 54528
rect 5592 54516 5598 54528
rect 13814 54516 13820 54528
rect 5592 54488 13820 54516
rect 5592 54476 5598 54488
rect 13814 54476 13820 54488
rect 13872 54476 13878 54528
rect 13814 53116 13820 53168
rect 13872 53156 13878 53168
rect 17862 53156 17868 53168
rect 13872 53128 17868 53156
rect 13872 53116 13878 53128
rect 17862 53116 17868 53128
rect 17920 53116 17926 53168
rect 12342 52980 12348 53032
rect 12400 53020 12406 53032
rect 15194 53020 15200 53032
rect 12400 52992 15200 53020
rect 12400 52980 12406 52992
rect 15194 52980 15200 52992
rect 15252 52980 15258 53032
rect 11974 52436 11980 52488
rect 12032 52476 12038 52488
rect 12032 52448 13860 52476
rect 12032 52436 12038 52448
rect 13832 52408 13860 52448
rect 18782 52408 18788 52420
rect 13832 52380 18788 52408
rect 18782 52368 18788 52380
rect 18840 52368 18846 52420
rect 361758 52368 361764 52420
rect 361816 52408 361822 52420
rect 407850 52408 407856 52420
rect 361816 52380 407856 52408
rect 361816 52368 361822 52380
rect 407850 52368 407856 52380
rect 407908 52368 407914 52420
rect 17862 51416 17868 51468
rect 17920 51456 17926 51468
rect 19518 51456 19524 51468
rect 17920 51428 19524 51456
rect 17920 51416 17926 51428
rect 19518 51416 19524 51428
rect 19576 51416 19582 51468
rect 540606 51076 540612 51128
rect 540664 51116 540670 51128
rect 543734 51116 543740 51128
rect 540664 51088 543740 51116
rect 540664 51076 540670 51088
rect 543734 51076 543740 51088
rect 543792 51076 543798 51128
rect 4982 50328 4988 50380
rect 5040 50368 5046 50380
rect 11698 50368 11704 50380
rect 5040 50340 11704 50368
rect 5040 50328 5046 50340
rect 11698 50328 11704 50340
rect 11756 50328 11762 50380
rect 12618 50328 12624 50380
rect 12676 50368 12682 50380
rect 20622 50368 20628 50380
rect 12676 50340 20628 50368
rect 12676 50328 12682 50340
rect 20622 50328 20628 50340
rect 20680 50328 20686 50380
rect 359550 50056 359556 50108
rect 359608 50096 359614 50108
rect 361206 50096 361212 50108
rect 359608 50068 361212 50096
rect 359608 50056 359614 50068
rect 361206 50056 361212 50068
rect 361264 50056 361270 50108
rect 15194 49716 15200 49768
rect 15252 49756 15258 49768
rect 15252 49728 16574 49756
rect 15252 49716 15258 49728
rect 16546 49688 16574 49728
rect 18046 49688 18052 49700
rect 16546 49660 18052 49688
rect 18046 49648 18052 49660
rect 18104 49648 18110 49700
rect 19518 48220 19524 48272
rect 19576 48260 19582 48272
rect 20714 48260 20720 48272
rect 19576 48232 20720 48260
rect 19576 48220 19582 48232
rect 20714 48220 20720 48232
rect 20772 48220 20778 48272
rect 18046 47880 18052 47932
rect 18104 47920 18110 47932
rect 20806 47920 20812 47932
rect 18104 47892 20812 47920
rect 18104 47880 18110 47892
rect 20806 47880 20812 47892
rect 20864 47880 20870 47932
rect 3142 46996 3148 47048
rect 3200 47036 3206 47048
rect 456150 47036 456156 47048
rect 3200 47008 456156 47036
rect 3200 46996 3206 47008
rect 456150 46996 456156 47008
rect 456208 46996 456214 47048
rect 3510 46860 3516 46912
rect 3568 46900 3574 46912
rect 460290 46900 460296 46912
rect 3568 46872 460296 46900
rect 3568 46860 3574 46872
rect 460290 46860 460296 46872
rect 460348 46860 460354 46912
rect 566458 46860 566464 46912
rect 566516 46900 566522 46912
rect 580166 46900 580172 46912
rect 566516 46872 580172 46900
rect 566516 46860 566522 46872
rect 580166 46860 580172 46872
rect 580224 46860 580230 46912
rect 3602 46792 3608 46844
rect 3660 46832 3666 46844
rect 460382 46832 460388 46844
rect 3660 46804 460388 46832
rect 3660 46792 3666 46804
rect 460382 46792 460388 46804
rect 460440 46792 460446 46844
rect 4062 46724 4068 46776
rect 4120 46764 4126 46776
rect 458910 46764 458916 46776
rect 4120 46736 458916 46764
rect 4120 46724 4126 46736
rect 458910 46724 458916 46736
rect 458968 46724 458974 46776
rect 3234 46656 3240 46708
rect 3292 46696 3298 46708
rect 456334 46696 456340 46708
rect 3292 46668 456340 46696
rect 3292 46656 3298 46668
rect 456334 46656 456340 46668
rect 456392 46656 456398 46708
rect 3326 46588 3332 46640
rect 3384 46628 3390 46640
rect 456242 46628 456248 46640
rect 3384 46600 456248 46628
rect 3384 46588 3390 46600
rect 456242 46588 456248 46600
rect 456300 46588 456306 46640
rect 3970 46520 3976 46572
rect 4028 46560 4034 46572
rect 456426 46560 456432 46572
rect 4028 46532 456432 46560
rect 4028 46520 4034 46532
rect 456426 46520 456432 46532
rect 456484 46520 456490 46572
rect 3786 46452 3792 46504
rect 3844 46492 3850 46504
rect 453482 46492 453488 46504
rect 3844 46464 453488 46492
rect 3844 46452 3850 46464
rect 453482 46452 453488 46464
rect 453540 46452 453546 46504
rect 3878 46384 3884 46436
rect 3936 46424 3942 46436
rect 453390 46424 453396 46436
rect 3936 46396 453396 46424
rect 3936 46384 3942 46396
rect 453390 46384 453396 46396
rect 453448 46384 453454 46436
rect 20898 46316 20904 46368
rect 20956 46356 20962 46368
rect 453574 46356 453580 46368
rect 20956 46328 453580 46356
rect 20956 46316 20962 46328
rect 453574 46316 453580 46328
rect 453632 46316 453638 46368
rect 21358 46248 21364 46300
rect 21416 46288 21422 46300
rect 450814 46288 450820 46300
rect 21416 46260 450820 46288
rect 21416 46248 21422 46260
rect 450814 46248 450820 46260
rect 450872 46248 450878 46300
rect 20806 46180 20812 46232
rect 20864 46220 20870 46232
rect 20864 46192 358032 46220
rect 20864 46180 20870 46192
rect 20714 46112 20720 46164
rect 20772 46152 20778 46164
rect 358004 46152 358032 46192
rect 359826 46180 359832 46232
rect 359884 46220 359890 46232
rect 362310 46220 362316 46232
rect 359884 46192 362316 46220
rect 359884 46180 359890 46192
rect 362310 46180 362316 46192
rect 362368 46180 362374 46232
rect 361390 46152 361396 46164
rect 20772 46124 354812 46152
rect 358004 46124 361396 46152
rect 20772 46112 20778 46124
rect 354784 46084 354812 46124
rect 361390 46112 361396 46124
rect 361448 46112 361454 46164
rect 361298 46084 361304 46096
rect 354784 46056 361304 46084
rect 361298 46044 361304 46056
rect 361356 46044 361362 46096
rect 3418 45500 3424 45552
rect 3476 45540 3482 45552
rect 453298 45540 453304 45552
rect 3476 45512 453304 45540
rect 3476 45500 3482 45512
rect 453298 45500 453304 45512
rect 453356 45500 453362 45552
rect 21450 45432 21456 45484
rect 21508 45472 21514 45484
rect 450998 45472 451004 45484
rect 21508 45444 451004 45472
rect 21508 45432 21514 45444
rect 450998 45432 451004 45444
rect 451056 45432 451062 45484
rect 3510 45364 3516 45416
rect 3568 45404 3574 45416
rect 396718 45404 396724 45416
rect 3568 45376 396724 45404
rect 3568 45364 3574 45376
rect 396718 45364 396724 45376
rect 396776 45364 396782 45416
rect 20714 45296 20720 45348
rect 20772 45336 20778 45348
rect 359826 45336 359832 45348
rect 20772 45308 359832 45336
rect 20772 45296 20778 45308
rect 359826 45296 359832 45308
rect 359884 45296 359890 45348
rect 65518 45228 65524 45280
rect 65576 45268 65582 45280
rect 403710 45268 403716 45280
rect 65576 45240 403716 45268
rect 65576 45228 65582 45240
rect 403710 45228 403716 45240
rect 403768 45228 403774 45280
rect 38378 45160 38384 45212
rect 38436 45200 38442 45212
rect 379238 45200 379244 45212
rect 38436 45172 379244 45200
rect 38436 45160 38442 45172
rect 379238 45160 379244 45172
rect 379296 45160 379302 45212
rect 62022 45092 62028 45144
rect 62080 45132 62086 45144
rect 403894 45132 403900 45144
rect 62080 45104 403900 45132
rect 62080 45092 62086 45104
rect 403894 45092 403900 45104
rect 403952 45092 403958 45144
rect 58434 45024 58440 45076
rect 58492 45064 58498 45076
rect 403618 45064 403624 45076
rect 58492 45036 403624 45064
rect 58492 45024 58498 45036
rect 403618 45024 403624 45036
rect 403676 45024 403682 45076
rect 54938 44956 54944 45008
rect 54996 44996 55002 45008
rect 403802 44996 403808 45008
rect 54996 44968 403808 44996
rect 54996 44956 55002 44968
rect 403802 44956 403808 44968
rect 403860 44956 403866 45008
rect 51350 44888 51356 44940
rect 51408 44928 51414 44940
rect 406470 44928 406476 44940
rect 51408 44900 406476 44928
rect 51408 44888 51414 44900
rect 406470 44888 406476 44900
rect 406528 44888 406534 44940
rect 47854 44820 47860 44872
rect 47912 44860 47918 44872
rect 406746 44860 406752 44872
rect 47912 44832 406752 44860
rect 47912 44820 47918 44832
rect 406746 44820 406752 44832
rect 406804 44820 406810 44872
rect 69106 44752 69112 44804
rect 69164 44792 69170 44804
rect 403986 44792 403992 44804
rect 69164 44764 403992 44792
rect 69164 44752 69170 44764
rect 403986 44752 403992 44764
rect 404044 44752 404050 44804
rect 84470 44684 84476 44736
rect 84528 44724 84534 44736
rect 387518 44724 387524 44736
rect 84528 44696 387524 44724
rect 84528 44684 84534 44696
rect 387518 44684 387524 44696
rect 387576 44684 387582 44736
rect 108114 44616 108120 44668
rect 108172 44656 108178 44668
rect 395798 44656 395804 44668
rect 108172 44628 395804 44656
rect 108172 44616 108178 44628
rect 395798 44616 395804 44628
rect 395856 44616 395862 44668
rect 93946 42712 93952 42764
rect 94004 42752 94010 42764
rect 398190 42752 398196 42764
rect 94004 42724 398196 42752
rect 94004 42712 94010 42724
rect 398190 42712 398196 42724
rect 398248 42712 398254 42764
rect 80882 42644 80888 42696
rect 80940 42684 80946 42696
rect 387426 42684 387432 42696
rect 80940 42656 387432 42684
rect 80940 42644 80946 42656
rect 387426 42644 387432 42656
rect 387484 42644 387490 42696
rect 90358 42576 90364 42628
rect 90416 42616 90422 42628
rect 398098 42616 398104 42628
rect 90416 42588 398104 42616
rect 90416 42576 90422 42588
rect 398098 42576 398104 42588
rect 398156 42576 398162 42628
rect 86862 42508 86868 42560
rect 86920 42548 86926 42560
rect 398374 42548 398380 42560
rect 86920 42520 398380 42548
rect 86920 42508 86926 42520
rect 398374 42508 398380 42520
rect 398432 42508 398438 42560
rect 83274 42440 83280 42492
rect 83332 42480 83338 42492
rect 401318 42480 401324 42492
rect 83332 42452 401324 42480
rect 83332 42440 83338 42452
rect 401318 42440 401324 42452
rect 401376 42440 401382 42492
rect 79686 42372 79692 42424
rect 79744 42412 79750 42424
rect 400950 42412 400956 42424
rect 79744 42384 400956 42412
rect 79744 42372 79750 42384
rect 400950 42372 400956 42384
rect 401008 42372 401014 42424
rect 76190 42304 76196 42356
rect 76248 42344 76254 42356
rect 401042 42344 401048 42356
rect 76248 42316 401048 42344
rect 76248 42304 76254 42316
rect 401042 42304 401048 42316
rect 401100 42304 401106 42356
rect 72602 42236 72608 42288
rect 72660 42276 72666 42288
rect 401134 42276 401140 42288
rect 72660 42248 401140 42276
rect 72660 42236 72666 42248
rect 401134 42236 401140 42248
rect 401192 42236 401198 42288
rect 111610 42168 111616 42220
rect 111668 42208 111674 42220
rect 460198 42208 460204 42220
rect 111668 42180 460204 42208
rect 111668 42168 111674 42180
rect 460198 42168 460204 42180
rect 460256 42168 460262 42220
rect 101030 42100 101036 42152
rect 101088 42140 101094 42152
rect 454678 42140 454684 42152
rect 101088 42112 454684 42140
rect 101088 42100 101094 42112
rect 454678 42100 454684 42112
rect 454736 42100 454742 42152
rect 12342 42032 12348 42084
rect 12400 42072 12406 42084
rect 401226 42072 401232 42084
rect 12400 42044 401232 42072
rect 12400 42032 12406 42044
rect 401226 42032 401232 42044
rect 401284 42032 401290 42084
rect 97442 41964 97448 42016
rect 97500 42004 97506 42016
rect 398282 42004 398288 42016
rect 97500 41976 398288 42004
rect 97500 41964 97506 41976
rect 398282 41964 398288 41976
rect 398340 41964 398346 42016
rect 106918 41896 106924 41948
rect 106976 41936 106982 41948
rect 370958 41936 370964 41948
rect 106976 41908 370964 41936
rect 106976 41896 106982 41908
rect 370958 41896 370964 41908
rect 371016 41896 371022 41948
rect 475378 41352 475384 41404
rect 475436 41392 475442 41404
rect 536834 41392 536840 41404
rect 475436 41364 536840 41392
rect 475436 41352 475442 41364
rect 536834 41352 536840 41364
rect 536892 41352 536898 41404
rect 102226 39992 102232 40044
rect 102284 40032 102290 40044
rect 384574 40032 384580 40044
rect 102284 40004 384580 40032
rect 102284 39992 102290 40004
rect 384574 39992 384580 40004
rect 384632 39992 384638 40044
rect 71498 39924 71504 39976
rect 71556 39964 71562 39976
rect 373534 39964 373540 39976
rect 71556 39936 373540 39964
rect 71556 39924 71562 39936
rect 373534 39924 373540 39936
rect 373592 39924 373598 39976
rect 59630 39856 59636 39908
rect 59688 39896 59694 39908
rect 390278 39896 390284 39908
rect 59688 39868 390284 39896
rect 59688 39856 59694 39868
rect 390278 39856 390284 39868
rect 390336 39856 390342 39908
rect 118786 39788 118792 39840
rect 118844 39828 118850 39840
rect 450630 39828 450636 39840
rect 118844 39800 450636 39828
rect 118844 39788 118850 39800
rect 450630 39788 450636 39800
rect 450688 39788 450694 39840
rect 56042 39720 56048 39772
rect 56100 39760 56106 39772
rect 390186 39760 390192 39772
rect 56100 39732 390192 39760
rect 56100 39720 56106 39732
rect 390186 39720 390192 39732
rect 390244 39720 390250 39772
rect 48958 39652 48964 39704
rect 49016 39692 49022 39704
rect 392854 39692 392860 39704
rect 49016 39664 392860 39692
rect 49016 39652 49022 39664
rect 392854 39652 392860 39664
rect 392912 39652 392918 39704
rect 104526 39584 104532 39636
rect 104584 39624 104590 39636
rect 451090 39624 451096 39636
rect 104584 39596 451096 39624
rect 104584 39584 104590 39596
rect 451090 39584 451096 39596
rect 451148 39584 451154 39636
rect 44266 39516 44272 39568
rect 44324 39556 44330 39568
rect 393038 39556 393044 39568
rect 44324 39528 393044 39556
rect 44324 39516 44330 39528
rect 393038 39516 393044 39528
rect 393096 39516 393102 39568
rect 40678 39448 40684 39500
rect 40736 39488 40742 39500
rect 392946 39488 392952 39500
rect 40736 39460 392952 39488
rect 40736 39448 40742 39460
rect 392946 39448 392952 39460
rect 393004 39448 393010 39500
rect 4062 39380 4068 39432
rect 4120 39420 4126 39432
rect 392762 39420 392768 39432
rect 4120 39392 392768 39420
rect 4120 39380 4126 39392
rect 392762 39380 392768 39392
rect 392820 39380 392826 39432
rect 26510 39312 26516 39364
rect 26568 39352 26574 39364
rect 450906 39352 450912 39364
rect 26568 39324 450912 39352
rect 26568 39312 26574 39324
rect 450906 39312 450912 39324
rect 450964 39312 450970 39364
rect 115198 39244 115204 39296
rect 115256 39284 115262 39296
rect 395614 39284 395620 39296
rect 115256 39256 395620 39284
rect 115256 39244 115262 39256
rect 395614 39244 395620 39256
rect 395672 39244 395678 39296
rect 122282 39176 122288 39228
rect 122340 39216 122346 39228
rect 395706 39216 395712 39228
rect 122340 39188 395712 39216
rect 122340 39176 122346 39188
rect 395706 39176 395712 39188
rect 395764 39176 395770 39228
rect 105722 37204 105728 37256
rect 105780 37244 105786 37256
rect 384482 37244 384488 37256
rect 105780 37216 384488 37244
rect 105780 37204 105786 37216
rect 384482 37204 384488 37216
rect 384540 37204 384546 37256
rect 98638 37136 98644 37188
rect 98696 37176 98702 37188
rect 384390 37176 384396 37188
rect 98696 37148 384396 37176
rect 98696 37136 98702 37148
rect 384390 37136 384396 37148
rect 384448 37136 384454 37188
rect 95142 37068 95148 37120
rect 95200 37108 95206 37120
rect 384298 37108 384304 37120
rect 95200 37080 384304 37108
rect 95200 37068 95206 37080
rect 384298 37068 384304 37080
rect 384356 37068 384362 37120
rect 91554 37000 91560 37052
rect 91612 37040 91618 37052
rect 387150 37040 387156 37052
rect 91612 37012 387156 37040
rect 91612 37000 91618 37012
rect 387150 37000 387156 37012
rect 387208 37000 387214 37052
rect 87966 36932 87972 36984
rect 88024 36972 88030 36984
rect 387242 36972 387248 36984
rect 88024 36944 387248 36972
rect 88024 36932 88030 36944
rect 387242 36932 387248 36944
rect 387300 36932 387306 36984
rect 77386 36864 77392 36916
rect 77444 36904 77450 36916
rect 387334 36904 387340 36916
rect 77444 36876 387340 36904
rect 77444 36864 77450 36876
rect 387334 36864 387340 36876
rect 387392 36864 387398 36916
rect 73798 36796 73804 36848
rect 73856 36836 73862 36848
rect 390002 36836 390008 36848
rect 73856 36808 390008 36836
rect 73856 36796 73862 36808
rect 390002 36796 390008 36808
rect 390060 36796 390066 36848
rect 70302 36728 70308 36780
rect 70360 36768 70366 36780
rect 390094 36768 390100 36780
rect 70360 36740 390100 36768
rect 70360 36728 70366 36740
rect 390094 36728 390100 36740
rect 390152 36728 390158 36780
rect 66714 36660 66720 36712
rect 66772 36700 66778 36712
rect 389910 36700 389916 36712
rect 66772 36672 389916 36700
rect 66772 36660 66778 36672
rect 389910 36660 389916 36672
rect 389968 36660 389974 36712
rect 63218 36592 63224 36644
rect 63276 36632 63282 36644
rect 389818 36632 389824 36644
rect 63276 36604 389824 36632
rect 63276 36592 63282 36604
rect 389818 36592 389824 36604
rect 389876 36592 389882 36644
rect 28902 36524 28908 36576
rect 28960 36564 28966 36576
rect 368198 36564 368204 36576
rect 28960 36536 368204 36564
rect 28960 36524 28966 36536
rect 368198 36524 368204 36536
rect 368256 36524 368262 36576
rect 109310 36456 109316 36508
rect 109368 36496 109374 36508
rect 381722 36496 381728 36508
rect 109368 36468 381728 36496
rect 109368 36456 109374 36468
rect 381722 36456 381728 36468
rect 381780 36456 381786 36508
rect 112806 36388 112812 36440
rect 112864 36428 112870 36440
rect 381998 36428 382004 36440
rect 112864 36400 382004 36428
rect 112864 36388 112870 36400
rect 381998 36388 382004 36400
rect 382056 36388 382062 36440
rect 119890 34416 119896 34468
rect 119948 34456 119954 34468
rect 381538 34456 381544 34468
rect 119948 34428 381544 34456
rect 119948 34416 119954 34428
rect 381538 34416 381544 34428
rect 381596 34416 381602 34468
rect 116394 34348 116400 34400
rect 116452 34388 116458 34400
rect 381814 34388 381820 34400
rect 116452 34360 381820 34388
rect 116452 34348 116458 34360
rect 381814 34348 381820 34360
rect 381872 34348 381878 34400
rect 60826 34280 60832 34332
rect 60884 34320 60890 34332
rect 376478 34320 376484 34332
rect 60884 34292 376484 34320
rect 60884 34280 60890 34292
rect 376478 34280 376484 34292
rect 376536 34280 376542 34332
rect 57238 34212 57244 34264
rect 57296 34252 57302 34264
rect 376386 34252 376392 34264
rect 57296 34224 376392 34252
rect 57296 34212 57302 34224
rect 376386 34212 376392 34224
rect 376444 34212 376450 34264
rect 50154 34144 50160 34196
rect 50212 34184 50218 34196
rect 376110 34184 376116 34196
rect 50212 34156 376116 34184
rect 50212 34144 50218 34156
rect 376110 34144 376116 34156
rect 376168 34144 376174 34196
rect 45462 34076 45468 34128
rect 45520 34116 45526 34128
rect 376202 34116 376208 34128
rect 45520 34088 376208 34116
rect 45520 34076 45526 34088
rect 376202 34076 376208 34088
rect 376260 34076 376266 34128
rect 41874 34008 41880 34060
rect 41932 34048 41938 34060
rect 376294 34048 376300 34060
rect 41932 34020 376300 34048
rect 41932 34008 41938 34020
rect 376294 34008 376300 34020
rect 376352 34008 376358 34060
rect 34790 33940 34796 33992
rect 34848 33980 34854 33992
rect 379054 33980 379060 33992
rect 34848 33952 379060 33980
rect 34848 33940 34854 33952
rect 379054 33940 379060 33952
rect 379112 33940 379118 33992
rect 31294 33872 31300 33924
rect 31352 33912 31358 33924
rect 379146 33912 379152 33924
rect 31352 33884 379152 33912
rect 31352 33872 31358 33884
rect 379146 33872 379152 33884
rect 379204 33872 379210 33924
rect 23014 33804 23020 33856
rect 23072 33844 23078 33856
rect 378962 33844 378968 33856
rect 23072 33816 378968 33844
rect 23072 33804 23078 33816
rect 378962 33804 378968 33816
rect 379020 33804 379026 33856
rect 18230 33736 18236 33788
rect 18288 33776 18294 33788
rect 381906 33776 381912 33788
rect 18288 33748 381912 33776
rect 18288 33736 18294 33748
rect 381906 33736 381912 33748
rect 381964 33736 381970 33788
rect 123478 33668 123484 33720
rect 123536 33708 123542 33720
rect 378778 33708 378784 33720
rect 123536 33680 378784 33708
rect 123536 33668 123542 33680
rect 378778 33668 378784 33680
rect 378836 33668 378842 33720
rect 111058 33600 111064 33652
rect 111116 33640 111122 33652
rect 365346 33640 365352 33652
rect 111116 33612 365352 33640
rect 111116 33600 111122 33612
rect 365346 33600 365352 33612
rect 365404 33600 365410 33652
rect 2866 33056 2872 33108
rect 2924 33096 2930 33108
rect 400858 33096 400864 33108
rect 2924 33068 400864 33096
rect 2924 33056 2930 33068
rect 400858 33056 400864 33068
rect 400916 33056 400922 33108
rect 569218 33056 569224 33108
rect 569276 33096 569282 33108
rect 580166 33096 580172 33108
rect 569276 33068 580172 33096
rect 569276 33056 569282 33068
rect 580166 33056 580172 33068
rect 580224 33056 580230 33108
rect 117590 31696 117596 31748
rect 117648 31736 117654 31748
rect 367738 31736 367744 31748
rect 117648 31708 367744 31736
rect 117648 31696 117654 31708
rect 367738 31696 367744 31708
rect 367796 31696 367802 31748
rect 114002 31628 114008 31680
rect 114060 31668 114066 31680
rect 368014 31668 368020 31680
rect 114060 31640 368020 31668
rect 114060 31628 114066 31640
rect 368014 31628 368020 31640
rect 368072 31628 368078 31680
rect 99834 31560 99840 31612
rect 99892 31600 99898 31612
rect 370774 31600 370780 31612
rect 99892 31572 370780 31600
rect 99892 31560 99898 31572
rect 370774 31560 370780 31572
rect 370832 31560 370838 31612
rect 96246 31492 96252 31544
rect 96304 31532 96310 31544
rect 370866 31532 370872 31544
rect 96304 31504 370872 31532
rect 96304 31492 96310 31504
rect 370866 31492 370872 31504
rect 370924 31492 370930 31544
rect 89162 31424 89168 31476
rect 89220 31464 89226 31476
rect 370498 31464 370504 31476
rect 89220 31436 370504 31464
rect 89220 31424 89226 31436
rect 370498 31424 370504 31436
rect 370556 31424 370562 31476
rect 78582 31356 78588 31408
rect 78640 31396 78646 31408
rect 370590 31396 370596 31408
rect 78640 31368 370596 31396
rect 78640 31356 78646 31368
rect 370590 31356 370596 31368
rect 370648 31356 370654 31408
rect 74994 31288 75000 31340
rect 75052 31328 75058 31340
rect 373258 31328 373264 31340
rect 75052 31300 373264 31328
rect 75052 31288 75058 31300
rect 373258 31288 373264 31300
rect 373316 31288 373322 31340
rect 67910 31220 67916 31272
rect 67968 31260 67974 31272
rect 373350 31260 373356 31272
rect 67968 31232 373356 31260
rect 67968 31220 67974 31232
rect 373350 31220 373356 31232
rect 373408 31220 373414 31272
rect 64322 31152 64328 31204
rect 64380 31192 64386 31204
rect 373442 31192 373448 31204
rect 64380 31164 373448 31192
rect 64380 31152 64386 31164
rect 373442 31152 373448 31164
rect 373500 31152 373506 31204
rect 19426 31084 19432 31136
rect 19484 31124 19490 31136
rect 368106 31124 368112 31136
rect 19484 31096 368112 31124
rect 19484 31084 19490 31096
rect 368106 31084 368112 31096
rect 368164 31084 368170 31136
rect 14734 31016 14740 31068
rect 14792 31056 14798 31068
rect 370682 31056 370688 31068
rect 14792 31028 370688 31056
rect 14792 31016 14798 31028
rect 370682 31016 370688 31028
rect 370740 31016 370746 31068
rect 121086 30948 121092 31000
rect 121144 30988 121150 31000
rect 367922 30988 367928 31000
rect 121144 30960 367928 30988
rect 121144 30948 121150 30960
rect 367922 30948 367928 30960
rect 367980 30948 367986 31000
rect 124674 30880 124680 30932
rect 124732 30920 124738 30932
rect 367830 30920 367836 30932
rect 124732 30892 367836 30920
rect 124732 30880 124738 30892
rect 367830 30880 367836 30892
rect 367888 30880 367894 30932
rect 46658 28432 46664 28484
rect 46716 28472 46722 28484
rect 365254 28472 365260 28484
rect 46716 28444 365260 28472
rect 46716 28432 46722 28444
rect 365254 28432 365260 28444
rect 365312 28432 365318 28484
rect 43070 28364 43076 28416
rect 43128 28404 43134 28416
rect 365070 28404 365076 28416
rect 43128 28376 365076 28404
rect 43128 28364 43134 28376
rect 365070 28364 365076 28376
rect 365128 28364 365134 28416
rect 35986 28296 35992 28348
rect 36044 28336 36050 28348
rect 364978 28336 364984 28348
rect 36044 28308 364984 28336
rect 36044 28296 36050 28308
rect 364978 28296 364984 28308
rect 365036 28296 365042 28348
rect 32398 28228 32404 28280
rect 32456 28268 32462 28280
rect 365162 28268 365168 28280
rect 32456 28240 365168 28268
rect 32456 28228 32462 28240
rect 365162 28228 365168 28240
rect 365220 28228 365226 28280
rect 3418 20612 3424 20664
rect 3476 20652 3482 20664
rect 381630 20652 381636 20664
rect 3476 20624 381636 20652
rect 3476 20612 3482 20624
rect 381630 20612 381636 20624
rect 381688 20612 381694 20664
rect 574738 20612 574744 20664
rect 574796 20652 574802 20664
rect 579982 20652 579988 20664
rect 574796 20624 579988 20652
rect 574796 20612 574802 20624
rect 579982 20612 579988 20624
rect 580040 20612 580046 20664
rect 3418 6808 3424 6860
rect 3476 6848 3482 6860
rect 395430 6848 395436 6860
rect 3476 6820 395436 6848
rect 3476 6808 3482 6820
rect 395430 6808 395436 6820
rect 395488 6808 395494 6860
rect 562318 6808 562324 6860
rect 562376 6848 562382 6860
rect 580166 6848 580172 6860
rect 562376 6820 580172 6848
rect 562376 6808 562382 6820
rect 580166 6808 580172 6820
rect 580224 6808 580230 6860
rect 85666 4088 85672 4140
rect 85724 4128 85730 4140
rect 363690 4128 363696 4140
rect 85724 4100 363696 4128
rect 85724 4088 85730 4100
rect 363690 4088 363696 4100
rect 363748 4088 363754 4140
rect 53742 4020 53748 4072
rect 53800 4060 53806 4072
rect 361114 4060 361120 4072
rect 53800 4032 361120 4060
rect 53800 4020 53806 4032
rect 361114 4020 361120 4032
rect 361172 4020 361178 4072
rect 39574 3952 39580 4004
rect 39632 3992 39638 4004
rect 360838 3992 360844 4004
rect 39632 3964 360844 3992
rect 39632 3952 39638 3964
rect 360838 3952 360844 3964
rect 360896 3952 360902 4004
rect 33594 3884 33600 3936
rect 33652 3924 33658 3936
rect 359458 3924 359464 3936
rect 33652 3896 359464 3924
rect 33652 3884 33658 3896
rect 359458 3884 359464 3896
rect 359516 3884 359522 3936
rect 27706 3816 27712 3868
rect 27764 3856 27770 3868
rect 378870 3856 378876 3868
rect 27764 3828 378876 3856
rect 27764 3816 27770 3828
rect 378870 3816 378876 3828
rect 378928 3816 378934 3868
rect 37182 3748 37188 3800
rect 37240 3788 37246 3800
rect 392670 3788 392676 3800
rect 37240 3760 392676 3788
rect 37240 3748 37246 3760
rect 392670 3748 392676 3760
rect 392728 3748 392734 3800
rect 82078 3680 82084 3732
rect 82136 3720 82142 3732
rect 450538 3720 450544 3732
rect 82136 3692 450544 3720
rect 82136 3680 82142 3692
rect 450538 3680 450544 3692
rect 450596 3680 450602 3732
rect 21818 3612 21824 3664
rect 21876 3652 21882 3664
rect 395522 3652 395528 3664
rect 21876 3624 395528 3652
rect 21876 3612 21882 3624
rect 395522 3612 395528 3624
rect 395580 3612 395586 3664
rect 24210 3544 24216 3596
rect 24268 3584 24274 3596
rect 407758 3584 407764 3596
rect 24268 3556 407764 3584
rect 24268 3544 24274 3556
rect 407758 3544 407764 3556
rect 407816 3544 407822 3596
rect 52546 3476 52552 3528
rect 52604 3516 52610 3528
rect 456058 3516 456064 3528
rect 52604 3488 456064 3516
rect 52604 3476 52610 3488
rect 456058 3476 456064 3488
rect 456116 3476 456122 3528
rect 17034 3408 17040 3460
rect 17092 3448 17098 3460
rect 450722 3448 450728 3460
rect 17092 3420 450728 3448
rect 17092 3408 17098 3420
rect 450722 3408 450728 3420
rect 450780 3408 450786 3460
rect 92750 3340 92756 3392
rect 92808 3380 92814 3392
rect 362218 3380 362224 3392
rect 92808 3352 362224 3380
rect 92808 3340 92814 3352
rect 362218 3340 362224 3352
rect 362276 3340 362282 3392
rect 103330 3272 103336 3324
rect 103388 3312 103394 3324
rect 361022 3312 361028 3324
rect 103388 3284 361028 3312
rect 103388 3272 103394 3284
rect 361022 3272 361028 3284
rect 361080 3272 361086 3324
rect 110506 3204 110512 3256
rect 110564 3244 110570 3256
rect 360930 3244 360936 3256
rect 110564 3216 360936 3244
rect 110564 3204 110570 3216
rect 360930 3204 360936 3216
rect 360988 3204 360994 3256
rect 6454 3136 6460 3188
rect 6512 3176 6518 3188
rect 111058 3176 111064 3188
rect 6512 3148 111064 3176
rect 6512 3136 6518 3148
rect 111058 3136 111064 3148
rect 111116 3136 111122 3188
rect 30098 2048 30104 2100
rect 30156 2088 30162 2100
rect 395338 2088 395344 2100
rect 30156 2060 395344 2088
rect 30156 2048 30162 2060
rect 395338 2048 395344 2060
rect 395396 2048 395402 2100
<< via1 >>
rect 267648 700816 267700 700868
rect 445116 700816 445168 700868
rect 235172 700748 235224 700800
rect 449256 700748 449308 700800
rect 218980 700680 219032 700732
rect 446496 700680 446548 700732
rect 154120 700612 154172 700664
rect 418804 700612 418856 700664
rect 429844 700612 429896 700664
rect 444104 700612 444156 700664
rect 170312 700544 170364 700596
rect 446404 700544 446456 700596
rect 137836 700476 137888 700528
rect 445208 700476 445260 700528
rect 105452 700408 105504 700460
rect 444196 700408 444248 700460
rect 447876 700408 447928 700460
rect 478512 700408 478564 700460
rect 40500 700340 40552 700392
rect 449164 700340 449216 700392
rect 8116 700272 8168 700324
rect 445024 700272 445076 700324
rect 447784 700272 447836 700324
rect 494796 700272 494848 700324
rect 348792 686536 348844 686588
rect 446588 686536 446640 686588
rect 283840 686468 283892 686520
rect 446680 686468 446732 686520
rect 332508 685312 332560 685364
rect 418896 685312 418948 685364
rect 202788 685244 202840 685296
rect 445300 685244 445352 685296
rect 89168 685176 89220 685228
rect 416044 685176 416096 685228
rect 72976 685108 73028 685160
rect 449348 685108 449400 685160
rect 19984 684564 20036 684616
rect 418988 684564 419040 684616
rect 3792 684496 3844 684548
rect 420184 684496 420236 684548
rect 18328 683748 18380 683800
rect 359464 683748 359516 683800
rect 21364 683680 21416 683732
rect 420736 683680 420788 683732
rect 4068 683612 4120 683664
rect 420276 683612 420328 683664
rect 3516 683544 3568 683596
rect 420368 683544 420420 683596
rect 3700 683476 3752 683528
rect 420644 683476 420696 683528
rect 3424 683408 3476 683460
rect 420552 683408 420604 683460
rect 3884 683340 3936 683392
rect 445484 683340 445536 683392
rect 3608 683272 3660 683324
rect 445392 683272 445444 683324
rect 3976 683204 4028 683256
rect 446864 683204 446916 683256
rect 3332 683136 3384 683188
rect 446312 683136 446364 683188
rect 576124 683136 576176 683188
rect 579620 683136 579672 683188
rect 3240 682660 3292 682712
rect 447048 682660 447100 682712
rect 17224 680348 17276 680400
rect 18328 680348 18380 680400
rect 359464 672052 359516 672104
rect 360844 672052 360896 672104
rect 361764 667904 361816 667956
rect 378876 667904 378928 667956
rect 14188 660968 14240 661020
rect 17224 661036 17276 661088
rect 3148 658180 3200 658232
rect 19984 658180 20036 658232
rect 361764 656888 361816 656940
rect 376024 656888 376076 656940
rect 11704 656616 11756 656668
rect 14188 656616 14240 656668
rect 361764 645872 361816 645924
rect 374644 645872 374696 645924
rect 10600 645804 10652 645856
rect 11704 645804 11756 645856
rect 5540 643696 5592 643748
rect 10600 643696 10652 643748
rect 4804 640296 4856 640348
rect 5540 640296 5592 640348
rect 361580 634788 361632 634840
rect 400864 634788 400916 634840
rect 3608 631320 3660 631372
rect 20904 631320 20956 631372
rect 361580 623772 361632 623824
rect 371884 623772 371936 623824
rect 570604 616836 570656 616888
rect 579620 616836 579672 616888
rect 361580 612824 361632 612876
rect 363604 612824 363656 612876
rect 458824 604120 458876 604172
rect 458824 603916 458876 603968
rect 459008 603712 459060 603764
rect 459468 603712 459520 603764
rect 459836 602080 459888 602132
rect 460112 602080 460164 602132
rect 361764 601672 361816 601724
rect 370504 601672 370556 601724
rect 460112 600244 460164 600296
rect 462320 600244 462372 600296
rect 457352 600176 457404 600228
rect 462964 600176 463016 600228
rect 457536 599768 457588 599820
rect 464344 599768 464396 599820
rect 459008 599700 459060 599752
rect 466460 599700 466512 599752
rect 458732 599632 458784 599684
rect 469220 599632 469272 599684
rect 457444 599564 457496 599616
rect 468484 599564 468536 599616
rect 515404 599564 515456 599616
rect 580540 599564 580592 599616
rect 457260 598680 457312 598732
rect 461584 598680 461636 598732
rect 459468 598408 459520 598460
rect 463700 598408 463752 598460
rect 458640 598272 458692 598324
rect 465080 598272 465132 598324
rect 488632 598272 488684 598324
rect 494336 598272 494388 598324
rect 360844 598204 360896 598256
rect 367744 598204 367796 598256
rect 457720 598204 457772 598256
rect 465724 598204 465776 598256
rect 493324 598204 493376 598256
rect 526720 598204 526772 598256
rect 459836 596844 459888 596896
rect 466552 596844 466604 596896
rect 450544 596776 450596 596828
rect 494980 596776 495032 596828
rect 457904 595892 457956 595944
rect 461676 595892 461728 595944
rect 460204 595484 460256 595536
rect 467932 595484 467984 595536
rect 457628 595416 457680 595468
rect 468576 595416 468628 595468
rect 460020 594124 460072 594176
rect 465172 594124 465224 594176
rect 457812 594056 457864 594108
rect 467104 594056 467156 594108
rect 361580 590792 361632 590844
rect 363696 590792 363748 590844
rect 511264 590656 511316 590708
rect 580172 590656 580224 590708
rect 367744 587800 367796 587852
rect 370596 587800 370648 587852
rect 361764 579640 361816 579692
rect 368020 579640 368072 579692
rect 370596 579572 370648 579624
rect 371976 579572 372028 579624
rect 511356 576852 511408 576904
rect 579988 576852 580040 576904
rect 371976 571276 372028 571328
rect 373264 571276 373316 571328
rect 361580 568760 361632 568812
rect 363788 568760 363840 568812
rect 373264 564340 373316 564392
rect 375288 564340 375340 564392
rect 515496 563048 515548 563100
rect 580172 563048 580224 563100
rect 361672 557540 361724 557592
rect 403624 557540 403676 557592
rect 375380 557132 375432 557184
rect 377772 557132 377824 557184
rect 377772 550604 377824 550656
rect 380164 550536 380216 550588
rect 361764 546456 361816 546508
rect 419080 546456 419132 546508
rect 459928 542988 459980 543040
rect 463792 542988 463844 543040
rect 380164 540880 380216 540932
rect 382280 540880 382332 540932
rect 519544 536800 519596 536852
rect 580172 536800 580224 536852
rect 361764 535440 361816 535492
rect 406384 535440 406436 535492
rect 382280 532652 382332 532704
rect 384304 532652 384356 532704
rect 361764 524424 361816 524476
rect 407764 524424 407816 524476
rect 518164 524424 518216 524476
rect 580172 524424 580224 524476
rect 384304 524084 384356 524136
rect 385684 524084 385736 524136
rect 457996 522316 458048 522368
rect 464436 522316 464488 522368
rect 459192 522248 459244 522300
rect 469404 522248 469456 522300
rect 459284 520888 459336 520940
rect 470600 520888 470652 520940
rect 482928 520888 482980 520940
rect 520280 520888 520332 520940
rect 458088 519596 458140 519648
rect 468668 519596 468720 519648
rect 459376 519528 459428 519580
rect 470876 519528 470928 519580
rect 449716 518168 449768 518220
rect 469864 518168 469916 518220
rect 494244 518168 494296 518220
rect 476028 517624 476080 517676
rect 494152 517624 494204 517676
rect 449808 517556 449860 517608
rect 488632 517556 488684 517608
rect 450360 517488 450412 517540
rect 494336 517488 494388 517540
rect 482284 517420 482336 517472
rect 450636 516808 450688 516860
rect 476028 516808 476080 516860
rect 449992 516740 450044 516792
rect 492128 516740 492180 516792
rect 385684 516128 385736 516180
rect 389180 516060 389232 516112
rect 3976 514768 4028 514820
rect 4804 514768 4856 514820
rect 502248 514020 502300 514072
rect 545120 514020 545172 514072
rect 361764 513340 361816 513392
rect 410524 513340 410576 513392
rect 492128 512592 492180 512644
rect 535460 512592 535512 512644
rect 389180 511912 389232 511964
rect 391204 511912 391256 511964
rect 516784 510620 516836 510672
rect 580172 510620 580224 510672
rect 494336 509872 494388 509924
rect 538220 509872 538272 509924
rect 494152 508512 494204 508564
rect 532700 508512 532752 508564
rect 391204 505792 391256 505844
rect 392584 505792 392636 505844
rect 495072 505724 495124 505776
rect 529940 505724 529992 505776
rect 361764 502324 361816 502376
rect 411904 502324 411956 502376
rect 463148 497700 463200 497752
rect 480260 497700 480312 497752
rect 458824 497632 458876 497684
rect 481640 497632 481692 497684
rect 457536 497564 457588 497616
rect 482652 497564 482704 497616
rect 457444 497496 457496 497548
rect 483848 497496 483900 497548
rect 454684 497428 454736 497480
rect 486240 497428 486292 497480
rect 455328 497020 455380 497072
rect 459560 497020 459612 497072
rect 456524 496952 456576 497004
rect 461032 496952 461084 497004
rect 453948 496884 454000 496936
rect 456616 496884 456668 496936
rect 452568 496816 452620 496868
rect 453672 496816 453724 496868
rect 455144 496816 455196 496868
rect 458088 496816 458140 496868
rect 483664 496816 483716 496868
rect 485044 496816 485096 496868
rect 361764 491308 361816 491360
rect 381636 491308 381688 491360
rect 518256 484372 518308 484424
rect 580172 484372 580224 484424
rect 361764 480224 361816 480276
rect 419172 480224 419224 480276
rect 361764 469208 361816 469260
rect 396724 469208 396776 469260
rect 494704 462476 494756 462528
rect 527640 462476 527692 462528
rect 453304 462408 453356 462460
rect 524696 462408 524748 462460
rect 450544 462340 450596 462392
rect 542360 462340 542412 462392
rect 467196 460980 467248 461032
rect 553860 460980 553912 461032
rect 458916 460912 458968 460964
rect 550916 460912 550968 460964
rect 447508 458804 447560 458856
rect 483664 458804 483716 458856
rect 361764 458192 361816 458244
rect 414664 458192 414716 458244
rect 569224 456764 569276 456816
rect 580172 456764 580224 456816
rect 392584 456696 392636 456748
rect 395344 456696 395396 456748
rect 488264 456016 488316 456068
rect 494704 456016 494756 456068
rect 461768 455472 461820 455524
rect 488264 455472 488316 455524
rect 452016 455404 452068 455456
rect 480996 455404 481048 455456
rect 449716 454724 449768 454776
rect 487160 454724 487212 454776
rect 449624 454656 449676 454708
rect 489920 454656 489972 454708
rect 459008 454044 459060 454096
rect 473728 454044 473780 454096
rect 447416 448468 447468 448520
rect 458916 448468 458968 448520
rect 447232 447856 447284 447908
rect 448336 447856 448388 447908
rect 459008 447856 459060 447908
rect 447140 447788 447192 447840
rect 447968 447788 448020 447840
rect 467196 447788 467248 447840
rect 422484 447380 422536 447432
rect 447232 447380 447284 447432
rect 437388 447312 437440 447364
rect 447140 447312 447192 447364
rect 432420 447244 432472 447296
rect 447416 447244 447468 447296
rect 427452 447176 427504 447228
rect 445668 447176 445720 447228
rect 361764 447108 361816 447160
rect 399484 447108 399536 447160
rect 442632 444320 442684 444372
rect 446220 444320 446272 444372
rect 361764 436092 361816 436144
rect 416136 436092 416188 436144
rect 395344 433236 395396 433288
rect 398104 433236 398156 433288
rect 458088 429972 458140 430024
rect 474280 429972 474332 430024
rect 459468 429904 459520 429956
rect 476948 429904 477000 429956
rect 459376 429836 459428 429888
rect 479616 429836 479668 429888
rect 480904 429156 480956 429208
rect 482284 429156 482336 429208
rect 483664 429156 483716 429208
rect 484952 429156 485004 429208
rect 457628 428408 457680 428460
rect 471612 428408 471664 428460
rect 361764 425076 361816 425128
rect 417424 425076 417476 425128
rect 503628 424328 503680 424380
rect 557540 424328 557592 424380
rect 398104 423580 398156 423632
rect 398840 423580 398892 423632
rect 529204 423580 529256 423632
rect 530216 423580 530268 423632
rect 530584 423580 530636 423632
rect 532792 423580 532844 423632
rect 511540 423512 511592 423564
rect 523776 423512 523828 423564
rect 522304 423444 522356 423496
rect 549536 423444 549588 423496
rect 502984 423376 503036 423428
rect 522488 423376 522540 423428
rect 523684 423376 523736 423428
rect 552112 423376 552164 423428
rect 487068 423308 487120 423360
rect 526352 423308 526404 423360
rect 526444 423308 526496 423360
rect 554688 423308 554740 423360
rect 488264 423240 488316 423292
rect 528928 423240 528980 423292
rect 489644 423172 489696 423224
rect 531504 423172 531556 423224
rect 498108 423104 498160 423156
rect 545672 423104 545724 423156
rect 499304 423036 499356 423088
rect 548248 423036 548300 423088
rect 444288 422968 444340 423020
rect 447876 422968 447928 423020
rect 500684 422968 500736 423020
rect 550824 422968 550876 423020
rect 502248 422900 502300 422952
rect 553400 422900 553452 422952
rect 484308 421540 484360 421592
rect 521200 421540 521252 421592
rect 495348 420180 495400 420232
rect 541808 420180 541860 420232
rect 398840 418820 398892 418872
rect 400680 418820 400732 418872
rect 425980 417732 426032 417784
rect 507952 417732 508004 417784
rect 425336 417664 425388 417716
rect 507860 417664 507912 417716
rect 422116 417596 422168 417648
rect 503996 417596 504048 417648
rect 421472 417528 421524 417580
rect 503720 417528 503772 417580
rect 424692 417460 424744 417512
rect 506480 417460 506532 417512
rect 424048 417392 424100 417444
rect 506572 417392 506624 417444
rect 423128 416304 423180 416356
rect 423588 416304 423640 416356
rect 486976 416032 487028 416084
rect 527640 416032 527692 416084
rect 361580 413992 361632 414044
rect 443644 413992 443696 414044
rect 400680 413924 400732 413976
rect 402336 413924 402388 413976
rect 402336 410524 402388 410576
rect 409144 410524 409196 410576
rect 511448 404336 511500 404388
rect 580172 404336 580224 404388
rect 361580 402976 361632 403028
rect 439504 402976 439556 403028
rect 497924 400868 497976 400920
rect 546500 400868 546552 400920
rect 494612 399440 494664 399492
rect 539600 399440 539652 399492
rect 493968 398080 494020 398132
rect 538220 398080 538272 398132
rect 493416 396720 493468 396772
rect 536840 396720 536892 396772
rect 409144 396040 409196 396092
rect 411628 395972 411680 396024
rect 460756 395292 460808 395344
rect 483664 395292 483716 395344
rect 492404 395292 492456 395344
rect 535460 395292 535512 395344
rect 496728 394000 496780 394052
rect 543740 394000 543792 394052
rect 423496 393932 423548 393984
rect 505560 393932 505612 393984
rect 463608 392572 463660 392624
rect 487160 392572 487212 392624
rect 491576 392572 491628 392624
rect 534172 392572 534224 392624
rect 361580 391960 361632 392012
rect 443736 391960 443788 392012
rect 495716 391280 495768 391332
rect 542360 391280 542412 391332
rect 411628 391212 411680 391264
rect 415400 391212 415452 391264
rect 423588 391212 423640 391264
rect 505284 391212 505336 391264
rect 459652 389852 459704 389904
rect 480904 389852 480956 389904
rect 448060 389784 448112 389836
rect 463148 389784 463200 389836
rect 464896 389784 464948 389836
rect 489920 389784 489972 389836
rect 490564 389784 490616 389836
rect 534080 389784 534132 389836
rect 458456 389240 458508 389292
rect 459468 389240 459520 389292
rect 465080 389240 465132 389292
rect 465908 389240 465960 389292
rect 466460 389240 466512 389292
rect 467380 389240 467432 389292
rect 486424 389240 486476 389292
rect 487068 389240 487120 389292
rect 497464 389240 497516 389292
rect 498108 389240 498160 389292
rect 506480 389240 506532 389292
rect 507124 389240 507176 389292
rect 415400 389104 415452 389156
rect 417516 389104 417568 389156
rect 453028 389104 453080 389156
rect 454040 389104 454092 389156
rect 456708 389104 456760 389156
rect 457628 389104 457680 389156
rect 468484 389036 468536 389088
rect 475844 389036 475896 389088
rect 468576 388968 468628 389020
rect 478052 388968 478104 389020
rect 502340 388968 502392 389020
rect 467104 388900 467156 388952
rect 478788 388900 478840 388952
rect 461584 388832 461636 388884
rect 473636 388832 473688 388884
rect 483940 388832 483992 388884
rect 502984 388832 503036 388884
rect 526444 388832 526496 388884
rect 461124 388764 461176 388816
rect 463608 388764 463660 388816
rect 464344 388764 464396 388816
rect 476580 388764 476632 388816
rect 500868 388764 500920 388816
rect 523684 388764 523736 388816
rect 462964 388696 463016 388748
rect 475108 388696 475160 388748
rect 499396 388696 499448 388748
rect 522304 388696 522356 388748
rect 468668 388628 468720 388680
rect 481732 388628 481784 388680
rect 484676 388628 484728 388680
rect 511540 388628 511592 388680
rect 447784 388560 447836 388612
rect 457444 388560 457496 388612
rect 465724 388560 465776 388612
rect 480260 388560 480312 388612
rect 485412 388560 485464 388612
rect 524420 388560 524472 388612
rect 447692 388492 447744 388544
rect 457536 388492 457588 388544
rect 464528 388492 464580 388544
rect 480996 388492 481048 388544
rect 488356 388492 488408 388544
rect 529204 388492 529256 388544
rect 450728 388424 450780 388476
rect 461768 388424 461820 388476
rect 463056 388424 463108 388476
rect 482468 388424 482520 388476
rect 489828 388424 489880 388476
rect 530584 388424 530636 388476
rect 461676 387880 461728 387932
rect 462596 387880 462648 387932
rect 461860 387812 461912 387864
rect 464896 387812 464948 387864
rect 447876 387200 447928 387252
rect 458824 387200 458876 387252
rect 448980 387132 449032 387184
rect 491300 387132 491352 387184
rect 449532 387064 449584 387116
rect 513380 387064 513432 387116
rect 448336 386656 448388 386708
rect 553952 386656 554004 386708
rect 381544 386588 381596 386640
rect 512092 386588 512144 386640
rect 378784 386520 378836 386572
rect 512552 386520 512604 386572
rect 367744 386452 367796 386504
rect 512000 386452 512052 386504
rect 367836 386384 367888 386436
rect 512276 386384 512328 386436
rect 448244 385976 448296 386028
rect 453304 385976 453356 386028
rect 448428 385636 448480 385688
rect 454408 385636 454460 385688
rect 448152 385364 448204 385416
rect 452016 385364 452068 385416
rect 449440 385092 449492 385144
rect 563428 385092 563480 385144
rect 367928 385024 367980 385076
rect 512368 385024 512420 385076
rect 513196 383732 513248 383784
rect 534724 383732 534776 383784
rect 513288 383664 513340 383716
rect 548524 383664 548576 383716
rect 362224 383596 362276 383648
rect 447140 383596 447192 383648
rect 378876 383528 378928 383580
rect 447232 383528 447284 383580
rect 512644 382916 512696 382968
rect 519728 382916 519780 382968
rect 513012 382712 513064 382764
rect 518348 382712 518400 382764
rect 512460 382440 512512 382492
rect 515588 382440 515640 382492
rect 374644 382168 374696 382220
rect 447232 382168 447284 382220
rect 376024 382100 376076 382152
rect 447140 382100 447192 382152
rect 361580 380876 361632 380928
rect 443828 380876 443880 380928
rect 512460 380876 512512 380928
rect 547144 380876 547196 380928
rect 363604 380808 363656 380860
rect 447416 380808 447468 380860
rect 371884 380740 371936 380792
rect 447140 380740 447192 380792
rect 400864 380672 400916 380724
rect 447232 380672 447284 380724
rect 512552 379720 512604 379772
rect 515680 379720 515732 379772
rect 513288 379516 513340 379568
rect 549904 379516 549956 379568
rect 363696 379448 363748 379500
rect 447324 379448 447376 379500
rect 370504 379380 370556 379432
rect 447140 379380 447192 379432
rect 417516 378904 417568 378956
rect 419264 378904 419316 378956
rect 513288 378292 513340 378344
rect 522304 378292 522356 378344
rect 512828 378224 512880 378276
rect 547236 378224 547288 378276
rect 514024 378156 514076 378208
rect 580172 378156 580224 378208
rect 363788 378088 363840 378140
rect 447232 378088 447284 378140
rect 368020 378020 368072 378072
rect 447140 378020 447192 378072
rect 513196 377408 513248 377460
rect 548616 377408 548668 377460
rect 513196 376728 513248 376780
rect 516968 376728 517020 376780
rect 403624 376660 403676 376712
rect 447140 376660 447192 376712
rect 419080 376592 419132 376644
rect 447232 376592 447284 376644
rect 513012 375980 513064 376032
rect 544384 375980 544436 376032
rect 406384 375300 406436 375352
rect 447140 375300 447192 375352
rect 407764 375232 407816 375284
rect 447232 375232 447284 375284
rect 513288 374144 513340 374196
rect 517520 374144 517572 374196
rect 410524 373940 410576 373992
rect 447140 373940 447192 373992
rect 411904 373872 411956 373924
rect 447232 373872 447284 373924
rect 513288 372648 513340 372700
rect 518900 372648 518952 372700
rect 512644 372580 512696 372632
rect 521660 372580 521712 372632
rect 381636 372512 381688 372564
rect 447140 372512 447192 372564
rect 419172 372444 419224 372496
rect 447232 372444 447284 372496
rect 512000 371696 512052 371748
rect 513840 371696 513892 371748
rect 396724 371152 396776 371204
rect 447140 371152 447192 371204
rect 414664 371084 414716 371136
rect 447232 371084 447284 371136
rect 512092 370200 512144 370252
rect 514760 370200 514812 370252
rect 513288 370064 513340 370116
rect 517612 370064 517664 370116
rect 361580 369860 361632 369912
rect 409880 369860 409932 369912
rect 513288 369860 513340 369912
rect 523040 369860 523092 369912
rect 399484 369792 399536 369844
rect 447140 369792 447192 369844
rect 416136 369724 416188 369776
rect 447232 369724 447284 369776
rect 419264 369316 419316 369368
rect 421564 369316 421616 369368
rect 512092 369112 512144 369164
rect 520280 369112 520332 369164
rect 512276 368568 512328 368620
rect 515128 368568 515180 368620
rect 417424 368432 417476 368484
rect 447140 368432 447192 368484
rect 443644 368364 443696 368416
rect 447232 368364 447284 368416
rect 513288 367344 513340 367396
rect 520372 367344 520424 367396
rect 439504 367004 439556 367056
rect 447140 367004 447192 367056
rect 443736 366936 443788 366988
rect 447232 366936 447284 366988
rect 513288 365712 513340 365764
rect 521752 365712 521804 365764
rect 409880 365644 409932 365696
rect 447140 365644 447192 365696
rect 443828 365576 443880 365628
rect 447232 365576 447284 365628
rect 512000 365576 512052 365628
rect 514208 365576 514260 365628
rect 513288 365032 513340 365084
rect 519084 365032 519136 365084
rect 512828 364352 512880 364404
rect 518992 364352 519044 364404
rect 573364 364352 573416 364404
rect 580172 364352 580224 364404
rect 512000 363196 512052 363248
rect 514852 363196 514904 363248
rect 432880 362992 432932 363044
rect 447232 362992 447284 363044
rect 432788 362924 432840 362976
rect 447140 362924 447192 362976
rect 421564 362448 421616 362500
rect 423588 362448 423640 362500
rect 512000 362312 512052 362364
rect 513656 362312 513708 362364
rect 442264 361632 442316 361684
rect 447232 361632 447284 361684
rect 513012 361632 513064 361684
rect 519176 361632 519228 361684
rect 432696 361564 432748 361616
rect 447140 361564 447192 361616
rect 513288 361564 513340 361616
rect 523132 361564 523184 361616
rect 512644 360680 512696 360732
rect 520556 360680 520608 360732
rect 512000 360408 512052 360460
rect 514944 360408 514996 360460
rect 439688 360272 439740 360324
rect 447232 360272 447284 360324
rect 436928 360204 436980 360256
rect 447140 360204 447192 360256
rect 547236 360136 547288 360188
rect 552020 360136 552072 360188
rect 534724 360068 534776 360120
rect 566740 360068 566792 360120
rect 549904 360000 549956 360052
rect 554964 360000 555016 360052
rect 548524 359932 548576 359984
rect 565268 359932 565320 359984
rect 547144 359864 547196 359916
rect 558184 359864 558236 359916
rect 515680 359796 515732 359848
rect 553768 359796 553820 359848
rect 522304 359728 522356 359780
rect 550824 359728 550876 359780
rect 443828 358844 443880 358896
rect 447232 358844 447284 358896
rect 435456 358776 435508 358828
rect 447140 358776 447192 358828
rect 513012 358776 513064 358828
rect 519268 358776 519320 358828
rect 548616 358708 548668 358760
rect 556712 358708 556764 358760
rect 519728 358640 519780 358692
rect 564072 358640 564124 358692
rect 518348 358572 518400 358624
rect 562600 358572 562652 358624
rect 544384 358504 544436 358556
rect 559656 358504 559708 358556
rect 515588 358436 515640 358488
rect 561128 358436 561180 358488
rect 423588 357416 423640 357468
rect 426348 357348 426400 357400
rect 512828 356328 512880 356380
rect 516232 356328 516284 356380
rect 513288 356192 513340 356244
rect 520464 356192 520516 356244
rect 513288 354968 513340 355020
rect 517704 354968 517756 355020
rect 513288 354696 513340 354748
rect 517888 354696 517940 354748
rect 512092 354152 512144 354204
rect 513748 354152 513800 354204
rect 445668 353948 445720 354000
rect 448428 353948 448480 354000
rect 513288 353472 513340 353524
rect 517796 353472 517848 353524
rect 446220 352520 446272 352572
rect 447784 352520 447836 352572
rect 512460 352248 512512 352300
rect 515220 352248 515272 352300
rect 426440 351908 426492 351960
rect 432972 351840 433024 351892
rect 512460 350820 512512 350872
rect 515588 350820 515640 350872
rect 512920 350616 512972 350668
rect 516324 350616 516376 350668
rect 407028 350548 407080 350600
rect 447140 350548 447192 350600
rect 364984 349800 365036 349852
rect 442356 349800 442408 349852
rect 512828 349664 512880 349716
rect 517980 349664 518032 349716
rect 432972 349528 433024 349580
rect 433984 349528 434036 349580
rect 513288 349392 513340 349444
rect 519360 349392 519412 349444
rect 512092 349256 512144 349308
rect 513932 349256 513984 349308
rect 513288 348440 513340 348492
rect 520648 348440 520700 348492
rect 513288 348168 513340 348220
rect 518072 348168 518124 348220
rect 361764 347760 361816 347812
rect 402244 347760 402296 347812
rect 362224 347692 362276 347744
rect 447140 347692 447192 347744
rect 512092 346740 512144 346792
rect 515036 346740 515088 346792
rect 512644 346536 512696 346588
rect 516508 346536 516560 346588
rect 512920 343680 512972 343732
rect 516416 343680 516468 343732
rect 513196 342592 513248 342644
rect 518348 342592 518400 342644
rect 513288 342252 513340 342304
rect 521844 342252 521896 342304
rect 512644 341232 512696 341284
rect 515312 341232 515364 341284
rect 444196 340960 444248 341012
rect 447232 340960 447284 341012
rect 512828 340960 512880 341012
rect 516600 340960 516652 341012
rect 361764 340892 361816 340944
rect 447140 340892 447192 340944
rect 513288 340008 513340 340060
rect 519452 340008 519504 340060
rect 431224 339532 431276 339584
rect 447140 339532 447192 339584
rect 371884 339464 371936 339516
rect 447232 339464 447284 339516
rect 513196 339464 513248 339516
rect 521936 339464 521988 339516
rect 513288 338512 513340 338564
rect 520740 338512 520792 338564
rect 436836 338172 436888 338224
rect 447140 338172 447192 338224
rect 435364 338104 435416 338156
rect 447232 338104 447284 338156
rect 402244 338036 402296 338088
rect 448428 338036 448480 338088
rect 449440 338036 449492 338088
rect 433984 337968 434036 338020
rect 436376 337968 436428 338020
rect 450084 337424 450136 337476
rect 450360 337424 450412 337476
rect 513288 337288 513340 337340
rect 519728 337288 519780 337340
rect 513104 337152 513156 337204
rect 516876 337152 516928 337204
rect 416780 336880 416832 336932
rect 450360 336880 450412 336932
rect 413100 336812 413152 336864
rect 450176 336812 450228 336864
rect 409420 336744 409472 336796
rect 450728 336744 450780 336796
rect 513196 336744 513248 336796
rect 522028 336744 522080 336796
rect 448428 336676 448480 336728
rect 449716 336676 449768 336728
rect 418804 336404 418856 336456
rect 439872 336404 439924 336456
rect 418896 336336 418948 336388
rect 442540 336336 442592 336388
rect 416044 336268 416096 336320
rect 439780 336268 439832 336320
rect 440884 336268 440936 336320
rect 447140 336268 447192 336320
rect 418988 336200 419040 336252
rect 449532 336200 449584 336252
rect 413652 336132 413704 336184
rect 449624 336132 449676 336184
rect 397460 336064 397512 336116
rect 447692 336064 447744 336116
rect 362224 335996 362276 336048
rect 444196 335996 444248 336048
rect 443736 335656 443788 335708
rect 447140 335656 447192 335708
rect 399484 335316 399536 335368
rect 447416 335316 447468 335368
rect 513288 335316 513340 335368
rect 522120 335316 522172 335368
rect 432604 334908 432656 334960
rect 447508 334908 447560 334960
rect 420552 334840 420604 334892
rect 442448 334840 442500 334892
rect 420736 334772 420788 334824
rect 442632 334772 442684 334824
rect 420184 334704 420236 334756
rect 444932 334704 444984 334756
rect 420276 334636 420328 334688
rect 445668 334636 445720 334688
rect 420644 334568 420696 334620
rect 449716 334568 449768 334620
rect 513288 334568 513340 334620
rect 520832 334568 520884 334620
rect 443644 334024 443696 334076
rect 447232 334024 447284 334076
rect 363788 333956 363840 334008
rect 447140 333956 447192 334008
rect 513288 333956 513340 334008
rect 522212 333956 522264 334008
rect 513012 333072 513064 333124
rect 516692 333072 516744 333124
rect 512644 332868 512696 332920
rect 514116 332868 514168 332920
rect 439596 332664 439648 332716
rect 447232 332664 447284 332716
rect 436744 332596 436796 332648
rect 447140 332596 447192 332648
rect 512644 331440 512696 331492
rect 516140 331440 516192 331492
rect 442908 330488 442960 330540
rect 447968 330488 448020 330540
rect 450084 330488 450136 330540
rect 450728 330488 450780 330540
rect 580724 330488 580776 330540
rect 580908 330488 580960 330540
rect 432880 330148 432932 330200
rect 439688 330148 439740 330200
rect 439504 329808 439556 329860
rect 447140 329808 447192 329860
rect 436376 329740 436428 329792
rect 438124 329740 438176 329792
rect 436008 328516 436060 328568
rect 449900 328516 449952 328568
rect 431868 328448 431920 328500
rect 450452 328448 450504 328500
rect 509516 326340 509568 326392
rect 510160 326340 510212 326392
rect 509332 326204 509384 326256
rect 509516 326204 509568 326256
rect 432880 324912 432932 324964
rect 442264 324912 442316 324964
rect 438124 323960 438176 324012
rect 439964 323960 440016 324012
rect 432696 322940 432748 322992
rect 436928 322940 436980 322992
rect 444104 322804 444156 322856
rect 570604 322872 570656 322924
rect 458272 322668 458324 322720
rect 458824 322668 458876 322720
rect 458548 322600 458600 322652
rect 580540 322804 580592 322856
rect 459100 322668 459152 322720
rect 468208 322668 468260 322720
rect 469036 322668 469088 322720
rect 469588 322668 469640 322720
rect 459376 322600 459428 322652
rect 468484 322600 468536 322652
rect 569224 322736 569276 322788
rect 471244 322668 471296 322720
rect 516784 322668 516836 322720
rect 471520 322600 471572 322652
rect 515496 322600 515548 322652
rect 444932 322532 444984 322584
rect 468760 322532 468812 322584
rect 470968 322532 471020 322584
rect 458824 322464 458876 322516
rect 459376 322464 459428 322516
rect 470140 322464 470192 322516
rect 484216 322532 484268 322584
rect 479800 322464 479852 322516
rect 518256 322464 518308 322516
rect 445668 322396 445720 322448
rect 483940 322396 483992 322448
rect 449716 322328 449768 322380
rect 455788 322328 455840 322380
rect 458272 322328 458324 322380
rect 460480 322328 460532 322380
rect 468484 322328 468536 322380
rect 471520 322328 471572 322380
rect 439872 322260 439924 322312
rect 472072 322260 472124 322312
rect 507860 322260 507912 322312
rect 580264 322260 580316 322312
rect 439964 322192 440016 322244
rect 466552 322192 466604 322244
rect 468208 322192 468260 322244
rect 471244 322192 471296 322244
rect 500224 322192 500276 322244
rect 580172 322192 580224 322244
rect 447692 322124 447744 322176
rect 481456 322124 481508 322176
rect 469312 322056 469364 322108
rect 469588 322056 469640 322108
rect 455788 321988 455840 322040
rect 463516 321988 463568 322040
rect 469036 321988 469088 322040
rect 470968 321988 471020 322040
rect 507308 321648 507360 321700
rect 509792 321648 509844 321700
rect 447048 321512 447100 321564
rect 463056 321512 463108 321564
rect 468576 321512 468628 321564
rect 573364 321512 573416 321564
rect 458364 321444 458416 321496
rect 511448 321444 511500 321496
rect 449256 321376 449308 321428
rect 461400 321376 461452 321428
rect 469404 321376 469456 321428
rect 518164 321376 518216 321428
rect 446404 321308 446456 321360
rect 461676 321308 461728 321360
rect 479064 321308 479116 321360
rect 514024 321308 514076 321360
rect 445024 321240 445076 321292
rect 483204 321240 483256 321292
rect 445484 321172 445536 321224
rect 473820 321172 473872 321224
rect 507400 321172 507452 321224
rect 513472 321172 513524 321224
rect 446496 321104 446548 321156
rect 471888 321104 471940 321156
rect 507216 321104 507268 321156
rect 516140 321104 516192 321156
rect 460204 321036 460256 321088
rect 513840 321036 513892 321088
rect 445116 320968 445168 321020
rect 482100 320968 482152 321020
rect 496820 320968 496872 321020
rect 580632 320968 580684 321020
rect 459928 320900 459980 320952
rect 580356 320900 580408 320952
rect 461860 320832 461912 320884
rect 580816 320832 580868 320884
rect 446956 320764 447008 320816
rect 473268 320764 473320 320816
rect 439780 320696 439832 320748
rect 472440 320696 472492 320748
rect 442540 320628 442592 320680
rect 481824 320628 481876 320680
rect 442356 320084 442408 320136
rect 446864 320016 446916 320068
rect 458088 320084 458140 320136
rect 461860 320084 461912 320136
rect 480720 320084 480772 320136
rect 507860 320084 507912 320136
rect 460848 320016 460900 320068
rect 466552 320016 466604 320068
rect 474372 320016 474424 320068
rect 479340 320016 479392 320068
rect 496820 320016 496872 320068
rect 463332 319948 463384 320000
rect 470232 319948 470284 320000
rect 576124 319948 576176 320000
rect 479892 319880 479944 319932
rect 519544 319880 519596 319932
rect 442632 319812 442684 319864
rect 463884 319812 463936 319864
rect 469680 319812 469732 319864
rect 511356 319812 511408 319864
rect 449624 319744 449676 319796
rect 471060 319744 471112 319796
rect 480996 319744 481048 319796
rect 519636 319744 519688 319796
rect 445392 319676 445444 319728
rect 462780 319676 462832 319728
rect 480444 319676 480496 319728
rect 515404 319676 515456 319728
rect 460388 319608 460440 319660
rect 465816 319608 465868 319660
rect 480168 319608 480220 319660
rect 511264 319608 511316 319660
rect 459008 319540 459060 319592
rect 465540 319540 465592 319592
rect 498660 319540 498712 319592
rect 534724 319540 534776 319592
rect 460296 319472 460348 319524
rect 476304 319472 476356 319524
rect 498108 319472 498160 319524
rect 533344 319472 533396 319524
rect 458824 319404 458876 319456
rect 476028 319404 476080 319456
rect 478788 319404 478840 319456
rect 500224 319404 500276 319456
rect 501696 319404 501748 319456
rect 538864 319404 538916 319456
rect 446588 319336 446640 319388
rect 471336 319336 471388 319388
rect 481272 319336 481324 319388
rect 510620 319336 510672 319388
rect 445300 319268 445352 319320
rect 482376 319268 482428 319320
rect 502800 319268 502852 319320
rect 530584 319268 530636 319320
rect 468852 319200 468904 319252
rect 580908 319200 580960 319252
rect 455788 319132 455840 319184
rect 456064 319132 456116 319184
rect 457168 319132 457220 319184
rect 457996 319132 458048 319184
rect 466828 319132 466880 319184
rect 467380 319132 467432 319184
rect 469956 319132 470008 319184
rect 580448 319132 580500 319184
rect 442448 319064 442500 319116
rect 484308 319064 484360 319116
rect 497464 319064 497516 319116
rect 498016 319064 498068 319116
rect 501604 319064 501656 319116
rect 502156 319064 502208 319116
rect 446680 318996 446732 319048
rect 466644 318928 466696 318980
rect 467380 318928 467432 318980
rect 471244 318996 471296 319048
rect 474648 318996 474700 319048
rect 471612 318928 471664 318980
rect 449532 318724 449584 318776
rect 483480 318724 483532 318776
rect 444288 318656 444340 318708
rect 470784 318656 470836 318708
rect 432052 318248 432104 318300
rect 435456 318248 435508 318300
rect 454776 318180 454828 318232
rect 491484 318180 491536 318232
rect 496176 318180 496228 318232
rect 539600 318180 539652 318232
rect 456064 318112 456116 318164
rect 512092 318112 512144 318164
rect 476856 318044 476908 318096
rect 569224 318044 569276 318096
rect 478512 317704 478564 317756
rect 479524 317704 479576 317756
rect 453396 317364 453448 317416
rect 464988 317364 465040 317416
rect 456340 317296 456392 317348
rect 475752 317296 475804 317348
rect 456432 317228 456484 317280
rect 475476 317228 475528 317280
rect 453304 317160 453356 317212
rect 475200 317160 475252 317212
rect 459192 317092 459244 317144
rect 486516 317092 486568 317144
rect 458916 317024 458968 317076
rect 485964 317024 486016 317076
rect 453488 316956 453540 317008
rect 485688 316956 485740 317008
rect 450636 316888 450688 316940
rect 457720 316888 457772 316940
rect 459100 316888 459152 316940
rect 491668 316956 491720 317008
rect 487252 316888 487304 316940
rect 488356 316888 488408 316940
rect 500316 316888 500368 316940
rect 539784 316888 539836 316940
rect 451924 316820 451976 316872
rect 495900 316820 495952 316872
rect 502524 316820 502576 316872
rect 542636 316820 542688 316872
rect 450636 316752 450688 316804
rect 509516 316752 509568 316804
rect 450820 316684 450872 316736
rect 474924 316684 474976 316736
rect 477960 316684 478012 316736
rect 547144 316684 547196 316736
rect 453580 316616 453632 316668
rect 464712 316616 464764 316668
rect 481732 316616 481784 316668
rect 484400 316616 484452 316668
rect 485872 316616 485924 316668
rect 486976 316616 487028 316668
rect 487528 316616 487580 316668
rect 487804 316616 487856 316668
rect 487896 316616 487948 316668
rect 488356 316616 488408 316668
rect 488632 316616 488684 316668
rect 489184 316616 489236 316668
rect 490288 316616 490340 316668
rect 490840 316616 490892 316668
rect 493324 316616 493376 316668
rect 493876 316616 493928 316668
rect 494152 316616 494204 316668
rect 495256 316616 495308 316668
rect 456248 316548 456300 316600
rect 465264 316548 465316 316600
rect 490012 316548 490064 316600
rect 491116 316548 491168 316600
rect 491392 316480 491444 316532
rect 492220 316480 492272 316532
rect 457812 316004 457864 316056
rect 461584 316004 461636 316056
rect 361764 315936 361816 315988
rect 371884 315936 371936 315988
rect 457444 315392 457496 315444
rect 489736 315392 489788 315444
rect 501604 315392 501656 315444
rect 539876 315392 539928 315444
rect 459284 315324 459336 315376
rect 492496 315324 492548 315376
rect 496636 315324 496688 315376
rect 539692 315324 539744 315376
rect 478144 315256 478196 315308
rect 551284 315256 551336 315308
rect 451004 314032 451056 314084
rect 484768 314032 484820 314084
rect 503168 314032 503220 314084
rect 543188 314032 543240 314084
rect 459376 313964 459428 314016
rect 493600 313964 493652 314016
rect 496728 313964 496780 314016
rect 540980 313964 541032 314016
rect 433156 313896 433208 313948
rect 443828 313896 443880 313948
rect 455788 313896 455840 313948
rect 566464 313896 566516 313948
rect 482100 313556 482152 313608
rect 484492 313556 484544 313608
rect 461676 313284 461728 313336
rect 463792 313284 463844 313336
rect 469036 313216 469088 313268
rect 580172 313216 580224 313268
rect 439688 312536 439740 312588
rect 471244 312536 471296 312588
rect 478880 312536 478932 312588
rect 481732 312536 481784 312588
rect 502064 312536 502116 312588
rect 542544 312536 542596 312588
rect 494612 311856 494664 311908
rect 494796 311856 494848 311908
rect 469864 311244 469916 311296
rect 482100 311244 482152 311296
rect 454868 311176 454920 311228
rect 494428 311176 494480 311228
rect 467380 311108 467432 311160
rect 548524 311108 548576 311160
rect 456524 309884 456576 309936
rect 495624 309884 495676 309936
rect 503536 309884 503588 309936
rect 538956 309884 539008 309936
rect 487712 309816 487764 309868
rect 530032 309816 530084 309868
rect 452016 309748 452068 309800
rect 494796 309748 494848 309800
rect 502156 309748 502208 309800
rect 541072 309748 541124 309800
rect 453672 308456 453724 308508
rect 489184 308456 489236 308508
rect 503260 308456 503312 308508
rect 539048 308456 539100 308508
rect 487804 308388 487856 308440
rect 529940 308388 529992 308440
rect 476764 308320 476816 308372
rect 478880 308320 478932 308372
rect 3516 307708 3568 307760
rect 4804 307708 4856 307760
rect 453764 307096 453816 307148
rect 490288 307096 490340 307148
rect 457352 307028 457404 307080
rect 576124 307028 576176 307080
rect 446128 306280 446180 306332
rect 469864 306280 469916 306332
rect 457536 306212 457588 306264
rect 491392 306212 491444 306264
rect 400864 306144 400916 306196
rect 465448 306144 465500 306196
rect 477316 306144 477368 306196
rect 544384 306144 544436 306196
rect 406660 306076 406712 306128
rect 509976 306076 510028 306128
rect 406476 306008 406528 306060
rect 509608 306008 509660 306060
rect 403808 305940 403860 305992
rect 511172 305940 511224 305992
rect 403624 305872 403676 305924
rect 511080 305872 511132 305924
rect 403900 305804 403952 305856
rect 513932 305804 513984 305856
rect 403716 305736 403768 305788
rect 515588 305736 515640 305788
rect 363604 305668 363656 305720
rect 512736 305668 512788 305720
rect 360844 305600 360896 305652
rect 512644 305600 512696 305652
rect 361764 304920 361816 304972
rect 431224 304920 431276 304972
rect 450452 304580 450504 304632
rect 455972 304580 456024 304632
rect 444748 304512 444800 304564
rect 461676 304512 461728 304564
rect 455880 304444 455932 304496
rect 562324 304444 562376 304496
rect 363696 304376 363748 304428
rect 512368 304376 512420 304428
rect 360936 304308 360988 304360
rect 512000 304308 512052 304360
rect 361028 304240 361080 304292
rect 512184 304240 512236 304292
rect 401048 303560 401100 303612
rect 510988 303560 511040 303612
rect 403992 303492 404044 303544
rect 515220 303492 515272 303544
rect 401140 303424 401192 303476
rect 513748 303424 513800 303476
rect 395620 303356 395672 303408
rect 510712 303356 510764 303408
rect 398288 303288 398340 303340
rect 514208 303288 514260 303340
rect 456616 303220 456668 303272
rect 571984 303220 572036 303272
rect 398104 303152 398156 303204
rect 513656 303152 513708 303204
rect 398380 303084 398432 303136
rect 514944 303084 514996 303136
rect 398196 303016 398248 303068
rect 514852 303016 514904 303068
rect 395804 302948 395856 303000
rect 517612 302948 517664 303000
rect 361120 302880 361172 302932
rect 512460 302880 512512 302932
rect 401324 302812 401376 302864
rect 510804 302812 510856 302864
rect 400956 302744 401008 302796
rect 509424 302744 509476 302796
rect 395436 302676 395488 302728
rect 485872 302676 485924 302728
rect 456708 301520 456760 301572
rect 573364 301520 573416 301572
rect 362224 301452 362276 301504
rect 512276 301452 512328 301504
rect 440976 300636 441028 300688
rect 446128 300636 446180 300688
rect 457996 300636 458048 300688
rect 533436 300636 533488 300688
rect 395712 300568 395764 300620
rect 516968 300568 517020 300620
rect 393044 300500 393096 300552
rect 516600 300500 516652 300552
rect 392676 300432 392728 300484
rect 516876 300432 516928 300484
rect 392860 300364 392912 300416
rect 518348 300364 518400 300416
rect 390192 300296 390244 300348
rect 516508 300296 516560 300348
rect 389916 300228 389968 300280
rect 516324 300228 516376 300280
rect 390284 300160 390336 300212
rect 518072 300160 518124 300212
rect 389824 300092 389876 300144
rect 517980 300092 518032 300144
rect 436928 299548 436980 299600
rect 439688 299548 439740 299600
rect 461584 299412 461636 299464
rect 580172 299412 580224 299464
rect 387432 298052 387484 298104
rect 513564 298052 513616 298104
rect 390008 297984 390060 298036
rect 517888 297984 517940 298036
rect 387340 297916 387392 297968
rect 516232 297916 516284 297968
rect 384396 297848 384448 297900
rect 513380 297848 513432 297900
rect 387524 297780 387576 297832
rect 519268 297780 519320 297832
rect 387156 297712 387208 297764
rect 519176 297712 519228 297764
rect 381728 297644 381780 297696
rect 514760 297644 514812 297696
rect 387248 297576 387300 297628
rect 520556 297576 520608 297628
rect 384304 297508 384356 297560
rect 519084 297508 519136 297560
rect 384488 297440 384540 297492
rect 520280 297440 520332 297492
rect 384580 297372 384632 297424
rect 520372 297372 520424 297424
rect 387064 297304 387116 297356
rect 509700 297304 509752 297356
rect 390100 297236 390152 297288
rect 510896 297236 510948 297288
rect 439688 297168 439740 297220
rect 444748 297168 444800 297220
rect 457628 297168 457680 297220
rect 574836 297168 574888 297220
rect 477408 295944 477460 295996
rect 570604 295944 570656 295996
rect 381912 295264 381964 295316
rect 510068 295264 510120 295316
rect 376024 295196 376076 295248
rect 507492 295196 507544 295248
rect 381820 295128 381872 295180
rect 517520 295128 517572 295180
rect 382004 295060 382056 295112
rect 518900 295060 518952 295112
rect 378876 294992 378928 295044
rect 516692 294992 516744 295044
rect 376208 294924 376260 294976
rect 515312 294924 515364 294976
rect 376116 294856 376168 294908
rect 516416 294856 516468 294908
rect 379060 294788 379112 294840
rect 519728 294788 519780 294840
rect 379244 294720 379296 294772
rect 520740 294720 520792 294772
rect 379152 294652 379204 294704
rect 520832 294652 520884 294704
rect 376300 294584 376352 294636
rect 519452 294584 519504 294636
rect 396724 294516 396776 294568
rect 486424 294516 486476 294568
rect 447876 294448 447928 294500
rect 536104 294448 536156 294500
rect 361764 293904 361816 293956
rect 435364 293904 435416 293956
rect 467288 293224 467340 293276
rect 555424 293224 555476 293276
rect 3424 292544 3476 292596
rect 4896 292544 4948 292596
rect 437480 292544 437532 292596
rect 440976 292544 441028 292596
rect 376392 292476 376444 292528
rect 515036 292476 515088 292528
rect 376484 292408 376536 292460
rect 520648 292408 520700 292460
rect 373540 292340 373592 292392
rect 517796 292340 517848 292392
rect 373264 292272 373316 292324
rect 517704 292272 517756 292324
rect 373448 292204 373500 292256
rect 519360 292204 519412 292256
rect 370872 292136 370924 292188
rect 518992 292136 519044 292188
rect 370596 292068 370648 292120
rect 520464 292068 520516 292120
rect 370780 292000 370832 292052
rect 521752 292000 521804 292052
rect 370964 291932 371016 291984
rect 523040 291932 523092 291984
rect 370504 291864 370556 291916
rect 523132 291864 523184 291916
rect 368020 291796 368072 291848
rect 521660 291796 521712 291848
rect 370688 291728 370740 291780
rect 507400 291728 507452 291780
rect 373356 291660 373408 291712
rect 507308 291660 507360 291712
rect 478420 291592 478472 291644
rect 559656 291592 559708 291644
rect 467012 290436 467064 290488
rect 558184 290436 558236 290488
rect 427084 289552 427136 289604
rect 437480 289552 437532 289604
rect 447784 289552 447836 289604
rect 464068 289552 464120 289604
rect 407764 289484 407816 289536
rect 507216 289484 507268 289536
rect 365352 289416 365404 289468
rect 507124 289416 507176 289468
rect 368204 289348 368256 289400
rect 522212 289348 522264 289400
rect 365260 289280 365312 289332
rect 521844 289280 521896 289332
rect 365076 289212 365128 289264
rect 521936 289212 521988 289264
rect 365168 289144 365220 289196
rect 522120 289144 522172 289196
rect 364984 289076 365036 289128
rect 522028 289076 522080 289128
rect 488356 287648 488408 287700
rect 531320 287648 531372 287700
rect 381636 286356 381688 286408
rect 476488 286356 476540 286408
rect 500132 286356 500184 286408
rect 541164 286356 541216 286408
rect 410524 286288 410576 286340
rect 436928 286288 436980 286340
rect 467656 286288 467708 286340
rect 580264 286288 580316 286340
rect 469220 284996 469272 285048
rect 476764 284996 476816 285048
rect 498844 284996 498896 285048
rect 539968 284996 540020 285048
rect 466828 284928 466880 284980
rect 559564 284928 559616 284980
rect 452292 283568 452344 283620
rect 494704 283568 494756 283620
rect 361764 282820 361816 282872
rect 436836 282820 436888 282872
rect 459468 282140 459520 282192
rect 489000 282140 489052 282192
rect 462964 281868 463016 281920
rect 469220 281868 469272 281920
rect 455052 280780 455104 280832
rect 493416 280780 493468 280832
rect 497648 280780 497700 280832
rect 542452 280780 542504 280832
rect 447876 279488 447928 279540
rect 462964 279488 463016 279540
rect 453948 279420 454000 279472
rect 490564 279420 490616 279472
rect 498016 279420 498068 279472
rect 543280 279420 543332 279472
rect 452384 277992 452436 278044
rect 494152 277992 494204 278044
rect 455236 276632 455288 276684
rect 494520 276632 494572 276684
rect 499948 276632 500000 276684
rect 540060 276632 540112 276684
rect 488080 275340 488132 275392
rect 530124 275340 530176 275392
rect 458640 275272 458692 275324
rect 493324 275272 493376 275324
rect 499028 275272 499080 275324
rect 541256 275272 541308 275324
rect 453856 273980 453908 274032
rect 488632 273980 488684 274032
rect 431224 273912 431276 273964
rect 439688 273912 439740 273964
rect 454960 273912 455012 273964
rect 491668 273912 491720 273964
rect 499396 273912 499448 273964
rect 541348 273912 541400 273964
rect 479524 273164 479576 273216
rect 579896 273164 579948 273216
rect 455144 272552 455196 272604
rect 492772 272552 492824 272604
rect 452108 272484 452160 272536
rect 490104 272484 490156 272536
rect 500776 272484 500828 272536
rect 541440 272484 541492 272536
rect 361764 271804 361816 271856
rect 432604 271804 432656 271856
rect 458732 271260 458784 271312
rect 488908 271260 488960 271312
rect 456616 271192 456668 271244
rect 490012 271192 490064 271244
rect 500500 271192 500552 271244
rect 540244 271192 540296 271244
rect 457628 271124 457680 271176
rect 493140 271124 493192 271176
rect 499120 271124 499172 271176
rect 540152 271124 540204 271176
rect 456708 269900 456760 269952
rect 487252 269900 487304 269952
rect 505008 269900 505060 269952
rect 543740 269900 543792 269952
rect 400128 269832 400180 269884
rect 410524 269832 410576 269884
rect 468760 269832 468812 269884
rect 580356 269832 580408 269884
rect 359464 269764 359516 269816
rect 512828 269764 512880 269816
rect 452200 268404 452252 268456
rect 490380 268404 490432 268456
rect 497740 268404 497792 268456
rect 542820 268404 542872 268456
rect 466368 268336 466420 268388
rect 574744 268336 574796 268388
rect 445024 264936 445076 264988
rect 447876 264936 447928 264988
rect 396816 263576 396868 263628
rect 400128 263576 400180 263628
rect 449808 263508 449860 263560
rect 456800 263508 456852 263560
rect 417424 262828 417476 262880
rect 427084 262828 427136 262880
rect 444656 262216 444708 262268
rect 447784 262216 447836 262268
rect 361764 260788 361816 260840
rect 440884 260788 440936 260840
rect 406844 260108 406896 260160
rect 417424 260108 417476 260160
rect 439688 258680 439740 258732
rect 444656 258680 444708 258732
rect 3976 253920 4028 253972
rect 5080 253920 5132 253972
rect 422944 253920 422996 253972
rect 431224 253920 431276 253972
rect 361764 249704 361816 249756
rect 399484 249704 399536 249756
rect 449440 249024 449492 249076
rect 457812 249024 457864 249076
rect 435640 245624 435692 245676
rect 439688 245624 439740 245676
rect 574836 245556 574888 245608
rect 580172 245556 580224 245608
rect 420184 245284 420236 245336
rect 422944 245284 422996 245336
rect 400220 244876 400272 244928
rect 406844 244876 406896 244928
rect 3792 243924 3844 243976
rect 4988 243924 5040 243976
rect 388444 242156 388496 242208
rect 400220 242156 400272 242208
rect 382924 239436 382976 239488
rect 388444 239436 388496 239488
rect 369124 239368 369176 239420
rect 396816 239368 396868 239420
rect 427084 239368 427136 239420
rect 435640 239368 435692 239420
rect 361764 238688 361816 238740
rect 443736 238688 443788 238740
rect 411904 235220 411956 235272
rect 420184 235220 420236 235272
rect 455972 234948 456024 235000
rect 457996 234948 458048 235000
rect 559656 233180 559708 233232
rect 580172 233180 580224 233232
rect 442264 232908 442316 232960
rect 445024 232908 445076 232960
rect 362316 229712 362368 229764
rect 369124 229712 369176 229764
rect 361764 227672 361816 227724
rect 443644 227672 443696 227724
rect 399484 225564 399536 225616
rect 411904 225564 411956 225616
rect 439688 223524 439740 223576
rect 442264 223524 442316 223576
rect 3884 222096 3936 222148
rect 5172 222096 5224 222148
rect 450360 221416 450412 221468
rect 457996 221416 458048 221468
rect 361212 220056 361264 220108
rect 382924 220056 382976 220108
rect 436100 218016 436152 218068
rect 439688 218016 439740 218068
rect 361580 216316 361632 216368
rect 363788 216316 363840 216368
rect 413100 214548 413152 214600
rect 436100 214548 436152 214600
rect 396264 213936 396316 213988
rect 399484 213936 399536 213988
rect 377404 211760 377456 211812
rect 396264 211760 396316 211812
rect 407856 210128 407908 210180
rect 413100 210128 413152 210180
rect 411904 209040 411956 209092
rect 427084 209040 427136 209092
rect 399484 207612 399536 207664
rect 407856 207612 407908 207664
rect 576124 206932 576176 206984
rect 579804 206932 579856 206984
rect 361764 205572 361816 205624
rect 439596 205572 439648 205624
rect 408500 198704 408552 198756
rect 411904 198704 411956 198756
rect 447324 197956 447376 198008
rect 475384 197956 475436 198008
rect 374644 195100 374696 195152
rect 377404 195100 377456 195152
rect 361672 194488 361724 194540
rect 436744 194488 436796 194540
rect 393964 194420 394016 194472
rect 399484 194420 399536 194472
rect 547144 193128 547196 193180
rect 580172 193128 580224 193180
rect 401600 191088 401652 191140
rect 408500 191088 408552 191140
rect 398472 186328 398524 186380
rect 401600 186328 401652 186380
rect 390652 186260 390704 186312
rect 393964 186260 394016 186312
rect 361672 183472 361724 183524
rect 447600 183472 447652 183524
rect 448060 183472 448112 183524
rect 447600 182792 447652 182844
rect 528560 182792 528612 182844
rect 388444 181568 388496 181620
rect 390652 181568 390704 181620
rect 362960 180072 363012 180124
rect 374644 180072 374696 180124
rect 559564 179324 559616 179376
rect 580172 179324 580224 179376
rect 361304 174632 361356 174684
rect 362960 174632 363012 174684
rect 361672 172456 361724 172508
rect 447600 172456 447652 172508
rect 448244 172456 448296 172508
rect 447600 171776 447652 171828
rect 524420 171776 524472 171828
rect 386052 168376 386104 168428
rect 388444 168376 388496 168428
rect 533436 166948 533488 167000
rect 580172 166948 580224 167000
rect 438584 163616 438636 163668
rect 439504 163616 439556 163668
rect 378692 162868 378744 162920
rect 386052 162868 386104 162920
rect 418712 162324 418764 162376
rect 457904 162324 457956 162376
rect 489920 162324 489972 162376
rect 414756 162256 414808 162308
rect 457996 162256 458048 162308
rect 485780 162256 485832 162308
rect 411628 162188 411680 162240
rect 458088 162188 458140 162240
rect 481640 162188 481692 162240
rect 445208 162120 445260 162172
rect 457812 162120 457864 162172
rect 533436 162120 533488 162172
rect 406844 161440 406896 161492
rect 414756 161440 414808 161492
rect 361764 161372 361816 161424
rect 448336 161372 448388 161424
rect 448336 160692 448388 160744
rect 521660 160692 521712 160744
rect 425336 160488 425388 160540
rect 426348 160488 426400 160540
rect 496820 160488 496872 160540
rect 428648 160420 428700 160472
rect 500960 160420 501012 160472
rect 422024 160352 422076 160404
rect 494060 160352 494112 160404
rect 431776 160284 431828 160336
rect 505100 160284 505152 160336
rect 404084 160216 404136 160268
rect 418160 160216 418212 160268
rect 435272 160216 435324 160268
rect 436008 160216 436060 160268
rect 509240 160216 509292 160268
rect 407856 160148 407908 160200
rect 411444 160148 411496 160200
rect 438584 160148 438636 160200
rect 513380 160148 513432 160200
rect 409696 160080 409748 160132
rect 441574 160080 441626 160132
rect 442908 160080 442960 160132
rect 517520 160080 517572 160132
rect 409144 159672 409196 159724
rect 421380 159672 421432 159724
rect 409236 159604 409288 159656
rect 425152 159604 425204 159656
rect 409328 159536 409380 159588
rect 428004 159536 428056 159588
rect 409420 159468 409472 159520
rect 431316 159468 431368 159520
rect 409512 159400 409564 159452
rect 434812 159400 434864 159452
rect 409604 159332 409656 159384
rect 437940 159332 437992 159384
rect 452568 158244 452620 158296
rect 456708 158244 456760 158296
rect 373632 156612 373684 156664
rect 378692 156612 378744 156664
rect 452568 155660 452620 155712
rect 456524 155660 456576 155712
rect 551284 153144 551336 153196
rect 580172 153144 580224 153196
rect 361764 150356 361816 150408
rect 409696 150356 409748 150408
rect 451556 150220 451608 150272
rect 455236 150220 455288 150272
rect 371240 149676 371292 149728
rect 398472 149676 398524 149728
rect 451740 148996 451792 149048
rect 454868 148996 454920 149048
rect 451740 147364 451792 147416
rect 458640 147364 458692 147416
rect 452568 146140 452620 146192
rect 459376 146140 459428 146192
rect 452568 144644 452620 144696
rect 455052 144644 455104 144696
rect 364248 144168 364300 144220
rect 371240 144168 371292 144220
rect 368388 143828 368440 143880
rect 373632 143828 373684 143880
rect 533436 143488 533488 143540
rect 533988 143488 534040 143540
rect 536104 143488 536156 143540
rect 537300 143488 537352 143540
rect 452568 143284 452620 143336
rect 457628 143284 457680 143336
rect 533988 142196 534040 142248
rect 540336 142196 540388 142248
rect 452568 141924 452620 141976
rect 455144 141924 455196 141976
rect 365444 140768 365496 140820
rect 368388 140768 368440 140820
rect 452568 140632 452620 140684
rect 459284 140632 459336 140684
rect 534724 140156 534776 140208
rect 542912 140156 542964 140208
rect 533344 140088 533396 140140
rect 542728 140088 542780 140140
rect 530584 140020 530636 140072
rect 543096 140020 543148 140072
rect 361764 139340 361816 139392
rect 409604 139340 409656 139392
rect 451556 139340 451608 139392
rect 457536 139340 457588 139392
rect 555424 139340 555476 139392
rect 580172 139340 580224 139392
rect 538864 138524 538916 138576
rect 543004 138524 543056 138576
rect 361396 137980 361448 138032
rect 364248 137980 364300 138032
rect 452568 137844 452620 137896
rect 454960 137844 455012 137896
rect 452568 136484 452620 136536
rect 459100 136484 459152 136536
rect 452568 135124 452620 135176
rect 454776 135124 454828 135176
rect 452568 133764 452620 133816
rect 456616 133764 456668 133816
rect 452476 132404 452528 132456
rect 453764 132404 453816 132456
rect 452568 131044 452620 131096
rect 453948 131044 454000 131096
rect 361488 130160 361540 130212
rect 365444 130160 365496 130212
rect 361580 128256 361632 128308
rect 409512 128256 409564 128308
rect 452568 126896 452620 126948
rect 457444 126896 457496 126948
rect 573364 126896 573416 126948
rect 580172 126896 580224 126948
rect 451924 126012 451976 126064
rect 453672 126012 453724 126064
rect 451924 124720 451976 124772
rect 453856 124720 453908 124772
rect 451924 123224 451976 123276
rect 459468 123224 459520 123276
rect 451740 122204 451792 122256
rect 458732 122204 458784 122256
rect 361580 117240 361632 117292
rect 409420 117240 409472 117292
rect 570604 113092 570656 113144
rect 579804 113092 579856 113144
rect 361580 106224 361632 106276
rect 409328 106224 409380 106276
rect 558184 100648 558236 100700
rect 580172 100648 580224 100700
rect 3700 98608 3752 98660
rect 20904 98608 20956 98660
rect 361764 95140 361816 95192
rect 409236 95140 409288 95192
rect 571984 86912 572036 86964
rect 580172 86912 580224 86964
rect 3608 86232 3660 86284
rect 20904 86232 20956 86284
rect 361764 84124 361816 84176
rect 409144 84124 409196 84176
rect 361764 73108 361816 73160
rect 404084 73108 404136 73160
rect 544384 73108 544436 73160
rect 580172 73108 580224 73160
rect 5080 70388 5132 70440
rect 7564 70320 7616 70372
rect 361764 62024 361816 62076
rect 406844 62024 406896 62076
rect 7564 60732 7616 60784
rect 10048 60664 10100 60716
rect 548524 60664 548576 60716
rect 580172 60664 580224 60716
rect 3516 59984 3568 60036
rect 20904 59984 20956 60036
rect 4804 59304 4856 59356
rect 5816 59304 5868 59356
rect 5816 57196 5868 57248
rect 9772 57196 9824 57248
rect 4896 56516 4948 56568
rect 7288 56516 7340 56568
rect 10048 56516 10100 56568
rect 12348 56516 12400 56568
rect 9772 56176 9824 56228
rect 12624 56176 12676 56228
rect 7288 54612 7340 54664
rect 11980 54612 12032 54664
rect 5540 54476 5592 54528
rect 13820 54476 13872 54528
rect 13820 53116 13872 53168
rect 17868 53116 17920 53168
rect 12348 52980 12400 53032
rect 15200 52980 15252 53032
rect 11980 52436 12032 52488
rect 18788 52368 18840 52420
rect 361764 52368 361816 52420
rect 407856 52368 407908 52420
rect 17868 51416 17920 51468
rect 19524 51416 19576 51468
rect 540612 51076 540664 51128
rect 543740 51076 543792 51128
rect 4988 50328 5040 50380
rect 11704 50328 11756 50380
rect 12624 50328 12676 50380
rect 20628 50328 20680 50380
rect 359556 50056 359608 50108
rect 361212 50056 361264 50108
rect 15200 49716 15252 49768
rect 18052 49648 18104 49700
rect 19524 48220 19576 48272
rect 20720 48220 20772 48272
rect 18052 47880 18104 47932
rect 20812 47880 20864 47932
rect 3148 46996 3200 47048
rect 456156 46996 456208 47048
rect 3516 46860 3568 46912
rect 460296 46860 460348 46912
rect 566464 46860 566516 46912
rect 580172 46860 580224 46912
rect 3608 46792 3660 46844
rect 460388 46792 460440 46844
rect 4068 46724 4120 46776
rect 458916 46724 458968 46776
rect 3240 46656 3292 46708
rect 456340 46656 456392 46708
rect 3332 46588 3384 46640
rect 456248 46588 456300 46640
rect 3976 46520 4028 46572
rect 456432 46520 456484 46572
rect 3792 46452 3844 46504
rect 453488 46452 453540 46504
rect 3884 46384 3936 46436
rect 453396 46384 453448 46436
rect 20904 46316 20956 46368
rect 453580 46316 453632 46368
rect 21364 46248 21416 46300
rect 450820 46248 450872 46300
rect 20812 46180 20864 46232
rect 20720 46112 20772 46164
rect 359832 46180 359884 46232
rect 362316 46180 362368 46232
rect 361396 46112 361448 46164
rect 361304 46044 361356 46096
rect 3424 45500 3476 45552
rect 453304 45500 453356 45552
rect 21456 45432 21508 45484
rect 451004 45432 451056 45484
rect 3516 45364 3568 45416
rect 396724 45364 396776 45416
rect 20720 45296 20772 45348
rect 359832 45296 359884 45348
rect 65524 45228 65576 45280
rect 403716 45228 403768 45280
rect 38384 45160 38436 45212
rect 379244 45160 379296 45212
rect 62028 45092 62080 45144
rect 403900 45092 403952 45144
rect 58440 45024 58492 45076
rect 403624 45024 403676 45076
rect 54944 44956 54996 45008
rect 403808 44956 403860 45008
rect 51356 44888 51408 44940
rect 406476 44888 406528 44940
rect 47860 44820 47912 44872
rect 406752 44820 406804 44872
rect 69112 44752 69164 44804
rect 403992 44752 404044 44804
rect 84476 44684 84528 44736
rect 387524 44684 387576 44736
rect 108120 44616 108172 44668
rect 395804 44616 395856 44668
rect 93952 42712 94004 42764
rect 398196 42712 398248 42764
rect 80888 42644 80940 42696
rect 387432 42644 387484 42696
rect 90364 42576 90416 42628
rect 398104 42576 398156 42628
rect 86868 42508 86920 42560
rect 398380 42508 398432 42560
rect 83280 42440 83332 42492
rect 401324 42440 401376 42492
rect 79692 42372 79744 42424
rect 400956 42372 401008 42424
rect 76196 42304 76248 42356
rect 401048 42304 401100 42356
rect 72608 42236 72660 42288
rect 401140 42236 401192 42288
rect 111616 42168 111668 42220
rect 460204 42168 460256 42220
rect 101036 42100 101088 42152
rect 454684 42100 454736 42152
rect 12348 42032 12400 42084
rect 401232 42032 401284 42084
rect 97448 41964 97500 42016
rect 398288 41964 398340 42016
rect 106924 41896 106976 41948
rect 370964 41896 371016 41948
rect 475384 41352 475436 41404
rect 536840 41352 536892 41404
rect 102232 39992 102284 40044
rect 384580 39992 384632 40044
rect 71504 39924 71556 39976
rect 373540 39924 373592 39976
rect 59636 39856 59688 39908
rect 390284 39856 390336 39908
rect 118792 39788 118844 39840
rect 450636 39788 450688 39840
rect 56048 39720 56100 39772
rect 390192 39720 390244 39772
rect 48964 39652 49016 39704
rect 392860 39652 392912 39704
rect 104532 39584 104584 39636
rect 451096 39584 451148 39636
rect 44272 39516 44324 39568
rect 393044 39516 393096 39568
rect 40684 39448 40736 39500
rect 392952 39448 393004 39500
rect 4068 39380 4120 39432
rect 392768 39380 392820 39432
rect 26516 39312 26568 39364
rect 450912 39312 450964 39364
rect 115204 39244 115256 39296
rect 395620 39244 395672 39296
rect 122288 39176 122340 39228
rect 395712 39176 395764 39228
rect 105728 37204 105780 37256
rect 384488 37204 384540 37256
rect 98644 37136 98696 37188
rect 384396 37136 384448 37188
rect 95148 37068 95200 37120
rect 384304 37068 384356 37120
rect 91560 37000 91612 37052
rect 387156 37000 387208 37052
rect 87972 36932 88024 36984
rect 387248 36932 387300 36984
rect 77392 36864 77444 36916
rect 387340 36864 387392 36916
rect 73804 36796 73856 36848
rect 390008 36796 390060 36848
rect 70308 36728 70360 36780
rect 390100 36728 390152 36780
rect 66720 36660 66772 36712
rect 389916 36660 389968 36712
rect 63224 36592 63276 36644
rect 389824 36592 389876 36644
rect 28908 36524 28960 36576
rect 368204 36524 368256 36576
rect 109316 36456 109368 36508
rect 381728 36456 381780 36508
rect 112812 36388 112864 36440
rect 382004 36388 382056 36440
rect 119896 34416 119948 34468
rect 381544 34416 381596 34468
rect 116400 34348 116452 34400
rect 381820 34348 381872 34400
rect 60832 34280 60884 34332
rect 376484 34280 376536 34332
rect 57244 34212 57296 34264
rect 376392 34212 376444 34264
rect 50160 34144 50212 34196
rect 376116 34144 376168 34196
rect 45468 34076 45520 34128
rect 376208 34076 376260 34128
rect 41880 34008 41932 34060
rect 376300 34008 376352 34060
rect 34796 33940 34848 33992
rect 379060 33940 379112 33992
rect 31300 33872 31352 33924
rect 379152 33872 379204 33924
rect 23020 33804 23072 33856
rect 378968 33804 379020 33856
rect 18236 33736 18288 33788
rect 381912 33736 381964 33788
rect 123484 33668 123536 33720
rect 378784 33668 378836 33720
rect 111064 33600 111116 33652
rect 365352 33600 365404 33652
rect 2872 33056 2924 33108
rect 400864 33056 400916 33108
rect 569224 33056 569276 33108
rect 580172 33056 580224 33108
rect 117596 31696 117648 31748
rect 367744 31696 367796 31748
rect 114008 31628 114060 31680
rect 368020 31628 368072 31680
rect 99840 31560 99892 31612
rect 370780 31560 370832 31612
rect 96252 31492 96304 31544
rect 370872 31492 370924 31544
rect 89168 31424 89220 31476
rect 370504 31424 370556 31476
rect 78588 31356 78640 31408
rect 370596 31356 370648 31408
rect 75000 31288 75052 31340
rect 373264 31288 373316 31340
rect 67916 31220 67968 31272
rect 373356 31220 373408 31272
rect 64328 31152 64380 31204
rect 373448 31152 373500 31204
rect 19432 31084 19484 31136
rect 368112 31084 368164 31136
rect 14740 31016 14792 31068
rect 370688 31016 370740 31068
rect 121092 30948 121144 31000
rect 367928 30948 367980 31000
rect 124680 30880 124732 30932
rect 367836 30880 367888 30932
rect 46664 28432 46716 28484
rect 365260 28432 365312 28484
rect 43076 28364 43128 28416
rect 365076 28364 365128 28416
rect 35992 28296 36044 28348
rect 364984 28296 365036 28348
rect 32404 28228 32456 28280
rect 365168 28228 365220 28280
rect 3424 20612 3476 20664
rect 381636 20612 381688 20664
rect 574744 20612 574796 20664
rect 579988 20612 580040 20664
rect 3424 6808 3476 6860
rect 395436 6808 395488 6860
rect 562324 6808 562376 6860
rect 580172 6808 580224 6860
rect 85672 4088 85724 4140
rect 363696 4088 363748 4140
rect 53748 4020 53800 4072
rect 361120 4020 361172 4072
rect 39580 3952 39632 4004
rect 360844 3952 360896 4004
rect 33600 3884 33652 3936
rect 359464 3884 359516 3936
rect 27712 3816 27764 3868
rect 378876 3816 378928 3868
rect 37188 3748 37240 3800
rect 392676 3748 392728 3800
rect 82084 3680 82136 3732
rect 450544 3680 450596 3732
rect 21824 3612 21876 3664
rect 395528 3612 395580 3664
rect 24216 3544 24268 3596
rect 407764 3544 407816 3596
rect 52552 3476 52604 3528
rect 456064 3476 456116 3528
rect 17040 3408 17092 3460
rect 450728 3408 450780 3460
rect 92756 3340 92808 3392
rect 362224 3340 362276 3392
rect 103336 3272 103388 3324
rect 361028 3272 361080 3324
rect 110512 3204 110564 3256
rect 360936 3204 360988 3256
rect 6460 3136 6512 3188
rect 111064 3136 111116 3188
rect 30104 2048 30156 2100
rect 395344 2048 395396 2100
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 8128 700330 8156 703520
rect 8116 700324 8168 700330
rect 8116 700266 8168 700272
rect 24320 686497 24348 703520
rect 40512 700398 40540 703520
rect 40500 700392 40552 700398
rect 40500 700334 40552 700340
rect 24306 686488 24362 686497
rect 24306 686423 24362 686432
rect 72988 685166 73016 703520
rect 89180 685234 89208 703520
rect 105464 700466 105492 703520
rect 137848 700534 137876 703520
rect 154132 700670 154160 703520
rect 154120 700664 154172 700670
rect 154120 700606 154172 700612
rect 170324 700602 170352 703520
rect 170312 700596 170364 700602
rect 170312 700538 170364 700544
rect 137836 700528 137888 700534
rect 137836 700470 137888 700476
rect 105452 700460 105504 700466
rect 105452 700402 105504 700408
rect 202800 685302 202828 703520
rect 218992 700738 219020 703520
rect 235184 700806 235212 703520
rect 267660 700874 267688 703520
rect 267648 700868 267700 700874
rect 267648 700810 267700 700816
rect 235172 700800 235224 700806
rect 235172 700742 235224 700748
rect 218980 700732 219032 700738
rect 218980 700674 219032 700680
rect 283852 686526 283880 703520
rect 300136 700369 300164 703520
rect 300122 700360 300178 700369
rect 300122 700295 300178 700304
rect 283840 686520 283892 686526
rect 283840 686462 283892 686468
rect 332520 685370 332548 703520
rect 348804 686594 348832 703520
rect 348792 686588 348844 686594
rect 348792 686530 348844 686536
rect 332508 685364 332560 685370
rect 332508 685306 332560 685312
rect 202788 685296 202840 685302
rect 202788 685238 202840 685244
rect 89168 685228 89220 685234
rect 89168 685170 89220 685176
rect 72976 685160 73028 685166
rect 72976 685102 73028 685108
rect 19984 684616 20036 684622
rect 19984 684558 20036 684564
rect 3792 684548 3844 684554
rect 3792 684490 3844 684496
rect 3516 683596 3568 683602
rect 3516 683538 3568 683544
rect 3424 683460 3476 683466
rect 3424 683402 3476 683408
rect 3332 683188 3384 683194
rect 3332 683130 3384 683136
rect 3240 682712 3292 682718
rect 3240 682654 3292 682660
rect 3148 658232 3200 658238
rect 3146 658200 3148 658209
rect 3200 658200 3202 658209
rect 3146 658135 3202 658144
rect 3252 580009 3280 682654
rect 3238 580000 3294 580009
rect 3238 579935 3294 579944
rect 3344 566953 3372 683130
rect 3330 566944 3386 566953
rect 3330 566879 3386 566888
rect 3436 449585 3464 683402
rect 3528 462641 3556 683538
rect 3700 683528 3752 683534
rect 3700 683470 3752 683476
rect 3608 683324 3660 683330
rect 3608 683266 3660 683272
rect 3620 632097 3648 683266
rect 3606 632088 3662 632097
rect 3606 632023 3662 632032
rect 3608 631372 3660 631378
rect 3608 631314 3660 631320
rect 3514 462632 3570 462641
rect 3514 462567 3570 462576
rect 3422 449576 3478 449585
rect 3422 449511 3478 449520
rect 3620 423609 3648 631314
rect 3712 475697 3740 683470
rect 3804 501809 3832 684490
rect 18328 683800 18380 683806
rect 18328 683742 18380 683748
rect 4068 683664 4120 683670
rect 4068 683606 4120 683612
rect 3884 683392 3936 683398
rect 3884 683334 3936 683340
rect 3896 514865 3924 683334
rect 3976 683256 4028 683262
rect 3976 683198 4028 683204
rect 3988 527921 4016 683198
rect 4080 553897 4108 683606
rect 18340 680406 18368 683742
rect 17224 680400 17276 680406
rect 17224 680342 17276 680348
rect 18328 680400 18380 680406
rect 18328 680342 18380 680348
rect 17236 661094 17264 680342
rect 17224 661088 17276 661094
rect 17224 661030 17276 661036
rect 14188 661020 14240 661026
rect 14188 660962 14240 660968
rect 14200 656674 14228 660962
rect 19996 658238 20024 684558
rect 359464 683800 359516 683806
rect 359464 683742 359516 683748
rect 21364 683732 21416 683738
rect 21364 683674 21416 683680
rect 19984 658232 20036 658238
rect 19984 658174 20036 658180
rect 11704 656668 11756 656674
rect 11704 656610 11756 656616
rect 14188 656668 14240 656674
rect 14188 656610 14240 656616
rect 11716 645862 11744 656610
rect 10600 645856 10652 645862
rect 10600 645798 10652 645804
rect 11704 645856 11756 645862
rect 11704 645798 11756 645804
rect 10612 643754 10640 645798
rect 5540 643748 5592 643754
rect 5540 643690 5592 643696
rect 10600 643748 10652 643754
rect 10600 643690 10652 643696
rect 5552 640354 5580 643690
rect 4804 640348 4856 640354
rect 4804 640290 4856 640296
rect 5540 640348 5592 640354
rect 5540 640290 5592 640296
rect 4066 553888 4122 553897
rect 4066 553823 4122 553832
rect 3974 527912 4030 527921
rect 3974 527847 4030 527856
rect 3882 514856 3938 514865
rect 4816 514826 4844 640290
rect 21376 634814 21404 683674
rect 359476 672110 359504 683742
rect 362222 679008 362278 679017
rect 362222 678943 362278 678952
rect 359464 672104 359516 672110
rect 359464 672046 359516 672052
rect 360844 672104 360896 672110
rect 360844 672046 360896 672052
rect 20916 634786 21404 634814
rect 20916 631378 20944 634786
rect 20904 631372 20956 631378
rect 20904 631314 20956 631320
rect 360856 598262 360884 672046
rect 361762 667992 361818 668001
rect 361762 667927 361764 667936
rect 361816 667927 361818 667936
rect 361764 667898 361816 667904
rect 361762 656976 361818 656985
rect 361762 656911 361764 656920
rect 361816 656911 361818 656920
rect 361764 656882 361816 656888
rect 361762 645960 361818 645969
rect 361762 645895 361764 645904
rect 361816 645895 361818 645904
rect 361764 645866 361816 645872
rect 361578 634944 361634 634953
rect 361578 634879 361634 634888
rect 361592 634846 361620 634879
rect 361580 634840 361632 634846
rect 361580 634782 361632 634788
rect 361578 623928 361634 623937
rect 361578 623863 361634 623872
rect 361592 623830 361620 623863
rect 361580 623824 361632 623830
rect 361580 623766 361632 623772
rect 361578 612912 361634 612921
rect 361578 612847 361580 612856
rect 361632 612847 361634 612856
rect 361580 612818 361632 612824
rect 361762 601896 361818 601905
rect 361762 601831 361818 601840
rect 361776 601730 361804 601831
rect 361764 601724 361816 601730
rect 361764 601666 361816 601672
rect 360844 598256 360896 598262
rect 360844 598198 360896 598204
rect 361578 590880 361634 590889
rect 361578 590815 361580 590824
rect 361632 590815 361634 590824
rect 361580 590786 361632 590792
rect 361762 579864 361818 579873
rect 361762 579799 361818 579808
rect 361776 579698 361804 579799
rect 361764 579692 361816 579698
rect 361764 579634 361816 579640
rect 361578 568848 361634 568857
rect 361578 568783 361580 568792
rect 361632 568783 361634 568792
rect 361580 568754 361632 568760
rect 361670 557832 361726 557841
rect 361670 557767 361726 557776
rect 361684 557598 361712 557767
rect 361672 557592 361724 557598
rect 361672 557534 361724 557540
rect 361762 546816 361818 546825
rect 361762 546751 361818 546760
rect 361776 546514 361804 546751
rect 361764 546508 361816 546514
rect 361764 546450 361816 546456
rect 361762 535800 361818 535809
rect 361762 535735 361818 535744
rect 361776 535498 361804 535735
rect 361764 535492 361816 535498
rect 361764 535434 361816 535440
rect 361762 524784 361818 524793
rect 361762 524719 361818 524728
rect 361776 524482 361804 524719
rect 361764 524476 361816 524482
rect 361764 524418 361816 524424
rect 3882 514791 3938 514800
rect 3976 514820 4028 514826
rect 3976 514762 4028 514768
rect 4804 514820 4856 514826
rect 4804 514762 4856 514768
rect 3790 501800 3846 501809
rect 3790 501735 3846 501744
rect 3698 475688 3754 475697
rect 3698 475623 3754 475632
rect 3606 423600 3662 423609
rect 3606 423535 3662 423544
rect 3988 410553 4016 514762
rect 361762 513768 361818 513777
rect 361762 513703 361818 513712
rect 361776 513398 361804 513703
rect 361764 513392 361816 513398
rect 361764 513334 361816 513340
rect 361762 502752 361818 502761
rect 361762 502687 361818 502696
rect 361776 502382 361804 502687
rect 361764 502376 361816 502382
rect 361764 502318 361816 502324
rect 361762 491736 361818 491745
rect 361762 491671 361818 491680
rect 361776 491366 361804 491671
rect 361764 491360 361816 491366
rect 361764 491302 361816 491308
rect 361762 480720 361818 480729
rect 361762 480655 361818 480664
rect 361776 480282 361804 480655
rect 361764 480276 361816 480282
rect 361764 480218 361816 480224
rect 361762 469704 361818 469713
rect 361762 469639 361818 469648
rect 361776 469266 361804 469639
rect 361764 469260 361816 469266
rect 361764 469202 361816 469208
rect 361762 458688 361818 458697
rect 361762 458623 361818 458632
rect 361776 458250 361804 458623
rect 361764 458244 361816 458250
rect 361764 458186 361816 458192
rect 361762 447672 361818 447681
rect 361762 447607 361818 447616
rect 361776 447166 361804 447607
rect 361764 447160 361816 447166
rect 361764 447102 361816 447108
rect 361762 436656 361818 436665
rect 361762 436591 361818 436600
rect 361776 436150 361804 436591
rect 361764 436144 361816 436150
rect 361764 436086 361816 436092
rect 361762 425640 361818 425649
rect 361762 425575 361818 425584
rect 361776 425134 361804 425575
rect 361764 425128 361816 425134
rect 361764 425070 361816 425076
rect 361578 414624 361634 414633
rect 361578 414559 361634 414568
rect 361592 414050 361620 414559
rect 361580 414044 361632 414050
rect 361580 413986 361632 413992
rect 3974 410544 4030 410553
rect 3974 410479 4030 410488
rect 361578 403608 361634 403617
rect 361578 403543 361634 403552
rect 361592 403034 361620 403543
rect 361580 403028 361632 403034
rect 361580 402970 361632 402976
rect 3790 397488 3846 397497
rect 3790 397423 3846 397432
rect 3514 358456 3570 358465
rect 3514 358391 3570 358400
rect 3422 345400 3478 345409
rect 3422 345335 3478 345344
rect 3436 292602 3464 345335
rect 3528 307766 3556 358391
rect 3516 307760 3568 307766
rect 3516 307702 3568 307708
rect 3698 306232 3754 306241
rect 3698 306167 3754 306176
rect 3606 293176 3662 293185
rect 3606 293111 3662 293120
rect 3424 292596 3476 292602
rect 3424 292538 3476 292544
rect 3514 267200 3570 267209
rect 3514 267135 3570 267144
rect 3422 254144 3478 254153
rect 3422 254079 3478 254088
rect 3330 162888 3386 162897
rect 3330 162823 3386 162832
rect 3238 149832 3294 149841
rect 3238 149767 3294 149776
rect 3146 98696 3202 98705
rect 3146 98631 3202 98640
rect 3160 47054 3188 98631
rect 3148 47048 3200 47054
rect 3148 46990 3200 46996
rect 3252 46714 3280 149767
rect 3240 46708 3292 46714
rect 3240 46650 3292 46656
rect 3344 46646 3372 162823
rect 3332 46640 3384 46646
rect 3332 46582 3384 46588
rect 3436 45558 3464 254079
rect 3528 60042 3556 267135
rect 3620 86290 3648 293111
rect 3712 98666 3740 306167
rect 3804 243982 3832 397423
rect 361578 392592 361634 392601
rect 361578 392527 361634 392536
rect 361592 392018 361620 392527
rect 361580 392012 361632 392018
rect 361580 391954 361632 391960
rect 362236 383654 362264 678943
rect 363604 612876 363656 612882
rect 363604 612818 363656 612824
rect 362224 383648 362276 383654
rect 362224 383590 362276 383596
rect 361578 381576 361634 381585
rect 361578 381511 361634 381520
rect 361592 380934 361620 381511
rect 361580 380928 361632 380934
rect 361580 380870 361632 380876
rect 363616 380866 363644 612818
rect 363696 590844 363748 590850
rect 363696 590786 363748 590792
rect 363604 380860 363656 380866
rect 363604 380802 363656 380808
rect 363708 379506 363736 590786
rect 363788 568812 363840 568818
rect 363788 568754 363840 568760
rect 363696 379500 363748 379506
rect 363696 379442 363748 379448
rect 363800 378146 363828 568754
rect 363788 378140 363840 378146
rect 363788 378082 363840 378088
rect 3882 371376 3938 371385
rect 3882 371311 3938 371320
rect 3792 243976 3844 243982
rect 3792 243918 3844 243924
rect 3790 241088 3846 241097
rect 3790 241023 3846 241032
rect 3700 98660 3752 98666
rect 3700 98602 3752 98608
rect 3608 86284 3660 86290
rect 3608 86226 3660 86232
rect 3606 71632 3662 71641
rect 3606 71567 3662 71576
rect 3516 60036 3568 60042
rect 3516 59978 3568 59984
rect 3514 58576 3570 58585
rect 3514 58511 3570 58520
rect 3528 46918 3556 58511
rect 3516 46912 3568 46918
rect 3516 46854 3568 46860
rect 3620 46850 3648 71567
rect 3608 46844 3660 46850
rect 3608 46786 3660 46792
rect 3804 46510 3832 241023
rect 3896 222154 3924 371311
rect 361578 370560 361634 370569
rect 361578 370495 361634 370504
rect 361592 369918 361620 370495
rect 361580 369912 361632 369918
rect 361580 369854 361632 369860
rect 362222 359544 362278 359553
rect 362222 359479 362278 359488
rect 361762 348528 361818 348537
rect 361762 348463 361818 348472
rect 361776 347818 361804 348463
rect 361764 347812 361816 347818
rect 361764 347754 361816 347760
rect 362236 347750 362264 359479
rect 364996 349858 365024 703520
rect 378876 667956 378928 667962
rect 378876 667898 378928 667904
rect 376024 656940 376076 656946
rect 376024 656882 376076 656888
rect 374644 645924 374696 645930
rect 374644 645866 374696 645872
rect 371884 623824 371936 623830
rect 371884 623766 371936 623772
rect 370504 601724 370556 601730
rect 370504 601666 370556 601672
rect 367744 598256 367796 598262
rect 367744 598198 367796 598204
rect 367756 587858 367784 598198
rect 367744 587852 367796 587858
rect 367744 587794 367796 587800
rect 368020 579692 368072 579698
rect 368020 579634 368072 579640
rect 367744 386504 367796 386510
rect 367744 386446 367796 386452
rect 364984 349852 365036 349858
rect 364984 349794 365036 349800
rect 362224 347744 362276 347750
rect 362224 347686 362276 347692
rect 361764 340944 361816 340950
rect 361764 340886 361816 340892
rect 361776 337521 361804 340886
rect 361762 337512 361818 337521
rect 361762 337447 361818 337456
rect 362224 336048 362276 336054
rect 362224 335990 362276 335996
rect 362236 326505 362264 335990
rect 363788 334008 363840 334014
rect 363788 333950 363840 333956
rect 362222 326496 362278 326505
rect 362222 326431 362278 326440
rect 3974 319288 4030 319297
rect 3974 319223 4030 319232
rect 3988 253978 4016 319223
rect 361764 315988 361816 315994
rect 361764 315930 361816 315936
rect 361776 315489 361804 315930
rect 361762 315480 361818 315489
rect 361762 315415 361818 315424
rect 4804 307760 4856 307766
rect 4804 307702 4856 307708
rect 3976 253972 4028 253978
rect 3976 253914 4028 253920
rect 3884 222148 3936 222154
rect 3884 222090 3936 222096
rect 3882 214976 3938 214985
rect 3882 214911 3938 214920
rect 3792 46504 3844 46510
rect 3792 46446 3844 46452
rect 3896 46442 3924 214911
rect 3974 201920 4030 201929
rect 3974 201855 4030 201864
rect 3988 46578 4016 201855
rect 4066 188864 4122 188873
rect 4066 188799 4122 188808
rect 4080 46782 4108 188799
rect 4816 59362 4844 307702
rect 363604 305720 363656 305726
rect 363604 305662 363656 305668
rect 360844 305652 360896 305658
rect 360844 305594 360896 305600
rect 4896 292596 4948 292602
rect 4896 292538 4948 292544
rect 4804 59356 4856 59362
rect 4804 59298 4856 59304
rect 4908 56574 4936 292538
rect 359464 269816 359516 269822
rect 359464 269758 359516 269764
rect 5080 253972 5132 253978
rect 5080 253914 5132 253920
rect 4988 243976 5040 243982
rect 4988 243918 5040 243924
rect 4896 56568 4948 56574
rect 4896 56510 4948 56516
rect 5000 50386 5028 243918
rect 5092 70446 5120 253914
rect 5172 222148 5224 222154
rect 5172 222090 5224 222096
rect 5080 70440 5132 70446
rect 5080 70382 5132 70388
rect 5184 55214 5212 222090
rect 20904 98660 20956 98666
rect 20904 98602 20956 98608
rect 20916 93854 20944 98602
rect 20916 93826 21404 93854
rect 20904 86284 20956 86290
rect 20904 86226 20956 86232
rect 20916 77217 20944 86226
rect 21376 77294 21404 93826
rect 21284 77266 21404 77294
rect 20902 77208 20958 77217
rect 20902 77143 20958 77152
rect 7564 70372 7616 70378
rect 7564 70314 7616 70320
rect 7576 60790 7604 70314
rect 21284 67634 21312 77266
rect 21454 77208 21510 77217
rect 21454 77143 21510 77152
rect 21284 67606 21404 67634
rect 7564 60784 7616 60790
rect 7564 60726 7616 60732
rect 10048 60716 10100 60722
rect 10048 60658 10100 60664
rect 5816 59356 5868 59362
rect 5816 59298 5868 59304
rect 5828 57254 5856 59298
rect 5816 57248 5868 57254
rect 5816 57190 5868 57196
rect 9772 57248 9824 57254
rect 9772 57190 9824 57196
rect 7288 56568 7340 56574
rect 7288 56510 7340 56516
rect 5184 55186 5580 55214
rect 5552 54534 5580 55186
rect 7300 54670 7328 56510
rect 9784 56234 9812 57190
rect 10060 56574 10088 60658
rect 20904 60036 20956 60042
rect 20904 59978 20956 59984
rect 10048 56568 10100 56574
rect 10048 56510 10100 56516
rect 12348 56568 12400 56574
rect 12348 56510 12400 56516
rect 9772 56228 9824 56234
rect 9772 56170 9824 56176
rect 7288 54664 7340 54670
rect 7288 54606 7340 54612
rect 11980 54664 12032 54670
rect 11980 54606 12032 54612
rect 5540 54528 5592 54534
rect 5540 54470 5592 54476
rect 11992 52494 12020 54606
rect 12360 53038 12388 56510
rect 12624 56228 12676 56234
rect 12624 56170 12676 56176
rect 12348 53032 12400 53038
rect 12348 52974 12400 52980
rect 11980 52488 12032 52494
rect 11980 52430 12032 52436
rect 12636 50386 12664 56170
rect 13820 54528 13872 54534
rect 13820 54470 13872 54476
rect 13832 53174 13860 54470
rect 13820 53168 13872 53174
rect 13820 53110 13872 53116
rect 17868 53168 17920 53174
rect 17868 53110 17920 53116
rect 15200 53032 15252 53038
rect 15200 52974 15252 52980
rect 4988 50380 5040 50386
rect 4988 50322 5040 50328
rect 11704 50380 11756 50386
rect 11704 50322 11756 50328
rect 12624 50380 12676 50386
rect 12624 50322 12676 50328
rect 11716 48929 11744 50322
rect 15212 49774 15240 52974
rect 17880 51474 17908 53110
rect 18788 52420 18840 52426
rect 18788 52362 18840 52368
rect 17868 51468 17920 51474
rect 17868 51410 17920 51416
rect 15200 49768 15252 49774
rect 15200 49710 15252 49716
rect 18052 49700 18104 49706
rect 18052 49642 18104 49648
rect 11702 48920 11758 48929
rect 11702 48855 11758 48864
rect 18064 47938 18092 49642
rect 18800 49337 18828 52362
rect 19524 51468 19576 51474
rect 19524 51410 19576 51416
rect 18786 49328 18842 49337
rect 18786 49263 18842 49272
rect 19536 48278 19564 51410
rect 20628 50380 20680 50386
rect 20628 50322 20680 50328
rect 19524 48272 19576 48278
rect 19524 48214 19576 48220
rect 18052 47932 18104 47938
rect 18052 47874 18104 47880
rect 4068 46776 4120 46782
rect 4068 46718 4120 46724
rect 3976 46572 4028 46578
rect 3976 46514 4028 46520
rect 3884 46436 3936 46442
rect 3884 46378 3936 46384
rect 3424 45552 3476 45558
rect 20640 45554 20668 50322
rect 20720 48272 20772 48278
rect 20720 48214 20772 48220
rect 20732 46170 20760 48214
rect 20812 47932 20864 47938
rect 20812 47874 20864 47880
rect 20824 46238 20852 47874
rect 20916 46374 20944 59978
rect 20904 46368 20956 46374
rect 20904 46310 20956 46316
rect 21376 46306 21404 67606
rect 21364 46300 21416 46306
rect 21364 46242 21416 46248
rect 20812 46232 20864 46238
rect 20812 46174 20864 46180
rect 20720 46164 20772 46170
rect 20720 46106 20772 46112
rect 3424 45494 3476 45500
rect 3514 45520 3570 45529
rect 20640 45526 20760 45554
rect 3514 45455 3570 45464
rect 3528 45422 3556 45455
rect 3516 45416 3568 45422
rect 3516 45358 3568 45364
rect 20732 45354 20760 45526
rect 21468 45490 21496 77143
rect 21456 45484 21508 45490
rect 21456 45426 21508 45432
rect 20720 45348 20772 45354
rect 20720 45290 20772 45296
rect 65524 45280 65576 45286
rect 65524 45222 65576 45228
rect 38384 45212 38436 45218
rect 38384 45154 38436 45160
rect 7654 44840 7710 44849
rect 7654 44775 7710 44784
rect 4068 39432 4120 39438
rect 4068 39374 4120 39380
rect 2872 33108 2924 33114
rect 2872 33050 2924 33056
rect 2884 32473 2912 33050
rect 2870 32464 2926 32473
rect 2870 32399 2926 32408
rect 3424 20664 3476 20670
rect 3424 20606 3476 20612
rect 3436 19417 3464 20606
rect 3422 19408 3478 19417
rect 3422 19343 3478 19352
rect 3424 6860 3476 6866
rect 3424 6802 3476 6808
rect 3436 6497 3464 6802
rect 3422 6488 3478 6497
rect 3422 6423 3478 6432
rect 2870 3632 2926 3641
rect 2870 3567 2926 3576
rect 1674 3496 1730 3505
rect 1674 3431 1730 3440
rect 570 3360 626 3369
rect 570 3295 626 3304
rect 584 480 612 3295
rect 1688 480 1716 3431
rect 2884 480 2912 3567
rect 4080 480 4108 39374
rect 5262 3224 5318 3233
rect 5262 3159 5318 3168
rect 6460 3188 6512 3194
rect 5276 480 5304 3159
rect 6460 3130 6512 3136
rect 6472 480 6500 3130
rect 7668 480 7696 44775
rect 12348 42084 12400 42090
rect 12348 42026 12400 42032
rect 9954 4040 10010 4049
rect 9954 3975 10010 3984
rect 8758 3768 8814 3777
rect 8758 3703 8814 3712
rect 8772 480 8800 3703
rect 9968 480 9996 3975
rect 12360 480 12388 42026
rect 26516 39364 26568 39370
rect 26516 39306 26568 39312
rect 23020 33856 23072 33862
rect 23020 33798 23072 33804
rect 18236 33788 18288 33794
rect 18236 33730 18288 33736
rect 14740 31068 14792 31074
rect 14740 31010 14792 31016
rect 13542 3904 13598 3913
rect 13542 3839 13598 3848
rect 13556 480 13584 3839
rect 14752 480 14780 31010
rect 17040 3460 17092 3466
rect 17040 3402 17092 3408
rect 17052 480 17080 3402
rect 18248 480 18276 33730
rect 19432 31136 19484 31142
rect 19432 31078 19484 31084
rect 19444 480 19472 31078
rect 21824 3664 21876 3670
rect 21824 3606 21876 3612
rect 21836 480 21864 3606
rect 23032 480 23060 33798
rect 24216 3596 24268 3602
rect 24216 3538 24268 3544
rect 24228 480 24256 3538
rect 26528 480 26556 39306
rect 28908 36576 28960 36582
rect 28908 36518 28960 36524
rect 27712 3868 27764 3874
rect 27712 3810 27764 3816
rect 27724 480 27752 3810
rect 28920 480 28948 36518
rect 34796 33992 34848 33998
rect 34796 33934 34848 33940
rect 31300 33924 31352 33930
rect 31300 33866 31352 33872
rect 30104 2100 30156 2106
rect 30104 2042 30156 2048
rect 30116 480 30144 2042
rect 31312 480 31340 33866
rect 32404 28280 32456 28286
rect 32404 28222 32456 28228
rect 32416 480 32444 28222
rect 33600 3936 33652 3942
rect 33600 3878 33652 3884
rect 33612 480 33640 3878
rect 34808 480 34836 33934
rect 35992 28348 36044 28354
rect 35992 28290 36044 28296
rect 36004 480 36032 28290
rect 37188 3800 37240 3806
rect 37188 3742 37240 3748
rect 37200 480 37228 3742
rect 38396 480 38424 45154
rect 62028 45144 62080 45150
rect 62028 45086 62080 45092
rect 58440 45076 58492 45082
rect 58440 45018 58492 45024
rect 54944 45008 54996 45014
rect 54944 44950 54996 44956
rect 51356 44940 51408 44946
rect 51356 44882 51408 44888
rect 47860 44872 47912 44878
rect 47860 44814 47912 44820
rect 44272 39568 44324 39574
rect 44272 39510 44324 39516
rect 40684 39500 40736 39506
rect 40684 39442 40736 39448
rect 39580 4004 39632 4010
rect 39580 3946 39632 3952
rect 39592 480 39620 3946
rect 40696 480 40724 39442
rect 41880 34060 41932 34066
rect 41880 34002 41932 34008
rect 41892 480 41920 34002
rect 43076 28416 43128 28422
rect 43076 28358 43128 28364
rect 43088 480 43116 28358
rect 44284 480 44312 39510
rect 45468 34128 45520 34134
rect 45468 34070 45520 34076
rect 45480 480 45508 34070
rect 46664 28484 46716 28490
rect 46664 28426 46716 28432
rect 46676 480 46704 28426
rect 47872 480 47900 44814
rect 48964 39704 49016 39710
rect 48964 39646 49016 39652
rect 48976 480 49004 39646
rect 50160 34196 50212 34202
rect 50160 34138 50212 34144
rect 50172 480 50200 34138
rect 51368 480 51396 44882
rect 53748 4072 53800 4078
rect 53748 4014 53800 4020
rect 52552 3528 52604 3534
rect 52552 3470 52604 3476
rect 52564 480 52592 3470
rect 53760 480 53788 4014
rect 54956 480 54984 44950
rect 56048 39772 56100 39778
rect 56048 39714 56100 39720
rect 56060 480 56088 39714
rect 57244 34264 57296 34270
rect 57244 34206 57296 34212
rect 57256 480 57284 34206
rect 58452 480 58480 45018
rect 59636 39908 59688 39914
rect 59636 39850 59688 39856
rect 59648 480 59676 39850
rect 60832 34332 60884 34338
rect 60832 34274 60884 34280
rect 60844 480 60872 34274
rect 62040 480 62068 45086
rect 63224 36644 63276 36650
rect 63224 36586 63276 36592
rect 63236 480 63264 36586
rect 64328 31204 64380 31210
rect 64328 31146 64380 31152
rect 64340 480 64368 31146
rect 65536 480 65564 45222
rect 69112 44804 69164 44810
rect 69112 44746 69164 44752
rect 66720 36712 66772 36718
rect 66720 36654 66772 36660
rect 66732 480 66760 36654
rect 67916 31272 67968 31278
rect 67916 31214 67968 31220
rect 67928 480 67956 31214
rect 69124 480 69152 44746
rect 84476 44736 84528 44742
rect 84476 44678 84528 44684
rect 80888 42696 80940 42702
rect 80888 42638 80940 42644
rect 79692 42424 79744 42430
rect 79692 42366 79744 42372
rect 76196 42356 76248 42362
rect 76196 42298 76248 42304
rect 72608 42288 72660 42294
rect 72608 42230 72660 42236
rect 71504 39976 71556 39982
rect 71504 39918 71556 39924
rect 70308 36780 70360 36786
rect 70308 36722 70360 36728
rect 70320 480 70348 36722
rect 71516 480 71544 39918
rect 72620 480 72648 42230
rect 73804 36848 73856 36854
rect 73804 36790 73856 36796
rect 73816 480 73844 36790
rect 75000 31340 75052 31346
rect 75000 31282 75052 31288
rect 75012 480 75040 31282
rect 76208 480 76236 42298
rect 77392 36916 77444 36922
rect 77392 36858 77444 36864
rect 77404 480 77432 36858
rect 78588 31408 78640 31414
rect 78588 31350 78640 31356
rect 78600 480 78628 31350
rect 79704 480 79732 42366
rect 80900 480 80928 42638
rect 83280 42492 83332 42498
rect 83280 42434 83332 42440
rect 82084 3732 82136 3738
rect 82084 3674 82136 3680
rect 82096 480 82124 3674
rect 83292 480 83320 42434
rect 84488 480 84516 44678
rect 108120 44668 108172 44674
rect 108120 44610 108172 44616
rect 93952 42764 94004 42770
rect 93952 42706 94004 42712
rect 90364 42628 90416 42634
rect 90364 42570 90416 42576
rect 86868 42560 86920 42566
rect 86868 42502 86920 42508
rect 85672 4140 85724 4146
rect 85672 4082 85724 4088
rect 85684 480 85712 4082
rect 86880 480 86908 42502
rect 87972 36984 88024 36990
rect 87972 36926 88024 36932
rect 87984 480 88012 36926
rect 89168 31476 89220 31482
rect 89168 31418 89220 31424
rect 89180 480 89208 31418
rect 90376 480 90404 42570
rect 91560 37052 91612 37058
rect 91560 36994 91612 37000
rect 91572 480 91600 36994
rect 92756 3392 92808 3398
rect 92756 3334 92808 3340
rect 92768 480 92796 3334
rect 93964 480 93992 42706
rect 101036 42152 101088 42158
rect 101036 42094 101088 42100
rect 97448 42016 97500 42022
rect 97448 41958 97500 41964
rect 95148 37120 95200 37126
rect 95148 37062 95200 37068
rect 95160 480 95188 37062
rect 96252 31544 96304 31550
rect 96252 31486 96304 31492
rect 96264 480 96292 31486
rect 97460 480 97488 41958
rect 98644 37188 98696 37194
rect 98644 37130 98696 37136
rect 98656 480 98684 37130
rect 99840 31612 99892 31618
rect 99840 31554 99892 31560
rect 99852 480 99880 31554
rect 101048 480 101076 42094
rect 106924 41948 106976 41954
rect 106924 41890 106976 41896
rect 102232 40044 102284 40050
rect 102232 39986 102284 39992
rect 102244 480 102272 39986
rect 104532 39636 104584 39642
rect 104532 39578 104584 39584
rect 103336 3324 103388 3330
rect 103336 3266 103388 3272
rect 103348 480 103376 3266
rect 104544 480 104572 39578
rect 105728 37256 105780 37262
rect 105728 37198 105780 37204
rect 105740 480 105768 37198
rect 106936 480 106964 41890
rect 108132 480 108160 44610
rect 111616 42220 111668 42226
rect 111616 42162 111668 42168
rect 109316 36508 109368 36514
rect 109316 36450 109368 36456
rect 109328 480 109356 36450
rect 111064 33652 111116 33658
rect 111064 33594 111116 33600
rect 110512 3256 110564 3262
rect 110512 3198 110564 3204
rect 110524 480 110552 3198
rect 111076 3194 111104 33594
rect 111064 3188 111116 3194
rect 111064 3130 111116 3136
rect 111628 480 111656 42162
rect 118792 39840 118844 39846
rect 118792 39782 118844 39788
rect 115204 39296 115256 39302
rect 115204 39238 115256 39244
rect 112812 36440 112864 36446
rect 112812 36382 112864 36388
rect 112824 480 112852 36382
rect 114008 31680 114060 31686
rect 114008 31622 114060 31628
rect 114020 480 114048 31622
rect 115216 480 115244 39238
rect 116400 34400 116452 34406
rect 116400 34342 116452 34348
rect 116412 480 116440 34342
rect 117596 31748 117648 31754
rect 117596 31690 117648 31696
rect 117608 480 117636 31690
rect 118804 480 118832 39782
rect 122288 39228 122340 39234
rect 122288 39170 122340 39176
rect 119896 34468 119948 34474
rect 119896 34410 119948 34416
rect 119908 480 119936 34410
rect 121092 31000 121144 31006
rect 121092 30942 121144 30948
rect 121104 480 121132 30942
rect 122300 480 122328 39170
rect 123484 33720 123536 33726
rect 123484 33662 123536 33668
rect 123496 480 123524 33662
rect 124680 30932 124732 30938
rect 124680 30874 124732 30880
rect 124692 480 124720 30874
rect 359476 3942 359504 269758
rect 359556 50108 359608 50114
rect 359556 50050 359608 50056
rect 359568 46345 359596 50050
rect 359554 46336 359610 46345
rect 359554 46271 359610 46280
rect 359832 46232 359884 46238
rect 359832 46174 359884 46180
rect 359844 45354 359872 46174
rect 359832 45348 359884 45354
rect 359832 45290 359884 45296
rect 360856 4010 360884 305594
rect 361764 304972 361816 304978
rect 361764 304914 361816 304920
rect 361776 304473 361804 304914
rect 361762 304464 361818 304473
rect 361762 304399 361818 304408
rect 360936 304360 360988 304366
rect 360936 304302 360988 304308
rect 360844 4004 360896 4010
rect 360844 3946 360896 3952
rect 359464 3936 359516 3942
rect 359464 3878 359516 3884
rect 360948 3262 360976 304302
rect 361028 304292 361080 304298
rect 361028 304234 361080 304240
rect 361040 3330 361068 304234
rect 361120 302932 361172 302938
rect 361120 302874 361172 302880
rect 361132 4078 361160 302874
rect 362224 301504 362276 301510
rect 362224 301446 362276 301452
rect 361764 293956 361816 293962
rect 361764 293898 361816 293904
rect 361776 293457 361804 293898
rect 361762 293448 361818 293457
rect 361762 293383 361818 293392
rect 361764 282872 361816 282878
rect 361764 282814 361816 282820
rect 361776 282441 361804 282814
rect 361762 282432 361818 282441
rect 361762 282367 361818 282376
rect 361764 271856 361816 271862
rect 361764 271798 361816 271804
rect 361776 271425 361804 271798
rect 361762 271416 361818 271425
rect 361762 271351 361818 271360
rect 361764 260840 361816 260846
rect 361764 260782 361816 260788
rect 361776 260409 361804 260782
rect 361762 260400 361818 260409
rect 361762 260335 361818 260344
rect 361764 249756 361816 249762
rect 361764 249698 361816 249704
rect 361776 249393 361804 249698
rect 361762 249384 361818 249393
rect 361762 249319 361818 249328
rect 361764 238740 361816 238746
rect 361764 238682 361816 238688
rect 361776 238377 361804 238682
rect 361762 238368 361818 238377
rect 361762 238303 361818 238312
rect 361764 227724 361816 227730
rect 361764 227666 361816 227672
rect 361776 227361 361804 227666
rect 361762 227352 361818 227361
rect 361762 227287 361818 227296
rect 361212 220108 361264 220114
rect 361212 220050 361264 220056
rect 361224 50114 361252 220050
rect 361580 216368 361632 216374
rect 361578 216336 361580 216345
rect 361632 216336 361634 216345
rect 361578 216271 361634 216280
rect 361764 205624 361816 205630
rect 361764 205566 361816 205572
rect 361776 205329 361804 205566
rect 361762 205320 361818 205329
rect 361762 205255 361818 205264
rect 361672 194540 361724 194546
rect 361672 194482 361724 194488
rect 361684 194313 361712 194482
rect 361670 194304 361726 194313
rect 361670 194239 361726 194248
rect 361672 183524 361724 183530
rect 361672 183466 361724 183472
rect 361684 183297 361712 183466
rect 361670 183288 361726 183297
rect 361670 183223 361726 183232
rect 361304 174684 361356 174690
rect 361304 174626 361356 174632
rect 361212 50108 361264 50114
rect 361212 50050 361264 50056
rect 361316 46102 361344 174626
rect 361672 172508 361724 172514
rect 361672 172450 361724 172456
rect 361684 172281 361712 172450
rect 361670 172272 361726 172281
rect 361670 172207 361726 172216
rect 361764 161424 361816 161430
rect 361764 161366 361816 161372
rect 361776 161265 361804 161366
rect 361762 161256 361818 161265
rect 361762 161191 361818 161200
rect 361764 150408 361816 150414
rect 361764 150350 361816 150356
rect 361776 150249 361804 150350
rect 361762 150240 361818 150249
rect 361762 150175 361818 150184
rect 361764 139392 361816 139398
rect 361764 139334 361816 139340
rect 361776 139233 361804 139334
rect 361762 139224 361818 139233
rect 361762 139159 361818 139168
rect 361396 138032 361448 138038
rect 361396 137974 361448 137980
rect 361408 46170 361436 137974
rect 361488 130212 361540 130218
rect 361488 130154 361540 130160
rect 361500 46481 361528 130154
rect 361580 128308 361632 128314
rect 361580 128250 361632 128256
rect 361592 128217 361620 128250
rect 361578 128208 361634 128217
rect 361578 128143 361634 128152
rect 361580 117292 361632 117298
rect 361580 117234 361632 117240
rect 361592 117201 361620 117234
rect 361578 117192 361634 117201
rect 361578 117127 361634 117136
rect 361580 106276 361632 106282
rect 361580 106218 361632 106224
rect 361592 106185 361620 106218
rect 361578 106176 361634 106185
rect 361578 106111 361634 106120
rect 361764 95192 361816 95198
rect 361762 95160 361764 95169
rect 361816 95160 361818 95169
rect 361762 95095 361818 95104
rect 361764 84176 361816 84182
rect 361762 84144 361764 84153
rect 361816 84144 361818 84153
rect 361762 84079 361818 84088
rect 361764 73160 361816 73166
rect 361762 73128 361764 73137
rect 361816 73128 361818 73137
rect 361762 73063 361818 73072
rect 361762 62112 361818 62121
rect 361762 62047 361764 62056
rect 361816 62047 361818 62056
rect 361764 62018 361816 62024
rect 361764 52420 361816 52426
rect 361764 52362 361816 52368
rect 361776 51105 361804 52362
rect 361762 51096 361818 51105
rect 361762 51031 361818 51040
rect 361486 46472 361542 46481
rect 361486 46407 361542 46416
rect 361396 46164 361448 46170
rect 361396 46106 361448 46112
rect 361304 46096 361356 46102
rect 361304 46038 361356 46044
rect 361120 4072 361172 4078
rect 361120 4014 361172 4020
rect 362236 3398 362264 301446
rect 362316 229764 362368 229770
rect 362316 229706 362368 229712
rect 362328 46238 362356 229706
rect 362960 180124 363012 180130
rect 362960 180066 363012 180072
rect 362972 174690 363000 180066
rect 362960 174684 363012 174690
rect 362960 174626 363012 174632
rect 362316 46232 362368 46238
rect 362316 46174 362368 46180
rect 362224 3392 362276 3398
rect 362224 3334 362276 3340
rect 361028 3324 361080 3330
rect 361028 3266 361080 3272
rect 360936 3256 360988 3262
rect 363616 3233 363644 305662
rect 363696 304428 363748 304434
rect 363696 304370 363748 304376
rect 363708 4146 363736 304370
rect 363800 216374 363828 333950
rect 365352 289468 365404 289474
rect 365352 289410 365404 289416
rect 365260 289332 365312 289338
rect 365260 289274 365312 289280
rect 365076 289264 365128 289270
rect 365076 289206 365128 289212
rect 364984 289128 365036 289134
rect 364984 289070 365036 289076
rect 363788 216368 363840 216374
rect 363788 216310 363840 216316
rect 364248 144220 364300 144226
rect 364248 144162 364300 144168
rect 364260 138038 364288 144162
rect 364248 138032 364300 138038
rect 364248 137974 364300 137980
rect 364996 28354 365024 289070
rect 365088 28422 365116 289206
rect 365168 289196 365220 289202
rect 365168 289138 365220 289144
rect 365076 28416 365128 28422
rect 365076 28358 365128 28364
rect 364984 28348 365036 28354
rect 364984 28290 365036 28296
rect 365180 28286 365208 289138
rect 365272 28490 365300 289274
rect 365364 33658 365392 289410
rect 365444 140820 365496 140826
rect 365444 140762 365496 140768
rect 365456 130218 365484 140762
rect 365444 130212 365496 130218
rect 365444 130154 365496 130160
rect 365352 33652 365404 33658
rect 365352 33594 365404 33600
rect 367756 31754 367784 386446
rect 367836 386436 367888 386442
rect 367836 386378 367888 386384
rect 367744 31748 367796 31754
rect 367744 31690 367796 31696
rect 367848 30938 367876 386378
rect 367928 385076 367980 385082
rect 367928 385018 367980 385024
rect 367940 31006 367968 385018
rect 368032 378078 368060 579634
rect 370516 379438 370544 601666
rect 370596 587852 370648 587858
rect 370596 587794 370648 587800
rect 370608 579630 370636 587794
rect 370596 579624 370648 579630
rect 370596 579566 370648 579572
rect 371896 380798 371924 623766
rect 371976 579624 372028 579630
rect 371976 579566 372028 579572
rect 371988 571334 372016 579566
rect 371976 571328 372028 571334
rect 371976 571270 372028 571276
rect 373264 571328 373316 571334
rect 373264 571270 373316 571276
rect 373276 564398 373304 571270
rect 373264 564392 373316 564398
rect 373264 564334 373316 564340
rect 374656 382226 374684 645866
rect 375288 564392 375340 564398
rect 375288 564334 375340 564340
rect 375300 557534 375328 564334
rect 375300 557506 375420 557534
rect 375392 557190 375420 557506
rect 375380 557184 375432 557190
rect 375380 557126 375432 557132
rect 374644 382220 374696 382226
rect 374644 382162 374696 382168
rect 376036 382158 376064 656882
rect 377772 557184 377824 557190
rect 377772 557126 377824 557132
rect 377784 550662 377812 557126
rect 377772 550656 377824 550662
rect 377772 550598 377824 550604
rect 378784 386572 378836 386578
rect 378784 386514 378836 386520
rect 376024 382152 376076 382158
rect 376024 382094 376076 382100
rect 371884 380792 371936 380798
rect 371884 380734 371936 380740
rect 370504 379432 370556 379438
rect 370504 379374 370556 379380
rect 368020 378072 368072 378078
rect 368020 378014 368072 378020
rect 371884 339516 371936 339522
rect 371884 339458 371936 339464
rect 371896 315994 371924 339458
rect 371884 315988 371936 315994
rect 371884 315930 371936 315936
rect 376024 295248 376076 295254
rect 376024 295190 376076 295196
rect 373540 292392 373592 292398
rect 373540 292334 373592 292340
rect 373264 292324 373316 292330
rect 373264 292266 373316 292272
rect 370872 292188 370924 292194
rect 370872 292130 370924 292136
rect 370596 292120 370648 292126
rect 370596 292062 370648 292068
rect 370504 291916 370556 291922
rect 370504 291858 370556 291864
rect 368020 291848 368072 291854
rect 368020 291790 368072 291796
rect 368110 291816 368166 291825
rect 368032 31686 368060 291790
rect 368110 291751 368166 291760
rect 368020 31680 368072 31686
rect 368020 31622 368072 31628
rect 368124 31142 368152 291751
rect 368204 289400 368256 289406
rect 368204 289342 368256 289348
rect 368216 36582 368244 289342
rect 369124 239420 369176 239426
rect 369124 239362 369176 239368
rect 369136 229770 369164 239362
rect 369124 229764 369176 229770
rect 369124 229706 369176 229712
rect 368388 143880 368440 143886
rect 368388 143822 368440 143828
rect 368400 140826 368428 143822
rect 368388 140820 368440 140826
rect 368388 140762 368440 140768
rect 368204 36576 368256 36582
rect 368204 36518 368256 36524
rect 370516 31482 370544 291858
rect 370504 31476 370556 31482
rect 370504 31418 370556 31424
rect 370608 31414 370636 292062
rect 370780 292052 370832 292058
rect 370780 291994 370832 292000
rect 370688 291780 370740 291786
rect 370688 291722 370740 291728
rect 370596 31408 370648 31414
rect 370596 31350 370648 31356
rect 368112 31136 368164 31142
rect 368112 31078 368164 31084
rect 370700 31074 370728 291722
rect 370792 31618 370820 291994
rect 370780 31612 370832 31618
rect 370780 31554 370832 31560
rect 370884 31550 370912 292130
rect 370964 291984 371016 291990
rect 370964 291926 371016 291932
rect 370976 41954 371004 291926
rect 371240 149728 371292 149734
rect 371240 149670 371292 149676
rect 371252 144226 371280 149670
rect 371240 144220 371292 144226
rect 371240 144162 371292 144168
rect 370964 41948 371016 41954
rect 370964 41890 371016 41896
rect 370872 31544 370924 31550
rect 370872 31486 370924 31492
rect 373276 31346 373304 292266
rect 373448 292256 373500 292262
rect 373448 292198 373500 292204
rect 373356 291712 373408 291718
rect 373356 291654 373408 291660
rect 373264 31340 373316 31346
rect 373264 31282 373316 31288
rect 373368 31278 373396 291654
rect 373356 31272 373408 31278
rect 373356 31214 373408 31220
rect 373460 31210 373488 292198
rect 373552 39982 373580 292334
rect 374644 195152 374696 195158
rect 374644 195094 374696 195100
rect 374656 180130 374684 195094
rect 374644 180124 374696 180130
rect 374644 180066 374696 180072
rect 373632 156664 373684 156670
rect 373632 156606 373684 156612
rect 373644 143886 373672 156606
rect 373632 143880 373684 143886
rect 373632 143822 373684 143828
rect 373540 39976 373592 39982
rect 373540 39918 373592 39924
rect 373448 31204 373500 31210
rect 373448 31146 373500 31152
rect 370688 31068 370740 31074
rect 370688 31010 370740 31016
rect 367928 31000 367980 31006
rect 367928 30942 367980 30948
rect 367836 30932 367888 30938
rect 367836 30874 367888 30880
rect 365260 28484 365312 28490
rect 365260 28426 365312 28432
rect 365168 28280 365220 28286
rect 365168 28222 365220 28228
rect 363696 4140 363748 4146
rect 363696 4082 363748 4088
rect 376036 4049 376064 295190
rect 376208 294976 376260 294982
rect 376208 294918 376260 294924
rect 376116 294908 376168 294914
rect 376116 294850 376168 294856
rect 376128 34202 376156 294850
rect 376116 34196 376168 34202
rect 376116 34138 376168 34144
rect 376220 34134 376248 294918
rect 376300 294636 376352 294642
rect 376300 294578 376352 294584
rect 376208 34128 376260 34134
rect 376208 34070 376260 34076
rect 376312 34066 376340 294578
rect 376392 292528 376444 292534
rect 376392 292470 376444 292476
rect 376404 34270 376432 292470
rect 376484 292460 376536 292466
rect 376484 292402 376536 292408
rect 376496 34338 376524 292402
rect 377404 211812 377456 211818
rect 377404 211754 377456 211760
rect 377416 195158 377444 211754
rect 377404 195152 377456 195158
rect 377404 195094 377456 195100
rect 378692 162920 378744 162926
rect 378692 162862 378744 162868
rect 378704 156670 378732 162862
rect 378692 156664 378744 156670
rect 378692 156606 378744 156612
rect 376484 34332 376536 34338
rect 376484 34274 376536 34280
rect 376392 34264 376444 34270
rect 376392 34206 376444 34212
rect 376300 34060 376352 34066
rect 376300 34002 376352 34008
rect 378796 33726 378824 386514
rect 378888 383586 378916 667898
rect 380164 550588 380216 550594
rect 380164 550530 380216 550536
rect 380176 540938 380204 550530
rect 380164 540932 380216 540938
rect 380164 540874 380216 540880
rect 382280 540932 382332 540938
rect 382280 540874 382332 540880
rect 382292 532710 382320 540874
rect 382280 532704 382332 532710
rect 382280 532646 382332 532652
rect 384304 532704 384356 532710
rect 384304 532646 384356 532652
rect 384316 524142 384344 532646
rect 384304 524136 384356 524142
rect 384304 524078 384356 524084
rect 385684 524136 385736 524142
rect 385684 524078 385736 524084
rect 385696 516186 385724 524078
rect 385684 516180 385736 516186
rect 385684 516122 385736 516128
rect 389180 516112 389232 516118
rect 389180 516054 389232 516060
rect 389192 511970 389220 516054
rect 389180 511964 389232 511970
rect 389180 511906 389232 511912
rect 391204 511964 391256 511970
rect 391204 511906 391256 511912
rect 391216 505850 391244 511906
rect 391204 505844 391256 505850
rect 391204 505786 391256 505792
rect 392584 505844 392636 505850
rect 392584 505786 392636 505792
rect 381636 491360 381688 491366
rect 381636 491302 381688 491308
rect 381544 386640 381596 386646
rect 381544 386582 381596 386588
rect 378876 383580 378928 383586
rect 378876 383522 378928 383528
rect 378876 295044 378928 295050
rect 378876 294986 378928 294992
rect 378784 33720 378836 33726
rect 378784 33662 378836 33668
rect 376022 4040 376078 4049
rect 376022 3975 376078 3984
rect 378888 3874 378916 294986
rect 379060 294840 379112 294846
rect 379060 294782 379112 294788
rect 378966 294536 379022 294545
rect 378966 294471 379022 294480
rect 378980 33862 379008 294471
rect 379072 33998 379100 294782
rect 379244 294772 379296 294778
rect 379244 294714 379296 294720
rect 379152 294704 379204 294710
rect 379152 294646 379204 294652
rect 379060 33992 379112 33998
rect 379060 33934 379112 33940
rect 379164 33930 379192 294646
rect 379256 45218 379284 294714
rect 379244 45212 379296 45218
rect 379244 45154 379296 45160
rect 381556 34474 381584 386582
rect 381648 372570 381676 491302
rect 392596 456754 392624 505786
rect 396724 469260 396776 469266
rect 396724 469202 396776 469208
rect 392584 456748 392636 456754
rect 392584 456690 392636 456696
rect 395344 456748 395396 456754
rect 395344 456690 395396 456696
rect 395356 433294 395384 456690
rect 395344 433288 395396 433294
rect 395344 433230 395396 433236
rect 381636 372564 381688 372570
rect 381636 372506 381688 372512
rect 396736 371210 396764 469202
rect 396724 371204 396776 371210
rect 396724 371146 396776 371152
rect 397472 336122 397500 703520
rect 400864 634840 400916 634846
rect 400864 634782 400916 634788
rect 399484 447160 399536 447166
rect 399484 447102 399536 447108
rect 398104 433288 398156 433294
rect 398104 433230 398156 433236
rect 398116 423638 398144 433230
rect 398104 423632 398156 423638
rect 398104 423574 398156 423580
rect 398840 423632 398892 423638
rect 398840 423574 398892 423580
rect 398852 418878 398880 423574
rect 398840 418872 398892 418878
rect 398840 418814 398892 418820
rect 399496 369850 399524 447102
rect 400680 418872 400732 418878
rect 400680 418814 400732 418820
rect 400692 413982 400720 418814
rect 400680 413976 400732 413982
rect 400680 413918 400732 413924
rect 400876 380730 400904 634782
rect 403624 557592 403676 557598
rect 403624 557534 403676 557540
rect 402336 413976 402388 413982
rect 402336 413918 402388 413924
rect 402348 410582 402376 413918
rect 402336 410576 402388 410582
rect 402336 410518 402388 410524
rect 400864 380724 400916 380730
rect 400864 380666 400916 380672
rect 403636 376718 403664 557534
rect 406384 535492 406436 535498
rect 406384 535434 406436 535440
rect 403624 376712 403676 376718
rect 403624 376654 403676 376660
rect 406396 375358 406424 535434
rect 407764 524476 407816 524482
rect 407764 524418 407816 524424
rect 406384 375352 406436 375358
rect 406384 375294 406436 375300
rect 407776 375290 407804 524418
rect 410524 513392 410576 513398
rect 410524 513334 410576 513340
rect 409144 410576 409196 410582
rect 409144 410518 409196 410524
rect 409156 396098 409184 410518
rect 409144 396092 409196 396098
rect 409144 396034 409196 396040
rect 407764 375284 407816 375290
rect 407764 375226 407816 375232
rect 410536 373998 410564 513334
rect 411904 502376 411956 502382
rect 411904 502318 411956 502324
rect 411628 396024 411680 396030
rect 411628 395966 411680 395972
rect 411640 391270 411668 395966
rect 411628 391264 411680 391270
rect 411628 391206 411680 391212
rect 410524 373992 410576 373998
rect 410524 373934 410576 373940
rect 411916 373930 411944 502318
rect 411904 373924 411956 373930
rect 411904 373866 411956 373872
rect 409880 369912 409932 369918
rect 409880 369854 409932 369860
rect 399484 369844 399536 369850
rect 399484 369786 399536 369792
rect 409892 365702 409920 369854
rect 409880 365696 409932 365702
rect 409880 365638 409932 365644
rect 407028 350600 407080 350606
rect 407028 350542 407080 350548
rect 402244 347812 402296 347818
rect 402244 347754 402296 347760
rect 402256 338094 402284 347754
rect 402244 338088 402296 338094
rect 402244 338030 402296 338036
rect 397460 336116 397512 336122
rect 397460 336058 397512 336064
rect 399484 335368 399536 335374
rect 399484 335310 399536 335316
rect 395620 303408 395672 303414
rect 395620 303350 395672 303356
rect 395436 302728 395488 302734
rect 395436 302670 395488 302676
rect 393044 300552 393096 300558
rect 392582 300520 392638 300529
rect 393044 300494 393096 300500
rect 392582 300455 392638 300464
rect 392676 300484 392728 300490
rect 390192 300348 390244 300354
rect 390192 300290 390244 300296
rect 389916 300280 389968 300286
rect 389916 300222 389968 300228
rect 389824 300144 389876 300150
rect 389824 300086 389876 300092
rect 387432 298104 387484 298110
rect 387432 298046 387484 298052
rect 387340 297968 387392 297974
rect 387340 297910 387392 297916
rect 384396 297900 384448 297906
rect 384396 297842 384448 297848
rect 381728 297696 381780 297702
rect 381728 297638 381780 297644
rect 381636 286408 381688 286414
rect 381636 286350 381688 286356
rect 381544 34468 381596 34474
rect 381544 34410 381596 34416
rect 379152 33924 379204 33930
rect 379152 33866 379204 33872
rect 378968 33856 379020 33862
rect 378968 33798 379020 33804
rect 381648 20670 381676 286350
rect 381740 36514 381768 297638
rect 384304 297560 384356 297566
rect 384304 297502 384356 297508
rect 381912 295316 381964 295322
rect 381912 295258 381964 295264
rect 381820 295180 381872 295186
rect 381820 295122 381872 295128
rect 381728 36508 381780 36514
rect 381728 36450 381780 36456
rect 381832 34406 381860 295122
rect 381820 34400 381872 34406
rect 381820 34342 381872 34348
rect 381924 33794 381952 295258
rect 382004 295112 382056 295118
rect 382004 295054 382056 295060
rect 382016 36446 382044 295054
rect 382924 239488 382976 239494
rect 382924 239430 382976 239436
rect 382936 220114 382964 239430
rect 382924 220108 382976 220114
rect 382924 220050 382976 220056
rect 384316 37126 384344 297502
rect 384408 37194 384436 297842
rect 387156 297764 387208 297770
rect 387156 297706 387208 297712
rect 384488 297492 384540 297498
rect 384488 297434 384540 297440
rect 384500 37262 384528 297434
rect 384580 297424 384632 297430
rect 384580 297366 384632 297372
rect 384592 40050 384620 297366
rect 387064 297356 387116 297362
rect 387064 297298 387116 297304
rect 386052 168428 386104 168434
rect 386052 168370 386104 168376
rect 386064 162926 386092 168370
rect 386052 162920 386104 162926
rect 386052 162862 386104 162868
rect 384580 40044 384632 40050
rect 384580 39986 384632 39992
rect 384488 37256 384540 37262
rect 384488 37198 384540 37204
rect 384396 37188 384448 37194
rect 384396 37130 384448 37136
rect 384304 37120 384356 37126
rect 384304 37062 384356 37068
rect 382004 36440 382056 36446
rect 382004 36382 382056 36388
rect 381912 33788 381964 33794
rect 381912 33730 381964 33736
rect 381636 20664 381688 20670
rect 381636 20606 381688 20612
rect 387076 3913 387104 297298
rect 387168 37058 387196 297706
rect 387248 297628 387300 297634
rect 387248 297570 387300 297576
rect 387156 37052 387208 37058
rect 387156 36994 387208 37000
rect 387260 36990 387288 297570
rect 387248 36984 387300 36990
rect 387248 36926 387300 36932
rect 387352 36922 387380 297910
rect 387444 42702 387472 298046
rect 387524 297832 387576 297838
rect 387524 297774 387576 297780
rect 387536 44742 387564 297774
rect 388444 242208 388496 242214
rect 388444 242150 388496 242156
rect 388456 239494 388484 242150
rect 388444 239488 388496 239494
rect 388444 239430 388496 239436
rect 388444 181620 388496 181626
rect 388444 181562 388496 181568
rect 388456 168434 388484 181562
rect 388444 168428 388496 168434
rect 388444 168370 388496 168376
rect 387524 44736 387576 44742
rect 387524 44678 387576 44684
rect 387432 42696 387484 42702
rect 387432 42638 387484 42644
rect 387340 36916 387392 36922
rect 387340 36858 387392 36864
rect 389836 36650 389864 300086
rect 389928 36718 389956 300222
rect 390008 298036 390060 298042
rect 390008 297978 390060 297984
rect 390020 36854 390048 297978
rect 390100 297288 390152 297294
rect 390100 297230 390152 297236
rect 390008 36848 390060 36854
rect 390008 36790 390060 36796
rect 390112 36786 390140 297230
rect 390204 39778 390232 300290
rect 390284 300212 390336 300218
rect 390284 300154 390336 300160
rect 390296 39914 390324 300154
rect 390652 186312 390704 186318
rect 390652 186254 390704 186260
rect 390664 181626 390692 186254
rect 390652 181620 390704 181626
rect 390652 181562 390704 181568
rect 390284 39908 390336 39914
rect 390284 39850 390336 39856
rect 390192 39772 390244 39778
rect 390192 39714 390244 39720
rect 390100 36780 390152 36786
rect 390100 36722 390152 36728
rect 389916 36712 389968 36718
rect 389916 36654 389968 36660
rect 389824 36644 389876 36650
rect 389824 36586 389876 36592
rect 387062 3904 387118 3913
rect 378876 3868 378928 3874
rect 387062 3839 387118 3848
rect 378876 3810 378928 3816
rect 392596 3777 392624 300455
rect 392676 300426 392728 300432
rect 392688 3806 392716 300426
rect 392860 300416 392912 300422
rect 392766 300384 392822 300393
rect 392860 300358 392912 300364
rect 392766 300319 392822 300328
rect 392780 39438 392808 300319
rect 392872 39710 392900 300358
rect 392950 300112 393006 300121
rect 392950 300047 393006 300056
rect 392860 39704 392912 39710
rect 392860 39646 392912 39652
rect 392964 39506 392992 300047
rect 393056 39574 393084 300494
rect 395342 300248 395398 300257
rect 395342 300183 395398 300192
rect 393964 194472 394016 194478
rect 393964 194414 394016 194420
rect 393976 186318 394004 194414
rect 393964 186312 394016 186318
rect 393964 186254 394016 186260
rect 393044 39568 393096 39574
rect 393044 39510 393096 39516
rect 392952 39500 393004 39506
rect 392952 39442 393004 39448
rect 392768 39432 392820 39438
rect 392768 39374 392820 39380
rect 392676 3800 392728 3806
rect 392582 3768 392638 3777
rect 392676 3742 392728 3748
rect 392582 3703 392638 3712
rect 360936 3198 360988 3204
rect 363602 3224 363658 3233
rect 363602 3159 363658 3168
rect 395356 2106 395384 300183
rect 395448 6866 395476 302670
rect 395526 300656 395582 300665
rect 395526 300591 395582 300600
rect 395436 6860 395488 6866
rect 395436 6802 395488 6808
rect 395540 3670 395568 300591
rect 395632 39302 395660 303350
rect 398288 303340 398340 303346
rect 398288 303282 398340 303288
rect 398104 303204 398156 303210
rect 398104 303146 398156 303152
rect 395804 303000 395856 303006
rect 395804 302942 395856 302948
rect 395712 300620 395764 300626
rect 395712 300562 395764 300568
rect 395620 39296 395672 39302
rect 395620 39238 395672 39244
rect 395724 39234 395752 300562
rect 395816 44674 395844 302942
rect 396724 294568 396776 294574
rect 396724 294510 396776 294516
rect 396264 213988 396316 213994
rect 396264 213930 396316 213936
rect 396276 211818 396304 213930
rect 396264 211812 396316 211818
rect 396264 211754 396316 211760
rect 396736 45422 396764 294510
rect 396816 263628 396868 263634
rect 396816 263570 396868 263576
rect 396828 239426 396856 263570
rect 396816 239420 396868 239426
rect 396816 239362 396868 239368
rect 396724 45416 396776 45422
rect 396724 45358 396776 45364
rect 395804 44668 395856 44674
rect 395804 44610 395856 44616
rect 398116 42634 398144 303146
rect 398196 303068 398248 303074
rect 398196 303010 398248 303016
rect 398208 42770 398236 303010
rect 398196 42764 398248 42770
rect 398196 42706 398248 42712
rect 398104 42628 398156 42634
rect 398104 42570 398156 42576
rect 398300 42022 398328 303282
rect 398380 303136 398432 303142
rect 398380 303078 398432 303084
rect 398392 42566 398420 303078
rect 399496 249762 399524 335310
rect 402256 334914 402284 338030
rect 407040 335354 407068 350542
rect 413100 336864 413152 336870
rect 413100 336806 413152 336812
rect 409420 336796 409472 336802
rect 409420 336738 409472 336744
rect 406120 335326 407068 335354
rect 406120 334914 406148 335326
rect 402086 334886 402284 334914
rect 405766 334886 406148 334914
rect 409432 334900 409460 336738
rect 413112 334900 413140 336806
rect 413664 336190 413692 703520
rect 429856 700670 429884 703520
rect 445116 700868 445168 700874
rect 445116 700810 445168 700816
rect 418804 700664 418856 700670
rect 418804 700606 418856 700612
rect 429844 700664 429896 700670
rect 429844 700606 429896 700612
rect 444104 700664 444156 700670
rect 444104 700606 444156 700612
rect 416044 685228 416096 685234
rect 416044 685170 416096 685176
rect 414664 458244 414716 458250
rect 414664 458186 414716 458192
rect 414676 371142 414704 458186
rect 415400 391264 415452 391270
rect 415400 391206 415452 391212
rect 415412 389162 415440 391206
rect 415400 389156 415452 389162
rect 415400 389098 415452 389104
rect 414664 371136 414716 371142
rect 414664 371078 414716 371084
rect 416056 336326 416084 685170
rect 416136 436144 416188 436150
rect 416136 436086 416188 436092
rect 416148 369782 416176 436086
rect 417424 425128 417476 425134
rect 417424 425070 417476 425076
rect 416136 369776 416188 369782
rect 416136 369718 416188 369724
rect 417436 368490 417464 425070
rect 417516 389156 417568 389162
rect 417516 389098 417568 389104
rect 417528 378962 417556 389098
rect 417516 378956 417568 378962
rect 417516 378898 417568 378904
rect 417424 368484 417476 368490
rect 417424 368426 417476 368432
rect 416780 336932 416832 336938
rect 416780 336874 416832 336880
rect 416044 336320 416096 336326
rect 416044 336262 416096 336268
rect 413652 336184 413704 336190
rect 413652 336126 413704 336132
rect 416792 334900 416820 336874
rect 418816 336462 418844 700606
rect 418896 685364 418948 685370
rect 418896 685306 418948 685312
rect 418804 336456 418856 336462
rect 418804 336398 418856 336404
rect 418908 336394 418936 685306
rect 418988 684616 419040 684622
rect 418988 684558 419040 684564
rect 418896 336388 418948 336394
rect 418896 336330 418948 336336
rect 419000 336258 419028 684558
rect 420184 684548 420236 684554
rect 420184 684490 420236 684496
rect 419080 546508 419132 546514
rect 419080 546450 419132 546456
rect 419092 376650 419120 546450
rect 419172 480276 419224 480282
rect 419172 480218 419224 480224
rect 419080 376644 419132 376650
rect 419080 376586 419132 376592
rect 419184 372502 419212 480218
rect 419264 378956 419316 378962
rect 419264 378898 419316 378904
rect 419172 372496 419224 372502
rect 419172 372438 419224 372444
rect 419276 369374 419304 378898
rect 419264 369368 419316 369374
rect 419264 369310 419316 369316
rect 418988 336252 419040 336258
rect 418988 336194 419040 336200
rect 420196 334762 420224 684490
rect 420736 683732 420788 683738
rect 420736 683674 420788 683680
rect 420276 683664 420328 683670
rect 420276 683606 420328 683612
rect 420184 334756 420236 334762
rect 420184 334698 420236 334704
rect 420288 334694 420316 683606
rect 420368 683596 420420 683602
rect 420368 683538 420420 683544
rect 420380 335209 420408 683538
rect 420644 683528 420696 683534
rect 420644 683470 420696 683476
rect 420552 683460 420604 683466
rect 420552 683402 420604 683408
rect 420366 335200 420422 335209
rect 420366 335135 420422 335144
rect 420564 334898 420592 683402
rect 420552 334892 420604 334898
rect 420552 334834 420604 334840
rect 420276 334688 420328 334694
rect 420276 334630 420328 334636
rect 420656 334626 420684 683470
rect 420748 334830 420776 683674
rect 422484 447432 422536 447438
rect 422484 447374 422536 447380
rect 422496 444924 422524 447374
rect 437388 447364 437440 447370
rect 437388 447306 437440 447312
rect 432420 447296 432472 447302
rect 432420 447238 432472 447244
rect 427452 447228 427504 447234
rect 427452 447170 427504 447176
rect 427464 444924 427492 447170
rect 432432 444924 432460 447238
rect 437400 444924 437428 447306
rect 442382 444378 442672 444394
rect 442382 444372 442684 444378
rect 442382 444366 442632 444372
rect 442632 444314 442684 444320
rect 421484 417586 421512 420036
rect 422128 417654 422156 420036
rect 422786 420022 423168 420050
rect 423430 420022 423536 420050
rect 422116 417648 422168 417654
rect 422116 417590 422168 417596
rect 421472 417580 421524 417586
rect 421472 417522 421524 417528
rect 423140 416362 423168 420022
rect 423128 416356 423180 416362
rect 423128 416298 423180 416304
rect 423508 393990 423536 420022
rect 424060 417450 424088 420036
rect 424704 417518 424732 420036
rect 425348 417722 425376 420036
rect 425992 417790 426020 420036
rect 425980 417784 426032 417790
rect 425980 417726 426032 417732
rect 425336 417716 425388 417722
rect 425336 417658 425388 417664
rect 424692 417512 424744 417518
rect 424692 417454 424744 417460
rect 424048 417444 424100 417450
rect 424048 417386 424100 417392
rect 423588 416356 423640 416362
rect 423588 416298 423640 416304
rect 423496 393984 423548 393990
rect 423496 393926 423548 393932
rect 423600 391270 423628 416298
rect 443644 414044 443696 414050
rect 443644 413986 443696 413992
rect 439504 403028 439556 403034
rect 439504 402970 439556 402976
rect 423588 391264 423640 391270
rect 423588 391206 423640 391212
rect 421564 369368 421616 369374
rect 421564 369310 421616 369316
rect 421576 362506 421604 369310
rect 439516 367062 439544 402970
rect 443656 368422 443684 413986
rect 443736 392012 443788 392018
rect 443736 391954 443788 391960
rect 443644 368416 443696 368422
rect 443644 368358 443696 368364
rect 439504 367056 439556 367062
rect 439504 366998 439556 367004
rect 443748 366994 443776 391954
rect 443828 380928 443880 380934
rect 443828 380870 443880 380876
rect 443736 366988 443788 366994
rect 443736 366930 443788 366936
rect 443840 365634 443868 380870
rect 443828 365628 443880 365634
rect 443828 365570 443880 365576
rect 432880 363044 432932 363050
rect 432880 362986 432932 362992
rect 432788 362976 432840 362982
rect 432788 362918 432840 362924
rect 421564 362500 421616 362506
rect 421564 362442 421616 362448
rect 423588 362500 423640 362506
rect 423588 362442 423640 362448
rect 423600 357474 423628 362442
rect 432696 361616 432748 361622
rect 432696 361558 432748 361564
rect 423588 357468 423640 357474
rect 423588 357410 423640 357416
rect 426348 357400 426400 357406
rect 426348 357342 426400 357348
rect 426360 354674 426388 357342
rect 426360 354646 426480 354674
rect 426452 351966 426480 354646
rect 426440 351960 426492 351966
rect 426440 351902 426492 351908
rect 431224 339584 431276 339590
rect 431224 339526 431276 339532
rect 427818 337104 427874 337113
rect 427818 337039 427874 337048
rect 420736 334824 420788 334830
rect 420736 334766 420788 334772
rect 427832 334642 427860 337039
rect 427832 334628 427952 334642
rect 420644 334620 420696 334626
rect 427846 334614 427952 334628
rect 420644 334562 420696 334568
rect 427924 334506 427952 334614
rect 428094 334520 428150 334529
rect 427846 334478 428094 334506
rect 428094 334455 428150 334464
rect 420458 334384 420514 334393
rect 420458 334319 420514 334328
rect 424138 334384 424194 334393
rect 424138 334319 424194 334328
rect 400864 306196 400916 306202
rect 400864 306138 400916 306144
rect 400128 269884 400180 269890
rect 400128 269826 400180 269832
rect 400140 263634 400168 269826
rect 400128 263628 400180 263634
rect 400128 263570 400180 263576
rect 399484 249756 399536 249762
rect 399484 249698 399536 249704
rect 400220 244928 400272 244934
rect 400220 244870 400272 244876
rect 400232 242214 400260 244870
rect 400220 242208 400272 242214
rect 400220 242150 400272 242156
rect 399484 225616 399536 225622
rect 399484 225558 399536 225564
rect 399496 213994 399524 225558
rect 399484 213988 399536 213994
rect 399484 213930 399536 213936
rect 399484 207664 399536 207670
rect 399484 207606 399536 207612
rect 399496 194478 399524 207606
rect 399484 194472 399536 194478
rect 399484 194414 399536 194420
rect 398472 186380 398524 186386
rect 398472 186322 398524 186328
rect 398484 149734 398512 186322
rect 398472 149728 398524 149734
rect 398472 149670 398524 149676
rect 398380 42560 398432 42566
rect 398380 42502 398432 42508
rect 398288 42016 398340 42022
rect 398288 41958 398340 41964
rect 395712 39228 395764 39234
rect 395712 39170 395764 39176
rect 400876 33114 400904 306138
rect 406660 306128 406712 306134
rect 406660 306070 406712 306076
rect 406476 306060 406528 306066
rect 406476 306002 406528 306008
rect 403808 305992 403860 305998
rect 403808 305934 403860 305940
rect 406382 305960 406438 305969
rect 403624 305924 403676 305930
rect 403624 305866 403676 305872
rect 401048 303612 401100 303618
rect 401048 303554 401100 303560
rect 400956 302796 401008 302802
rect 400956 302738 401008 302744
rect 400968 42430 400996 302738
rect 400956 42424 401008 42430
rect 400956 42366 401008 42372
rect 401060 42362 401088 303554
rect 401140 303476 401192 303482
rect 401140 303418 401192 303424
rect 401048 42356 401100 42362
rect 401048 42298 401100 42304
rect 401152 42294 401180 303418
rect 401324 302864 401376 302870
rect 401230 302832 401286 302841
rect 401324 302806 401376 302812
rect 401230 302767 401286 302776
rect 401140 42288 401192 42294
rect 401140 42230 401192 42236
rect 401244 42090 401272 302767
rect 401336 42498 401364 302806
rect 401600 191140 401652 191146
rect 401600 191082 401652 191088
rect 401612 186386 401640 191082
rect 401600 186380 401652 186386
rect 401600 186322 401652 186328
rect 403636 45082 403664 305866
rect 403716 305788 403768 305794
rect 403716 305730 403768 305736
rect 403728 45286 403756 305730
rect 403716 45280 403768 45286
rect 403716 45222 403768 45228
rect 403624 45076 403676 45082
rect 403624 45018 403676 45024
rect 403820 45014 403848 305934
rect 406382 305895 406438 305904
rect 403900 305856 403952 305862
rect 403900 305798 403952 305804
rect 403912 45150 403940 305798
rect 403992 303544 404044 303550
rect 403992 303486 404044 303492
rect 403900 45144 403952 45150
rect 403900 45086 403952 45092
rect 403808 45008 403860 45014
rect 403808 44950 403860 44956
rect 404004 44810 404032 303486
rect 404084 160268 404136 160274
rect 404084 160210 404136 160216
rect 404096 73166 404124 160210
rect 404084 73160 404136 73166
rect 404084 73102 404136 73108
rect 403992 44804 404044 44810
rect 403992 44746 404044 44752
rect 401324 42492 401376 42498
rect 401324 42434 401376 42440
rect 401232 42084 401284 42090
rect 401232 42026 401284 42032
rect 400864 33108 400916 33114
rect 400864 33050 400916 33056
rect 395528 3664 395580 3670
rect 395528 3606 395580 3612
rect 406396 3505 406424 305895
rect 406488 44946 406516 306002
rect 406566 305688 406622 305697
rect 406566 305623 406622 305632
rect 406476 44940 406528 44946
rect 406476 44882 406528 44888
rect 406580 3641 406608 305623
rect 406672 44849 406700 306070
rect 406750 305824 406806 305833
rect 406750 305759 406806 305768
rect 406764 44878 406792 305759
rect 431236 304978 431264 339526
rect 432604 334960 432656 334966
rect 432604 334902 432656 334908
rect 431868 328500 431920 328506
rect 431868 328442 431920 328448
rect 431224 304972 431276 304978
rect 431224 304914 431276 304920
rect 427084 289604 427136 289610
rect 427084 289546 427136 289552
rect 407764 289536 407816 289542
rect 407764 289478 407816 289484
rect 406844 260160 406896 260166
rect 406844 260102 406896 260108
rect 406856 244934 406884 260102
rect 406844 244928 406896 244934
rect 406844 244870 406896 244876
rect 406844 161492 406896 161498
rect 406844 161434 406896 161440
rect 406856 62082 406884 161434
rect 406844 62076 406896 62082
rect 406844 62018 406896 62024
rect 406752 44872 406804 44878
rect 406658 44840 406714 44849
rect 406752 44814 406804 44820
rect 406658 44775 406714 44784
rect 406566 3632 406622 3641
rect 407776 3602 407804 289478
rect 410524 286340 410576 286346
rect 410524 286282 410576 286288
rect 410536 269890 410564 286282
rect 410524 269884 410576 269890
rect 410524 269826 410576 269832
rect 427096 262886 427124 289546
rect 431224 273964 431276 273970
rect 431224 273906 431276 273912
rect 417424 262880 417476 262886
rect 417424 262822 417476 262828
rect 427084 262880 427136 262886
rect 427084 262822 427136 262828
rect 417436 260166 417464 262822
rect 417424 260160 417476 260166
rect 417424 260102 417476 260108
rect 431236 253978 431264 273906
rect 422944 253972 422996 253978
rect 422944 253914 422996 253920
rect 431224 253972 431276 253978
rect 431224 253914 431276 253920
rect 422956 245342 422984 253914
rect 420184 245336 420236 245342
rect 420184 245278 420236 245284
rect 422944 245336 422996 245342
rect 422944 245278 422996 245284
rect 420196 235278 420224 245278
rect 427084 239420 427136 239426
rect 427084 239362 427136 239368
rect 411904 235272 411956 235278
rect 411904 235214 411956 235220
rect 420184 235272 420236 235278
rect 420184 235214 420236 235220
rect 411916 225622 411944 235214
rect 411904 225616 411956 225622
rect 411904 225558 411956 225564
rect 413100 214600 413152 214606
rect 413100 214542 413152 214548
rect 413112 210186 413140 214542
rect 407856 210180 407908 210186
rect 407856 210122 407908 210128
rect 413100 210180 413152 210186
rect 413100 210122 413152 210128
rect 407868 207670 407896 210122
rect 427096 209098 427124 239362
rect 411904 209092 411956 209098
rect 411904 209034 411956 209040
rect 427084 209092 427136 209098
rect 427084 209034 427136 209040
rect 407856 207664 407908 207670
rect 407856 207606 407908 207612
rect 411916 198762 411944 209034
rect 408500 198756 408552 198762
rect 408500 198698 408552 198704
rect 411904 198756 411956 198762
rect 411904 198698 411956 198704
rect 408512 191146 408540 198698
rect 408500 191140 408552 191146
rect 408500 191082 408552 191088
rect 422022 162752 422078 162761
rect 422022 162687 422078 162696
rect 426346 162752 426402 162761
rect 426346 162687 426402 162696
rect 428646 162752 428702 162761
rect 428646 162687 428702 162696
rect 418712 162376 418764 162382
rect 418712 162318 418764 162324
rect 414756 162308 414808 162314
rect 414756 162250 414808 162256
rect 411628 162240 411680 162246
rect 411628 162182 411680 162188
rect 407856 160200 407908 160206
rect 407856 160142 407908 160148
rect 411444 160200 411496 160206
rect 411444 160142 411496 160148
rect 407868 52426 407896 160142
rect 409696 160132 409748 160138
rect 409696 160074 409748 160080
rect 409144 159724 409196 159730
rect 409144 159666 409196 159672
rect 409156 84182 409184 159666
rect 409236 159656 409288 159662
rect 409236 159598 409288 159604
rect 409248 95198 409276 159598
rect 409328 159588 409380 159594
rect 409328 159530 409380 159536
rect 409340 106282 409368 159530
rect 409420 159520 409472 159526
rect 409420 159462 409472 159468
rect 409432 117298 409460 159462
rect 409512 159452 409564 159458
rect 409512 159394 409564 159400
rect 409524 128314 409552 159394
rect 409604 159384 409656 159390
rect 409604 159326 409656 159332
rect 409616 139398 409644 159326
rect 409708 150414 409736 160074
rect 411456 159882 411484 160142
rect 411640 159882 411668 162182
rect 414768 161498 414796 162250
rect 414756 161492 414808 161498
rect 414756 161434 414808 161440
rect 414768 159882 414796 161434
rect 418160 160268 418212 160274
rect 418160 160210 418212 160216
rect 418172 159882 418200 160210
rect 418724 159882 418752 162318
rect 422036 160410 422064 162687
rect 426360 160546 426388 162687
rect 425336 160540 425388 160546
rect 425336 160482 425388 160488
rect 426348 160540 426400 160546
rect 426348 160482 426400 160488
rect 422024 160404 422076 160410
rect 422024 160346 422076 160352
rect 411456 159854 411792 159882
rect 414768 159854 415104 159882
rect 418172 159854 418752 159882
rect 422036 159746 422064 160346
rect 425348 159882 425376 160482
rect 428660 160478 428688 162687
rect 431880 161474 431908 328442
rect 432052 318300 432104 318306
rect 432052 318242 432104 318248
rect 432064 310865 432092 318242
rect 432050 310856 432106 310865
rect 432050 310791 432106 310800
rect 432616 271862 432644 334902
rect 432708 325553 432736 361558
rect 432800 329225 432828 362918
rect 432892 332897 432920 362986
rect 442264 361684 442316 361690
rect 442264 361626 442316 361632
rect 439688 360324 439740 360330
rect 439688 360266 439740 360272
rect 436928 360256 436980 360262
rect 436928 360198 436980 360204
rect 435456 358828 435508 358834
rect 435456 358770 435508 358776
rect 432972 351892 433024 351898
rect 432972 351834 433024 351840
rect 432984 349586 433012 351834
rect 432972 349580 433024 349586
rect 432972 349522 433024 349528
rect 433984 349580 434036 349586
rect 433984 349522 434036 349528
rect 433996 338026 434024 349522
rect 435364 338156 435416 338162
rect 435364 338098 435416 338104
rect 433984 338020 434036 338026
rect 433984 337962 434036 337968
rect 432878 332888 432934 332897
rect 432878 332823 432934 332832
rect 432880 330200 432932 330206
rect 432880 330142 432932 330148
rect 432786 329216 432842 329225
rect 432786 329151 432842 329160
rect 432892 325694 432920 330142
rect 432800 325666 432920 325694
rect 432694 325544 432750 325553
rect 432694 325479 432750 325488
rect 432696 322992 432748 322998
rect 432696 322934 432748 322940
rect 432708 314537 432736 322934
rect 432800 318209 432828 325666
rect 432880 324964 432932 324970
rect 432880 324906 432932 324912
rect 432892 321881 432920 324906
rect 432878 321872 432934 321881
rect 432878 321807 432934 321816
rect 432786 318200 432842 318209
rect 432786 318135 432842 318144
rect 432694 314528 432750 314537
rect 432694 314463 432750 314472
rect 433156 313948 433208 313954
rect 433156 313890 433208 313896
rect 433168 307193 433196 313890
rect 433154 307184 433210 307193
rect 433154 307119 433210 307128
rect 435376 293962 435404 338098
rect 435468 318306 435496 358770
rect 436836 338224 436888 338230
rect 436836 338166 436888 338172
rect 436376 338020 436428 338026
rect 436376 337962 436428 337968
rect 436388 329798 436416 337962
rect 436744 332648 436796 332654
rect 436744 332590 436796 332596
rect 436376 329792 436428 329798
rect 436376 329734 436428 329740
rect 436008 328568 436060 328574
rect 436008 328510 436060 328516
rect 435456 318300 435508 318306
rect 435456 318242 435508 318248
rect 435364 293956 435416 293962
rect 435364 293898 435416 293904
rect 432604 271856 432656 271862
rect 432604 271798 432656 271804
rect 435640 245676 435692 245682
rect 435640 245618 435692 245624
rect 435652 239426 435680 245618
rect 435640 239420 435692 239426
rect 435640 239362 435692 239368
rect 431788 161446 431908 161474
rect 428648 160472 428700 160478
rect 428648 160414 428700 160420
rect 425040 159854 425376 159882
rect 421392 159730 422064 159746
rect 421380 159724 422064 159730
rect 421432 159718 422064 159724
rect 421380 159666 421432 159672
rect 425164 159662 425192 159854
rect 425152 159656 425204 159662
rect 428660 159610 428688 160414
rect 431788 160342 431816 161446
rect 431776 160336 431828 160342
rect 431776 160278 431828 160284
rect 425152 159598 425204 159604
rect 428016 159594 428688 159610
rect 428004 159588 428688 159594
rect 428056 159582 428688 159588
rect 428004 159530 428056 159536
rect 431316 159520 431368 159526
rect 431316 159462 431368 159468
rect 431328 159338 431356 159462
rect 431788 159338 431816 160278
rect 436020 160274 436048 328510
rect 436100 218068 436152 218074
rect 436100 218010 436152 218016
rect 436112 214606 436140 218010
rect 436100 214600 436152 214606
rect 436100 214542 436152 214548
rect 436756 194546 436784 332590
rect 436848 282878 436876 338166
rect 436940 322998 436968 360198
rect 439596 332716 439648 332722
rect 439596 332658 439648 332664
rect 439504 329860 439556 329866
rect 439504 329802 439556 329808
rect 438124 329792 438176 329798
rect 438124 329734 438176 329740
rect 438136 324018 438164 329734
rect 438124 324012 438176 324018
rect 438124 323954 438176 323960
rect 436928 322992 436980 322998
rect 436928 322934 436980 322940
rect 436928 299600 436980 299606
rect 436928 299542 436980 299548
rect 436940 286346 436968 299542
rect 437480 292596 437532 292602
rect 437480 292538 437532 292544
rect 437492 289610 437520 292538
rect 437480 289604 437532 289610
rect 437480 289546 437532 289552
rect 436928 286340 436980 286346
rect 436928 286282 436980 286288
rect 436836 282872 436888 282878
rect 436836 282814 436888 282820
rect 436744 194540 436796 194546
rect 436744 194482 436796 194488
rect 439516 163674 439544 329802
rect 439608 205630 439636 332658
rect 439700 330206 439728 360266
rect 439872 336456 439924 336462
rect 439872 336398 439924 336404
rect 439780 336320 439832 336326
rect 439780 336262 439832 336268
rect 439688 330200 439740 330206
rect 439688 330142 439740 330148
rect 439792 320754 439820 336262
rect 439884 322318 439912 336398
rect 440884 336320 440936 336326
rect 440884 336262 440936 336268
rect 439964 324012 440016 324018
rect 439964 323954 440016 323960
rect 439872 322312 439924 322318
rect 439872 322254 439924 322260
rect 439976 322250 440004 323954
rect 439964 322244 440016 322250
rect 439964 322186 440016 322192
rect 439780 320748 439832 320754
rect 439780 320690 439832 320696
rect 439688 312588 439740 312594
rect 439688 312530 439740 312536
rect 439700 299606 439728 312530
rect 439688 299600 439740 299606
rect 439688 299542 439740 299548
rect 439688 297220 439740 297226
rect 439688 297162 439740 297168
rect 439700 273970 439728 297162
rect 439688 273964 439740 273970
rect 439688 273906 439740 273912
rect 440896 260846 440924 336262
rect 442276 324970 442304 361626
rect 443828 358896 443880 358902
rect 443828 358838 443880 358844
rect 442356 349852 442408 349858
rect 442356 349794 442408 349800
rect 442264 324964 442316 324970
rect 442264 324906 442316 324912
rect 442368 320142 442396 349794
rect 442540 336388 442592 336394
rect 442540 336330 442592 336336
rect 442448 334892 442500 334898
rect 442448 334834 442500 334840
rect 442356 320136 442408 320142
rect 442356 320078 442408 320084
rect 442460 319122 442488 334834
rect 442552 320686 442580 336330
rect 443736 335708 443788 335714
rect 443736 335650 443788 335656
rect 442632 334824 442684 334830
rect 442632 334766 442684 334772
rect 442540 320680 442592 320686
rect 442540 320622 442592 320628
rect 442644 319870 442672 334766
rect 443644 334076 443696 334082
rect 443644 334018 443696 334024
rect 442908 330540 442960 330546
rect 442908 330482 442960 330488
rect 442632 319864 442684 319870
rect 442632 319806 442684 319812
rect 442448 319116 442500 319122
rect 442448 319058 442500 319064
rect 440976 300688 441028 300694
rect 440976 300630 441028 300636
rect 440988 292602 441016 300630
rect 440976 292596 441028 292602
rect 440976 292538 441028 292544
rect 440884 260840 440936 260846
rect 440884 260782 440936 260788
rect 439688 258732 439740 258738
rect 439688 258674 439740 258680
rect 439700 245682 439728 258674
rect 439688 245676 439740 245682
rect 439688 245618 439740 245624
rect 442264 232960 442316 232966
rect 442264 232902 442316 232908
rect 442276 223582 442304 232902
rect 439688 223576 439740 223582
rect 439688 223518 439740 223524
rect 442264 223576 442316 223582
rect 442264 223518 442316 223524
rect 439700 218074 439728 223518
rect 439688 218068 439740 218074
rect 439688 218010 439740 218016
rect 439596 205624 439648 205630
rect 439596 205566 439648 205572
rect 438584 163668 438636 163674
rect 438584 163610 438636 163616
rect 439504 163668 439556 163674
rect 439504 163610 439556 163616
rect 435272 160268 435324 160274
rect 435272 160210 435324 160216
rect 436008 160268 436060 160274
rect 436008 160210 436060 160216
rect 435284 159882 435312 160210
rect 438596 160206 438624 163610
rect 438584 160200 438636 160206
rect 438584 160142 438636 160148
rect 434824 159854 435312 159882
rect 434824 159458 434852 159854
rect 434812 159452 434864 159458
rect 434812 159394 434864 159400
rect 431328 159310 431816 159338
rect 437940 159384 437992 159390
rect 438596 159338 438624 160142
rect 442920 160138 442948 330482
rect 443656 227730 443684 334018
rect 443748 238746 443776 335650
rect 443840 313954 443868 358838
rect 444116 322862 444144 700606
rect 444196 700460 444248 700466
rect 444196 700402 444248 700408
rect 444208 421977 444236 700402
rect 445024 700324 445076 700330
rect 445024 700266 445076 700272
rect 444288 423020 444340 423026
rect 444288 422962 444340 422968
rect 444194 421968 444250 421977
rect 444194 421903 444250 421912
rect 444196 341012 444248 341018
rect 444196 340954 444248 340960
rect 444208 336054 444236 340954
rect 444196 336048 444248 336054
rect 444196 335990 444248 335996
rect 444104 322856 444156 322862
rect 444104 322798 444156 322804
rect 444300 318714 444328 422962
rect 444932 334756 444984 334762
rect 444932 334698 444984 334704
rect 444944 322590 444972 334698
rect 444932 322584 444984 322590
rect 444932 322526 444984 322532
rect 445036 321298 445064 700266
rect 445024 321292 445076 321298
rect 445024 321234 445076 321240
rect 445128 321026 445156 700810
rect 449256 700800 449308 700806
rect 449256 700742 449308 700748
rect 446496 700732 446548 700738
rect 446496 700674 446548 700680
rect 446404 700596 446456 700602
rect 446404 700538 446456 700544
rect 445208 700528 445260 700534
rect 445208 700470 445260 700476
rect 445220 322697 445248 700470
rect 445300 685296 445352 685302
rect 445300 685238 445352 685244
rect 445206 322688 445262 322697
rect 445206 322623 445262 322632
rect 445116 321020 445168 321026
rect 445116 320962 445168 320968
rect 445312 319326 445340 685238
rect 445484 683392 445536 683398
rect 445484 683334 445536 683340
rect 445392 683324 445444 683330
rect 445392 683266 445444 683272
rect 445404 319734 445432 683266
rect 445496 321230 445524 683334
rect 446312 683188 446364 683194
rect 446312 683130 446364 683136
rect 445574 682816 445630 682825
rect 445574 682751 445630 682760
rect 445588 322833 445616 682751
rect 445668 447228 445720 447234
rect 445668 447170 445720 447176
rect 445680 354006 445708 447170
rect 446220 444372 446272 444378
rect 446220 444314 446272 444320
rect 445668 354000 445720 354006
rect 445668 353942 445720 353948
rect 446232 352578 446260 444314
rect 446220 352572 446272 352578
rect 446220 352514 446272 352520
rect 445668 334688 445720 334694
rect 445668 334630 445720 334636
rect 445574 322824 445630 322833
rect 445574 322759 445630 322768
rect 445680 322454 445708 334630
rect 446324 322561 446352 683130
rect 446310 322552 446366 322561
rect 446310 322487 446366 322496
rect 445668 322448 445720 322454
rect 445668 322390 445720 322396
rect 446416 321366 446444 700538
rect 446404 321360 446456 321366
rect 446404 321302 446456 321308
rect 445484 321224 445536 321230
rect 445484 321166 445536 321172
rect 446508 321162 446536 700674
rect 447876 700460 447928 700466
rect 447876 700402 447928 700408
rect 447784 700324 447836 700330
rect 447784 700266 447836 700272
rect 446588 686588 446640 686594
rect 446588 686530 446640 686536
rect 446496 321156 446548 321162
rect 446496 321098 446548 321104
rect 445392 319728 445444 319734
rect 445392 319670 445444 319676
rect 446600 319394 446628 686530
rect 446680 686520 446732 686526
rect 446680 686462 446732 686468
rect 446588 319388 446640 319394
rect 446588 319330 446640 319336
rect 445300 319320 445352 319326
rect 445300 319262 445352 319268
rect 446692 319054 446720 686462
rect 446770 683360 446826 683369
rect 446770 683295 446826 683304
rect 446784 319705 446812 683295
rect 446864 683256 446916 683262
rect 446864 683198 446916 683204
rect 446954 683224 447010 683233
rect 446876 320074 446904 683198
rect 446954 683159 447010 683168
rect 446968 320822 446996 683159
rect 447048 682712 447100 682718
rect 447048 682654 447100 682660
rect 447060 321570 447088 682654
rect 447508 458856 447560 458862
rect 447508 458798 447560 458804
rect 447416 448520 447468 448526
rect 447416 448462 447468 448468
rect 447232 447908 447284 447914
rect 447232 447850 447284 447856
rect 447140 447840 447192 447846
rect 447140 447782 447192 447788
rect 447152 447370 447180 447782
rect 447244 447438 447272 447850
rect 447232 447432 447284 447438
rect 447232 447374 447284 447380
rect 447140 447364 447192 447370
rect 447140 447306 447192 447312
rect 447428 447302 447456 448462
rect 447416 447296 447468 447302
rect 447414 447264 447416 447273
rect 447468 447264 447470 447273
rect 447414 447199 447470 447208
rect 447140 383648 447192 383654
rect 447138 383616 447140 383625
rect 447192 383616 447194 383625
rect 447138 383551 447194 383560
rect 447232 383580 447284 383586
rect 447232 383522 447284 383528
rect 447244 382945 447272 383522
rect 447230 382936 447286 382945
rect 447230 382871 447286 382880
rect 447138 382256 447194 382265
rect 447138 382191 447194 382200
rect 447232 382220 447284 382226
rect 447152 382158 447180 382191
rect 447232 382162 447284 382168
rect 447140 382152 447192 382158
rect 447140 382094 447192 382100
rect 447244 381585 447272 382162
rect 447230 381576 447286 381585
rect 447230 381511 447286 381520
rect 447230 380896 447286 380905
rect 447230 380831 447286 380840
rect 447416 380860 447468 380866
rect 447140 380792 447192 380798
rect 447140 380734 447192 380740
rect 447152 380225 447180 380734
rect 447244 380730 447272 380831
rect 447416 380802 447468 380808
rect 447232 380724 447284 380730
rect 447232 380666 447284 380672
rect 447138 380216 447194 380225
rect 447138 380151 447194 380160
rect 447428 379545 447456 380802
rect 447414 379536 447470 379545
rect 447324 379500 447376 379506
rect 447414 379471 447470 379480
rect 447324 379442 447376 379448
rect 447140 379432 447192 379438
rect 447140 379374 447192 379380
rect 447152 378865 447180 379374
rect 447138 378856 447194 378865
rect 447138 378791 447194 378800
rect 447336 378185 447364 379442
rect 447322 378176 447378 378185
rect 447232 378140 447284 378146
rect 447322 378111 447378 378120
rect 447232 378082 447284 378088
rect 447140 378072 447192 378078
rect 447140 378014 447192 378020
rect 447152 377505 447180 378014
rect 447138 377496 447194 377505
rect 447138 377431 447194 377440
rect 447244 376825 447272 378082
rect 447230 376816 447286 376825
rect 447230 376751 447286 376760
rect 447140 376712 447192 376718
rect 447140 376654 447192 376660
rect 447152 376145 447180 376654
rect 447232 376644 447284 376650
rect 447232 376586 447284 376592
rect 447138 376136 447194 376145
rect 447138 376071 447194 376080
rect 447244 375465 447272 376586
rect 447230 375456 447286 375465
rect 447230 375391 447286 375400
rect 447140 375352 447192 375358
rect 447140 375294 447192 375300
rect 447152 374785 447180 375294
rect 447232 375284 447284 375290
rect 447232 375226 447284 375232
rect 447138 374776 447194 374785
rect 447138 374711 447194 374720
rect 447244 374105 447272 375226
rect 447230 374096 447286 374105
rect 447230 374031 447286 374040
rect 447140 373992 447192 373998
rect 447140 373934 447192 373940
rect 447152 373425 447180 373934
rect 447232 373924 447284 373930
rect 447232 373866 447284 373872
rect 447138 373416 447194 373425
rect 447138 373351 447194 373360
rect 447244 372745 447272 373866
rect 447230 372736 447286 372745
rect 447230 372671 447286 372680
rect 447140 372564 447192 372570
rect 447140 372506 447192 372512
rect 447152 372065 447180 372506
rect 447232 372496 447284 372502
rect 447232 372438 447284 372444
rect 447138 372056 447194 372065
rect 447138 371991 447194 372000
rect 447244 371385 447272 372438
rect 447230 371376 447286 371385
rect 447230 371311 447286 371320
rect 447140 371204 447192 371210
rect 447140 371146 447192 371152
rect 447152 370705 447180 371146
rect 447232 371136 447284 371142
rect 447232 371078 447284 371084
rect 447138 370696 447194 370705
rect 447138 370631 447194 370640
rect 447244 370025 447272 371078
rect 447230 370016 447286 370025
rect 447230 369951 447286 369960
rect 447140 369844 447192 369850
rect 447140 369786 447192 369792
rect 447152 369345 447180 369786
rect 447232 369776 447284 369782
rect 447232 369718 447284 369724
rect 447138 369336 447194 369345
rect 447138 369271 447194 369280
rect 447244 368665 447272 369718
rect 447230 368656 447286 368665
rect 447230 368591 447286 368600
rect 447140 368484 447192 368490
rect 447140 368426 447192 368432
rect 447152 367985 447180 368426
rect 447232 368416 447284 368422
rect 447232 368358 447284 368364
rect 447138 367976 447194 367985
rect 447138 367911 447194 367920
rect 447244 367305 447272 368358
rect 447230 367296 447286 367305
rect 447230 367231 447286 367240
rect 447140 367056 447192 367062
rect 447140 366998 447192 367004
rect 447152 366625 447180 366998
rect 447232 366988 447284 366994
rect 447232 366930 447284 366936
rect 447138 366616 447194 366625
rect 447138 366551 447194 366560
rect 447244 365945 447272 366930
rect 447230 365936 447286 365945
rect 447230 365871 447286 365880
rect 447140 365696 447192 365702
rect 447140 365638 447192 365644
rect 447152 364585 447180 365638
rect 447232 365628 447284 365634
rect 447232 365570 447284 365576
rect 447244 365265 447272 365570
rect 447230 365256 447286 365265
rect 447230 365191 447286 365200
rect 447138 364576 447194 364585
rect 447138 364511 447194 364520
rect 447230 363896 447286 363905
rect 447230 363831 447286 363840
rect 447138 363216 447194 363225
rect 447138 363151 447194 363160
rect 447152 362982 447180 363151
rect 447244 363050 447272 363831
rect 447232 363044 447284 363050
rect 447232 362986 447284 362992
rect 447140 362976 447192 362982
rect 447140 362918 447192 362924
rect 447138 362536 447194 362545
rect 447138 362471 447194 362480
rect 447152 361622 447180 362471
rect 447230 361856 447286 361865
rect 447230 361791 447286 361800
rect 447244 361690 447272 361791
rect 447232 361684 447284 361690
rect 447232 361626 447284 361632
rect 447140 361616 447192 361622
rect 447140 361558 447192 361564
rect 447230 361176 447286 361185
rect 447230 361111 447286 361120
rect 447138 360496 447194 360505
rect 447138 360431 447194 360440
rect 447152 360262 447180 360431
rect 447244 360330 447272 361111
rect 447232 360324 447284 360330
rect 447232 360266 447284 360272
rect 447140 360256 447192 360262
rect 447140 360198 447192 360204
rect 447138 359816 447194 359825
rect 447138 359751 447194 359760
rect 447152 358834 447180 359751
rect 447230 359136 447286 359145
rect 447230 359071 447286 359080
rect 447244 358902 447272 359071
rect 447232 358896 447284 358902
rect 447232 358838 447284 358844
rect 447140 358828 447192 358834
rect 447140 358770 447192 358776
rect 447520 355065 447548 458798
rect 447796 422385 447824 700266
rect 447888 423026 447916 700402
rect 449164 700392 449216 700398
rect 449164 700334 449216 700340
rect 448336 447908 448388 447914
rect 448336 447850 448388 447856
rect 447968 447840 448020 447846
rect 447968 447782 448020 447788
rect 447876 423020 447928 423026
rect 447876 422962 447928 422968
rect 447782 422376 447838 422385
rect 447782 422311 447838 422320
rect 447784 388612 447836 388618
rect 447784 388554 447836 388560
rect 447692 388544 447744 388550
rect 447692 388486 447744 388492
rect 447506 355056 447562 355065
rect 447506 354991 447562 355000
rect 447704 353705 447732 388486
rect 447796 354385 447824 388554
rect 447876 387252 447928 387258
rect 447876 387194 447928 387200
rect 447782 354376 447838 354385
rect 447782 354311 447838 354320
rect 447690 353696 447746 353705
rect 447690 353631 447746 353640
rect 447888 353025 447916 387194
rect 447874 353016 447930 353025
rect 447874 352951 447930 352960
rect 447784 352572 447836 352578
rect 447784 352514 447836 352520
rect 447322 351656 447378 351665
rect 447322 351591 447378 351600
rect 447138 350976 447194 350985
rect 447138 350911 447194 350920
rect 447152 350606 447180 350911
rect 447140 350600 447192 350606
rect 447140 350542 447192 350548
rect 447140 347744 447192 347750
rect 447140 347686 447192 347692
rect 447152 347585 447180 347686
rect 447138 347576 447194 347585
rect 447138 347511 447194 347520
rect 447138 342136 447194 342145
rect 447138 342071 447194 342080
rect 447152 340950 447180 342071
rect 447230 341456 447286 341465
rect 447230 341391 447286 341400
rect 447244 341018 447272 341391
rect 447232 341012 447284 341018
rect 447232 340954 447284 340960
rect 447140 340944 447192 340950
rect 447140 340886 447192 340892
rect 447230 340776 447286 340785
rect 447230 340711 447286 340720
rect 447138 340096 447194 340105
rect 447138 340031 447194 340040
rect 447152 339590 447180 340031
rect 447140 339584 447192 339590
rect 447140 339526 447192 339532
rect 447244 339522 447272 340711
rect 447232 339516 447284 339522
rect 447232 339458 447284 339464
rect 447230 339416 447286 339425
rect 447230 339351 447286 339360
rect 447138 338736 447194 338745
rect 447138 338671 447194 338680
rect 447152 338230 447180 338671
rect 447140 338224 447192 338230
rect 447140 338166 447192 338172
rect 447244 338162 447272 339351
rect 447232 338156 447284 338162
rect 447232 338098 447284 338104
rect 447138 337376 447194 337385
rect 447138 337311 447194 337320
rect 447152 336326 447180 337311
rect 447140 336320 447192 336326
rect 447140 336262 447192 336268
rect 447138 336016 447194 336025
rect 447138 335951 447194 335960
rect 447152 335714 447180 335951
rect 447140 335708 447192 335714
rect 447140 335650 447192 335656
rect 447230 335336 447286 335345
rect 447230 335271 447286 335280
rect 447138 334656 447194 334665
rect 447138 334591 447194 334600
rect 447152 334014 447180 334591
rect 447244 334082 447272 335271
rect 447232 334076 447284 334082
rect 447232 334018 447284 334024
rect 447140 334008 447192 334014
rect 447140 333950 447192 333956
rect 447230 333976 447286 333985
rect 447230 333911 447286 333920
rect 447138 333296 447194 333305
rect 447138 333231 447194 333240
rect 447152 332654 447180 333231
rect 447244 332722 447272 333911
rect 447232 332716 447284 332722
rect 447232 332658 447284 332664
rect 447140 332648 447192 332654
rect 447140 332590 447192 332596
rect 447138 329896 447194 329905
rect 447138 329831 447140 329840
rect 447192 329831 447194 329840
rect 447140 329802 447192 329808
rect 447048 321564 447100 321570
rect 447048 321506 447100 321512
rect 446956 320816 447008 320822
rect 446956 320758 447008 320764
rect 446864 320068 446916 320074
rect 446864 320010 446916 320016
rect 446770 319696 446826 319705
rect 446770 319631 446826 319640
rect 446680 319048 446732 319054
rect 446680 318990 446732 318996
rect 444288 318708 444340 318714
rect 444288 318650 444340 318656
rect 443828 313948 443880 313954
rect 443828 313890 443880 313896
rect 446128 306332 446180 306338
rect 446128 306274 446180 306280
rect 444748 304564 444800 304570
rect 444748 304506 444800 304512
rect 444760 297226 444788 304506
rect 446140 300694 446168 306274
rect 446128 300688 446180 300694
rect 446128 300630 446180 300636
rect 444748 297220 444800 297226
rect 444748 297162 444800 297168
rect 445024 264988 445076 264994
rect 445024 264930 445076 264936
rect 444656 262268 444708 262274
rect 444656 262210 444708 262216
rect 444668 258738 444696 262210
rect 444656 258732 444708 258738
rect 444656 258674 444708 258680
rect 443736 238740 443788 238746
rect 443736 238682 443788 238688
rect 445036 232966 445064 264930
rect 445024 232960 445076 232966
rect 445024 232902 445076 232908
rect 443644 227724 443696 227730
rect 443644 227666 443696 227672
rect 447336 198014 447364 351591
rect 447506 338056 447562 338065
rect 447506 337991 447562 338000
rect 447414 336696 447470 336705
rect 447414 336631 447470 336640
rect 447428 335374 447456 336631
rect 447416 335368 447468 335374
rect 447416 335310 447468 335316
rect 447520 334966 447548 337991
rect 447692 336116 447744 336122
rect 447692 336058 447744 336064
rect 447508 334960 447560 334966
rect 447508 334902 447560 334908
rect 447704 322182 447732 336058
rect 447796 331265 447824 352514
rect 447874 345536 447930 345545
rect 447874 345471 447930 345480
rect 447782 331256 447838 331265
rect 447782 331191 447838 331200
rect 447692 322176 447744 322182
rect 447692 322118 447744 322124
rect 447888 294506 447916 345471
rect 447980 330585 448008 447782
rect 448060 389836 448112 389842
rect 448060 389778 448112 389784
rect 448072 352345 448100 389778
rect 448348 386714 448376 447850
rect 448980 387184 449032 387190
rect 448980 387126 449032 387132
rect 448336 386708 448388 386714
rect 448336 386650 448388 386656
rect 448244 386028 448296 386034
rect 448244 385970 448296 385976
rect 448152 385416 448204 385422
rect 448152 385358 448204 385364
rect 448058 352336 448114 352345
rect 448058 352271 448114 352280
rect 448164 348945 448192 385358
rect 448150 348936 448206 348945
rect 448150 348871 448206 348880
rect 448256 346905 448284 385970
rect 448242 346896 448298 346905
rect 448242 346831 448298 346840
rect 448348 343482 448376 386650
rect 448428 385688 448480 385694
rect 448428 385630 448480 385636
rect 448440 355745 448468 385630
rect 448992 358465 449020 387126
rect 449070 387016 449126 387025
rect 449070 386951 449126 386960
rect 448978 358456 449034 358465
rect 448978 358391 449034 358400
rect 449084 357105 449112 386951
rect 449070 357096 449126 357105
rect 449070 357031 449126 357040
rect 448426 355736 448482 355745
rect 448426 355671 448482 355680
rect 448428 354000 448480 354006
rect 448428 353942 448480 353948
rect 448440 344865 448468 353942
rect 448426 344856 448482 344865
rect 448426 344791 448482 344800
rect 448426 343496 448482 343505
rect 448348 343454 448426 343482
rect 448426 343431 448482 343440
rect 448440 338094 448468 343431
rect 448428 338088 448480 338094
rect 448428 338030 448480 338036
rect 448428 336728 448480 336734
rect 448428 336670 448480 336676
rect 448058 332616 448114 332625
rect 448058 332551 448114 332560
rect 447966 330576 448022 330585
rect 447966 330511 447968 330520
rect 448020 330511 448022 330520
rect 447968 330482 448020 330488
rect 447876 294500 447928 294506
rect 447876 294442 447928 294448
rect 447784 289604 447836 289610
rect 447784 289546 447836 289552
rect 447796 262274 447824 289546
rect 447876 279540 447928 279546
rect 447876 279482 447928 279488
rect 447888 264994 447916 279482
rect 447876 264988 447928 264994
rect 447876 264930 447928 264936
rect 447784 262268 447836 262274
rect 447784 262210 447836 262216
rect 447324 198008 447376 198014
rect 447324 197950 447376 197956
rect 448072 183530 448100 332551
rect 448242 331936 448298 331945
rect 448242 331871 448298 331880
rect 447600 183524 447652 183530
rect 447600 183466 447652 183472
rect 448060 183524 448112 183530
rect 448060 183466 448112 183472
rect 447612 182850 447640 183466
rect 447600 182844 447652 182850
rect 447600 182786 447652 182792
rect 448256 172514 448284 331871
rect 448334 331256 448390 331265
rect 448334 331191 448390 331200
rect 447600 172508 447652 172514
rect 447600 172450 447652 172456
rect 448244 172508 448296 172514
rect 448244 172450 448296 172456
rect 447612 171834 447640 172450
rect 447600 171828 447652 171834
rect 447600 171770 447652 171776
rect 445208 162172 445260 162178
rect 445208 162114 445260 162120
rect 441574 160132 441626 160138
rect 441574 160074 441626 160080
rect 442908 160132 442960 160138
rect 442908 160074 442960 160080
rect 441586 159868 441614 160074
rect 445220 159882 445248 162114
rect 448348 161430 448376 331191
rect 448336 161424 448388 161430
rect 448336 161366 448388 161372
rect 448348 160750 448376 161366
rect 448336 160744 448388 160750
rect 448336 160686 448388 160692
rect 448440 159882 448468 336670
rect 449176 321473 449204 700334
rect 449162 321464 449218 321473
rect 449268 321434 449296 700742
rect 449348 685160 449400 685166
rect 449348 685102 449400 685108
rect 449162 321399 449218 321408
rect 449256 321428 449308 321434
rect 449256 321370 449308 321376
rect 449360 319569 449388 685102
rect 462332 670585 462360 703520
rect 478524 700466 478552 703520
rect 478512 700460 478564 700466
rect 478512 700402 478564 700408
rect 494808 700330 494836 703520
rect 494796 700324 494848 700330
rect 494796 700266 494848 700272
rect 527192 699825 527220 703520
rect 543476 700369 543504 703520
rect 543462 700360 543518 700369
rect 543462 700295 543518 700304
rect 559668 699825 559696 703520
rect 527178 699816 527234 699825
rect 527178 699751 527234 699760
rect 559654 699816 559710 699825
rect 559654 699751 559710 699760
rect 580262 697232 580318 697241
rect 580262 697167 580318 697176
rect 579618 683904 579674 683913
rect 579618 683839 579674 683848
rect 579632 683194 579660 683839
rect 576124 683188 576176 683194
rect 576124 683130 576176 683136
rect 579620 683188 579672 683194
rect 579620 683130 579672 683136
rect 462318 670576 462374 670585
rect 462318 670511 462374 670520
rect 457902 667992 457958 668001
rect 457902 667927 457958 667936
rect 457718 657520 457774 657529
rect 457718 657455 457774 657464
rect 457626 650176 457682 650185
rect 457626 650111 457682 650120
rect 457534 645960 457590 645969
rect 457534 645895 457590 645904
rect 457442 643240 457498 643249
rect 457442 643175 457498 643184
rect 457350 640384 457406 640393
rect 457350 640319 457406 640328
rect 457258 635488 457314 635497
rect 457258 635423 457314 635432
rect 457272 598738 457300 635423
rect 457364 600234 457392 640319
rect 457352 600228 457404 600234
rect 457352 600170 457404 600176
rect 457456 599622 457484 643175
rect 457548 599826 457576 645895
rect 457536 599820 457588 599826
rect 457536 599762 457588 599768
rect 457444 599616 457496 599622
rect 457444 599558 457496 599564
rect 457260 598732 457312 598738
rect 457260 598674 457312 598680
rect 450544 596828 450596 596834
rect 450544 596770 450596 596776
rect 449716 518220 449768 518226
rect 449716 518162 449768 518168
rect 449728 503509 449756 518162
rect 449808 517608 449860 517614
rect 449808 517550 449860 517556
rect 449714 503500 449770 503509
rect 449714 503435 449770 503444
rect 449716 454776 449768 454782
rect 449716 454718 449768 454724
rect 449624 454708 449676 454714
rect 449624 454650 449676 454656
rect 449532 387116 449584 387122
rect 449532 387058 449584 387064
rect 449440 385144 449492 385150
rect 449440 385086 449492 385092
rect 449452 348265 449480 385086
rect 449438 348256 449494 348265
rect 449438 348191 449494 348200
rect 449544 342825 449572 387058
rect 449636 357785 449664 454650
rect 449622 357776 449678 357785
rect 449622 357711 449678 357720
rect 449728 356425 449756 454718
rect 449714 356416 449770 356425
rect 449714 356351 449770 356360
rect 449714 350296 449770 350305
rect 449714 350231 449770 350240
rect 449728 345014 449756 350231
rect 449820 349625 449848 517550
rect 450360 517540 450412 517546
rect 450360 517482 450412 517488
rect 449992 516792 450044 516798
rect 449992 516734 450044 516740
rect 450004 507657 450032 516734
rect 450372 510241 450400 517482
rect 450450 516896 450506 516905
rect 450450 516831 450506 516840
rect 450464 514729 450492 516831
rect 450450 514720 450506 514729
rect 450450 514655 450506 514664
rect 450556 512417 450584 596770
rect 457640 595474 457668 650111
rect 457732 598262 457760 657455
rect 457810 652896 457866 652905
rect 457810 652831 457866 652840
rect 457720 598256 457772 598262
rect 457720 598198 457772 598204
rect 457628 595468 457680 595474
rect 457628 595410 457680 595416
rect 457824 594114 457852 652831
rect 457916 595950 457944 667927
rect 458086 662552 458142 662561
rect 458086 662487 458142 662496
rect 457994 659968 458050 659977
rect 457994 659903 458050 659912
rect 457904 595944 457956 595950
rect 457904 595886 457956 595892
rect 457812 594108 457864 594114
rect 457812 594050 457864 594056
rect 458008 522374 458036 659903
rect 457996 522368 458048 522374
rect 457996 522310 458048 522316
rect 458100 519654 458128 662487
rect 459098 637936 459154 637945
rect 459098 637871 459154 637880
rect 459006 633448 459062 633457
rect 459006 633383 459062 633392
rect 458822 630728 458878 630737
rect 458822 630663 458878 630672
rect 458638 611416 458694 611425
rect 458638 611351 458694 611360
rect 458652 598330 458680 611351
rect 458836 604178 458864 630663
rect 458914 621072 458970 621081
rect 458914 621007 458970 621016
rect 458824 604172 458876 604178
rect 458824 604114 458876 604120
rect 458928 604058 458956 621007
rect 458744 604030 458956 604058
rect 458744 599690 458772 604030
rect 458824 603968 458876 603974
rect 459020 603922 459048 633383
rect 458824 603910 458876 603916
rect 458732 599684 458784 599690
rect 458732 599626 458784 599632
rect 458640 598324 458692 598330
rect 458640 598266 458692 598272
rect 458088 519648 458140 519654
rect 458088 519590 458140 519596
rect 458836 518265 458864 603910
rect 458928 603894 459048 603922
rect 458928 599593 458956 603894
rect 459008 603764 459060 603770
rect 459008 603706 459060 603712
rect 459020 599758 459048 603706
rect 459008 599752 459060 599758
rect 459008 599694 459060 599700
rect 458914 599584 458970 599593
rect 458914 599519 458970 599528
rect 459112 543017 459140 637871
rect 459374 628144 459430 628153
rect 459374 628079 459430 628088
rect 459282 625832 459338 625841
rect 459282 625767 459338 625776
rect 459190 623928 459246 623937
rect 459190 623863 459246 623872
rect 459098 543008 459154 543017
rect 459098 542943 459154 542952
rect 459204 522306 459232 623863
rect 459192 522300 459244 522306
rect 459192 522242 459244 522248
rect 459296 520946 459324 625767
rect 459284 520940 459336 520946
rect 459284 520882 459336 520888
rect 459388 519586 459416 628079
rect 460202 618352 460258 618361
rect 460202 618287 460258 618296
rect 459466 616040 459522 616049
rect 459466 615975 459522 615984
rect 459480 603770 459508 615975
rect 460110 613864 460166 613873
rect 460110 613799 460166 613808
rect 460018 608696 460074 608705
rect 460018 608631 460074 608640
rect 459926 606384 459982 606393
rect 459926 606319 459982 606328
rect 459468 603764 459520 603770
rect 459468 603706 459520 603712
rect 459466 603664 459522 603673
rect 459466 603599 459522 603608
rect 459480 598466 459508 603599
rect 459836 602132 459888 602138
rect 459836 602074 459888 602080
rect 459468 598460 459520 598466
rect 459468 598402 459520 598408
rect 459848 596902 459876 602074
rect 459836 596896 459888 596902
rect 459836 596838 459888 596844
rect 459940 543046 459968 606319
rect 460032 594182 460060 608631
rect 460124 602138 460152 613799
rect 460112 602132 460164 602138
rect 460112 602074 460164 602080
rect 460110 602032 460166 602041
rect 460110 601967 460166 601976
rect 460124 600302 460152 601967
rect 460112 600296 460164 600302
rect 460112 600238 460164 600244
rect 460216 595542 460244 618287
rect 570604 616888 570656 616894
rect 570604 616830 570656 616836
rect 462320 600296 462372 600302
rect 462320 600238 462372 600244
rect 461584 598732 461636 598738
rect 461584 598674 461636 598680
rect 460204 595536 460256 595542
rect 460204 595478 460256 595484
rect 460020 594176 460072 594182
rect 460020 594118 460072 594124
rect 459928 543040 459980 543046
rect 459928 542982 459980 542988
rect 459376 519580 459428 519586
rect 459376 519522 459428 519528
rect 458822 518256 458878 518265
rect 458822 518191 458878 518200
rect 450636 516860 450688 516866
rect 450636 516802 450688 516808
rect 450542 512408 450598 512417
rect 450542 512343 450598 512352
rect 450358 510232 450414 510241
rect 450358 510167 450414 510176
rect 450372 509234 450400 510167
rect 450372 509206 450492 509234
rect 449990 507648 450046 507657
rect 449990 507583 450046 507592
rect 449806 349616 449862 349625
rect 449806 349551 449862 349560
rect 449728 344986 449848 345014
rect 449714 344176 449770 344185
rect 449714 344111 449770 344120
rect 449530 342816 449586 342825
rect 449530 342751 449586 342760
rect 449440 338088 449492 338094
rect 449440 338030 449492 338036
rect 449346 319560 449402 319569
rect 449346 319495 449402 319504
rect 449452 249082 449480 338030
rect 449728 336734 449756 344111
rect 449716 336728 449768 336734
rect 449716 336670 449768 336676
rect 449532 336252 449584 336258
rect 449532 336194 449584 336200
rect 449544 318782 449572 336194
rect 449624 336184 449676 336190
rect 449624 336126 449676 336132
rect 449636 319802 449664 336126
rect 449716 334620 449768 334626
rect 449716 334562 449768 334568
rect 449728 322386 449756 334562
rect 449716 322380 449768 322386
rect 449716 322322 449768 322328
rect 449624 319796 449676 319802
rect 449624 319738 449676 319744
rect 449532 318776 449584 318782
rect 449532 318718 449584 318724
rect 449820 263566 449848 344986
rect 450004 334121 450032 507583
rect 450082 505472 450138 505481
rect 450082 505407 450138 505416
rect 450096 337482 450124 505407
rect 450174 503296 450230 503305
rect 450174 503231 450230 503240
rect 450084 337476 450136 337482
rect 450084 337418 450136 337424
rect 450188 336870 450216 503231
rect 450266 337784 450322 337793
rect 450266 337719 450322 337728
rect 450280 337113 450308 337719
rect 450360 337476 450412 337482
rect 450360 337418 450412 337424
rect 450266 337104 450322 337113
rect 450266 337039 450322 337048
rect 450176 336864 450228 336870
rect 450176 336806 450228 336812
rect 449990 334112 450046 334121
rect 449990 334047 450046 334056
rect 449898 328944 449954 328953
rect 449898 328879 449954 328888
rect 449912 328574 449940 328879
rect 449900 328568 449952 328574
rect 449900 328510 449952 328516
rect 450004 326641 450032 334047
rect 450084 330540 450136 330546
rect 450084 330482 450136 330488
rect 449990 326632 450046 326641
rect 449990 326567 450046 326576
rect 450096 324601 450124 330482
rect 450188 324850 450216 336806
rect 450280 328001 450308 337039
rect 450372 336938 450400 337418
rect 450360 336932 450412 336938
rect 450360 336874 450412 336880
rect 450266 327992 450322 328001
rect 450266 327927 450322 327936
rect 450372 325694 450400 336874
rect 450464 335354 450492 509206
rect 450556 462398 450584 512343
rect 450648 505481 450676 516802
rect 450634 505472 450690 505481
rect 450634 505407 450690 505416
rect 450648 500126 450754 500154
rect 451936 500126 452226 500154
rect 450544 462392 450596 462398
rect 450544 462334 450596 462340
rect 450556 337793 450584 462334
rect 450648 402974 450676 500126
rect 450648 402946 450860 402974
rect 450728 388476 450780 388482
rect 450728 388418 450780 388424
rect 450542 337784 450598 337793
rect 450542 337719 450598 337728
rect 450740 336802 450768 388418
rect 450832 385900 450860 402946
rect 451936 385914 451964 500126
rect 453684 496874 453712 500140
rect 454052 500126 455170 500154
rect 453948 496936 454000 496942
rect 453948 496878 454000 496884
rect 452568 496868 452620 496874
rect 452568 496810 452620 496816
rect 453672 496868 453724 496874
rect 453672 496810 453724 496816
rect 452016 455456 452068 455462
rect 452016 455398 452068 455404
rect 451582 385886 451964 385914
rect 452028 385422 452056 455398
rect 452580 385914 452608 496810
rect 453304 462460 453356 462466
rect 453304 462402 453356 462408
rect 453028 389156 453080 389162
rect 453028 389098 453080 389104
rect 452318 385886 452608 385914
rect 453040 385900 453068 389098
rect 453316 386034 453344 462402
rect 453304 386028 453356 386034
rect 453304 385970 453356 385976
rect 453960 385914 453988 496878
rect 454052 389162 454080 500126
rect 454684 497480 454736 497486
rect 454684 497422 454736 497428
rect 454696 393314 454724 497422
rect 455328 497072 455380 497078
rect 455328 497014 455380 497020
rect 455144 496868 455196 496874
rect 455144 496810 455196 496816
rect 455156 393314 455184 496810
rect 455340 393314 455368 497014
rect 456524 497004 456576 497010
rect 456524 496946 456576 496952
rect 456536 393314 456564 496946
rect 456628 496942 456656 500140
rect 457536 497616 457588 497622
rect 457536 497558 457588 497564
rect 457444 497548 457496 497554
rect 457444 497490 457496 497496
rect 456616 496936 456668 496942
rect 456616 496878 456668 496884
rect 454420 393286 454724 393314
rect 454880 393286 455184 393314
rect 455248 393286 455368 393314
rect 456352 393286 456564 393314
rect 454040 389156 454092 389162
rect 454040 389098 454092 389104
rect 453790 385886 453988 385914
rect 454420 385694 454448 393286
rect 454880 385914 454908 393286
rect 454526 385886 454908 385914
rect 455248 385900 455276 393286
rect 456352 385914 456380 393286
rect 456708 389156 456760 389162
rect 456708 389098 456760 389104
rect 455998 385886 456380 385914
rect 456720 385900 456748 389098
rect 457456 388618 457484 497490
rect 457444 388612 457496 388618
rect 457444 388554 457496 388560
rect 457548 388550 457576 497558
rect 458100 496874 458128 500140
rect 458824 497684 458876 497690
rect 458824 497626 458876 497632
rect 458088 496868 458140 496874
rect 458088 496810 458140 496816
rect 458088 430024 458140 430030
rect 458088 429966 458140 429972
rect 457628 428460 457680 428466
rect 457628 428402 457680 428408
rect 457640 389162 457668 428402
rect 458100 393314 458128 429966
rect 457824 393286 458128 393314
rect 457628 389156 457680 389162
rect 457628 389098 457680 389104
rect 457536 388544 457588 388550
rect 457536 388486 457588 388492
rect 457824 385914 457852 393286
rect 458456 389292 458508 389298
rect 458456 389234 458508 389240
rect 458468 385914 458496 389234
rect 458836 387258 458864 497626
rect 459572 497078 459600 500140
rect 459560 497072 459612 497078
rect 459560 497014 459612 497020
rect 461044 497010 461072 500140
rect 461032 497004 461084 497010
rect 461032 496946 461084 496952
rect 458916 460964 458968 460970
rect 458916 460906 458968 460912
rect 458928 448526 458956 460906
rect 459008 454096 459060 454102
rect 459008 454038 459060 454044
rect 458916 448520 458968 448526
rect 458916 448462 458968 448468
rect 459020 447914 459048 454038
rect 459008 447908 459060 447914
rect 459008 447850 459060 447856
rect 459468 429956 459520 429962
rect 459468 429898 459520 429904
rect 459376 429888 459428 429894
rect 459376 429830 459428 429836
rect 459388 393314 459416 429830
rect 459296 393286 459416 393314
rect 458824 387252 458876 387258
rect 458824 387194 458876 387200
rect 459296 385914 459324 393286
rect 459480 389298 459508 429898
rect 460756 395344 460808 395350
rect 460756 395286 460808 395292
rect 459652 389904 459704 389910
rect 459652 389846 459704 389852
rect 459468 389292 459520 389298
rect 459468 389234 459520 389240
rect 457470 385886 457852 385914
rect 458206 385886 458496 385914
rect 458942 385886 459324 385914
rect 459664 385900 459692 389846
rect 460768 385914 460796 395286
rect 461596 388890 461624 598674
rect 461676 595944 461728 595950
rect 461676 595886 461728 595892
rect 461584 388884 461636 388890
rect 461584 388826 461636 388832
rect 461124 388816 461176 388822
rect 461124 388758 461176 388764
rect 460414 385886 460796 385914
rect 461136 385900 461164 388758
rect 461688 387938 461716 595886
rect 461768 455524 461820 455530
rect 461768 455466 461820 455472
rect 461780 388482 461808 455466
rect 462332 402974 462360 600238
rect 462964 600228 463016 600234
rect 462964 600170 463016 600176
rect 462332 402946 462912 402974
rect 461768 388476 461820 388482
rect 461768 388418 461820 388424
rect 461676 387932 461728 387938
rect 461676 387874 461728 387880
rect 462596 387932 462648 387938
rect 462596 387874 462648 387880
rect 461860 387864 461912 387870
rect 461860 387806 461912 387812
rect 461872 385900 461900 387806
rect 462608 385900 462636 387874
rect 462884 385914 462912 402946
rect 462976 388754 463004 600170
rect 463160 600086 463266 600114
rect 469614 600086 469904 600114
rect 475962 600086 476068 600114
rect 463054 517576 463110 517585
rect 463054 517511 463110 517520
rect 462964 388748 463016 388754
rect 462964 388690 463016 388696
rect 463068 388482 463096 517511
rect 463160 501129 463188 600086
rect 464344 599820 464396 599826
rect 464344 599762 464396 599768
rect 463700 598460 463752 598466
rect 463700 598402 463752 598408
rect 463146 501120 463202 501129
rect 463146 501055 463202 501064
rect 463148 497752 463200 497758
rect 463148 497694 463200 497700
rect 463160 389842 463188 497694
rect 463608 392624 463660 392630
rect 463608 392566 463660 392572
rect 463148 389836 463200 389842
rect 463148 389778 463200 389784
rect 463620 388822 463648 392566
rect 463608 388816 463660 388822
rect 463608 388758 463660 388764
rect 463056 388476 463108 388482
rect 463056 388418 463108 388424
rect 463712 385914 463740 598402
rect 463792 543040 463844 543046
rect 463792 542982 463844 542988
rect 463804 402974 463832 542982
rect 463804 402946 464292 402974
rect 464264 386050 464292 402946
rect 464356 388822 464384 599762
rect 466460 599752 466512 599758
rect 466460 599694 466512 599700
rect 465080 598324 465132 598330
rect 465080 598266 465132 598272
rect 464436 522368 464488 522374
rect 464436 522310 464488 522316
rect 464448 402974 464476 522310
rect 464448 402946 464568 402974
rect 464344 388816 464396 388822
rect 464344 388758 464396 388764
rect 464540 388550 464568 402946
rect 464896 389836 464948 389842
rect 464896 389778 464948 389784
rect 464528 388544 464580 388550
rect 464528 388486 464580 388492
rect 464908 387870 464936 389778
rect 465092 389298 465120 598266
rect 465724 598256 465776 598262
rect 465724 598198 465776 598204
rect 465172 594176 465224 594182
rect 465172 594118 465224 594124
rect 465080 389292 465132 389298
rect 465080 389234 465132 389240
rect 464896 387864 464948 387870
rect 464896 387806 464948 387812
rect 464264 386022 464384 386050
rect 464356 385914 464384 386022
rect 465184 385914 465212 594118
rect 465736 388618 465764 598198
rect 466472 389298 466500 599694
rect 469220 599684 469272 599690
rect 469220 599626 469272 599632
rect 468484 599616 468536 599622
rect 468484 599558 468536 599564
rect 466552 596896 466604 596902
rect 466552 596838 466604 596844
rect 465908 389292 465960 389298
rect 465908 389234 465960 389240
rect 466460 389292 466512 389298
rect 466460 389234 466512 389240
rect 465724 388612 465776 388618
rect 465724 388554 465776 388560
rect 465920 385914 465948 389234
rect 466564 385914 466592 596838
rect 467932 595536 467984 595542
rect 467932 595478 467984 595484
rect 467104 594108 467156 594114
rect 467104 594050 467156 594056
rect 467116 388958 467144 594050
rect 467196 461032 467248 461038
rect 467196 460974 467248 460980
rect 467208 447846 467236 460974
rect 467196 447840 467248 447846
rect 467196 447782 467248 447788
rect 467944 402974 467972 595478
rect 467944 402946 468064 402974
rect 467380 389292 467432 389298
rect 467380 389234 467432 389240
rect 467104 388952 467156 388958
rect 467104 388894 467156 388900
rect 467392 385914 467420 389234
rect 468036 385914 468064 402946
rect 468496 389094 468524 599558
rect 468576 595468 468628 595474
rect 468576 595410 468628 595416
rect 468484 389088 468536 389094
rect 468484 389030 468536 389036
rect 468588 389026 468616 595410
rect 468668 519648 468720 519654
rect 468668 519590 468720 519596
rect 468576 389020 468628 389026
rect 468576 388962 468628 388968
rect 468680 388686 468708 519590
rect 468668 388680 468720 388686
rect 468668 388622 468720 388628
rect 462884 385886 463358 385914
rect 463712 385886 464094 385914
rect 464356 385886 464830 385914
rect 465184 385886 465566 385914
rect 465920 385886 466302 385914
rect 466564 385886 467038 385914
rect 467392 385886 467774 385914
rect 468036 385886 468510 385914
rect 469232 385900 469260 599626
rect 469404 522300 469456 522306
rect 469404 522242 469456 522248
rect 469416 402974 469444 522242
rect 469876 518226 469904 600086
rect 470600 520940 470652 520946
rect 470600 520882 470652 520888
rect 469864 518220 469916 518226
rect 469864 518162 469916 518168
rect 469416 402946 469536 402974
rect 469508 385914 469536 402946
rect 470612 385914 470640 520882
rect 470876 519580 470928 519586
rect 470876 519522 470928 519528
rect 470888 402974 470916 519522
rect 476040 517682 476068 600086
rect 476028 517676 476080 517682
rect 476028 517618 476080 517624
rect 476040 516866 476068 517618
rect 482296 517478 482324 600100
rect 488644 598330 488672 600100
rect 488632 598324 488684 598330
rect 488632 598266 488684 598272
rect 494336 598324 494388 598330
rect 494336 598266 494388 598272
rect 493324 598256 493376 598262
rect 493324 598198 493376 598204
rect 482928 520940 482980 520946
rect 482928 520882 482980 520888
rect 482742 517576 482798 517585
rect 482940 517562 482968 520882
rect 488632 517608 488684 517614
rect 482798 517534 483000 517562
rect 488684 517556 488980 517562
rect 488632 517550 488980 517556
rect 488644 517534 488980 517550
rect 482742 517511 482798 517520
rect 482284 517472 482336 517478
rect 482284 517414 482336 517420
rect 476028 516860 476080 516866
rect 476028 516802 476080 516808
rect 492128 516792 492180 516798
rect 492128 516734 492180 516740
rect 492140 512650 492168 516734
rect 492128 512644 492180 512650
rect 492128 512586 492180 512592
rect 492140 512485 492168 512586
rect 492126 512476 492182 512485
rect 492126 512411 492182 512420
rect 480272 500126 480608 500154
rect 481652 500126 481804 500154
rect 482664 500126 483000 500154
rect 483860 500126 484196 500154
rect 485056 500126 485392 500154
rect 486252 500126 486588 500154
rect 487172 500126 487784 500154
rect 488980 500126 489224 500154
rect 480272 497758 480300 500126
rect 480260 497752 480312 497758
rect 480260 497694 480312 497700
rect 481652 497690 481680 500126
rect 481640 497684 481692 497690
rect 481640 497626 481692 497632
rect 482664 497622 482692 500126
rect 482652 497616 482704 497622
rect 482652 497558 482704 497564
rect 483860 497554 483888 500126
rect 483848 497548 483900 497554
rect 483848 497490 483900 497496
rect 485056 496874 485084 500126
rect 486252 497486 486280 500126
rect 486240 497480 486292 497486
rect 486240 497422 486292 497428
rect 483664 496868 483716 496874
rect 483664 496810 483716 496816
rect 485044 496868 485096 496874
rect 485044 496810 485096 496816
rect 473726 462904 473782 462913
rect 473726 462839 473782 462848
rect 473740 454102 473768 462839
rect 483676 458862 483704 496810
rect 483664 458856 483716 458862
rect 483664 458798 483716 458804
rect 480996 455456 481048 455462
rect 480996 455398 481048 455404
rect 473728 454096 473780 454102
rect 473728 454038 473780 454044
rect 473740 453900 473768 454038
rect 481008 453900 481036 455398
rect 487172 454782 487200 500126
rect 489196 496913 489224 500126
rect 489932 500126 490176 500154
rect 491312 500126 491372 500154
rect 489182 496904 489238 496913
rect 489182 496839 489238 496848
rect 488264 456068 488316 456074
rect 488264 456010 488316 456016
rect 488276 455530 488304 456010
rect 488264 455524 488316 455530
rect 488264 455466 488316 455472
rect 487160 454776 487212 454782
rect 487160 454718 487212 454724
rect 488276 453900 488304 455466
rect 489932 454714 489960 500126
rect 489920 454708 489972 454714
rect 489920 454650 489972 454656
rect 471624 428466 471652 432140
rect 474292 430030 474320 432140
rect 474280 430024 474332 430030
rect 474280 429966 474332 429972
rect 476960 429962 476988 432140
rect 476948 429956 477000 429962
rect 476948 429898 477000 429904
rect 479628 429894 479656 432140
rect 479616 429888 479668 429894
rect 479616 429830 479668 429836
rect 482296 429214 482324 432140
rect 484964 429214 484992 432140
rect 487172 432126 487646 432154
rect 489932 432126 490314 432154
rect 480904 429208 480956 429214
rect 480904 429150 480956 429156
rect 482284 429208 482336 429214
rect 482284 429150 482336 429156
rect 483664 429208 483716 429214
rect 483664 429150 483716 429156
rect 484952 429208 485004 429214
rect 484952 429150 485004 429156
rect 476118 428496 476174 428505
rect 471612 428460 471664 428466
rect 476118 428431 476174 428440
rect 471612 428402 471664 428408
rect 476132 402974 476160 428431
rect 470888 402946 471008 402974
rect 476132 402946 476896 402974
rect 470980 385914 471008 402946
rect 475844 389088 475896 389094
rect 472162 389056 472218 389065
rect 472162 388991 472218 389000
rect 474370 389056 474426 389065
rect 475844 389030 475896 389036
rect 474370 388991 474426 389000
rect 469508 385886 469982 385914
rect 470612 385886 470718 385914
rect 470980 385886 471454 385914
rect 472176 385900 472204 388991
rect 472898 388920 472954 388929
rect 472898 388855 472954 388864
rect 473636 388884 473688 388890
rect 472912 385900 472940 388855
rect 473636 388826 473688 388832
rect 473648 385900 473676 388826
rect 474384 385900 474412 388991
rect 475108 388748 475160 388754
rect 475108 388690 475160 388696
rect 475120 385900 475148 388690
rect 475856 385900 475884 389030
rect 476580 388816 476632 388822
rect 476580 388758 476632 388764
rect 476592 385900 476620 388758
rect 476868 385914 476896 402946
rect 480916 389910 480944 429150
rect 483676 395350 483704 429150
rect 487068 423360 487120 423366
rect 487068 423302 487120 423308
rect 484308 421592 484360 421598
rect 484308 421534 484360 421540
rect 483664 395344 483716 395350
rect 483664 395286 483716 395292
rect 484320 393314 484348 421534
rect 486976 416084 487028 416090
rect 486976 416026 487028 416032
rect 486988 393314 487016 416026
rect 483584 393286 484348 393314
rect 486896 393286 487016 393314
rect 480904 389904 480956 389910
rect 480904 389846 480956 389852
rect 479522 389056 479578 389065
rect 478052 389020 478104 389026
rect 479522 388991 479578 389000
rect 478052 388962 478104 388968
rect 476868 385886 477342 385914
rect 478064 385900 478092 388962
rect 478788 388952 478840 388958
rect 478788 388894 478840 388900
rect 478800 385900 478828 388894
rect 479536 385900 479564 388991
rect 481732 388680 481784 388686
rect 481732 388622 481784 388628
rect 480260 388612 480312 388618
rect 480260 388554 480312 388560
rect 480272 385900 480300 388554
rect 480996 388544 481048 388550
rect 480996 388486 481048 388492
rect 481008 385900 481036 388486
rect 481744 385900 481772 388622
rect 482468 388476 482520 388482
rect 482468 388418 482520 388424
rect 482480 385900 482508 388418
rect 483584 385914 483612 393286
rect 486424 389292 486476 389298
rect 486424 389234 486476 389240
rect 483940 388884 483992 388890
rect 483940 388826 483992 388832
rect 483230 385886 483612 385914
rect 483952 385900 483980 388826
rect 484676 388680 484728 388686
rect 484676 388622 484728 388628
rect 484688 385900 484716 388622
rect 485412 388612 485464 388618
rect 485412 388554 485464 388560
rect 485424 385900 485452 388554
rect 486436 385914 486464 389234
rect 486174 385886 486464 385914
rect 486896 385900 486924 393286
rect 487080 389298 487108 423302
rect 487172 392630 487200 432126
rect 488264 423292 488316 423298
rect 488264 423234 488316 423240
rect 488276 393314 488304 423234
rect 489644 423224 489696 423230
rect 489644 423166 489696 423172
rect 489656 393314 489684 423166
rect 488000 393286 488304 393314
rect 489472 393286 489684 393314
rect 487160 392624 487212 392630
rect 487160 392566 487212 392572
rect 487068 389292 487120 389298
rect 487068 389234 487120 389240
rect 488000 385914 488028 393286
rect 488356 388544 488408 388550
rect 488356 388486 488408 388492
rect 487646 385886 488028 385914
rect 488368 385900 488396 388486
rect 489472 385914 489500 393286
rect 489932 389842 489960 432126
rect 489920 389836 489972 389842
rect 489920 389778 489972 389784
rect 490564 389836 490616 389842
rect 490564 389778 490616 389784
rect 489828 388476 489880 388482
rect 489828 388418 489880 388424
rect 489118 385886 489500 385914
rect 489840 385900 489868 388418
rect 490576 385900 490604 389778
rect 491312 387190 491340 500126
rect 492404 395344 492456 395350
rect 492404 395286 492456 395292
rect 491576 392624 491628 392630
rect 491576 392566 491628 392572
rect 491300 387184 491352 387190
rect 491300 387126 491352 387132
rect 491588 385914 491616 392566
rect 492416 385914 492444 395286
rect 493336 392601 493364 598198
rect 494244 518220 494296 518226
rect 494244 518162 494296 518168
rect 494152 517676 494204 517682
rect 494152 517618 494204 517624
rect 494164 508881 494192 517618
rect 494150 508872 494206 508881
rect 494150 508807 494206 508816
rect 494164 508570 494192 508807
rect 494152 508564 494204 508570
rect 494152 508506 494204 508512
rect 494256 505753 494284 518162
rect 494348 517546 494376 598266
rect 494992 596834 495020 600100
rect 500972 600086 501354 600114
rect 507136 600086 507702 600114
rect 513392 600086 514050 600114
rect 520292 600086 520398 600114
rect 494980 596828 495032 596834
rect 494980 596770 495032 596776
rect 494336 517540 494388 517546
rect 494336 517482 494388 517488
rect 494348 515953 494376 517482
rect 500972 516905 501000 600086
rect 500958 516896 501014 516905
rect 500958 516831 501014 516840
rect 502246 516896 502302 516905
rect 502246 516831 502302 516840
rect 494334 515944 494390 515953
rect 494334 515879 494390 515888
rect 494348 509930 494376 515879
rect 502260 514078 502288 516831
rect 507136 516769 507164 600086
rect 511264 590708 511316 590714
rect 511264 590650 511316 590656
rect 510618 518120 510674 518129
rect 510618 518055 510674 518064
rect 507122 516760 507178 516769
rect 507122 516695 507178 516704
rect 502248 514072 502300 514078
rect 502248 514014 502300 514020
rect 494336 509924 494388 509930
rect 494336 509866 494388 509872
rect 495072 505776 495124 505782
rect 494242 505744 494298 505753
rect 494242 505679 494298 505688
rect 495070 505744 495072 505753
rect 495124 505744 495126 505753
rect 495070 505679 495126 505688
rect 494702 501256 494758 501265
rect 494702 501191 494758 501200
rect 494716 462534 494744 501191
rect 494704 462528 494756 462534
rect 494704 462470 494756 462476
rect 494716 456074 494744 462470
rect 494704 456068 494756 456074
rect 494704 456010 494756 456016
rect 503628 424380 503680 424386
rect 503628 424322 503680 424328
rect 502984 423428 503036 423434
rect 502984 423370 503036 423376
rect 498108 423156 498160 423162
rect 498108 423098 498160 423104
rect 495348 420232 495400 420238
rect 495348 420174 495400 420180
rect 494612 399492 494664 399498
rect 494612 399434 494664 399440
rect 493968 398132 494020 398138
rect 493968 398074 494020 398080
rect 493416 396772 493468 396778
rect 493416 396714 493468 396720
rect 493322 392592 493378 392601
rect 493322 392527 493378 392536
rect 493428 386050 493456 396714
rect 493152 386022 493456 386050
rect 493152 385914 493180 386022
rect 493980 385914 494008 398074
rect 494624 385914 494652 399434
rect 495360 385914 495388 420174
rect 497924 400920 497976 400926
rect 497924 400862 497976 400868
rect 496728 394052 496780 394058
rect 496728 393994 496780 394000
rect 495716 391332 495768 391338
rect 495716 391274 495768 391280
rect 491326 385886 491616 385914
rect 492062 385886 492444 385914
rect 492798 385886 493180 385914
rect 493534 385886 494008 385914
rect 494270 385886 494652 385914
rect 495006 385886 495388 385914
rect 495728 385900 495756 391274
rect 496740 385914 496768 393994
rect 497464 389292 497516 389298
rect 497464 389234 497516 389240
rect 497476 385914 497504 389234
rect 496478 385886 496768 385914
rect 497214 385886 497504 385914
rect 497936 385900 497964 400862
rect 498120 389298 498148 423098
rect 499304 423088 499356 423094
rect 499304 423030 499356 423036
rect 499316 393314 499344 423030
rect 500684 423020 500736 423026
rect 500684 422962 500736 422968
rect 500696 393314 500724 422962
rect 502248 422952 502300 422958
rect 502248 422894 502300 422900
rect 502260 393314 502288 422894
rect 499040 393286 499344 393314
rect 500512 393286 500724 393314
rect 501984 393286 502288 393314
rect 498108 389292 498160 389298
rect 498108 389234 498160 389240
rect 499040 385914 499068 393286
rect 499396 388748 499448 388754
rect 499396 388690 499448 388696
rect 498686 385886 499068 385914
rect 499408 385900 499436 388690
rect 500512 385914 500540 393286
rect 500868 388816 500920 388822
rect 500868 388758 500920 388764
rect 500158 385886 500540 385914
rect 500880 385900 500908 388758
rect 501984 385914 502012 393286
rect 502340 389020 502392 389026
rect 502340 388962 502392 388968
rect 501630 385886 502012 385914
rect 502352 385900 502380 388962
rect 502996 388890 503024 423370
rect 503640 393314 503668 424322
rect 507952 417784 508004 417790
rect 507952 417726 508004 417732
rect 507860 417716 507912 417722
rect 507860 417658 507912 417664
rect 503996 417648 504048 417654
rect 503996 417590 504048 417596
rect 503720 417580 503772 417586
rect 503720 417522 503772 417528
rect 503456 393286 503668 393314
rect 502984 388884 503036 388890
rect 502984 388826 503036 388832
rect 503456 385914 503484 393286
rect 503102 385886 503484 385914
rect 503732 385914 503760 417522
rect 504008 402974 504036 417590
rect 506480 417512 506532 417518
rect 506480 417454 506532 417460
rect 504008 402946 504128 402974
rect 504100 385914 504128 402946
rect 505560 393984 505612 393990
rect 505560 393926 505612 393932
rect 505284 391264 505336 391270
rect 505284 391206 505336 391212
rect 503732 385886 503838 385914
rect 504100 385886 504574 385914
rect 505296 385900 505324 391206
rect 505572 385914 505600 393926
rect 506492 389298 506520 417454
rect 506572 417444 506624 417450
rect 506572 417386 506624 417392
rect 506480 389292 506532 389298
rect 506480 389234 506532 389240
rect 506584 385914 506612 417386
rect 507124 389292 507176 389298
rect 507124 389234 507176 389240
rect 507136 385914 507164 389234
rect 507872 385914 507900 417658
rect 507964 402974 507992 417726
rect 507964 402946 508544 402974
rect 508516 385914 508544 402946
rect 505572 385886 506046 385914
rect 506584 385886 506782 385914
rect 507136 385886 507518 385914
rect 507872 385886 508254 385914
rect 508516 385886 508990 385914
rect 454408 385688 454460 385694
rect 454408 385630 454460 385636
rect 452016 385416 452068 385422
rect 452016 385358 452068 385364
rect 509330 375592 509386 375601
rect 509330 375527 509386 375536
rect 450728 336796 450780 336802
rect 450728 336738 450780 336744
rect 450464 335326 450584 335354
rect 450556 334257 450584 335326
rect 450542 334248 450598 334257
rect 450542 334183 450598 334192
rect 450450 328672 450506 328681
rect 450450 328607 450506 328616
rect 450464 328506 450492 328607
rect 450452 328500 450504 328506
rect 450452 328442 450504 328448
rect 450556 327321 450584 334183
rect 450740 330546 450768 336738
rect 450728 330540 450780 330546
rect 450728 330482 450780 330488
rect 450542 327312 450598 327321
rect 450542 327247 450598 327256
rect 509344 326262 509372 375527
rect 509514 367024 509570 367033
rect 509514 366959 509570 366968
rect 509422 357640 509478 357649
rect 509422 357575 509478 357584
rect 509332 326256 509384 326262
rect 509332 326198 509384 326204
rect 450372 325666 450492 325694
rect 450464 325553 450492 325666
rect 450450 325544 450506 325553
rect 450450 325479 450506 325488
rect 450358 324864 450414 324873
rect 450188 324822 450358 324850
rect 450358 324799 450414 324808
rect 450082 324592 450138 324601
rect 450082 324527 450138 324536
rect 449808 263560 449860 263566
rect 449808 263502 449860 263508
rect 449440 249076 449492 249082
rect 449440 249018 449492 249024
rect 450372 221474 450400 324799
rect 450464 304638 450492 325479
rect 450634 324184 450690 324193
rect 450634 324119 450690 324128
rect 450542 317112 450598 317121
rect 450542 317047 450598 317056
rect 450452 304632 450504 304638
rect 450452 304574 450504 304580
rect 450360 221468 450412 221474
rect 450360 221410 450412 221416
rect 444912 159854 445248 159882
rect 448224 159854 448468 159882
rect 437992 159332 438624 159338
rect 437940 159326 438624 159332
rect 437952 159310 438624 159326
rect 409696 150408 409748 150414
rect 409696 150350 409748 150356
rect 409604 139392 409656 139398
rect 409604 139334 409656 139340
rect 409512 128308 409564 128314
rect 409512 128250 409564 128256
rect 409420 117292 409472 117298
rect 409420 117234 409472 117240
rect 409328 106276 409380 106282
rect 409328 106218 409380 106224
rect 409236 95192 409288 95198
rect 409236 95134 409288 95140
rect 409144 84176 409196 84182
rect 409144 84118 409196 84124
rect 407856 52420 407908 52426
rect 407856 52362 407908 52368
rect 450556 3738 450584 317047
rect 450648 316946 450676 324119
rect 509330 322960 509386 322969
rect 509330 322895 509386 322904
rect 458272 322720 458324 322726
rect 458824 322720 458876 322726
rect 458272 322662 458324 322668
rect 458284 322386 458312 322662
rect 458560 322658 458666 322674
rect 459100 322720 459152 322726
rect 458824 322662 458876 322668
rect 458942 322668 459100 322674
rect 468208 322720 468260 322726
rect 458942 322662 459152 322668
rect 458548 322652 458666 322658
rect 458600 322646 458666 322652
rect 458548 322594 458600 322600
rect 458836 322522 458864 322662
rect 458942 322646 459140 322662
rect 459218 322658 459416 322674
rect 468208 322662 468260 322668
rect 469036 322720 469088 322726
rect 469036 322662 469088 322668
rect 469588 322720 469640 322726
rect 469588 322662 469640 322668
rect 471244 322720 471296 322726
rect 471244 322662 471296 322668
rect 482650 322688 482706 322697
rect 459218 322652 459428 322658
rect 459218 322646 459376 322652
rect 459376 322594 459428 322600
rect 459388 322522 459494 322538
rect 458824 322516 458876 322522
rect 458824 322458 458876 322464
rect 459376 322516 459494 322522
rect 459428 322510 459494 322516
rect 459376 322458 459428 322464
rect 460492 322386 460598 322402
rect 455788 322380 455840 322386
rect 455788 322322 455840 322328
rect 458272 322380 458324 322386
rect 458272 322322 458324 322328
rect 460480 322380 460598 322386
rect 460532 322374 460598 322380
rect 460480 322322 460532 322328
rect 455800 322046 455828 322322
rect 468220 322250 468248 322662
rect 468484 322652 468536 322658
rect 468484 322594 468536 322600
rect 468496 322386 468524 322594
rect 468760 322584 468812 322590
rect 468760 322526 468812 322532
rect 468772 322425 468800 322526
rect 468758 322416 468814 322425
rect 468484 322380 468536 322386
rect 468758 322351 468814 322360
rect 468484 322322 468536 322328
rect 466552 322244 466604 322250
rect 466552 322186 466604 322192
rect 468208 322244 468260 322250
rect 468208 322186 468260 322192
rect 455788 322040 455840 322046
rect 455788 321982 455840 321988
rect 455788 319184 455840 319190
rect 455788 319126 455840 319132
rect 454776 318232 454828 318238
rect 454776 318174 454828 318180
rect 453396 317416 453448 317422
rect 453396 317358 453448 317364
rect 453304 317212 453356 317218
rect 453304 317154 453356 317160
rect 450910 316976 450966 316985
rect 450636 316940 450688 316946
rect 450910 316911 450966 316920
rect 450636 316882 450688 316888
rect 450636 316804 450688 316810
rect 450636 316746 450688 316752
rect 450648 39846 450676 316746
rect 450820 316736 450872 316742
rect 450726 316704 450782 316713
rect 450820 316678 450872 316684
rect 450726 316639 450782 316648
rect 450636 39840 450688 39846
rect 450636 39782 450688 39788
rect 450544 3732 450596 3738
rect 450544 3674 450596 3680
rect 406566 3567 406622 3576
rect 407764 3596 407816 3602
rect 407764 3538 407816 3544
rect 406382 3496 406438 3505
rect 450740 3466 450768 316639
rect 450832 46306 450860 316678
rect 450820 46300 450872 46306
rect 450820 46242 450872 46248
rect 450924 39370 450952 316911
rect 451924 316872 451976 316878
rect 451094 316840 451150 316849
rect 451924 316814 451976 316820
rect 451094 316775 451150 316784
rect 451004 314084 451056 314090
rect 451004 314026 451056 314032
rect 451016 45490 451044 314026
rect 451004 45484 451056 45490
rect 451004 45426 451056 45432
rect 451108 39642 451136 316775
rect 451936 156913 451964 316814
rect 452016 309800 452068 309806
rect 452016 309742 452068 309748
rect 451922 156904 451978 156913
rect 451922 156839 451978 156848
rect 452028 151473 452056 309742
rect 452292 283620 452344 283626
rect 452292 283562 452344 283568
rect 452108 272536 452160 272542
rect 452108 272478 452160 272484
rect 452014 151464 452070 151473
rect 452014 151399 452070 151408
rect 451556 150272 451608 150278
rect 451556 150214 451608 150220
rect 451568 150113 451596 150214
rect 451554 150104 451610 150113
rect 451554 150039 451610 150048
rect 451740 149048 451792 149054
rect 451740 148990 451792 148996
rect 451752 148753 451780 148990
rect 451738 148744 451794 148753
rect 451738 148679 451794 148688
rect 451740 147416 451792 147422
rect 451738 147384 451740 147393
rect 451792 147384 451794 147393
rect 451738 147319 451794 147328
rect 451556 139392 451608 139398
rect 451556 139334 451608 139340
rect 451568 139233 451596 139334
rect 451554 139224 451610 139233
rect 451554 139159 451610 139168
rect 452120 128353 452148 272478
rect 452200 268456 452252 268462
rect 452200 268398 452252 268404
rect 452212 129713 452240 268398
rect 452304 152833 452332 283562
rect 452384 278044 452436 278050
rect 452384 277986 452436 277992
rect 452396 154193 452424 277986
rect 452568 158296 452620 158302
rect 452566 158264 452568 158273
rect 452620 158264 452622 158273
rect 452566 158199 452622 158208
rect 452568 155712 452620 155718
rect 452568 155654 452620 155660
rect 452580 155553 452608 155654
rect 452566 155544 452622 155553
rect 452566 155479 452622 155488
rect 452382 154184 452438 154193
rect 452382 154119 452438 154128
rect 452290 152824 452346 152833
rect 452290 152759 452346 152768
rect 452568 146192 452620 146198
rect 452568 146134 452620 146140
rect 452580 146033 452608 146134
rect 452566 146024 452622 146033
rect 452566 145959 452622 145968
rect 452568 144696 452620 144702
rect 452566 144664 452568 144673
rect 452620 144664 452622 144673
rect 452566 144599 452622 144608
rect 452568 143336 452620 143342
rect 452566 143304 452568 143313
rect 452620 143304 452622 143313
rect 452566 143239 452622 143248
rect 452568 141976 452620 141982
rect 452566 141944 452568 141953
rect 452620 141944 452622 141953
rect 452566 141879 452622 141888
rect 452568 140684 452620 140690
rect 452568 140626 452620 140632
rect 452580 140593 452608 140626
rect 452566 140584 452622 140593
rect 452566 140519 452622 140528
rect 452568 137896 452620 137902
rect 452566 137864 452568 137873
rect 452620 137864 452622 137873
rect 452566 137799 452622 137808
rect 452568 136536 452620 136542
rect 452566 136504 452568 136513
rect 452620 136504 452622 136513
rect 452566 136439 452622 136448
rect 452568 135176 452620 135182
rect 452566 135144 452568 135153
rect 452620 135144 452622 135153
rect 452566 135079 452622 135088
rect 452568 133816 452620 133822
rect 452566 133784 452568 133793
rect 452620 133784 452622 133793
rect 452566 133719 452622 133728
rect 452476 132456 452528 132462
rect 452474 132424 452476 132433
rect 452528 132424 452530 132433
rect 452474 132359 452530 132368
rect 452568 131096 452620 131102
rect 452566 131064 452568 131073
rect 452620 131064 452622 131073
rect 452566 130999 452622 131008
rect 452198 129704 452254 129713
rect 452198 129639 452254 129648
rect 452106 128344 452162 128353
rect 452106 128279 452162 128288
rect 452566 126984 452622 126993
rect 452566 126919 452568 126928
rect 452620 126919 452622 126928
rect 452568 126890 452620 126896
rect 451924 126064 451976 126070
rect 451924 126006 451976 126012
rect 451936 125633 451964 126006
rect 451922 125624 451978 125633
rect 451922 125559 451978 125568
rect 451924 124772 451976 124778
rect 451924 124714 451976 124720
rect 451936 124273 451964 124714
rect 451922 124264 451978 124273
rect 451922 124199 451978 124208
rect 451924 123276 451976 123282
rect 451924 123218 451976 123224
rect 451936 122913 451964 123218
rect 451922 122904 451978 122913
rect 451922 122839 451978 122848
rect 451740 122256 451792 122262
rect 451740 122198 451792 122204
rect 451752 121553 451780 122198
rect 451738 121544 451794 121553
rect 451738 121479 451794 121488
rect 453316 45558 453344 317154
rect 453408 46442 453436 317358
rect 454682 317248 454738 317257
rect 454682 317183 454738 317192
rect 453488 317008 453540 317014
rect 453488 316950 453540 316956
rect 453500 46510 453528 316950
rect 453580 316668 453632 316674
rect 453580 316610 453632 316616
rect 453488 46504 453540 46510
rect 453488 46446 453540 46452
rect 453396 46436 453448 46442
rect 453396 46378 453448 46384
rect 453592 46374 453620 316610
rect 453672 308508 453724 308514
rect 453672 308450 453724 308456
rect 453684 126070 453712 308450
rect 453764 307148 453816 307154
rect 453764 307090 453816 307096
rect 453776 132462 453804 307090
rect 453948 279472 454000 279478
rect 453948 279414 454000 279420
rect 453856 274032 453908 274038
rect 453856 273974 453908 273980
rect 453764 132456 453816 132462
rect 453764 132398 453816 132404
rect 453672 126064 453724 126070
rect 453672 126006 453724 126012
rect 453868 124778 453896 273974
rect 453960 131102 453988 279414
rect 453948 131096 454000 131102
rect 453948 131038 454000 131044
rect 453856 124772 453908 124778
rect 453856 124714 453908 124720
rect 453580 46368 453632 46374
rect 453580 46310 453632 46316
rect 453304 45552 453356 45558
rect 453304 45494 453356 45500
rect 454696 42158 454724 317183
rect 454788 135182 454816 318174
rect 455800 313954 455828 319126
rect 455788 313948 455840 313954
rect 455788 313890 455840 313896
rect 454868 311228 454920 311234
rect 454868 311170 454920 311176
rect 454880 149054 454908 311170
rect 455892 304502 455920 322116
rect 456076 322102 456182 322130
rect 456458 322102 456656 322130
rect 456076 319190 456104 322102
rect 456154 319424 456210 319433
rect 456154 319359 456210 319368
rect 456064 319184 456116 319190
rect 456064 319126 456116 319132
rect 456064 318164 456116 318170
rect 456064 318106 456116 318112
rect 455972 304632 456024 304638
rect 455972 304574 456024 304580
rect 455880 304496 455932 304502
rect 455880 304438 455932 304444
rect 455052 280832 455104 280838
rect 455052 280774 455104 280780
rect 454960 273964 455012 273970
rect 454960 273906 455012 273912
rect 454868 149048 454920 149054
rect 454868 148990 454920 148996
rect 454972 137902 455000 273906
rect 455064 144702 455092 280774
rect 455236 276684 455288 276690
rect 455236 276626 455288 276632
rect 455144 272604 455196 272610
rect 455144 272546 455196 272552
rect 455052 144696 455104 144702
rect 455052 144638 455104 144644
rect 455156 141982 455184 272546
rect 455248 150278 455276 276626
rect 455984 235006 456012 304574
rect 455972 235000 456024 235006
rect 455972 234942 456024 234948
rect 455236 150272 455288 150278
rect 455236 150214 455288 150220
rect 455144 141976 455196 141982
rect 455144 141918 455196 141924
rect 454960 137896 455012 137902
rect 454960 137838 455012 137844
rect 454776 135176 454828 135182
rect 454776 135118 454828 135124
rect 454684 42152 454736 42158
rect 454684 42094 454736 42100
rect 451096 39636 451148 39642
rect 451096 39578 451148 39584
rect 450912 39364 450964 39370
rect 450912 39306 450964 39312
rect 456076 3534 456104 318106
rect 456168 47054 456196 319359
rect 456340 317348 456392 317354
rect 456340 317290 456392 317296
rect 456248 316600 456300 316606
rect 456248 316542 456300 316548
rect 456156 47048 456208 47054
rect 456156 46990 456208 46996
rect 456260 46646 456288 316542
rect 456352 46714 456380 317290
rect 456432 317280 456484 317286
rect 456432 317222 456484 317228
rect 456340 46708 456392 46714
rect 456340 46650 456392 46656
rect 456248 46640 456300 46646
rect 456248 46582 456300 46588
rect 456444 46578 456472 317222
rect 456524 309936 456576 309942
rect 456524 309878 456576 309884
rect 456536 155718 456564 309878
rect 456628 303278 456656 322102
rect 456616 303272 456668 303278
rect 456616 303214 456668 303220
rect 456720 301578 456748 322116
rect 457010 322102 457208 322130
rect 457180 319190 457208 322102
rect 457168 319184 457220 319190
rect 457168 319126 457220 319132
rect 457272 316034 457300 322116
rect 457548 316034 457576 322116
rect 457720 316940 457772 316946
rect 457720 316882 457772 316888
rect 457272 316006 457392 316034
rect 457548 316006 457668 316034
rect 457364 307086 457392 316006
rect 457444 315444 457496 315450
rect 457444 315386 457496 315392
rect 457352 307080 457404 307086
rect 457352 307022 457404 307028
rect 456708 301572 456760 301578
rect 456708 301514 456760 301520
rect 456616 271244 456668 271250
rect 456616 271186 456668 271192
rect 456524 155712 456576 155718
rect 456524 155654 456576 155660
rect 456628 133822 456656 271186
rect 456708 269952 456760 269958
rect 456708 269894 456760 269900
rect 456720 158302 456748 269894
rect 456800 263560 456852 263566
rect 456800 263502 456852 263508
rect 456812 262721 456840 263502
rect 456798 262712 456854 262721
rect 456798 262647 456854 262656
rect 456708 158296 456760 158302
rect 456708 158238 456760 158244
rect 456616 133816 456668 133822
rect 456616 133758 456668 133764
rect 457456 126954 457484 315386
rect 457536 306264 457588 306270
rect 457536 306206 457588 306212
rect 457548 139398 457576 306206
rect 457640 297226 457668 316006
rect 457628 297220 457680 297226
rect 457628 297162 457680 297168
rect 457628 271176 457680 271182
rect 457628 271118 457680 271124
rect 457640 143342 457668 271118
rect 457732 207233 457760 316882
rect 457824 316062 457852 322116
rect 458100 320142 458128 322116
rect 458376 321502 458404 322116
rect 459770 322102 459968 322130
rect 458364 321496 458416 321502
rect 458364 321438 458416 321444
rect 459940 320958 459968 322102
rect 459928 320952 459980 320958
rect 459928 320894 459980 320900
rect 460032 320657 460060 322116
rect 460204 321088 460256 321094
rect 460204 321030 460256 321036
rect 460018 320648 460074 320657
rect 460018 320583 460074 320592
rect 458088 320136 458140 320142
rect 458088 320078 458140 320084
rect 459008 319592 459060 319598
rect 459008 319534 459060 319540
rect 458824 319456 458876 319462
rect 458824 319398 458876 319404
rect 457996 319184 458048 319190
rect 457996 319126 458048 319132
rect 457812 316056 457864 316062
rect 457812 315998 457864 316004
rect 458008 300694 458036 319126
rect 457996 300688 458048 300694
rect 457996 300630 458048 300636
rect 458640 275324 458692 275330
rect 458640 275266 458692 275272
rect 457812 249076 457864 249082
rect 457812 249018 457864 249024
rect 457824 248849 457852 249018
rect 457810 248840 457866 248849
rect 457810 248775 457866 248784
rect 457718 207224 457774 207233
rect 457718 207159 457774 207168
rect 457824 162178 457852 248775
rect 457996 235000 458048 235006
rect 457994 234968 457996 234977
rect 458048 234968 458050 234977
rect 457994 234903 458050 234912
rect 458008 229094 458036 234903
rect 457916 229066 458036 229094
rect 457916 162382 457944 229066
rect 457996 221468 458048 221474
rect 457996 221410 458048 221416
rect 458008 221105 458036 221410
rect 457994 221096 458050 221105
rect 457994 221031 458050 221040
rect 457904 162376 457956 162382
rect 457904 162318 457956 162324
rect 458008 162314 458036 221031
rect 458086 207224 458142 207233
rect 458086 207159 458142 207168
rect 457996 162308 458048 162314
rect 457996 162250 458048 162256
rect 458100 162246 458128 207159
rect 458088 162240 458140 162246
rect 458088 162182 458140 162188
rect 457812 162172 457864 162178
rect 457812 162114 457864 162120
rect 458652 147422 458680 275266
rect 458732 271312 458784 271318
rect 458732 271254 458784 271260
rect 458640 147416 458692 147422
rect 458640 147358 458692 147364
rect 457628 143336 457680 143342
rect 457628 143278 457680 143284
rect 457536 139392 457588 139398
rect 457536 139334 457588 139340
rect 457444 126948 457496 126954
rect 457444 126890 457496 126896
rect 458744 122262 458772 271254
rect 458732 122256 458784 122262
rect 458732 122198 458784 122204
rect 458836 46617 458864 319398
rect 458916 317076 458968 317082
rect 458916 317018 458968 317024
rect 458928 46782 458956 317018
rect 459020 46889 459048 319534
rect 459192 317144 459244 317150
rect 459192 317086 459244 317092
rect 459100 316940 459152 316946
rect 459100 316882 459152 316888
rect 459112 136542 459140 316882
rect 459100 136536 459152 136542
rect 459100 136478 459152 136484
rect 459006 46880 459062 46889
rect 459006 46815 459062 46824
rect 458916 46776 458968 46782
rect 459204 46753 459232 317086
rect 459284 315376 459336 315382
rect 459284 315318 459336 315324
rect 459296 140690 459324 315318
rect 459376 314016 459428 314022
rect 459376 313958 459428 313964
rect 459388 146198 459416 313958
rect 459468 282192 459520 282198
rect 459468 282134 459520 282140
rect 459376 146192 459428 146198
rect 459376 146134 459428 146140
rect 459284 140684 459336 140690
rect 459284 140626 459336 140632
rect 459480 123282 459508 282134
rect 459468 123276 459520 123282
rect 459468 123218 459520 123224
rect 458916 46718 458968 46724
rect 459190 46744 459246 46753
rect 459190 46679 459246 46688
rect 458822 46608 458878 46617
rect 456432 46572 456484 46578
rect 458822 46543 458878 46552
rect 456432 46514 456484 46520
rect 460216 42226 460244 321030
rect 460308 320113 460336 322116
rect 460294 320104 460350 320113
rect 460860 320074 460888 322116
rect 461136 321337 461164 322116
rect 461412 321434 461440 322116
rect 461400 321428 461452 321434
rect 461400 321370 461452 321376
rect 461688 321366 461716 322116
rect 461676 321360 461728 321366
rect 461122 321328 461178 321337
rect 461676 321302 461728 321308
rect 461122 321263 461178 321272
rect 461964 321065 461992 322116
rect 462240 321473 462268 322116
rect 462226 321464 462282 321473
rect 462226 321399 462282 321408
rect 462516 321201 462544 322116
rect 462502 321192 462558 321201
rect 462502 321127 462558 321136
rect 461950 321056 462006 321065
rect 461950 320991 462006 321000
rect 461860 320884 461912 320890
rect 461860 320826 461912 320832
rect 461872 320142 461900 320826
rect 461860 320136 461912 320142
rect 461860 320078 461912 320084
rect 460294 320039 460350 320048
rect 460848 320068 460900 320074
rect 460848 320010 460900 320016
rect 462792 319734 462820 322116
rect 463068 321570 463096 322116
rect 463056 321564 463108 321570
rect 463056 321506 463108 321512
rect 463344 320006 463372 322116
rect 463528 322102 463634 322130
rect 463528 322046 463556 322102
rect 463516 322040 463568 322046
rect 463516 321982 463568 321988
rect 463332 320000 463384 320006
rect 463332 319942 463384 319948
rect 463896 319870 463924 322116
rect 464080 322102 464186 322130
rect 464356 322102 464462 322130
rect 463884 319864 463936 319870
rect 463884 319806 463936 319812
rect 462780 319728 462832 319734
rect 462780 319670 462832 319676
rect 460388 319660 460440 319666
rect 460388 319602 460440 319608
rect 460296 319524 460348 319530
rect 460296 319466 460348 319472
rect 460308 46918 460336 319466
rect 460296 46912 460348 46918
rect 460296 46854 460348 46860
rect 460400 46850 460428 319602
rect 464080 319138 464108 322102
rect 463804 319110 464108 319138
rect 461584 316056 461636 316062
rect 461584 315998 461636 316004
rect 461596 299470 461624 315998
rect 463804 313342 463832 319110
rect 464356 316034 464384 322102
rect 464724 316674 464752 322116
rect 465000 317422 465028 322116
rect 464988 317416 465040 317422
rect 464988 317358 465040 317364
rect 464712 316668 464764 316674
rect 464712 316610 464764 316616
rect 465276 316606 465304 322116
rect 465552 319598 465580 322116
rect 465828 319666 465856 322116
rect 466012 322102 466118 322130
rect 465816 319660 465868 319666
rect 465816 319602 465868 319608
rect 465540 319592 465592 319598
rect 465540 319534 465592 319540
rect 465264 316600 465316 316606
rect 465264 316542 465316 316548
rect 466012 316034 466040 322102
rect 464080 316006 464384 316034
rect 465460 316006 466040 316034
rect 461676 313336 461728 313342
rect 461676 313278 461728 313284
rect 463792 313336 463844 313342
rect 463792 313278 463844 313284
rect 461688 304570 461716 313278
rect 461676 304564 461728 304570
rect 461676 304506 461728 304512
rect 461584 299464 461636 299470
rect 461584 299406 461636 299412
rect 464080 289610 464108 316006
rect 465460 306202 465488 316006
rect 465448 306196 465500 306202
rect 465448 306138 465500 306144
rect 464068 289604 464120 289610
rect 464068 289546 464120 289552
rect 462964 281920 463016 281926
rect 462964 281862 463016 281868
rect 462976 279546 463004 281862
rect 462964 279540 463016 279546
rect 462964 279482 463016 279488
rect 466380 268394 466408 322116
rect 466564 320074 466592 322186
rect 466552 320068 466604 320074
rect 466552 320010 466604 320016
rect 466656 318986 466684 322116
rect 466828 319184 466880 319190
rect 466828 319126 466880 319132
rect 466644 318980 466696 318986
rect 466644 318922 466696 318928
rect 466840 284986 466868 319126
rect 466932 316034 466960 322116
rect 467208 316034 467236 322116
rect 467392 322102 467498 322130
rect 467668 322102 467774 322130
rect 468050 322102 468248 322130
rect 468326 322102 468524 322130
rect 467392 319190 467420 322102
rect 467380 319184 467432 319190
rect 467380 319126 467432 319132
rect 467380 318980 467432 318986
rect 467380 318922 467432 318928
rect 466932 316006 467052 316034
rect 467208 316006 467328 316034
rect 467024 290494 467052 316006
rect 467300 293282 467328 316006
rect 467392 311166 467420 318922
rect 467380 311160 467432 311166
rect 467380 311102 467432 311108
rect 467288 293276 467340 293282
rect 467288 293218 467340 293224
rect 467012 290488 467064 290494
rect 467012 290430 467064 290436
rect 467668 286346 467696 322102
rect 468220 316034 468248 322102
rect 468496 319138 468524 322102
rect 468588 321570 468616 322116
rect 468576 321564 468628 321570
rect 468576 321506 468628 321512
rect 468864 319258 468892 322116
rect 469048 322046 469076 322662
rect 469154 322114 469352 322130
rect 469154 322108 469364 322114
rect 469154 322102 469312 322108
rect 469312 322050 469364 322056
rect 469036 322040 469088 322046
rect 469036 321982 469088 321988
rect 469416 321434 469444 322116
rect 469600 322114 469628 322662
rect 470968 322584 471020 322590
rect 470968 322526 471020 322532
rect 470140 322516 470192 322522
rect 470140 322458 470192 322464
rect 470152 322425 470180 322458
rect 470138 322416 470194 322425
rect 470138 322351 470194 322360
rect 469588 322108 469640 322114
rect 469588 322050 469640 322056
rect 469404 321428 469456 321434
rect 469404 321370 469456 321376
rect 469692 319870 469720 322116
rect 469680 319864 469732 319870
rect 469680 319806 469732 319812
rect 468852 319252 468904 319258
rect 468852 319194 468904 319200
rect 469968 319190 469996 322116
rect 470244 320006 470272 322116
rect 470520 321337 470548 322116
rect 470506 321328 470562 321337
rect 470506 321263 470562 321272
rect 470232 320000 470284 320006
rect 470232 319942 470284 319948
rect 469956 319184 470008 319190
rect 468496 319110 469076 319138
rect 469956 319126 470008 319132
rect 468220 316006 468800 316034
rect 467656 286340 467708 286346
rect 467656 286282 467708 286288
rect 466828 284980 466880 284986
rect 466828 284922 466880 284928
rect 468772 269890 468800 316006
rect 469048 313274 469076 319110
rect 470796 318714 470824 322116
rect 470980 322046 471008 322526
rect 471256 322250 471284 322662
rect 471520 322652 471572 322658
rect 482650 322623 482706 322632
rect 483754 322688 483810 322697
rect 483754 322623 483810 322632
rect 507122 322688 507178 322697
rect 507122 322623 507178 322632
rect 471520 322594 471572 322600
rect 471532 322386 471560 322594
rect 484216 322584 484268 322590
rect 473542 322552 473598 322561
rect 479642 322522 479840 322538
rect 484268 322532 484334 322538
rect 484216 322526 484334 322532
rect 479642 322516 479852 322522
rect 479642 322510 479800 322516
rect 473542 322487 473598 322496
rect 484228 322510 484334 322526
rect 479800 322458 479852 322464
rect 483940 322448 483992 322454
rect 483992 322396 484058 322402
rect 483940 322390 484058 322396
rect 471520 322380 471572 322386
rect 483952 322374 484058 322390
rect 471520 322322 471572 322328
rect 472072 322312 472124 322318
rect 472124 322260 472190 322266
rect 472072 322254 472190 322260
rect 471244 322244 471296 322250
rect 472084 322238 472190 322254
rect 500224 322244 500276 322250
rect 471244 322186 471296 322192
rect 500224 322186 500276 322192
rect 481456 322176 481508 322182
rect 470968 322040 471020 322046
rect 470968 321982 471020 321988
rect 471072 319802 471100 322116
rect 471060 319796 471112 319802
rect 471060 319738 471112 319744
rect 471348 319394 471376 322116
rect 471336 319388 471388 319394
rect 471336 319330 471388 319336
rect 471244 319048 471296 319054
rect 471244 318990 471296 318996
rect 470784 318708 470836 318714
rect 470784 318650 470836 318656
rect 469036 313268 469088 313274
rect 469036 313210 469088 313216
rect 471256 312594 471284 318990
rect 471624 318986 471652 322116
rect 471900 321162 471928 322116
rect 471888 321156 471940 321162
rect 471888 321098 471940 321104
rect 472452 320754 472480 322116
rect 472440 320748 472492 320754
rect 472440 320690 472492 320696
rect 472728 319977 472756 322116
rect 472714 319968 472770 319977
rect 472714 319903 472770 319912
rect 473004 319705 473032 322116
rect 473280 320822 473308 322116
rect 473832 321230 473860 322116
rect 473820 321224 473872 321230
rect 473820 321166 473872 321172
rect 473268 320816 473320 320822
rect 473268 320758 473320 320764
rect 474108 319841 474136 322116
rect 474384 320074 474412 322116
rect 474372 320068 474424 320074
rect 474372 320010 474424 320016
rect 474094 319832 474150 319841
rect 474094 319767 474150 319776
rect 472990 319696 473046 319705
rect 472990 319631 473046 319640
rect 474660 319054 474688 322116
rect 474648 319048 474700 319054
rect 474648 318990 474700 318996
rect 471612 318980 471664 318986
rect 471612 318922 471664 318928
rect 474936 316742 474964 322116
rect 475212 317218 475240 322116
rect 475488 317286 475516 322116
rect 475764 317354 475792 322116
rect 476040 319462 476068 322116
rect 476316 319530 476344 322116
rect 476500 322102 476606 322130
rect 476304 319524 476356 319530
rect 476304 319466 476356 319472
rect 476028 319456 476080 319462
rect 476028 319398 476080 319404
rect 475752 317348 475804 317354
rect 475752 317290 475804 317296
rect 475476 317280 475528 317286
rect 475476 317222 475528 317228
rect 475200 317212 475252 317218
rect 475200 317154 475252 317160
rect 474924 316736 474976 316742
rect 474924 316678 474976 316684
rect 471244 312588 471296 312594
rect 471244 312530 471296 312536
rect 469864 311296 469916 311302
rect 469864 311238 469916 311244
rect 469876 306338 469904 311238
rect 469864 306332 469916 306338
rect 469864 306274 469916 306280
rect 476500 286414 476528 322102
rect 476868 318102 476896 322116
rect 477158 322102 477356 322130
rect 476856 318096 476908 318102
rect 476856 318038 476908 318044
rect 476764 308372 476816 308378
rect 476764 308314 476816 308320
rect 476488 286408 476540 286414
rect 476488 286350 476540 286356
rect 476776 285054 476804 308314
rect 477328 306202 477356 322102
rect 477316 306196 477368 306202
rect 477316 306138 477368 306144
rect 477420 296002 477448 322116
rect 477710 322102 477908 322130
rect 477880 316034 477908 322102
rect 477972 316742 478000 322116
rect 478262 322102 478460 322130
rect 481508 322124 481574 322130
rect 481456 322118 481574 322124
rect 477960 316736 478012 316742
rect 477960 316678 478012 316684
rect 477880 316006 478184 316034
rect 478156 315314 478184 316006
rect 478144 315308 478196 315314
rect 478144 315250 478196 315256
rect 477408 295996 477460 296002
rect 477408 295938 477460 295944
rect 478432 291650 478460 322102
rect 478524 317762 478552 322116
rect 478800 319462 478828 322116
rect 479076 321366 479104 322116
rect 479064 321360 479116 321366
rect 479064 321302 479116 321308
rect 479352 320074 479380 322116
rect 479340 320068 479392 320074
rect 479340 320010 479392 320016
rect 479904 319938 479932 322116
rect 479892 319932 479944 319938
rect 479892 319874 479944 319880
rect 480180 319666 480208 322116
rect 480456 319734 480484 322116
rect 480732 320142 480760 322116
rect 480720 320136 480772 320142
rect 480720 320078 480772 320084
rect 481008 319802 481036 322116
rect 480996 319796 481048 319802
rect 480996 319738 481048 319744
rect 480444 319728 480496 319734
rect 480444 319670 480496 319676
rect 480168 319660 480220 319666
rect 480168 319602 480220 319608
rect 478788 319456 478840 319462
rect 478788 319398 478840 319404
rect 481284 319394 481312 322116
rect 481468 322102 481574 322118
rect 481836 320686 481864 322116
rect 482112 321026 482140 322116
rect 482100 321020 482152 321026
rect 482100 320962 482152 320968
rect 481824 320680 481876 320686
rect 481824 320622 481876 320628
rect 481272 319388 481324 319394
rect 481272 319330 481324 319336
rect 482388 319326 482416 322116
rect 482940 319569 482968 322116
rect 483216 321298 483244 322116
rect 483204 321292 483256 321298
rect 483204 321234 483256 321240
rect 482926 319560 482982 319569
rect 482926 319495 482982 319504
rect 482376 319320 482428 319326
rect 482376 319262 482428 319268
rect 483492 318782 483520 322116
rect 484504 322102 484610 322130
rect 484780 322102 484886 322130
rect 485056 322102 485162 322130
rect 485332 322102 485438 322130
rect 484504 320090 484532 322102
rect 484412 320062 484532 320090
rect 484412 319410 484440 320062
rect 484320 319382 484440 319410
rect 484320 319122 484348 319382
rect 484780 319274 484808 322102
rect 484412 319246 484808 319274
rect 484308 319116 484360 319122
rect 484308 319058 484360 319064
rect 483480 318776 483532 318782
rect 483480 318718 483532 318724
rect 478512 317756 478564 317762
rect 478512 317698 478564 317704
rect 479524 317756 479576 317762
rect 479524 317698 479576 317704
rect 478880 312588 478932 312594
rect 478880 312530 478932 312536
rect 478892 308378 478920 312530
rect 478880 308372 478932 308378
rect 478880 308314 478932 308320
rect 478420 291644 478472 291650
rect 478420 291586 478472 291592
rect 469220 285048 469272 285054
rect 469220 284990 469272 284996
rect 476764 285048 476816 285054
rect 476764 284990 476816 284996
rect 469232 281926 469260 284990
rect 469220 281920 469272 281926
rect 469220 281862 469272 281868
rect 479536 273222 479564 317698
rect 484412 316674 484440 319246
rect 485056 319138 485084 322102
rect 484504 319110 485084 319138
rect 481732 316668 481784 316674
rect 481732 316610 481784 316616
rect 484400 316668 484452 316674
rect 484400 316610 484452 316616
rect 481744 312594 481772 316610
rect 484504 313614 484532 319110
rect 485332 316034 485360 322102
rect 485700 317014 485728 322116
rect 485976 317082 486004 322116
rect 486252 319433 486280 322116
rect 486238 319424 486294 319433
rect 486238 319359 486294 319368
rect 486528 317150 486556 322116
rect 486712 322102 486818 322130
rect 486988 322102 487094 322130
rect 487370 322102 487568 322130
rect 486516 317144 486568 317150
rect 486516 317086 486568 317092
rect 485964 317076 486016 317082
rect 485964 317018 486016 317024
rect 485688 317008 485740 317014
rect 485688 316950 485740 316956
rect 485872 316668 485924 316674
rect 485872 316610 485924 316616
rect 484780 316006 485360 316034
rect 484780 314090 484808 316006
rect 484768 314084 484820 314090
rect 484768 314026 484820 314032
rect 482100 313608 482152 313614
rect 482100 313550 482152 313556
rect 484492 313608 484544 313614
rect 484492 313550 484544 313556
rect 481732 312588 481784 312594
rect 481732 312530 481784 312536
rect 482112 311302 482140 313550
rect 482100 311296 482152 311302
rect 482100 311238 482152 311244
rect 485884 302734 485912 316610
rect 486712 311894 486740 322102
rect 486988 316674 487016 322102
rect 487252 316940 487304 316946
rect 487252 316882 487304 316888
rect 486976 316668 487028 316674
rect 486976 316610 487028 316616
rect 486436 311866 486740 311894
rect 485872 302728 485924 302734
rect 485872 302670 485924 302676
rect 486436 294574 486464 311866
rect 486424 294568 486476 294574
rect 486424 294510 486476 294516
rect 479524 273216 479576 273222
rect 479524 273158 479576 273164
rect 487264 269958 487292 316882
rect 487540 316674 487568 322102
rect 487632 321554 487660 322116
rect 487632 321526 487752 321554
rect 487528 316668 487580 316674
rect 487528 316610 487580 316616
rect 487724 309874 487752 321526
rect 487908 316674 487936 322116
rect 488092 322102 488198 322130
rect 488368 322102 488474 322130
rect 488750 322102 488948 322130
rect 487804 316668 487856 316674
rect 487804 316610 487856 316616
rect 487896 316668 487948 316674
rect 487896 316610 487948 316616
rect 487712 309868 487764 309874
rect 487712 309810 487764 309816
rect 487816 308446 487844 316610
rect 487804 308440 487856 308446
rect 487804 308382 487856 308388
rect 488092 275398 488120 322102
rect 488368 316946 488396 322102
rect 488356 316940 488408 316946
rect 488356 316882 488408 316888
rect 488356 316668 488408 316674
rect 488356 316610 488408 316616
rect 488632 316668 488684 316674
rect 488632 316610 488684 316616
rect 488368 287706 488396 316610
rect 488356 287700 488408 287706
rect 488356 287642 488408 287648
rect 488080 275392 488132 275398
rect 488080 275334 488132 275340
rect 488644 274038 488672 316610
rect 488632 274032 488684 274038
rect 488632 273974 488684 273980
rect 488920 271318 488948 322102
rect 489012 282198 489040 322116
rect 489196 322102 489302 322130
rect 489472 322102 489578 322130
rect 489748 322102 489854 322130
rect 489196 316674 489224 322102
rect 489184 316668 489236 316674
rect 489184 316610 489236 316616
rect 489472 311894 489500 322102
rect 489748 315450 489776 322102
rect 490012 316600 490064 316606
rect 490012 316542 490064 316548
rect 489736 315444 489788 315450
rect 489736 315386 489788 315392
rect 489196 311866 489500 311894
rect 489196 308514 489224 311866
rect 489184 308508 489236 308514
rect 489184 308450 489236 308456
rect 489000 282192 489052 282198
rect 489000 282134 489052 282140
rect 488908 271312 488960 271318
rect 488908 271254 488960 271260
rect 490024 271250 490052 316542
rect 490116 272542 490144 322116
rect 490288 316668 490340 316674
rect 490288 316610 490340 316616
rect 490300 307154 490328 316610
rect 490288 307148 490340 307154
rect 490288 307090 490340 307096
rect 490104 272536 490156 272542
rect 490104 272478 490156 272484
rect 490012 271244 490064 271250
rect 490012 271186 490064 271192
rect 487252 269952 487304 269958
rect 487252 269894 487304 269900
rect 468760 269884 468812 269890
rect 468760 269826 468812 269832
rect 490392 268462 490420 322116
rect 490576 322102 490682 322130
rect 490852 322102 490958 322130
rect 491128 322102 491234 322130
rect 490576 279478 490604 322102
rect 490852 316674 490880 322102
rect 490840 316668 490892 316674
rect 490840 316610 490892 316616
rect 491128 316606 491156 322102
rect 491496 318238 491524 322116
rect 491680 322102 491786 322130
rect 491956 322102 492062 322130
rect 492232 322102 492338 322130
rect 492508 322102 492614 322130
rect 492784 322102 492890 322130
rect 491484 318232 491536 318238
rect 491484 318174 491536 318180
rect 491680 317014 491708 322102
rect 491668 317008 491720 317014
rect 491668 316950 491720 316956
rect 491116 316600 491168 316606
rect 491116 316542 491168 316548
rect 491392 316532 491444 316538
rect 491392 316474 491444 316480
rect 491404 306270 491432 316474
rect 491956 311894 491984 322102
rect 492232 316538 492260 322102
rect 492220 316532 492272 316538
rect 492220 316474 492272 316480
rect 492508 315382 492536 322102
rect 492496 315376 492548 315382
rect 492496 315318 492548 315324
rect 491680 311866 491984 311894
rect 491392 306264 491444 306270
rect 491392 306206 491444 306212
rect 490564 279472 490616 279478
rect 490564 279414 490616 279420
rect 491680 273970 491708 311866
rect 491668 273964 491720 273970
rect 491668 273906 491720 273912
rect 492784 272610 492812 322102
rect 492772 272604 492824 272610
rect 492772 272546 492824 272552
rect 493152 271182 493180 322116
rect 493324 316668 493376 316674
rect 493324 316610 493376 316616
rect 493336 275330 493364 316610
rect 493428 280838 493456 322116
rect 493612 322102 493718 322130
rect 493888 322102 493994 322130
rect 494270 322102 494468 322130
rect 493612 314022 493640 322102
rect 493888 316674 493916 322102
rect 493876 316668 493928 316674
rect 493876 316610 493928 316616
rect 494152 316668 494204 316674
rect 494152 316610 494204 316616
rect 493600 314016 493652 314022
rect 493600 313958 493652 313964
rect 493416 280832 493468 280838
rect 493416 280774 493468 280780
rect 494164 278050 494192 316610
rect 494440 311234 494468 322102
rect 494428 311228 494480 311234
rect 494428 311170 494480 311176
rect 494152 278044 494204 278050
rect 494152 277986 494204 277992
rect 494532 276690 494560 322116
rect 494716 322102 494822 322130
rect 494992 322102 495098 322130
rect 495268 322102 495374 322130
rect 494716 321554 494744 322102
rect 494992 321554 495020 322102
rect 494624 321526 494744 321554
rect 494808 321526 495020 321554
rect 494624 311914 494652 321526
rect 494808 316826 494836 321526
rect 494716 316798 494836 316826
rect 494612 311908 494664 311914
rect 494612 311850 494664 311856
rect 494716 283626 494744 316798
rect 495268 316674 495296 322102
rect 495256 316668 495308 316674
rect 495256 316610 495308 316616
rect 494796 311908 494848 311914
rect 494796 311850 494848 311856
rect 494808 309806 494836 311850
rect 495636 309942 495664 322116
rect 495912 316878 495940 322116
rect 496188 318238 496216 322116
rect 496478 322102 496676 322130
rect 496176 318232 496228 318238
rect 496176 318174 496228 318180
rect 495900 316872 495952 316878
rect 495900 316814 495952 316820
rect 496648 315382 496676 322102
rect 496636 315376 496688 315382
rect 496636 315318 496688 315324
rect 496740 314022 496768 322116
rect 497030 322102 497228 322130
rect 497306 322102 497504 322130
rect 496820 321020 496872 321026
rect 496820 320962 496872 320968
rect 496832 320074 496860 320962
rect 496820 320068 496872 320074
rect 496820 320010 496872 320016
rect 496728 314016 496780 314022
rect 496728 313958 496780 313964
rect 497200 311137 497228 322102
rect 497476 319122 497504 322102
rect 497464 319116 497516 319122
rect 497464 319058 497516 319064
rect 497568 316034 497596 322116
rect 497752 322102 497858 322130
rect 497568 316006 497688 316034
rect 497186 311128 497242 311137
rect 497186 311063 497242 311072
rect 495624 309936 495676 309942
rect 495624 309878 495676 309884
rect 494796 309800 494848 309806
rect 494796 309742 494848 309748
rect 494704 283620 494756 283626
rect 494704 283562 494756 283568
rect 497660 280838 497688 316006
rect 497648 280832 497700 280838
rect 497648 280774 497700 280780
rect 494520 276684 494572 276690
rect 494520 276626 494572 276632
rect 493324 275324 493376 275330
rect 493324 275266 493376 275272
rect 493140 271176 493192 271182
rect 493140 271118 493192 271124
rect 497752 268462 497780 322102
rect 498120 319530 498148 322116
rect 498410 322102 498608 322130
rect 498108 319524 498160 319530
rect 498108 319466 498160 319472
rect 498016 319116 498068 319122
rect 498016 319058 498068 319064
rect 498028 279478 498056 319058
rect 498580 316034 498608 322102
rect 498672 319598 498700 322116
rect 498660 319592 498712 319598
rect 498660 319534 498712 319540
rect 498948 316034 498976 322116
rect 499132 322102 499238 322130
rect 499408 322102 499514 322130
rect 499790 322102 499988 322130
rect 498580 316006 498884 316034
rect 498948 316006 499068 316034
rect 498856 285054 498884 316006
rect 498844 285048 498896 285054
rect 498844 284990 498896 284996
rect 498016 279472 498068 279478
rect 498016 279414 498068 279420
rect 499040 275330 499068 316006
rect 499028 275324 499080 275330
rect 499028 275266 499080 275272
rect 499132 271182 499160 322102
rect 499408 273970 499436 322102
rect 499960 276690 499988 322102
rect 500052 316034 500080 322116
rect 500236 319462 500264 322186
rect 500224 319456 500276 319462
rect 500224 319398 500276 319404
rect 500328 316946 500356 322116
rect 500512 322102 500618 322130
rect 500788 322102 500894 322130
rect 501170 322102 501368 322130
rect 501446 322102 501644 322130
rect 500316 316940 500368 316946
rect 500316 316882 500368 316888
rect 500052 316006 500172 316034
rect 500144 286414 500172 316006
rect 500132 286408 500184 286414
rect 500132 286350 500184 286356
rect 499948 276684 500000 276690
rect 499948 276626 500000 276632
rect 499396 273964 499448 273970
rect 499396 273906 499448 273912
rect 500512 271250 500540 322102
rect 500788 272542 500816 322102
rect 501340 316034 501368 322102
rect 501616 319122 501644 322102
rect 501708 319462 501736 322116
rect 501696 319456 501748 319462
rect 501696 319398 501748 319404
rect 501604 319116 501656 319122
rect 501604 319058 501656 319064
rect 501984 316034 502012 322116
rect 502156 319116 502208 319122
rect 502156 319058 502208 319064
rect 501340 316006 501644 316034
rect 501984 316006 502104 316034
rect 501616 315450 501644 316006
rect 501604 315444 501656 315450
rect 501604 315386 501656 315392
rect 502076 312594 502104 316006
rect 502064 312588 502116 312594
rect 502064 312530 502116 312536
rect 502168 309806 502196 319058
rect 502156 309800 502208 309806
rect 502156 309742 502208 309748
rect 502260 278089 502288 322116
rect 502536 316878 502564 322116
rect 502812 319326 502840 322116
rect 502800 319320 502852 319326
rect 502800 319262 502852 319268
rect 502524 316872 502576 316878
rect 502524 316814 502576 316820
rect 503088 316034 503116 322116
rect 503272 322102 503378 322130
rect 503548 322102 503654 322130
rect 503930 322102 505048 322130
rect 503088 316006 503208 316034
rect 503180 314090 503208 316006
rect 503168 314084 503220 314090
rect 503168 314026 503220 314032
rect 503272 308514 503300 322102
rect 503548 309942 503576 322102
rect 503536 309936 503588 309942
rect 503536 309878 503588 309884
rect 503260 308508 503312 308514
rect 503260 308450 503312 308456
rect 502246 278080 502302 278089
rect 502246 278015 502302 278024
rect 500776 272536 500828 272542
rect 500776 272478 500828 272484
rect 500500 271244 500552 271250
rect 500500 271186 500552 271192
rect 499120 271176 499172 271182
rect 499120 271118 499172 271124
rect 505020 269958 505048 322102
rect 507136 289474 507164 322623
rect 507860 322312 507912 322318
rect 507860 322254 507912 322260
rect 507308 321700 507360 321706
rect 507308 321642 507360 321648
rect 507216 321156 507268 321162
rect 507216 321098 507268 321104
rect 507228 289542 507256 321098
rect 507320 291718 507348 321642
rect 507490 321464 507546 321473
rect 507490 321399 507546 321408
rect 507400 321224 507452 321230
rect 507400 321166 507452 321172
rect 507412 291786 507440 321166
rect 507504 295254 507532 321399
rect 507872 320142 507900 322254
rect 509344 320793 509372 322895
rect 509330 320784 509386 320793
rect 509330 320719 509386 320728
rect 507860 320136 507912 320142
rect 507860 320078 507912 320084
rect 509436 302802 509464 357575
rect 509528 326398 509556 366959
rect 509790 351792 509846 351801
rect 509790 351727 509846 351736
rect 509606 344040 509662 344049
rect 509606 343975 509662 343984
rect 509516 326392 509568 326398
rect 509516 326334 509568 326340
rect 509516 326256 509568 326262
rect 509516 326198 509568 326204
rect 509528 316810 509556 326198
rect 509516 316804 509568 316810
rect 509516 316746 509568 316752
rect 509620 306066 509648 343975
rect 509698 328400 509754 328409
rect 509698 328335 509754 328344
rect 509608 306060 509660 306066
rect 509608 306002 509660 306008
rect 509424 302796 509476 302802
rect 509424 302738 509476 302744
rect 509712 297362 509740 328335
rect 509804 321706 509832 351727
rect 510066 330304 510122 330313
rect 510066 330239 510122 330248
rect 509882 327720 509938 327729
rect 509882 327655 509938 327664
rect 509792 321700 509844 321706
rect 509792 321642 509844 321648
rect 509896 302841 509924 327655
rect 509974 326088 510030 326097
rect 509974 326023 510030 326032
rect 509988 306134 510016 326023
rect 509976 306128 510028 306134
rect 509976 306070 510028 306076
rect 509882 302832 509938 302841
rect 509882 302767 509938 302776
rect 509700 297356 509752 297362
rect 509700 297298 509752 297304
rect 510080 295322 510108 330239
rect 510160 326392 510212 326398
rect 510160 326334 510212 326340
rect 510172 317257 510200 326334
rect 510632 319394 510660 518055
rect 510710 373824 510766 373833
rect 510710 373759 510766 373768
rect 510620 319388 510672 319394
rect 510620 319330 510672 319336
rect 510158 317248 510214 317257
rect 510158 317183 510214 317192
rect 510724 303414 510752 373759
rect 510802 359136 510858 359145
rect 510802 359071 510858 359080
rect 510712 303408 510764 303414
rect 510712 303350 510764 303356
rect 510816 302870 510844 359071
rect 510986 355872 511042 355881
rect 510986 355807 511042 355816
rect 510894 353152 510950 353161
rect 510894 353087 510950 353096
rect 510804 302864 510856 302870
rect 510804 302806 510856 302812
rect 510908 297294 510936 353087
rect 511000 303618 511028 355807
rect 511078 347712 511134 347721
rect 511078 347647 511134 347656
rect 511092 305930 511120 347647
rect 511170 346080 511226 346089
rect 511170 346015 511226 346024
rect 511184 305998 511212 346015
rect 511276 319666 511304 590650
rect 511356 576904 511408 576910
rect 511356 576846 511408 576852
rect 511368 319870 511396 576846
rect 511540 423564 511592 423570
rect 511540 423506 511592 423512
rect 511448 404388 511500 404394
rect 511448 404330 511500 404336
rect 511460 321502 511488 404330
rect 511552 388686 511580 423506
rect 511540 388680 511592 388686
rect 511540 388622 511592 388628
rect 513392 387122 513420 600086
rect 515404 599616 515456 599622
rect 515404 599558 515456 599564
rect 513380 387116 513432 387122
rect 513380 387058 513432 387064
rect 512092 386640 512144 386646
rect 512092 386582 512144 386588
rect 512000 386504 512052 386510
rect 512000 386446 512052 386452
rect 512012 374921 512040 386446
rect 512104 376009 512132 386582
rect 512552 386572 512604 386578
rect 512552 386514 512604 386520
rect 512276 386436 512328 386442
rect 512276 386378 512328 386384
rect 512288 378185 512316 386378
rect 512368 385076 512420 385082
rect 512368 385018 512420 385024
rect 512274 378176 512330 378185
rect 512274 378111 512330 378120
rect 512380 376553 512408 385018
rect 512458 382528 512514 382537
rect 512458 382463 512460 382472
rect 512512 382463 512514 382472
rect 512460 382434 512512 382440
rect 512458 381440 512514 381449
rect 512458 381375 512514 381384
rect 512472 380934 512500 381375
rect 512460 380928 512512 380934
rect 512460 380870 512512 380876
rect 512564 379930 512592 386514
rect 513194 384704 513250 384713
rect 513194 384639 513250 384648
rect 513208 383790 513236 384639
rect 513286 384160 513342 384169
rect 513286 384095 513342 384104
rect 513196 383784 513248 383790
rect 513196 383726 513248 383732
rect 513300 383722 513328 384095
rect 513288 383716 513340 383722
rect 513288 383658 513340 383664
rect 512642 383616 512698 383625
rect 512642 383551 512698 383560
rect 512656 382974 512684 383551
rect 513010 383072 513066 383081
rect 513010 383007 513066 383016
rect 512644 382968 512696 382974
rect 512644 382910 512696 382916
rect 513024 382770 513052 383007
rect 513012 382764 513064 382770
rect 513012 382706 513064 382712
rect 513010 381984 513066 381993
rect 513010 381919 513066 381928
rect 512472 379902 512592 379930
rect 512472 377641 512500 379902
rect 512550 379808 512606 379817
rect 512550 379743 512552 379752
rect 512604 379743 512606 379752
rect 512552 379714 512604 379720
rect 512826 379264 512882 379273
rect 512826 379199 512882 379208
rect 512840 378282 512868 379199
rect 512828 378276 512880 378282
rect 512828 378218 512880 378224
rect 512458 377632 512514 377641
rect 512458 377567 512514 377576
rect 512366 376544 512422 376553
rect 512366 376479 512422 376488
rect 513024 376038 513052 381919
rect 513194 380896 513250 380905
rect 513194 380831 513250 380840
rect 513208 377466 513236 380831
rect 513286 380352 513342 380361
rect 513286 380287 513342 380296
rect 513300 379574 513328 380287
rect 513288 379568 513340 379574
rect 513288 379510 513340 379516
rect 513286 378720 513342 378729
rect 513286 378655 513342 378664
rect 513300 378350 513328 378655
rect 513288 378344 513340 378350
rect 513288 378286 513340 378292
rect 514024 378208 514076 378214
rect 514024 378150 514076 378156
rect 513196 377460 513248 377466
rect 513196 377402 513248 377408
rect 513194 377088 513250 377097
rect 513194 377023 513250 377032
rect 513208 376786 513236 377023
rect 513196 376780 513248 376786
rect 513196 376722 513248 376728
rect 513012 376032 513064 376038
rect 512090 376000 512146 376009
rect 513012 375974 513064 375980
rect 512090 375935 512146 375944
rect 511998 374912 512054 374921
rect 511998 374847 512054 374856
rect 513286 374368 513342 374377
rect 513286 374303 513342 374312
rect 513300 374202 513328 374303
rect 513288 374196 513340 374202
rect 513288 374138 513340 374144
rect 512642 373280 512698 373289
rect 512642 373215 512698 373224
rect 512656 372638 512684 373215
rect 513286 372736 513342 372745
rect 513286 372671 513288 372680
rect 513340 372671 513342 372680
rect 513288 372642 513340 372648
rect 512644 372632 512696 372638
rect 512644 372574 512696 372580
rect 511998 372192 512054 372201
rect 511998 372127 512054 372136
rect 512012 371754 512040 372127
rect 512000 371748 512052 371754
rect 512000 371690 512052 371696
rect 513840 371748 513892 371754
rect 513840 371690 513892 371696
rect 511998 371648 512054 371657
rect 511998 371583 512054 371592
rect 512012 369050 512040 371583
rect 512090 371104 512146 371113
rect 512090 371039 512146 371048
rect 512104 370258 512132 371039
rect 513286 370560 513342 370569
rect 513286 370495 513342 370504
rect 512092 370252 512144 370258
rect 512092 370194 512144 370200
rect 513300 370122 513328 370495
rect 513288 370116 513340 370122
rect 513288 370058 513340 370064
rect 513286 370016 513342 370025
rect 513286 369951 513342 369960
rect 513300 369918 513328 369951
rect 513288 369912 513340 369918
rect 513288 369854 513340 369860
rect 512090 369472 512146 369481
rect 512090 369407 512146 369416
rect 512104 369170 512132 369407
rect 512092 369164 512144 369170
rect 512092 369106 512144 369112
rect 512012 369022 512132 369050
rect 511998 365664 512054 365673
rect 511998 365599 512000 365608
rect 512052 365599 512054 365608
rect 512000 365570 512052 365576
rect 511998 364032 512054 364041
rect 511998 363967 512054 363976
rect 512012 363254 512040 363967
rect 512000 363248 512052 363254
rect 512000 363190 512052 363196
rect 511998 362400 512054 362409
rect 511998 362335 512000 362344
rect 512052 362335 512054 362344
rect 512000 362306 512052 362312
rect 511998 360768 512054 360777
rect 511998 360703 512054 360712
rect 512012 360466 512040 360703
rect 512000 360460 512052 360466
rect 512000 360402 512052 360408
rect 512104 354674 512132 369022
rect 512274 368928 512330 368937
rect 512274 368863 512330 368872
rect 512288 368626 512316 368863
rect 512276 368620 512328 368626
rect 512276 368562 512328 368568
rect 512182 368384 512238 368393
rect 512182 368319 512238 368328
rect 512012 354646 512132 354674
rect 511448 321496 511500 321502
rect 511448 321438 511500 321444
rect 511356 319864 511408 319870
rect 511356 319806 511408 319812
rect 511264 319660 511316 319666
rect 511264 319602 511316 319608
rect 511172 305992 511224 305998
rect 511172 305934 511224 305940
rect 511080 305924 511132 305930
rect 511080 305866 511132 305872
rect 512012 304366 512040 354646
rect 512090 354240 512146 354249
rect 512090 354175 512092 354184
rect 512144 354175 512146 354184
rect 512092 354146 512144 354152
rect 512090 349344 512146 349353
rect 512090 349279 512092 349288
rect 512144 349279 512146 349288
rect 512092 349250 512144 349256
rect 512090 347168 512146 347177
rect 512090 347103 512146 347112
rect 512104 346798 512132 347103
rect 512092 346792 512144 346798
rect 512092 346734 512144 346740
rect 512090 344992 512146 345001
rect 512090 344927 512146 344936
rect 512104 318170 512132 344927
rect 512092 318164 512144 318170
rect 512092 318106 512144 318112
rect 512000 304360 512052 304366
rect 512000 304302 512052 304308
rect 512196 304298 512224 368319
rect 513286 367840 513342 367849
rect 513286 367775 513342 367784
rect 513300 367402 513328 367775
rect 513288 367396 513340 367402
rect 513288 367338 513340 367344
rect 513286 366752 513342 366761
rect 513286 366687 513342 366696
rect 513300 365770 513328 366687
rect 513378 366208 513434 366217
rect 513378 366143 513434 366152
rect 513288 365764 513340 365770
rect 513288 365706 513340 365712
rect 512826 365120 512882 365129
rect 512826 365055 512882 365064
rect 513288 365084 513340 365090
rect 512840 364410 512868 365055
rect 513288 365026 513340 365032
rect 513300 364585 513328 365026
rect 513286 364576 513342 364585
rect 513286 364511 513342 364520
rect 512828 364404 512880 364410
rect 512828 364346 512880 364352
rect 512274 363488 512330 363497
rect 512274 363423 512330 363432
rect 512184 304292 512236 304298
rect 512184 304234 512236 304240
rect 510988 303612 511040 303618
rect 510988 303554 511040 303560
rect 512288 301510 512316 363423
rect 513010 362944 513066 362953
rect 513010 362879 513066 362888
rect 513024 361690 513052 362879
rect 513286 361856 513342 361865
rect 513286 361791 513342 361800
rect 513012 361684 513064 361690
rect 513012 361626 513064 361632
rect 513300 361622 513328 361791
rect 513288 361616 513340 361622
rect 513288 361558 513340 361564
rect 512642 361312 512698 361321
rect 512642 361247 512698 361256
rect 512656 360738 512684 361247
rect 512644 360732 512696 360738
rect 512644 360674 512696 360680
rect 512366 360224 512422 360233
rect 512366 360159 512422 360168
rect 512380 304434 512408 360159
rect 513010 359680 513066 359689
rect 513010 359615 513066 359624
rect 513024 358834 513052 359615
rect 513012 358828 513064 358834
rect 513012 358770 513064 358776
rect 512550 358592 512606 358601
rect 512550 358527 512606 358536
rect 512458 352608 512514 352617
rect 512458 352543 512514 352552
rect 512472 352306 512500 352543
rect 512460 352300 512512 352306
rect 512460 352242 512512 352248
rect 512458 350976 512514 350985
rect 512458 350911 512514 350920
rect 512472 350878 512500 350911
rect 512460 350872 512512 350878
rect 512460 350814 512512 350820
rect 512458 345536 512514 345545
rect 512458 345471 512514 345480
rect 512368 304428 512420 304434
rect 512368 304370 512420 304376
rect 512472 302938 512500 345471
rect 512564 317121 512592 358527
rect 513286 356960 513342 356969
rect 513286 356895 513342 356904
rect 512826 356416 512882 356425
rect 512826 356351 512828 356360
rect 512880 356351 512882 356360
rect 512828 356322 512880 356328
rect 513300 356250 513328 356895
rect 513288 356244 513340 356250
rect 513288 356186 513340 356192
rect 513286 355328 513342 355337
rect 513286 355263 513342 355272
rect 513300 355026 513328 355263
rect 513288 355020 513340 355026
rect 513288 354962 513340 354968
rect 513286 354784 513342 354793
rect 513286 354719 513288 354728
rect 513340 354719 513342 354728
rect 513288 354690 513340 354696
rect 513286 353696 513342 353705
rect 513286 353631 513342 353640
rect 513300 353530 513328 353631
rect 513288 353524 513340 353530
rect 513288 353466 513340 353472
rect 512918 351520 512974 351529
rect 512918 351455 512974 351464
rect 512932 350674 512960 351455
rect 512920 350668 512972 350674
rect 512920 350610 512972 350616
rect 513286 350432 513342 350441
rect 513286 350367 513342 350376
rect 512826 349888 512882 349897
rect 512826 349823 512882 349832
rect 512840 349722 512868 349823
rect 512828 349716 512880 349722
rect 512828 349658 512880 349664
rect 513300 349450 513328 350367
rect 513288 349444 513340 349450
rect 513288 349386 513340 349392
rect 513286 348800 513342 348809
rect 513286 348735 513342 348744
rect 513300 348498 513328 348735
rect 513288 348492 513340 348498
rect 513288 348434 513340 348440
rect 513286 348256 513342 348265
rect 513286 348191 513288 348200
rect 513340 348191 513342 348200
rect 513288 348162 513340 348168
rect 512642 346624 512698 346633
rect 512642 346559 512644 346568
rect 512696 346559 512698 346568
rect 512644 346530 512696 346536
rect 512918 343904 512974 343913
rect 512918 343839 512974 343848
rect 512932 343738 512960 343839
rect 512920 343732 512972 343738
rect 512920 343674 512972 343680
rect 513194 343360 513250 343369
rect 513194 343295 513250 343304
rect 513208 342650 513236 343295
rect 513196 342644 513248 342650
rect 513196 342586 513248 342592
rect 513288 342304 513340 342310
rect 513286 342272 513288 342281
rect 513340 342272 513342 342281
rect 513286 342207 513342 342216
rect 512642 341728 512698 341737
rect 512642 341663 512698 341672
rect 512656 341290 512684 341663
rect 512644 341284 512696 341290
rect 512644 341226 512696 341232
rect 512826 341184 512882 341193
rect 512826 341119 512882 341128
rect 512840 341018 512868 341119
rect 512828 341012 512880 341018
rect 512828 340954 512880 340960
rect 513194 340640 513250 340649
rect 513194 340575 513250 340584
rect 513208 339522 513236 340575
rect 513286 340096 513342 340105
rect 513286 340031 513288 340040
rect 513340 340031 513342 340040
rect 513288 340002 513340 340008
rect 513196 339516 513248 339522
rect 513196 339458 513248 339464
rect 512734 339008 512790 339017
rect 512734 338943 512790 338952
rect 512642 333024 512698 333033
rect 512642 332959 512698 332968
rect 512656 332926 512684 332959
rect 512644 332920 512696 332926
rect 512644 332862 512696 332868
rect 512642 332480 512698 332489
rect 512642 332415 512698 332424
rect 512656 331498 512684 332415
rect 512644 331492 512696 331498
rect 512644 331434 512696 331440
rect 512748 331214 512776 338943
rect 513288 338564 513340 338570
rect 513288 338506 513340 338512
rect 513300 338473 513328 338506
rect 513286 338464 513342 338473
rect 513286 338399 513342 338408
rect 513102 337920 513158 337929
rect 513102 337855 513158 337864
rect 513116 337210 513144 337855
rect 513194 337376 513250 337385
rect 513194 337311 513250 337320
rect 513288 337340 513340 337346
rect 513104 337204 513156 337210
rect 513104 337146 513156 337152
rect 513208 336802 513236 337311
rect 513288 337282 513340 337288
rect 513300 336841 513328 337282
rect 513286 336832 513342 336841
rect 513196 336796 513248 336802
rect 513286 336767 513342 336776
rect 513196 336738 513248 336744
rect 512826 336288 512882 336297
rect 512826 336223 512882 336232
rect 512656 331186 512776 331214
rect 512550 317112 512606 317121
rect 512550 317047 512606 317056
rect 512656 305658 512684 331186
rect 512734 325408 512790 325417
rect 512734 325343 512790 325352
rect 512748 305726 512776 325343
rect 512736 305720 512788 305726
rect 512736 305662 512788 305668
rect 512644 305652 512696 305658
rect 512644 305594 512696 305600
rect 512460 302932 512512 302938
rect 512460 302874 512512 302880
rect 512276 301504 512328 301510
rect 512276 301446 512328 301452
rect 510896 297288 510948 297294
rect 510896 297230 510948 297236
rect 510068 295316 510120 295322
rect 510068 295258 510120 295264
rect 507492 295248 507544 295254
rect 507492 295190 507544 295196
rect 507400 291780 507452 291786
rect 507400 291722 507452 291728
rect 507308 291712 507360 291718
rect 507308 291654 507360 291660
rect 507216 289536 507268 289542
rect 507216 289478 507268 289484
rect 507124 289468 507176 289474
rect 507124 289410 507176 289416
rect 505008 269952 505060 269958
rect 505008 269894 505060 269900
rect 512840 269822 512868 336223
rect 513286 335744 513342 335753
rect 513286 335679 513342 335688
rect 513300 335374 513328 335679
rect 513288 335368 513340 335374
rect 513288 335310 513340 335316
rect 513286 335200 513342 335209
rect 513286 335135 513342 335144
rect 513300 334626 513328 335135
rect 513288 334620 513340 334626
rect 513288 334562 513340 334568
rect 513286 334112 513342 334121
rect 513286 334047 513342 334056
rect 513300 334014 513328 334047
rect 513288 334008 513340 334014
rect 513288 333950 513340 333956
rect 513010 333568 513066 333577
rect 513010 333503 513066 333512
rect 513024 333130 513052 333503
rect 513012 333124 513064 333130
rect 513012 333066 513064 333072
rect 513392 297906 513420 366143
rect 513656 362364 513708 362370
rect 513656 362306 513708 362312
rect 513562 358048 513618 358057
rect 513562 357983 513618 357992
rect 513470 329216 513526 329225
rect 513470 329151 513526 329160
rect 513484 321230 513512 329151
rect 513472 321224 513524 321230
rect 513472 321166 513524 321172
rect 513576 298110 513604 357983
rect 513668 303210 513696 362306
rect 513748 354204 513800 354210
rect 513748 354146 513800 354152
rect 513760 303482 513788 354146
rect 513852 321094 513880 371690
rect 513932 349308 513984 349314
rect 513932 349250 513984 349256
rect 513840 321088 513892 321094
rect 513840 321030 513892 321036
rect 513944 305862 513972 349250
rect 514036 321366 514064 378150
rect 514760 370252 514812 370258
rect 514760 370194 514812 370200
rect 514208 365628 514260 365634
rect 514208 365570 514260 365576
rect 514116 332920 514168 332926
rect 514116 332862 514168 332868
rect 514024 321360 514076 321366
rect 514024 321302 514076 321308
rect 514128 316985 514156 332862
rect 514114 316976 514170 316985
rect 514114 316911 514170 316920
rect 513932 305856 513984 305862
rect 513932 305798 513984 305804
rect 513748 303476 513800 303482
rect 513748 303418 513800 303424
rect 514220 303346 514248 365570
rect 514208 303340 514260 303346
rect 514208 303282 514260 303288
rect 513656 303204 513708 303210
rect 513656 303146 513708 303152
rect 513564 298104 513616 298110
rect 513564 298046 513616 298052
rect 513380 297900 513432 297906
rect 513380 297842 513432 297848
rect 514772 297702 514800 370194
rect 515128 368620 515180 368626
rect 515128 368562 515180 368568
rect 514852 363248 514904 363254
rect 514852 363190 514904 363196
rect 514864 303074 514892 363190
rect 514944 360460 514996 360466
rect 514944 360402 514996 360408
rect 514956 303142 514984 360402
rect 515036 346792 515088 346798
rect 515036 346734 515088 346740
rect 514944 303136 514996 303142
rect 514944 303078 514996 303084
rect 514852 303068 514904 303074
rect 514852 303010 514904 303016
rect 514760 297696 514812 297702
rect 514760 297638 514812 297644
rect 515048 292534 515076 346734
rect 515140 316849 515168 368562
rect 515220 352300 515272 352306
rect 515220 352242 515272 352248
rect 515126 316840 515182 316849
rect 515126 316775 515182 316784
rect 515232 303550 515260 352242
rect 515312 341284 515364 341290
rect 515312 341226 515364 341232
rect 515220 303544 515272 303550
rect 515220 303486 515272 303492
rect 515324 294982 515352 341226
rect 515416 319734 515444 599558
rect 515496 563100 515548 563106
rect 515496 563042 515548 563048
rect 515508 322658 515536 563042
rect 519544 536852 519596 536858
rect 519544 536794 519596 536800
rect 518164 524476 518216 524482
rect 518164 524418 518216 524424
rect 516784 510672 516836 510678
rect 516784 510614 516836 510620
rect 515588 382492 515640 382498
rect 515588 382434 515640 382440
rect 515600 358494 515628 382434
rect 515680 379772 515732 379778
rect 515680 379714 515732 379720
rect 515692 359854 515720 379714
rect 515680 359848 515732 359854
rect 515680 359790 515732 359796
rect 515588 358488 515640 358494
rect 515588 358430 515640 358436
rect 516232 356380 516284 356386
rect 516232 356322 516284 356328
rect 515588 350872 515640 350878
rect 515588 350814 515640 350820
rect 515496 322652 515548 322658
rect 515496 322594 515548 322600
rect 515404 319728 515456 319734
rect 515404 319670 515456 319676
rect 515600 305794 515628 350814
rect 516140 331492 516192 331498
rect 516140 331434 516192 331440
rect 516152 321162 516180 331434
rect 516140 321156 516192 321162
rect 516140 321098 516192 321104
rect 515588 305788 515640 305794
rect 515588 305730 515640 305736
rect 516244 297974 516272 356322
rect 516324 350668 516376 350674
rect 516324 350610 516376 350616
rect 516336 300286 516364 350610
rect 516508 346588 516560 346594
rect 516508 346530 516560 346536
rect 516416 343732 516468 343738
rect 516416 343674 516468 343680
rect 516324 300280 516376 300286
rect 516324 300222 516376 300228
rect 516232 297968 516284 297974
rect 516232 297910 516284 297916
rect 515312 294976 515364 294982
rect 515312 294918 515364 294924
rect 516428 294914 516456 343674
rect 516520 300354 516548 346530
rect 516600 341012 516652 341018
rect 516600 340954 516652 340960
rect 516612 300558 516640 340954
rect 516692 333124 516744 333130
rect 516692 333066 516744 333072
rect 516600 300552 516652 300558
rect 516600 300494 516652 300500
rect 516508 300348 516560 300354
rect 516508 300290 516560 300296
rect 516704 295050 516732 333066
rect 516796 322726 516824 510614
rect 516968 376780 517020 376786
rect 516968 376722 517020 376728
rect 516876 337204 516928 337210
rect 516876 337146 516928 337152
rect 516784 322720 516836 322726
rect 516784 322662 516836 322668
rect 516888 300490 516916 337146
rect 516980 300626 517008 376722
rect 517520 374196 517572 374202
rect 517520 374138 517572 374144
rect 516968 300620 517020 300626
rect 516968 300562 517020 300568
rect 516876 300484 516928 300490
rect 516876 300426 516928 300432
rect 517532 295186 517560 374138
rect 517612 370116 517664 370122
rect 517612 370058 517664 370064
rect 517624 303006 517652 370058
rect 517704 355020 517756 355026
rect 517704 354962 517756 354968
rect 517612 303000 517664 303006
rect 517612 302942 517664 302948
rect 517520 295180 517572 295186
rect 517520 295122 517572 295128
rect 516692 295044 516744 295050
rect 516692 294986 516744 294992
rect 516416 294908 516468 294914
rect 516416 294850 516468 294856
rect 515036 292528 515088 292534
rect 515036 292470 515088 292476
rect 517716 292330 517744 354962
rect 517888 354748 517940 354754
rect 517888 354690 517940 354696
rect 517796 353524 517848 353530
rect 517796 353466 517848 353472
rect 517808 292398 517836 353466
rect 517900 298042 517928 354690
rect 517980 349716 518032 349722
rect 517980 349658 518032 349664
rect 517992 300150 518020 349658
rect 518072 348220 518124 348226
rect 518072 348162 518124 348168
rect 518084 300218 518112 348162
rect 518176 321434 518204 524418
rect 518256 484424 518308 484430
rect 518256 484366 518308 484372
rect 518268 322522 518296 484366
rect 518348 382764 518400 382770
rect 518348 382706 518400 382712
rect 518360 358630 518388 382706
rect 518900 372700 518952 372706
rect 518900 372642 518952 372648
rect 518348 358624 518400 358630
rect 518348 358566 518400 358572
rect 518348 342644 518400 342650
rect 518348 342586 518400 342592
rect 518256 322516 518308 322522
rect 518256 322458 518308 322464
rect 518164 321428 518216 321434
rect 518164 321370 518216 321376
rect 518360 300422 518388 342586
rect 518348 300416 518400 300422
rect 518348 300358 518400 300364
rect 518072 300212 518124 300218
rect 518072 300154 518124 300160
rect 517980 300144 518032 300150
rect 517980 300086 518032 300092
rect 517888 298036 517940 298042
rect 517888 297978 517940 297984
rect 518912 295118 518940 372642
rect 519084 365084 519136 365090
rect 519084 365026 519136 365032
rect 518992 364404 519044 364410
rect 518992 364346 519044 364352
rect 518900 295112 518952 295118
rect 518900 295054 518952 295060
rect 517796 292392 517848 292398
rect 517796 292334 517848 292340
rect 517704 292324 517756 292330
rect 517704 292266 517756 292272
rect 519004 292194 519032 364346
rect 519096 297566 519124 365026
rect 519176 361684 519228 361690
rect 519176 361626 519228 361632
rect 519188 297770 519216 361626
rect 519268 358828 519320 358834
rect 519268 358770 519320 358776
rect 519280 297838 519308 358770
rect 519360 349444 519412 349450
rect 519360 349386 519412 349392
rect 519268 297832 519320 297838
rect 519268 297774 519320 297780
rect 519176 297764 519228 297770
rect 519176 297706 519228 297712
rect 519084 297560 519136 297566
rect 519084 297502 519136 297508
rect 519372 292262 519400 349386
rect 519452 340060 519504 340066
rect 519452 340002 519504 340008
rect 519464 294642 519492 340002
rect 519556 319938 519584 536794
rect 520292 520946 520320 600086
rect 526732 598262 526760 600100
rect 526720 598256 526772 598262
rect 526720 598198 526772 598204
rect 520280 520940 520332 520946
rect 520280 520882 520332 520888
rect 547878 516760 547934 516769
rect 547878 516695 547934 516704
rect 545120 514072 545172 514078
rect 545120 514014 545172 514020
rect 535460 512644 535512 512650
rect 535460 512586 535512 512592
rect 532700 508564 532752 508570
rect 532700 508506 532752 508512
rect 529940 505776 529992 505782
rect 529940 505718 529992 505724
rect 519634 502344 519690 502353
rect 519634 502279 519690 502288
rect 519544 319932 519596 319938
rect 519544 319874 519596 319880
rect 519648 319802 519676 502279
rect 529952 480254 529980 505718
rect 532712 480254 532740 508506
rect 535472 480254 535500 512586
rect 538220 509924 538272 509930
rect 538220 509866 538272 509872
rect 538232 480254 538260 509866
rect 529952 480226 530256 480254
rect 532712 480226 533200 480254
rect 535472 480226 536144 480254
rect 538232 480226 539088 480254
rect 521750 462904 521806 462913
rect 521750 462839 521806 462848
rect 521764 460972 521792 462839
rect 527640 462528 527692 462534
rect 527640 462470 527692 462476
rect 524696 462460 524748 462466
rect 524696 462402 524748 462408
rect 524708 460972 524736 462402
rect 527652 460972 527680 462470
rect 530228 460986 530256 480226
rect 533172 460986 533200 480226
rect 536116 460986 536144 480226
rect 539060 460986 539088 480226
rect 542360 462392 542412 462398
rect 542360 462334 542412 462340
rect 530228 460958 530610 460986
rect 533172 460958 533554 460986
rect 536116 460958 536498 460986
rect 539060 460958 539442 460986
rect 542372 460972 542400 462334
rect 545132 460986 545160 514014
rect 547892 460986 547920 516695
rect 553860 461032 553912 461038
rect 545132 460958 545330 460986
rect 547892 460958 548274 460986
rect 550928 460970 551218 460986
rect 553912 460980 554162 460986
rect 553860 460974 554162 460980
rect 550916 460964 551218 460970
rect 550968 460958 551218 460964
rect 553872 460958 554162 460974
rect 550916 460906 550968 460912
rect 569224 456816 569276 456822
rect 569224 456758 569276 456764
rect 557538 442912 557594 442921
rect 557538 442847 557594 442856
rect 521212 421598 521240 425068
rect 522304 423496 522356 423502
rect 522304 423438 522356 423444
rect 521200 421592 521252 421598
rect 521200 421534 521252 421540
rect 522316 388754 522344 423438
rect 522500 423434 522528 425068
rect 523788 423570 523816 425068
rect 524708 425054 525090 425082
rect 523776 423564 523828 423570
rect 523776 423506 523828 423512
rect 522488 423428 522540 423434
rect 522488 423370 522540 423376
rect 523684 423428 523736 423434
rect 523684 423370 523736 423376
rect 523696 388822 523724 423370
rect 524708 412634 524736 425054
rect 526364 423366 526392 425068
rect 526352 423360 526404 423366
rect 526352 423302 526404 423308
rect 526444 423360 526496 423366
rect 526444 423302 526496 423308
rect 524432 412606 524736 412634
rect 523684 388816 523736 388822
rect 523684 388758 523736 388764
rect 522304 388748 522356 388754
rect 522304 388690 522356 388696
rect 524432 388618 524460 412606
rect 526456 388890 526484 423302
rect 527652 416090 527680 425068
rect 528940 423298 528968 425068
rect 530228 423638 530256 425068
rect 529204 423632 529256 423638
rect 529204 423574 529256 423580
rect 530216 423632 530268 423638
rect 530216 423574 530268 423580
rect 530584 423632 530636 423638
rect 530584 423574 530636 423580
rect 528928 423292 528980 423298
rect 528928 423234 528980 423240
rect 527640 416084 527692 416090
rect 527640 416026 527692 416032
rect 526444 388884 526496 388890
rect 526444 388826 526496 388832
rect 524420 388612 524472 388618
rect 524420 388554 524472 388560
rect 529216 388550 529244 423574
rect 529204 388544 529256 388550
rect 529204 388486 529256 388492
rect 530596 388482 530624 423574
rect 531516 423230 531544 425068
rect 532804 423638 532832 425068
rect 532792 423632 532844 423638
rect 532792 423574 532844 423580
rect 531504 423224 531556 423230
rect 531504 423166 531556 423172
rect 534092 389842 534120 425068
rect 535012 425054 535394 425082
rect 536300 425054 536682 425082
rect 537588 425054 537970 425082
rect 538876 425054 539258 425082
rect 540164 425054 540546 425082
rect 535012 412634 535040 425054
rect 536300 412634 536328 425054
rect 537588 412634 537616 425054
rect 538876 412634 538904 425054
rect 540164 412634 540192 425054
rect 541820 420238 541848 425068
rect 542740 425054 543122 425082
rect 544028 425054 544410 425082
rect 541808 420232 541860 420238
rect 541808 420174 541860 420180
rect 542740 412634 542768 425054
rect 544028 412634 544056 425054
rect 545684 423162 545712 425068
rect 546604 425054 546986 425082
rect 545672 423156 545724 423162
rect 545672 423098 545724 423104
rect 546604 412634 546632 425054
rect 548260 423094 548288 425068
rect 549548 423502 549576 425068
rect 549536 423496 549588 423502
rect 549536 423438 549588 423444
rect 548248 423088 548300 423094
rect 548248 423030 548300 423036
rect 550836 423026 550864 425068
rect 552124 423434 552152 425068
rect 552112 423428 552164 423434
rect 552112 423370 552164 423376
rect 550824 423020 550876 423026
rect 550824 422962 550876 422968
rect 553412 422958 553440 425068
rect 554700 423366 554728 425068
rect 557552 424386 557580 442847
rect 557540 424380 557592 424386
rect 557540 424322 557592 424328
rect 554688 423360 554740 423366
rect 554688 423302 554740 423308
rect 553400 422952 553452 422958
rect 553400 422894 553452 422900
rect 534184 412606 535040 412634
rect 535472 412606 536328 412634
rect 536852 412606 537616 412634
rect 538232 412606 538904 412634
rect 539612 412606 540192 412634
rect 542372 412606 542768 412634
rect 543752 412606 544056 412634
rect 546512 412606 546632 412634
rect 534184 392630 534212 412606
rect 535472 395350 535500 412606
rect 536852 396778 536880 412606
rect 538232 398138 538260 412606
rect 539612 399498 539640 412606
rect 539600 399492 539652 399498
rect 539600 399434 539652 399440
rect 538220 398132 538272 398138
rect 538220 398074 538272 398080
rect 536840 396772 536892 396778
rect 536840 396714 536892 396720
rect 535460 395344 535512 395350
rect 535460 395286 535512 395292
rect 534172 392624 534224 392630
rect 534172 392566 534224 392572
rect 542372 391338 542400 412606
rect 543752 394058 543780 412606
rect 546512 400926 546540 412606
rect 546500 400920 546552 400926
rect 546500 400862 546552 400868
rect 543740 394052 543792 394058
rect 543740 393994 543792 394000
rect 542360 391332 542412 391338
rect 542360 391274 542412 391280
rect 534080 389836 534132 389842
rect 534080 389778 534132 389784
rect 530584 388476 530636 388482
rect 530584 388418 530636 388424
rect 553952 386708 554004 386714
rect 553952 386650 554004 386656
rect 534724 383784 534776 383790
rect 534724 383726 534776 383732
rect 519728 382968 519780 382974
rect 519728 382910 519780 382916
rect 519740 358698 519768 382910
rect 522304 378344 522356 378350
rect 522304 378286 522356 378292
rect 521660 372632 521712 372638
rect 521660 372574 521712 372580
rect 520280 369164 520332 369170
rect 520280 369106 520332 369112
rect 519728 358692 519780 358698
rect 519728 358634 519780 358640
rect 519728 337340 519780 337346
rect 519728 337282 519780 337288
rect 519636 319796 519688 319802
rect 519636 319738 519688 319744
rect 519740 294846 519768 337282
rect 520292 297498 520320 369106
rect 520372 367396 520424 367402
rect 520372 367338 520424 367344
rect 520280 297492 520332 297498
rect 520280 297434 520332 297440
rect 520384 297430 520412 367338
rect 520556 360732 520608 360738
rect 520556 360674 520608 360680
rect 520464 356244 520516 356250
rect 520464 356186 520516 356192
rect 520372 297424 520424 297430
rect 520372 297366 520424 297372
rect 519728 294840 519780 294846
rect 519728 294782 519780 294788
rect 519452 294636 519504 294642
rect 519452 294578 519504 294584
rect 519360 292256 519412 292262
rect 519360 292198 519412 292204
rect 518992 292188 519044 292194
rect 518992 292130 519044 292136
rect 520476 292126 520504 356186
rect 520568 297634 520596 360674
rect 520648 348492 520700 348498
rect 520648 348434 520700 348440
rect 520556 297628 520608 297634
rect 520556 297570 520608 297576
rect 520660 292466 520688 348434
rect 520740 338564 520792 338570
rect 520740 338506 520792 338512
rect 520752 294778 520780 338506
rect 520832 334620 520884 334626
rect 520832 334562 520884 334568
rect 520740 294772 520792 294778
rect 520740 294714 520792 294720
rect 520844 294710 520872 334562
rect 520832 294704 520884 294710
rect 520832 294646 520884 294652
rect 520648 292460 520700 292466
rect 520648 292402 520700 292408
rect 520464 292120 520516 292126
rect 520464 292062 520516 292068
rect 521672 291854 521700 372574
rect 521752 365764 521804 365770
rect 521752 365706 521804 365712
rect 521764 292058 521792 365706
rect 522316 359786 522344 378286
rect 523040 369912 523092 369918
rect 523040 369854 523092 369860
rect 522304 359780 522356 359786
rect 522304 359722 522356 359728
rect 521844 342304 521896 342310
rect 521844 342246 521896 342252
rect 521752 292052 521804 292058
rect 521752 291994 521804 292000
rect 521660 291848 521712 291854
rect 521660 291790 521712 291796
rect 521856 289338 521884 342246
rect 521936 339516 521988 339522
rect 521936 339458 521988 339464
rect 521844 289332 521896 289338
rect 521844 289274 521896 289280
rect 521948 289270 521976 339458
rect 522028 336796 522080 336802
rect 522028 336738 522080 336744
rect 521936 289264 521988 289270
rect 521936 289206 521988 289212
rect 522040 289134 522068 336738
rect 522120 335368 522172 335374
rect 522120 335310 522172 335316
rect 522132 289202 522160 335310
rect 522212 334008 522264 334014
rect 522212 333950 522264 333956
rect 522224 289406 522252 333950
rect 523052 291990 523080 369854
rect 523132 361616 523184 361622
rect 523132 361558 523184 361564
rect 523040 291984 523092 291990
rect 523040 291926 523092 291932
rect 523144 291922 523172 361558
rect 534736 360126 534764 383726
rect 548524 383716 548576 383722
rect 548524 383658 548576 383664
rect 547144 380928 547196 380934
rect 547144 380870 547196 380876
rect 544384 376032 544436 376038
rect 544384 375974 544436 375980
rect 534724 360120 534776 360126
rect 534724 360062 534776 360068
rect 544396 358562 544424 375974
rect 547156 359922 547184 380870
rect 547236 378276 547288 378282
rect 547236 378218 547288 378224
rect 547248 360194 547276 378218
rect 547236 360188 547288 360194
rect 547236 360130 547288 360136
rect 548536 359990 548564 383658
rect 549904 379568 549956 379574
rect 549904 379510 549956 379516
rect 548616 377460 548668 377466
rect 548616 377402 548668 377408
rect 548524 359984 548576 359990
rect 548524 359926 548576 359932
rect 547144 359916 547196 359922
rect 547144 359858 547196 359864
rect 548628 358766 548656 377402
rect 549916 360058 549944 379510
rect 553964 377890 553992 386650
rect 563428 385144 563480 385150
rect 563428 385086 563480 385092
rect 553964 377862 554438 377890
rect 563440 377876 563468 385086
rect 552032 360194 552322 360210
rect 552020 360188 552322 360194
rect 552072 360182 552322 360188
rect 552020 360130 552072 360136
rect 566740 360120 566792 360126
rect 549904 360052 549956 360058
rect 549904 359994 549956 360000
rect 550836 359786 550864 360060
rect 553780 359854 553808 360060
rect 554976 360058 555266 360074
rect 554964 360052 555266 360058
rect 555016 360046 555266 360052
rect 554964 359994 555016 360000
rect 553768 359848 553820 359854
rect 553768 359790 553820 359796
rect 550824 359780 550876 359786
rect 550824 359722 550876 359728
rect 556724 358766 556752 360060
rect 558196 359922 558224 360060
rect 558184 359916 558236 359922
rect 558184 359858 558236 359864
rect 548616 358760 548668 358766
rect 548616 358702 548668 358708
rect 556712 358760 556764 358766
rect 556712 358702 556764 358708
rect 559668 358562 559696 360060
rect 544384 358556 544436 358562
rect 544384 358498 544436 358504
rect 559656 358556 559708 358562
rect 559656 358498 559708 358504
rect 561140 358494 561168 360060
rect 562612 358630 562640 360060
rect 564084 358698 564112 360060
rect 565280 360046 565570 360074
rect 566792 360068 567042 360074
rect 566740 360062 567042 360068
rect 566752 360046 567042 360062
rect 565280 359990 565308 360046
rect 565268 359984 565320 359990
rect 565268 359926 565320 359932
rect 564072 358692 564124 358698
rect 564072 358634 564124 358640
rect 562600 358624 562652 358630
rect 562600 358566 562652 358572
rect 561128 358488 561180 358494
rect 561128 358430 561180 358436
rect 569236 322794 569264 456758
rect 570616 322930 570644 616830
rect 573364 364404 573416 364410
rect 573364 364346 573416 364352
rect 570604 322924 570656 322930
rect 570604 322866 570656 322872
rect 569224 322788 569276 322794
rect 569224 322730 569276 322736
rect 573376 321570 573404 364346
rect 573364 321564 573416 321570
rect 573364 321506 573416 321512
rect 576136 320006 576164 683130
rect 579618 617536 579674 617545
rect 579618 617471 579674 617480
rect 579632 616894 579660 617471
rect 579620 616888 579672 616894
rect 579620 616830 579672 616836
rect 580170 591016 580226 591025
rect 580170 590951 580226 590960
rect 580184 590714 580212 590951
rect 580172 590708 580224 590714
rect 580172 590650 580224 590656
rect 579986 577688 580042 577697
rect 579986 577623 580042 577632
rect 580000 576910 580028 577623
rect 579988 576904 580040 576910
rect 579988 576846 580040 576852
rect 580170 564360 580226 564369
rect 580170 564295 580226 564304
rect 580184 563106 580212 564295
rect 580172 563100 580224 563106
rect 580172 563042 580224 563048
rect 580170 537840 580226 537849
rect 580170 537775 580226 537784
rect 580184 536858 580212 537775
rect 580172 536852 580224 536858
rect 580172 536794 580224 536800
rect 580170 524512 580226 524521
rect 580170 524447 580172 524456
rect 580224 524447 580226 524456
rect 580172 524418 580224 524424
rect 580170 511320 580226 511329
rect 580170 511255 580226 511264
rect 580184 510678 580212 511255
rect 580172 510672 580224 510678
rect 580172 510614 580224 510620
rect 580170 484664 580226 484673
rect 580170 484599 580226 484608
rect 580184 484430 580212 484599
rect 580172 484424 580224 484430
rect 580172 484366 580224 484372
rect 580170 458144 580226 458153
rect 580170 458079 580226 458088
rect 580184 456822 580212 458079
rect 580172 456816 580224 456822
rect 580172 456758 580224 456764
rect 580170 404968 580226 404977
rect 580170 404903 580226 404912
rect 580184 404394 580212 404903
rect 580172 404388 580224 404394
rect 580172 404330 580224 404336
rect 580170 378448 580226 378457
rect 580170 378383 580226 378392
rect 580184 378214 580212 378383
rect 580172 378208 580224 378214
rect 580172 378150 580224 378156
rect 580170 365120 580226 365129
rect 580170 365055 580226 365064
rect 580184 364410 580212 365055
rect 580172 364404 580224 364410
rect 580172 364346 580224 364352
rect 580170 325272 580226 325281
rect 580170 325207 580226 325216
rect 580184 322250 580212 325207
rect 580276 322318 580304 697167
rect 580354 670712 580410 670721
rect 580354 670647 580410 670656
rect 580264 322312 580316 322318
rect 580264 322254 580316 322260
rect 580172 322244 580224 322250
rect 580172 322186 580224 322192
rect 580368 320958 580396 670647
rect 580538 644056 580594 644065
rect 580538 643991 580594 644000
rect 580446 630864 580502 630873
rect 580446 630799 580502 630808
rect 580356 320952 580408 320958
rect 580356 320894 580408 320900
rect 576124 320000 576176 320006
rect 576124 319942 576176 319948
rect 534724 319592 534776 319598
rect 534724 319534 534776 319540
rect 533344 319524 533396 319530
rect 533344 319466 533396 319472
rect 530584 319320 530636 319326
rect 530584 319262 530636 319268
rect 530032 309868 530084 309874
rect 530032 309810 530084 309816
rect 529940 308440 529992 308446
rect 529940 308382 529992 308388
rect 523132 291916 523184 291922
rect 523132 291858 523184 291864
rect 522212 289400 522264 289406
rect 522212 289342 522264 289348
rect 522120 289196 522172 289202
rect 522120 289138 522172 289144
rect 522028 289128 522080 289134
rect 522028 289070 522080 289076
rect 512828 269816 512880 269822
rect 512828 269758 512880 269764
rect 490380 268456 490432 268462
rect 490380 268398 490432 268404
rect 497740 268456 497792 268462
rect 497740 268398 497792 268404
rect 466368 268388 466420 268394
rect 466368 268330 466420 268336
rect 529952 209273 529980 308382
rect 530044 226250 530072 309810
rect 530124 275392 530176 275398
rect 530124 275334 530176 275340
rect 530136 261089 530164 275334
rect 530122 261080 530178 261089
rect 530122 261015 530178 261024
rect 530122 226264 530178 226273
rect 530044 226222 530122 226250
rect 530122 226199 530178 226208
rect 529938 209264 529994 209273
rect 529938 209199 529994 209208
rect 475384 198008 475436 198014
rect 475384 197950 475436 197956
rect 460388 46844 460440 46850
rect 460388 46786 460440 46792
rect 460204 42220 460256 42226
rect 460204 42162 460256 42168
rect 475396 41410 475424 197950
rect 528560 182844 528612 182850
rect 528560 182786 528612 182792
rect 524420 171828 524472 171834
rect 524420 171770 524472 171776
rect 489920 162376 489972 162382
rect 489920 162318 489972 162324
rect 485780 162308 485832 162314
rect 485780 162250 485832 162256
rect 481640 162240 481692 162246
rect 481640 162182 481692 162188
rect 481652 151814 481680 162182
rect 481652 151786 481864 151814
rect 481836 139890 481864 151786
rect 485792 139890 485820 162250
rect 489932 139890 489960 162318
rect 521660 160744 521712 160750
rect 521660 160686 521712 160692
rect 496820 160540 496872 160546
rect 496820 160482 496872 160488
rect 494060 160404 494112 160410
rect 494060 160346 494112 160352
rect 494072 139890 494100 160346
rect 496832 151814 496860 160482
rect 500960 160472 501012 160478
rect 500960 160414 501012 160420
rect 500972 151814 501000 160414
rect 505100 160336 505152 160342
rect 505100 160278 505152 160284
rect 505112 151814 505140 160278
rect 509240 160268 509292 160274
rect 509240 160210 509292 160216
rect 509252 151814 509280 160210
rect 513380 160200 513432 160206
rect 513380 160142 513432 160148
rect 513392 151814 513420 160142
rect 517520 160132 517572 160138
rect 517520 160074 517572 160080
rect 496832 151786 497688 151814
rect 500972 151786 501644 151814
rect 505112 151786 505600 151814
rect 509252 151786 509556 151814
rect 513392 151786 513512 151814
rect 497660 139890 497688 151786
rect 501616 139890 501644 151786
rect 505572 139890 505600 151786
rect 509528 139890 509556 151786
rect 513484 139890 513512 151786
rect 517532 139890 517560 160074
rect 521672 139890 521700 160686
rect 524432 151814 524460 171770
rect 528572 151814 528600 182786
rect 524432 151786 525380 151814
rect 528572 151786 529336 151814
rect 525352 139890 525380 151786
rect 529308 139890 529336 151786
rect 530596 140078 530624 319262
rect 531320 287700 531372 287706
rect 531320 287642 531372 287648
rect 531332 243681 531360 287642
rect 531318 243672 531374 243681
rect 531318 243607 531374 243616
rect 533356 140146 533384 319466
rect 533436 300688 533488 300694
rect 533436 300630 533488 300636
rect 533448 167006 533476 300630
rect 533436 167000 533488 167006
rect 533436 166942 533488 166948
rect 533436 162172 533488 162178
rect 533436 162114 533488 162120
rect 533448 143546 533476 162114
rect 533436 143540 533488 143546
rect 533436 143482 533488 143488
rect 533988 143540 534040 143546
rect 533988 143482 534040 143488
rect 534000 142254 534028 143482
rect 533988 142248 534040 142254
rect 533988 142190 534040 142196
rect 533344 140140 533396 140146
rect 533344 140082 533396 140088
rect 530584 140072 530636 140078
rect 530584 140014 530636 140020
rect 534000 139890 534028 142190
rect 534736 140214 534764 319534
rect 538864 319456 538916 319462
rect 538864 319398 538916 319404
rect 536104 294500 536156 294506
rect 536104 294442 536156 294448
rect 536116 143546 536144 294442
rect 536104 143540 536156 143546
rect 536104 143482 536156 143488
rect 537300 143540 537352 143546
rect 537300 143482 537352 143488
rect 534724 140208 534776 140214
rect 534724 140150 534776 140156
rect 481836 139862 482264 139890
rect 485792 139862 486220 139890
rect 489932 139862 490176 139890
rect 494072 139862 494132 139890
rect 497660 139862 498088 139890
rect 501616 139862 502044 139890
rect 505572 139862 506000 139890
rect 509528 139862 509956 139890
rect 513484 139862 513912 139890
rect 517532 139862 517868 139890
rect 521672 139862 521824 139890
rect 525352 139862 525780 139890
rect 529308 139862 529736 139890
rect 533692 139862 534028 139890
rect 537312 139890 537340 143482
rect 537312 139862 537648 139890
rect 538876 138582 538904 319398
rect 580460 319190 580488 630799
rect 580552 599622 580580 643991
rect 580540 599616 580592 599622
rect 580540 599558 580592 599564
rect 580538 471472 580594 471481
rect 580538 471407 580594 471416
rect 580552 322862 580580 471407
rect 580630 431624 580686 431633
rect 580630 431559 580686 431568
rect 580540 322856 580592 322862
rect 580540 322798 580592 322804
rect 580644 321026 580672 431559
rect 580722 418296 580778 418305
rect 580722 418231 580778 418240
rect 580736 330546 580764 418231
rect 580814 351928 580870 351937
rect 580814 351863 580870 351872
rect 580724 330540 580776 330546
rect 580724 330482 580776 330488
rect 580632 321020 580684 321026
rect 580632 320962 580684 320968
rect 580828 320890 580856 351863
rect 580908 330540 580960 330546
rect 580908 330482 580960 330488
rect 580816 320884 580868 320890
rect 580816 320826 580868 320832
rect 580920 319258 580948 330482
rect 580908 319252 580960 319258
rect 580908 319194 580960 319200
rect 580448 319184 580500 319190
rect 580448 319126 580500 319132
rect 539600 318232 539652 318238
rect 539600 318174 539652 318180
rect 538956 309936 539008 309942
rect 538956 309878 539008 309884
rect 538864 138576 538916 138582
rect 538864 138518 538916 138524
rect 538968 138009 538996 309878
rect 539048 308508 539100 308514
rect 539048 308450 539100 308456
rect 539060 151814 539088 308450
rect 539060 151786 539364 151814
rect 538954 138000 539010 138009
rect 538954 137935 539010 137944
rect 539336 135697 539364 151786
rect 539322 135688 539378 135697
rect 539322 135623 539378 135632
rect 539612 82793 539640 318174
rect 569224 318096 569276 318102
rect 569224 318038 569276 318044
rect 539784 316940 539836 316946
rect 539784 316882 539836 316888
rect 539692 315376 539744 315382
rect 539692 315318 539744 315324
rect 539704 84969 539732 315318
rect 539796 113257 539824 316882
rect 542636 316872 542688 316878
rect 542636 316814 542688 316820
rect 539876 315444 539928 315450
rect 539876 315386 539928 315392
rect 539888 119649 539916 315386
rect 540980 314016 541032 314022
rect 540980 313958 541032 313964
rect 539968 285048 540020 285054
rect 539968 284990 540020 284996
rect 539874 119640 539930 119649
rect 539874 119575 539930 119584
rect 539782 113248 539838 113257
rect 539782 113183 539838 113192
rect 539980 99249 540008 284990
rect 540060 276684 540112 276690
rect 540060 276626 540112 276632
rect 540072 108769 540100 276626
rect 540244 271244 540296 271250
rect 540244 271186 540296 271192
rect 540152 271176 540204 271182
rect 540152 271118 540204 271124
rect 540058 108760 540114 108769
rect 540058 108695 540114 108704
rect 540164 104825 540192 271118
rect 540256 115025 540284 271186
rect 540336 142248 540388 142254
rect 540336 142190 540388 142196
rect 540242 115016 540298 115025
rect 540242 114951 540298 114960
rect 540150 104816 540206 104825
rect 540150 104751 540206 104760
rect 539966 99240 540022 99249
rect 539966 99175 540022 99184
rect 539690 84960 539746 84969
rect 539690 84895 539746 84904
rect 539598 82784 539654 82793
rect 539598 82719 539654 82728
rect 475384 41404 475436 41410
rect 475384 41346 475436 41352
rect 536840 41404 536892 41410
rect 536840 41346 536892 41352
rect 536852 41041 536880 41346
rect 536838 41032 536894 41041
rect 536838 40967 536894 40976
rect 540348 34241 540376 142190
rect 540992 86465 541020 313958
rect 542544 312588 542596 312594
rect 542544 312530 542596 312536
rect 541072 309800 541124 309806
rect 541072 309742 541124 309748
rect 541084 121145 541112 309742
rect 541164 286408 541216 286414
rect 541164 286350 541216 286356
rect 541070 121136 541126 121145
rect 541070 121071 541126 121080
rect 541176 110945 541204 286350
rect 542452 280832 542504 280838
rect 542452 280774 542504 280780
rect 541256 275324 541308 275330
rect 541256 275266 541308 275272
rect 541162 110936 541218 110945
rect 541162 110871 541218 110880
rect 541268 102785 541296 275266
rect 541348 273964 541400 273970
rect 541348 273906 541400 273912
rect 541360 106865 541388 273906
rect 541440 272536 541492 272542
rect 541440 272478 541492 272484
rect 541452 117065 541480 272478
rect 541438 117056 541494 117065
rect 541438 116991 541494 117000
rect 541346 106856 541402 106865
rect 541346 106791 541402 106800
rect 541254 102776 541310 102785
rect 541254 102711 541310 102720
rect 542464 92585 542492 280774
rect 542556 125225 542584 312530
rect 542648 129305 542676 316814
rect 547144 316736 547196 316742
rect 547144 316678 547196 316684
rect 543188 314084 543240 314090
rect 543188 314026 543240 314032
rect 542820 268456 542872 268462
rect 542820 268398 542872 268404
rect 542728 140140 542780 140146
rect 542728 140082 542780 140088
rect 542634 129296 542690 129305
rect 542634 129231 542690 129240
rect 542542 125216 542598 125225
rect 542542 125151 542598 125160
rect 542740 96665 542768 140082
rect 542726 96656 542782 96665
rect 542726 96591 542782 96600
rect 542832 94625 542860 268398
rect 542912 140208 542964 140214
rect 542912 140150 542964 140156
rect 542924 100745 542952 140150
rect 543096 140072 543148 140078
rect 543096 140014 543148 140020
rect 543004 138576 543056 138582
rect 543004 138518 543056 138524
rect 543016 123185 543044 138518
rect 543108 131345 543136 140014
rect 543200 133385 543228 314026
rect 544384 306196 544436 306202
rect 544384 306138 544436 306144
rect 543280 279472 543332 279478
rect 543280 279414 543332 279420
rect 543186 133376 543242 133385
rect 543186 133311 543242 133320
rect 543094 131336 543150 131345
rect 543094 131271 543150 131280
rect 543002 123176 543058 123185
rect 543002 123111 543058 123120
rect 542910 100736 542966 100745
rect 542910 100671 542966 100680
rect 542818 94616 542874 94625
rect 542818 94551 542874 94560
rect 542450 92576 542506 92585
rect 542450 92511 542506 92520
rect 543292 90545 543320 279414
rect 543740 269952 543792 269958
rect 543740 269894 543792 269900
rect 543278 90536 543334 90545
rect 543278 90471 543334 90480
rect 540978 86456 541034 86465
rect 540978 86391 541034 86400
rect 543752 51134 543780 269894
rect 544396 73166 544424 306138
rect 547156 193186 547184 316678
rect 551284 315308 551336 315314
rect 551284 315250 551336 315256
rect 548524 311160 548576 311166
rect 548524 311102 548576 311108
rect 547144 193180 547196 193186
rect 547144 193122 547196 193128
rect 544384 73160 544436 73166
rect 544384 73102 544436 73108
rect 548536 60722 548564 311102
rect 551296 153202 551324 315250
rect 566464 313948 566516 313954
rect 566464 313890 566516 313896
rect 562324 304496 562376 304502
rect 562324 304438 562376 304444
rect 555424 293276 555476 293282
rect 555424 293218 555476 293224
rect 551284 153196 551336 153202
rect 551284 153138 551336 153144
rect 555436 139398 555464 293218
rect 559656 291644 559708 291650
rect 559656 291586 559708 291592
rect 558184 290488 558236 290494
rect 558184 290430 558236 290436
rect 555424 139392 555476 139398
rect 555424 139334 555476 139340
rect 558196 100706 558224 290430
rect 559564 284980 559616 284986
rect 559564 284922 559616 284928
rect 559576 179382 559604 284922
rect 559668 233238 559696 291586
rect 559656 233232 559708 233238
rect 559656 233174 559708 233180
rect 559564 179376 559616 179382
rect 559564 179318 559616 179324
rect 558184 100700 558236 100706
rect 558184 100642 558236 100648
rect 548524 60716 548576 60722
rect 548524 60658 548576 60664
rect 540612 51128 540664 51134
rect 540612 51070 540664 51076
rect 543740 51128 543792 51134
rect 543740 51070 543792 51076
rect 540624 48929 540652 51070
rect 540610 48920 540666 48929
rect 540610 48855 540666 48864
rect 540334 34232 540390 34241
rect 540334 34167 540390 34176
rect 562336 6866 562364 304438
rect 566476 46918 566504 313890
rect 566464 46912 566516 46918
rect 566464 46854 566516 46860
rect 569236 33114 569264 318038
rect 580172 313268 580224 313274
rect 580172 313210 580224 313216
rect 580184 312089 580212 313210
rect 580170 312080 580226 312089
rect 580170 312015 580226 312024
rect 576124 307080 576176 307086
rect 576124 307022 576176 307028
rect 571984 303272 572036 303278
rect 571984 303214 572036 303220
rect 570604 295996 570656 296002
rect 570604 295938 570656 295944
rect 570616 113150 570644 295938
rect 570604 113144 570656 113150
rect 570604 113086 570656 113092
rect 571996 86970 572024 303214
rect 573364 301572 573416 301578
rect 573364 301514 573416 301520
rect 573376 126954 573404 301514
rect 574836 297220 574888 297226
rect 574836 297162 574888 297168
rect 574744 268388 574796 268394
rect 574744 268330 574796 268336
rect 573364 126948 573416 126954
rect 573364 126890 573416 126896
rect 571984 86964 572036 86970
rect 571984 86906 572036 86912
rect 569224 33108 569276 33114
rect 569224 33050 569276 33056
rect 574756 20670 574784 268330
rect 574848 245614 574876 297162
rect 574836 245608 574888 245614
rect 574836 245550 574888 245556
rect 576136 206990 576164 307022
rect 580172 299464 580224 299470
rect 580172 299406 580224 299412
rect 580184 298761 580212 299406
rect 580170 298752 580226 298761
rect 580170 298687 580226 298696
rect 580264 286340 580316 286346
rect 580264 286282 580316 286288
rect 579896 273216 579948 273222
rect 579896 273158 579948 273164
rect 579908 272241 579936 273158
rect 579894 272232 579950 272241
rect 579894 272167 579950 272176
rect 580172 245608 580224 245614
rect 580170 245576 580172 245585
rect 580224 245576 580226 245585
rect 580170 245511 580226 245520
rect 580172 233232 580224 233238
rect 580172 233174 580224 233180
rect 580184 232393 580212 233174
rect 580170 232384 580226 232393
rect 580170 232319 580226 232328
rect 580276 219065 580304 286282
rect 580356 269884 580408 269890
rect 580356 269826 580408 269832
rect 580368 258913 580396 269826
rect 580354 258904 580410 258913
rect 580354 258839 580410 258848
rect 580262 219056 580318 219065
rect 580262 218991 580318 219000
rect 576124 206984 576176 206990
rect 576124 206926 576176 206932
rect 579804 206984 579856 206990
rect 579804 206926 579856 206932
rect 579816 205737 579844 206926
rect 579802 205728 579858 205737
rect 579802 205663 579858 205672
rect 580172 193180 580224 193186
rect 580172 193122 580224 193128
rect 580184 192545 580212 193122
rect 580170 192536 580226 192545
rect 580170 192471 580226 192480
rect 580172 179376 580224 179382
rect 580172 179318 580224 179324
rect 580184 179217 580212 179318
rect 580170 179208 580226 179217
rect 580170 179143 580226 179152
rect 580172 167000 580224 167006
rect 580172 166942 580224 166948
rect 580184 165889 580212 166942
rect 580170 165880 580226 165889
rect 580170 165815 580226 165824
rect 580172 153196 580224 153202
rect 580172 153138 580224 153144
rect 580184 152697 580212 153138
rect 580170 152688 580226 152697
rect 580170 152623 580226 152632
rect 580172 139392 580224 139398
rect 580170 139360 580172 139369
rect 580224 139360 580226 139369
rect 580170 139295 580226 139304
rect 580172 126948 580224 126954
rect 580172 126890 580224 126896
rect 580184 126041 580212 126890
rect 580170 126032 580226 126041
rect 580170 125967 580226 125976
rect 579804 113144 579856 113150
rect 579804 113086 579856 113092
rect 579816 112849 579844 113086
rect 579802 112840 579858 112849
rect 579802 112775 579858 112784
rect 580172 100700 580224 100706
rect 580172 100642 580224 100648
rect 580184 99521 580212 100642
rect 580170 99512 580226 99521
rect 580170 99447 580226 99456
rect 580172 86964 580224 86970
rect 580172 86906 580224 86912
rect 580184 86193 580212 86906
rect 580170 86184 580226 86193
rect 580170 86119 580226 86128
rect 580172 73160 580224 73166
rect 580172 73102 580224 73108
rect 580184 73001 580212 73102
rect 580170 72992 580226 73001
rect 580170 72927 580226 72936
rect 580172 60716 580224 60722
rect 580172 60658 580224 60664
rect 580184 59673 580212 60658
rect 580170 59664 580226 59673
rect 580170 59599 580226 59608
rect 580172 46912 580224 46918
rect 580172 46854 580224 46860
rect 580184 46345 580212 46854
rect 580170 46336 580226 46345
rect 580170 46271 580226 46280
rect 580170 33144 580226 33153
rect 580170 33079 580172 33088
rect 580224 33079 580226 33088
rect 580172 33050 580224 33056
rect 574744 20664 574796 20670
rect 574744 20606 574796 20612
rect 579988 20664 580040 20670
rect 579988 20606 580040 20612
rect 580000 19825 580028 20606
rect 579986 19816 580042 19825
rect 579986 19751 580042 19760
rect 562324 6860 562376 6866
rect 562324 6802 562376 6808
rect 580172 6860 580224 6866
rect 580172 6802 580224 6808
rect 580184 6633 580212 6802
rect 580170 6624 580226 6633
rect 580170 6559 580226 6568
rect 456064 3528 456116 3534
rect 456064 3470 456116 3476
rect 406382 3431 406438 3440
rect 450728 3460 450780 3466
rect 450728 3402 450780 3408
rect 395344 2100 395396 2106
rect 395344 2042 395396 2048
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9926 -960 10038 480
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14710 -960 14822 480
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 18206 -960 18318 480
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22990 -960 23102 480
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26486 -960 26598 480
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 31270 -960 31382 480
rect 32374 -960 32486 480
rect 33570 -960 33682 480
rect 34766 -960 34878 480
rect 35962 -960 36074 480
rect 37158 -960 37270 480
rect 38354 -960 38466 480
rect 39550 -960 39662 480
rect 40654 -960 40766 480
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45438 -960 45550 480
rect 46634 -960 46746 480
rect 47830 -960 47942 480
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53718 -960 53830 480
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 57214 -960 57326 480
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61998 -960 62110 480
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67886 -960 67998 480
rect 69082 -960 69194 480
rect 70278 -960 70390 480
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 76166 -960 76278 480
rect 77362 -960 77474 480
rect 78558 -960 78670 480
rect 79662 -960 79774 480
rect 80858 -960 80970 480
rect 82054 -960 82166 480
rect 83250 -960 83362 480
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 86838 -960 86950 480
rect 87942 -960 88054 480
rect 89138 -960 89250 480
rect 90334 -960 90446 480
rect 91530 -960 91642 480
rect 92726 -960 92838 480
rect 93922 -960 94034 480
rect 95118 -960 95230 480
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98614 -960 98726 480
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104502 -960 104614 480
rect 105698 -960 105810 480
rect 106894 -960 107006 480
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112782 -960 112894 480
rect 113978 -960 114090 480
rect 115174 -960 115286 480
rect 116370 -960 116482 480
rect 117566 -960 117678 480
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 123454 -960 123566 480
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 148294 -960 148406 480
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 174238 -960 174350 480
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 179022 -960 179134 480
rect 180218 -960 180330 480
rect 181414 -960 181526 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 199078 -960 199190 480
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220422 -960 220534 480
rect 221526 -960 221638 480
rect 222722 -960 222834 480
rect 223918 -960 224030 480
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236982 -960 237094 480
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248758 -960 248870 480
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273598 -960 273710 480
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 279486 -960 279598 480
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293654 -960 293766 480
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 304326 -960 304438 480
rect 305522 -960 305634 480
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318494 -960 318606 480
rect 319690 -960 319802 480
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 354006 -960 354118 480
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370566 -960 370678 480
rect 371670 -960 371782 480
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 378846 -960 378958 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 387126 -960 387238 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396510 -960 396622 480
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409574 -960 409686 480
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 413070 -960 413182 480
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417854 -960 417966 480
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 421350 -960 421462 480
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 427238 -960 427350 480
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435518 -960 435630 480
rect 436714 -960 436826 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 446190 -960 446302 480
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 460358 -960 460470 480
rect 461554 -960 461666 480
rect 462750 -960 462862 480
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 471030 -960 471142 480
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474526 -960 474638 480
rect 475722 -960 475834 480
rect 476918 -960 477030 480
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482806 -960 482918 480
rect 484002 -960 484114 480
rect 485198 -960 485310 480
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 491086 -960 491198 480
rect 492282 -960 492394 480
rect 493478 -960 493590 480
rect 494674 -960 494786 480
rect 495870 -960 495982 480
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499366 -960 499478 480
rect 500562 -960 500674 480
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 504150 -960 504262 480
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507646 -960 507758 480
rect 508842 -960 508954 480
rect 510038 -960 510150 480
rect 511234 -960 511346 480
rect 512430 -960 512542 480
rect 513534 -960 513646 480
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 518318 -960 518430 480
rect 519514 -960 519626 480
rect 520710 -960 520822 480
rect 521814 -960 521926 480
rect 523010 -960 523122 480
rect 524206 -960 524318 480
rect 525402 -960 525514 480
rect 526598 -960 526710 480
rect 527794 -960 527906 480
rect 528990 -960 529102 480
rect 530094 -960 530206 480
rect 531290 -960 531402 480
rect 532486 -960 532598 480
rect 533682 -960 533794 480
rect 534878 -960 534990 480
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538374 -960 538486 480
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 543158 -960 543270 480
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546654 -960 546766 480
rect 547850 -960 547962 480
rect 549046 -960 549158 480
rect 550242 -960 550354 480
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 557326 -960 557438 480
rect 558522 -960 558634 480
rect 559718 -960 559830 480
rect 560822 -960 560934 480
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564410 -960 564522 480
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 24306 686432 24362 686488
rect 300122 700304 300178 700360
rect 3146 658180 3148 658200
rect 3148 658180 3200 658200
rect 3200 658180 3202 658200
rect 3146 658144 3202 658180
rect 3238 579944 3294 580000
rect 3330 566888 3386 566944
rect 3606 632032 3662 632088
rect 3514 462576 3570 462632
rect 3422 449520 3478 449576
rect 4066 553832 4122 553888
rect 3974 527856 4030 527912
rect 3882 514800 3938 514856
rect 362222 678952 362278 679008
rect 361762 667956 361818 667992
rect 361762 667936 361764 667956
rect 361764 667936 361816 667956
rect 361816 667936 361818 667956
rect 361762 656940 361818 656976
rect 361762 656920 361764 656940
rect 361764 656920 361816 656940
rect 361816 656920 361818 656940
rect 361762 645924 361818 645960
rect 361762 645904 361764 645924
rect 361764 645904 361816 645924
rect 361816 645904 361818 645924
rect 361578 634888 361634 634944
rect 361578 623872 361634 623928
rect 361578 612876 361634 612912
rect 361578 612856 361580 612876
rect 361580 612856 361632 612876
rect 361632 612856 361634 612876
rect 361762 601840 361818 601896
rect 361578 590844 361634 590880
rect 361578 590824 361580 590844
rect 361580 590824 361632 590844
rect 361632 590824 361634 590844
rect 361762 579808 361818 579864
rect 361578 568812 361634 568848
rect 361578 568792 361580 568812
rect 361580 568792 361632 568812
rect 361632 568792 361634 568812
rect 361670 557776 361726 557832
rect 361762 546760 361818 546816
rect 361762 535744 361818 535800
rect 361762 524728 361818 524784
rect 3790 501744 3846 501800
rect 3698 475632 3754 475688
rect 3606 423544 3662 423600
rect 361762 513712 361818 513768
rect 361762 502696 361818 502752
rect 361762 491680 361818 491736
rect 361762 480664 361818 480720
rect 361762 469648 361818 469704
rect 361762 458632 361818 458688
rect 361762 447616 361818 447672
rect 361762 436600 361818 436656
rect 361762 425584 361818 425640
rect 361578 414568 361634 414624
rect 3974 410488 4030 410544
rect 361578 403552 361634 403608
rect 3790 397432 3846 397488
rect 3514 358400 3570 358456
rect 3422 345344 3478 345400
rect 3698 306176 3754 306232
rect 3606 293120 3662 293176
rect 3514 267144 3570 267200
rect 3422 254088 3478 254144
rect 3330 162832 3386 162888
rect 3238 149776 3294 149832
rect 3146 98640 3202 98696
rect 361578 392536 361634 392592
rect 361578 381520 361634 381576
rect 3882 371320 3938 371376
rect 3790 241032 3846 241088
rect 3606 71576 3662 71632
rect 3514 58520 3570 58576
rect 361578 370504 361634 370560
rect 362222 359488 362278 359544
rect 361762 348472 361818 348528
rect 361762 337456 361818 337512
rect 362222 326440 362278 326496
rect 3974 319232 4030 319288
rect 361762 315424 361818 315480
rect 3882 214920 3938 214976
rect 3974 201864 4030 201920
rect 4066 188808 4122 188864
rect 20902 77152 20958 77208
rect 21454 77152 21510 77208
rect 11702 48864 11758 48920
rect 18786 49272 18842 49328
rect 3514 45464 3570 45520
rect 7654 44784 7710 44840
rect 2870 32408 2926 32464
rect 3422 19352 3478 19408
rect 3422 6432 3478 6488
rect 2870 3576 2926 3632
rect 1674 3440 1730 3496
rect 570 3304 626 3360
rect 5262 3168 5318 3224
rect 9954 3984 10010 4040
rect 8758 3712 8814 3768
rect 13542 3848 13598 3904
rect 359554 46280 359610 46336
rect 361762 304408 361818 304464
rect 361762 293392 361818 293448
rect 361762 282376 361818 282432
rect 361762 271360 361818 271416
rect 361762 260344 361818 260400
rect 361762 249328 361818 249384
rect 361762 238312 361818 238368
rect 361762 227296 361818 227352
rect 361578 216316 361580 216336
rect 361580 216316 361632 216336
rect 361632 216316 361634 216336
rect 361578 216280 361634 216316
rect 361762 205264 361818 205320
rect 361670 194248 361726 194304
rect 361670 183232 361726 183288
rect 361670 172216 361726 172272
rect 361762 161200 361818 161256
rect 361762 150184 361818 150240
rect 361762 139168 361818 139224
rect 361578 128152 361634 128208
rect 361578 117136 361634 117192
rect 361578 106120 361634 106176
rect 361762 95140 361764 95160
rect 361764 95140 361816 95160
rect 361816 95140 361818 95160
rect 361762 95104 361818 95140
rect 361762 84124 361764 84144
rect 361764 84124 361816 84144
rect 361816 84124 361818 84144
rect 361762 84088 361818 84124
rect 361762 73108 361764 73128
rect 361764 73108 361816 73128
rect 361816 73108 361818 73128
rect 361762 73072 361818 73108
rect 361762 62076 361818 62112
rect 361762 62056 361764 62076
rect 361764 62056 361816 62076
rect 361816 62056 361818 62076
rect 361762 51040 361818 51096
rect 361486 46416 361542 46472
rect 368110 291760 368166 291816
rect 376022 3984 376078 4040
rect 378966 294480 379022 294536
rect 392582 300464 392638 300520
rect 387062 3848 387118 3904
rect 392766 300328 392822 300384
rect 392950 300056 393006 300112
rect 395342 300192 395398 300248
rect 392582 3712 392638 3768
rect 363602 3168 363658 3224
rect 395526 300600 395582 300656
rect 420366 335144 420422 335200
rect 427818 337048 427874 337104
rect 428094 334464 428150 334520
rect 420458 334328 420514 334384
rect 424138 334328 424194 334384
rect 401230 302776 401286 302832
rect 406382 305904 406438 305960
rect 406566 305632 406622 305688
rect 406750 305768 406806 305824
rect 406658 44784 406714 44840
rect 406566 3576 406622 3632
rect 422022 162696 422078 162752
rect 426346 162696 426402 162752
rect 428646 162696 428702 162752
rect 432050 310800 432106 310856
rect 432878 332832 432934 332888
rect 432786 329160 432842 329216
rect 432694 325488 432750 325544
rect 432878 321816 432934 321872
rect 432786 318144 432842 318200
rect 432694 314472 432750 314528
rect 433154 307128 433210 307184
rect 444194 421912 444250 421968
rect 445206 322632 445262 322688
rect 445574 682760 445630 682816
rect 445574 322768 445630 322824
rect 446310 322496 446366 322552
rect 446770 683304 446826 683360
rect 446954 683168 447010 683224
rect 447414 447244 447416 447264
rect 447416 447244 447468 447264
rect 447468 447244 447470 447264
rect 447414 447208 447470 447244
rect 447138 383596 447140 383616
rect 447140 383596 447192 383616
rect 447192 383596 447194 383616
rect 447138 383560 447194 383596
rect 447230 382880 447286 382936
rect 447138 382200 447194 382256
rect 447230 381520 447286 381576
rect 447230 380840 447286 380896
rect 447138 380160 447194 380216
rect 447414 379480 447470 379536
rect 447138 378800 447194 378856
rect 447322 378120 447378 378176
rect 447138 377440 447194 377496
rect 447230 376760 447286 376816
rect 447138 376080 447194 376136
rect 447230 375400 447286 375456
rect 447138 374720 447194 374776
rect 447230 374040 447286 374096
rect 447138 373360 447194 373416
rect 447230 372680 447286 372736
rect 447138 372000 447194 372056
rect 447230 371320 447286 371376
rect 447138 370640 447194 370696
rect 447230 369960 447286 370016
rect 447138 369280 447194 369336
rect 447230 368600 447286 368656
rect 447138 367920 447194 367976
rect 447230 367240 447286 367296
rect 447138 366560 447194 366616
rect 447230 365880 447286 365936
rect 447230 365200 447286 365256
rect 447138 364520 447194 364576
rect 447230 363840 447286 363896
rect 447138 363160 447194 363216
rect 447138 362480 447194 362536
rect 447230 361800 447286 361856
rect 447230 361120 447286 361176
rect 447138 360440 447194 360496
rect 447138 359760 447194 359816
rect 447230 359080 447286 359136
rect 447782 422320 447838 422376
rect 447506 355000 447562 355056
rect 447782 354320 447838 354376
rect 447690 353640 447746 353696
rect 447874 352960 447930 353016
rect 447322 351600 447378 351656
rect 447138 350920 447194 350976
rect 447138 347520 447194 347576
rect 447138 342080 447194 342136
rect 447230 341400 447286 341456
rect 447230 340720 447286 340776
rect 447138 340040 447194 340096
rect 447230 339360 447286 339416
rect 447138 338680 447194 338736
rect 447138 337320 447194 337376
rect 447138 335960 447194 336016
rect 447230 335280 447286 335336
rect 447138 334600 447194 334656
rect 447230 333920 447286 333976
rect 447138 333240 447194 333296
rect 447138 329860 447194 329896
rect 447138 329840 447140 329860
rect 447140 329840 447192 329860
rect 447192 329840 447194 329860
rect 446770 319640 446826 319696
rect 447506 338000 447562 338056
rect 447414 336640 447470 336696
rect 447874 345480 447930 345536
rect 447782 331200 447838 331256
rect 448058 352280 448114 352336
rect 448150 348880 448206 348936
rect 448242 346840 448298 346896
rect 449070 386960 449126 387016
rect 448978 358400 449034 358456
rect 449070 357040 449126 357096
rect 448426 355680 448482 355736
rect 448426 344800 448482 344856
rect 448426 343440 448482 343496
rect 448058 332560 448114 332616
rect 447966 330540 448022 330576
rect 447966 330520 447968 330540
rect 447968 330520 448020 330540
rect 448020 330520 448022 330540
rect 448242 331880 448298 331936
rect 448334 331200 448390 331256
rect 449162 321408 449218 321464
rect 543462 700304 543518 700360
rect 527178 699760 527234 699816
rect 559654 699760 559710 699816
rect 580262 697176 580318 697232
rect 579618 683848 579674 683904
rect 462318 670520 462374 670576
rect 457902 667936 457958 667992
rect 457718 657464 457774 657520
rect 457626 650120 457682 650176
rect 457534 645904 457590 645960
rect 457442 643184 457498 643240
rect 457350 640328 457406 640384
rect 457258 635432 457314 635488
rect 449714 503444 449770 503500
rect 449438 348200 449494 348256
rect 449622 357720 449678 357776
rect 449714 356360 449770 356416
rect 449714 350240 449770 350296
rect 450450 516840 450506 516896
rect 450450 514664 450506 514720
rect 457810 652840 457866 652896
rect 458086 662496 458142 662552
rect 457994 659912 458050 659968
rect 459098 637880 459154 637936
rect 459006 633392 459062 633448
rect 458822 630672 458878 630728
rect 458638 611360 458694 611416
rect 458914 621016 458970 621072
rect 458914 599528 458970 599584
rect 459374 628088 459430 628144
rect 459282 625776 459338 625832
rect 459190 623872 459246 623928
rect 459098 542952 459154 543008
rect 460202 618296 460258 618352
rect 459466 615984 459522 616040
rect 460110 613808 460166 613864
rect 460018 608640 460074 608696
rect 459926 606328 459982 606384
rect 459466 603608 459522 603664
rect 460110 601976 460166 602032
rect 458822 518200 458878 518256
rect 450542 512352 450598 512408
rect 450358 510176 450414 510232
rect 449990 507592 450046 507648
rect 449806 349560 449862 349616
rect 449714 344120 449770 344176
rect 449530 342760 449586 342816
rect 449346 319504 449402 319560
rect 450082 505416 450138 505472
rect 450174 503240 450230 503296
rect 450266 337728 450322 337784
rect 450266 337048 450322 337104
rect 449990 334056 450046 334112
rect 449898 328888 449954 328944
rect 449990 326576 450046 326632
rect 450266 327936 450322 327992
rect 450634 505416 450690 505472
rect 450542 337728 450598 337784
rect 463054 517520 463110 517576
rect 463146 501064 463202 501120
rect 482742 517520 482798 517576
rect 492126 512420 492182 512476
rect 473726 462848 473782 462904
rect 489182 496848 489238 496904
rect 476118 428440 476174 428496
rect 472162 389000 472218 389056
rect 474370 389000 474426 389056
rect 472898 388864 472954 388920
rect 479522 389000 479578 389056
rect 494150 508816 494206 508872
rect 500958 516840 501014 516896
rect 502246 516840 502302 516896
rect 494334 515888 494390 515944
rect 510618 518064 510674 518120
rect 507122 516704 507178 516760
rect 494242 505688 494298 505744
rect 495070 505724 495072 505744
rect 495072 505724 495124 505744
rect 495124 505724 495126 505744
rect 495070 505688 495126 505724
rect 494702 501200 494758 501256
rect 493322 392536 493378 392592
rect 509330 375536 509386 375592
rect 450542 334192 450598 334248
rect 450450 328616 450506 328672
rect 450542 327256 450598 327312
rect 509514 366968 509570 367024
rect 509422 357584 509478 357640
rect 450450 325488 450506 325544
rect 450358 324808 450414 324864
rect 450082 324536 450138 324592
rect 450634 324128 450690 324184
rect 450542 317056 450598 317112
rect 509330 322904 509386 322960
rect 468758 322360 468814 322416
rect 450910 316920 450966 316976
rect 450726 316648 450782 316704
rect 406382 3440 406438 3496
rect 451094 316784 451150 316840
rect 451922 156848 451978 156904
rect 452014 151408 452070 151464
rect 451554 150048 451610 150104
rect 451738 148688 451794 148744
rect 451738 147364 451740 147384
rect 451740 147364 451792 147384
rect 451792 147364 451794 147384
rect 451738 147328 451794 147364
rect 451554 139168 451610 139224
rect 452566 158244 452568 158264
rect 452568 158244 452620 158264
rect 452620 158244 452622 158264
rect 452566 158208 452622 158244
rect 452566 155488 452622 155544
rect 452382 154128 452438 154184
rect 452290 152768 452346 152824
rect 452566 145968 452622 146024
rect 452566 144644 452568 144664
rect 452568 144644 452620 144664
rect 452620 144644 452622 144664
rect 452566 144608 452622 144644
rect 452566 143284 452568 143304
rect 452568 143284 452620 143304
rect 452620 143284 452622 143304
rect 452566 143248 452622 143284
rect 452566 141924 452568 141944
rect 452568 141924 452620 141944
rect 452620 141924 452622 141944
rect 452566 141888 452622 141924
rect 452566 140528 452622 140584
rect 452566 137844 452568 137864
rect 452568 137844 452620 137864
rect 452620 137844 452622 137864
rect 452566 137808 452622 137844
rect 452566 136484 452568 136504
rect 452568 136484 452620 136504
rect 452620 136484 452622 136504
rect 452566 136448 452622 136484
rect 452566 135124 452568 135144
rect 452568 135124 452620 135144
rect 452620 135124 452622 135144
rect 452566 135088 452622 135124
rect 452566 133764 452568 133784
rect 452568 133764 452620 133784
rect 452620 133764 452622 133784
rect 452566 133728 452622 133764
rect 452474 132404 452476 132424
rect 452476 132404 452528 132424
rect 452528 132404 452530 132424
rect 452474 132368 452530 132404
rect 452566 131044 452568 131064
rect 452568 131044 452620 131064
rect 452620 131044 452622 131064
rect 452566 131008 452622 131044
rect 452198 129648 452254 129704
rect 452106 128288 452162 128344
rect 452566 126948 452622 126984
rect 452566 126928 452568 126948
rect 452568 126928 452620 126948
rect 452620 126928 452622 126948
rect 451922 125568 451978 125624
rect 451922 124208 451978 124264
rect 451922 122848 451978 122904
rect 451738 121488 451794 121544
rect 454682 317192 454738 317248
rect 456154 319368 456210 319424
rect 456798 262656 456854 262712
rect 460018 320592 460074 320648
rect 457810 248784 457866 248840
rect 457718 207168 457774 207224
rect 457994 234948 457996 234968
rect 457996 234948 458048 234968
rect 458048 234948 458050 234968
rect 457994 234912 458050 234948
rect 457994 221040 458050 221096
rect 458086 207168 458142 207224
rect 459006 46824 459062 46880
rect 459190 46688 459246 46744
rect 458822 46552 458878 46608
rect 460294 320048 460350 320104
rect 461122 321272 461178 321328
rect 462226 321408 462282 321464
rect 462502 321136 462558 321192
rect 461950 321000 462006 321056
rect 470138 322360 470194 322416
rect 470506 321272 470562 321328
rect 482650 322632 482706 322688
rect 483754 322632 483810 322688
rect 507122 322632 507178 322688
rect 473542 322496 473598 322552
rect 472714 319912 472770 319968
rect 474094 319776 474150 319832
rect 472990 319640 473046 319696
rect 482926 319504 482982 319560
rect 486238 319368 486294 319424
rect 497186 311072 497242 311128
rect 502246 278024 502302 278080
rect 507490 321408 507546 321464
rect 509330 320728 509386 320784
rect 509790 351736 509846 351792
rect 509606 343984 509662 344040
rect 509698 328344 509754 328400
rect 510066 330248 510122 330304
rect 509882 327664 509938 327720
rect 509974 326032 510030 326088
rect 509882 302776 509938 302832
rect 510710 373768 510766 373824
rect 510158 317192 510214 317248
rect 510802 359080 510858 359136
rect 510986 355816 511042 355872
rect 510894 353096 510950 353152
rect 511078 347656 511134 347712
rect 511170 346024 511226 346080
rect 512274 378120 512330 378176
rect 512458 382492 512514 382528
rect 512458 382472 512460 382492
rect 512460 382472 512512 382492
rect 512512 382472 512514 382492
rect 512458 381384 512514 381440
rect 513194 384648 513250 384704
rect 513286 384104 513342 384160
rect 512642 383560 512698 383616
rect 513010 383016 513066 383072
rect 513010 381928 513066 381984
rect 512550 379772 512606 379808
rect 512550 379752 512552 379772
rect 512552 379752 512604 379772
rect 512604 379752 512606 379772
rect 512826 379208 512882 379264
rect 512458 377576 512514 377632
rect 512366 376488 512422 376544
rect 513194 380840 513250 380896
rect 513286 380296 513342 380352
rect 513286 378664 513342 378720
rect 513194 377032 513250 377088
rect 512090 375944 512146 376000
rect 511998 374856 512054 374912
rect 513286 374312 513342 374368
rect 512642 373224 512698 373280
rect 513286 372700 513342 372736
rect 513286 372680 513288 372700
rect 513288 372680 513340 372700
rect 513340 372680 513342 372700
rect 511998 372136 512054 372192
rect 511998 371592 512054 371648
rect 512090 371048 512146 371104
rect 513286 370504 513342 370560
rect 513286 369960 513342 370016
rect 512090 369416 512146 369472
rect 511998 365628 512054 365664
rect 511998 365608 512000 365628
rect 512000 365608 512052 365628
rect 512052 365608 512054 365628
rect 511998 363976 512054 364032
rect 511998 362364 512054 362400
rect 511998 362344 512000 362364
rect 512000 362344 512052 362364
rect 512052 362344 512054 362364
rect 511998 360712 512054 360768
rect 512274 368872 512330 368928
rect 512182 368328 512238 368384
rect 512090 354204 512146 354240
rect 512090 354184 512092 354204
rect 512092 354184 512144 354204
rect 512144 354184 512146 354204
rect 512090 349308 512146 349344
rect 512090 349288 512092 349308
rect 512092 349288 512144 349308
rect 512144 349288 512146 349308
rect 512090 347112 512146 347168
rect 512090 344936 512146 344992
rect 513286 367784 513342 367840
rect 513286 366696 513342 366752
rect 513378 366152 513434 366208
rect 512826 365064 512882 365120
rect 513286 364520 513342 364576
rect 512274 363432 512330 363488
rect 513010 362888 513066 362944
rect 513286 361800 513342 361856
rect 512642 361256 512698 361312
rect 512366 360168 512422 360224
rect 513010 359624 513066 359680
rect 512550 358536 512606 358592
rect 512458 352552 512514 352608
rect 512458 350920 512514 350976
rect 512458 345480 512514 345536
rect 513286 356904 513342 356960
rect 512826 356380 512882 356416
rect 512826 356360 512828 356380
rect 512828 356360 512880 356380
rect 512880 356360 512882 356380
rect 513286 355272 513342 355328
rect 513286 354748 513342 354784
rect 513286 354728 513288 354748
rect 513288 354728 513340 354748
rect 513340 354728 513342 354748
rect 513286 353640 513342 353696
rect 512918 351464 512974 351520
rect 513286 350376 513342 350432
rect 512826 349832 512882 349888
rect 513286 348744 513342 348800
rect 513286 348220 513342 348256
rect 513286 348200 513288 348220
rect 513288 348200 513340 348220
rect 513340 348200 513342 348220
rect 512642 346588 512698 346624
rect 512642 346568 512644 346588
rect 512644 346568 512696 346588
rect 512696 346568 512698 346588
rect 512918 343848 512974 343904
rect 513194 343304 513250 343360
rect 513286 342252 513288 342272
rect 513288 342252 513340 342272
rect 513340 342252 513342 342272
rect 513286 342216 513342 342252
rect 512642 341672 512698 341728
rect 512826 341128 512882 341184
rect 513194 340584 513250 340640
rect 513286 340060 513342 340096
rect 513286 340040 513288 340060
rect 513288 340040 513340 340060
rect 513340 340040 513342 340060
rect 512734 338952 512790 339008
rect 512642 332968 512698 333024
rect 512642 332424 512698 332480
rect 513286 338408 513342 338464
rect 513102 337864 513158 337920
rect 513194 337320 513250 337376
rect 513286 336776 513342 336832
rect 512826 336232 512882 336288
rect 512550 317056 512606 317112
rect 512734 325352 512790 325408
rect 513286 335688 513342 335744
rect 513286 335144 513342 335200
rect 513286 334056 513342 334112
rect 513010 333512 513066 333568
rect 513562 357992 513618 358048
rect 513470 329160 513526 329216
rect 514114 316920 514170 316976
rect 515126 316784 515182 316840
rect 547878 516704 547934 516760
rect 519634 502288 519690 502344
rect 521750 462848 521806 462904
rect 557538 442856 557594 442912
rect 579618 617480 579674 617536
rect 580170 590960 580226 591016
rect 579986 577632 580042 577688
rect 580170 564304 580226 564360
rect 580170 537784 580226 537840
rect 580170 524476 580226 524512
rect 580170 524456 580172 524476
rect 580172 524456 580224 524476
rect 580224 524456 580226 524476
rect 580170 511264 580226 511320
rect 580170 484608 580226 484664
rect 580170 458088 580226 458144
rect 580170 404912 580226 404968
rect 580170 378392 580226 378448
rect 580170 365064 580226 365120
rect 580170 325216 580226 325272
rect 580354 670656 580410 670712
rect 580538 644000 580594 644056
rect 580446 630808 580502 630864
rect 530122 261024 530178 261080
rect 530122 226208 530178 226264
rect 529938 209208 529994 209264
rect 531318 243616 531374 243672
rect 580538 471416 580594 471472
rect 580630 431568 580686 431624
rect 580722 418240 580778 418296
rect 580814 351872 580870 351928
rect 538954 137944 539010 138000
rect 539322 135632 539378 135688
rect 539874 119584 539930 119640
rect 539782 113192 539838 113248
rect 540058 108704 540114 108760
rect 540242 114960 540298 115016
rect 540150 104760 540206 104816
rect 539966 99184 540022 99240
rect 539690 84904 539746 84960
rect 539598 82728 539654 82784
rect 536838 40976 536894 41032
rect 541070 121080 541126 121136
rect 541162 110880 541218 110936
rect 541438 117000 541494 117056
rect 541346 106800 541402 106856
rect 541254 102720 541310 102776
rect 542634 129240 542690 129296
rect 542542 125160 542598 125216
rect 542726 96600 542782 96656
rect 543186 133320 543242 133376
rect 543094 131280 543150 131336
rect 543002 123120 543058 123176
rect 542910 100680 542966 100736
rect 542818 94560 542874 94616
rect 542450 92520 542506 92576
rect 543278 90480 543334 90536
rect 540978 86400 541034 86456
rect 540610 48864 540666 48920
rect 540334 34176 540390 34232
rect 580170 312024 580226 312080
rect 580170 298696 580226 298752
rect 579894 272176 579950 272232
rect 580170 245556 580172 245576
rect 580172 245556 580224 245576
rect 580224 245556 580226 245576
rect 580170 245520 580226 245556
rect 580170 232328 580226 232384
rect 580354 258848 580410 258904
rect 580262 219000 580318 219056
rect 579802 205672 579858 205728
rect 580170 192480 580226 192536
rect 580170 179152 580226 179208
rect 580170 165824 580226 165880
rect 580170 152632 580226 152688
rect 580170 139340 580172 139360
rect 580172 139340 580224 139360
rect 580224 139340 580226 139360
rect 580170 139304 580226 139340
rect 580170 125976 580226 126032
rect 579802 112784 579858 112840
rect 580170 99456 580226 99512
rect 580170 86128 580226 86184
rect 580170 72936 580226 72992
rect 580170 59608 580226 59664
rect 580170 46280 580226 46336
rect 580170 33108 580226 33144
rect 580170 33088 580172 33108
rect 580172 33088 580224 33108
rect 580224 33088 580226 33108
rect 579986 19760 580042 19816
rect 580170 6568 580226 6624
<< metal3 >>
rect 300117 700362 300183 700365
rect 444230 700362 444236 700364
rect 300117 700360 444236 700362
rect 300117 700304 300122 700360
rect 300178 700304 444236 700360
rect 300117 700302 444236 700304
rect 300117 700299 300183 700302
rect 444230 700300 444236 700302
rect 444300 700300 444306 700364
rect 530526 700300 530532 700364
rect 530596 700362 530602 700364
rect 543457 700362 543523 700365
rect 530596 700360 543523 700362
rect 530596 700304 543462 700360
rect 543518 700304 543523 700360
rect 530596 700302 543523 700304
rect 530596 700300 530602 700302
rect 543457 700299 543523 700302
rect 527173 699820 527239 699821
rect 527173 699818 527220 699820
rect 527128 699816 527220 699818
rect 527128 699760 527178 699816
rect 527128 699758 527220 699760
rect 527173 699756 527220 699758
rect 527284 699756 527290 699820
rect 558126 699756 558132 699820
rect 558196 699818 558202 699820
rect 559649 699818 559715 699821
rect 558196 699816 559715 699818
rect 558196 699760 559654 699816
rect 559710 699760 559715 699816
rect 558196 699758 559715 699760
rect 558196 699756 558202 699758
rect 527173 699755 527239 699756
rect 559649 699755 559715 699758
rect -960 697220 480 697460
rect 580257 697234 580323 697237
rect 583520 697234 584960 697324
rect 580257 697232 584960 697234
rect 580257 697176 580262 697232
rect 580318 697176 584960 697232
rect 580257 697174 584960 697176
rect 580257 697171 580323 697174
rect 583520 697084 584960 697174
rect 24301 686490 24367 686493
rect 446254 686490 446260 686492
rect 24301 686488 446260 686490
rect 24301 686432 24306 686488
rect 24362 686432 446260 686488
rect 24301 686430 446260 686432
rect 24301 686427 24367 686430
rect 446254 686428 446260 686430
rect 446324 686428 446330 686492
rect -960 684314 480 684404
rect 447726 684314 447732 684316
rect -960 684254 447732 684314
rect -960 684164 480 684254
rect 447726 684252 447732 684254
rect 447796 684252 447802 684316
rect 579613 683906 579679 683909
rect 583520 683906 584960 683996
rect 579613 683904 584960 683906
rect 579613 683848 579618 683904
rect 579674 683848 584960 683904
rect 579613 683846 584960 683848
rect 579613 683843 579679 683846
rect 583520 683756 584960 683846
rect 3734 683300 3740 683364
rect 3804 683362 3810 683364
rect 446765 683362 446831 683365
rect 3804 683360 446831 683362
rect 3804 683304 446770 683360
rect 446826 683304 446831 683360
rect 3804 683302 446831 683304
rect 3804 683300 3810 683302
rect 446765 683299 446831 683302
rect 3550 683164 3556 683228
rect 3620 683226 3626 683228
rect 446949 683226 447015 683229
rect 3620 683224 447015 683226
rect 3620 683168 446954 683224
rect 447010 683168 447015 683224
rect 3620 683166 447015 683168
rect 3620 683164 3626 683166
rect 446949 683163 447015 683166
rect 3366 682756 3372 682820
rect 3436 682818 3442 682820
rect 445569 682818 445635 682821
rect 3436 682816 445635 682818
rect 3436 682760 445574 682816
rect 445630 682760 445635 682816
rect 3436 682758 445635 682760
rect 3436 682756 3442 682758
rect 445569 682755 445635 682758
rect 362217 679010 362283 679013
rect 359812 679008 362283 679010
rect 359812 678952 362222 679008
rect 362278 678952 362283 679008
rect 359812 678950 362283 678952
rect 362217 678947 362283 678950
rect -960 671258 480 671348
rect 3734 671258 3740 671260
rect -960 671198 3740 671258
rect -960 671108 480 671198
rect 3734 671196 3740 671198
rect 3804 671196 3810 671260
rect 580349 670714 580415 670717
rect 583520 670714 584960 670804
rect 580349 670712 584960 670714
rect 580349 670656 580354 670712
rect 580410 670656 584960 670712
rect 580349 670654 584960 670656
rect 580349 670651 580415 670654
rect 459502 670516 459508 670580
rect 459572 670578 459578 670580
rect 462313 670578 462379 670581
rect 459572 670576 462379 670578
rect 459572 670520 462318 670576
rect 462374 670520 462379 670576
rect 583520 670564 584960 670654
rect 459572 670518 462379 670520
rect 459572 670516 459578 670518
rect 462313 670515 462379 670518
rect 361757 667994 361823 667997
rect 359812 667992 361823 667994
rect 359812 667936 361762 667992
rect 361818 667936 361823 667992
rect 359812 667934 361823 667936
rect 361757 667931 361823 667934
rect 457897 667994 457963 667997
rect 457897 667992 460092 667994
rect 457897 667936 457902 667992
rect 457958 667936 460092 667992
rect 457897 667934 460092 667936
rect 457897 667931 457963 667934
rect 458030 665212 458036 665276
rect 458100 665274 458106 665276
rect 460062 665274 460122 665448
rect 458100 665214 460122 665274
rect 458100 665212 458106 665214
rect 458081 662554 458147 662557
rect 460062 662554 460122 663000
rect 458081 662552 460122 662554
rect 458081 662496 458086 662552
rect 458142 662496 460122 662552
rect 458081 662494 460122 662496
rect 458081 662491 458147 662494
rect 457989 659970 458055 659973
rect 460062 659970 460122 660552
rect 457989 659968 460122 659970
rect 457989 659912 457994 659968
rect 458050 659912 460122 659968
rect 457989 659910 460122 659912
rect 457989 659907 458055 659910
rect -960 658202 480 658292
rect 3141 658202 3207 658205
rect -960 658200 3207 658202
rect -960 658144 3146 658200
rect 3202 658144 3207 658200
rect -960 658142 3207 658144
rect -960 658052 480 658142
rect 3141 658139 3207 658142
rect 457713 657522 457779 657525
rect 460062 657522 460122 658104
rect 457713 657520 460122 657522
rect 457713 657464 457718 657520
rect 457774 657464 460122 657520
rect 457713 657462 460122 657464
rect 457713 657459 457779 657462
rect 583520 657236 584960 657476
rect 361757 656978 361823 656981
rect 359812 656976 361823 656978
rect 359812 656920 361762 656976
rect 361818 656920 361823 656976
rect 359812 656918 361823 656920
rect 361757 656915 361823 656918
rect 459134 655692 459140 655756
rect 459204 655754 459210 655756
rect 459204 655694 460092 655754
rect 459204 655692 459210 655694
rect 457805 652898 457871 652901
rect 460062 652898 460122 653208
rect 457805 652896 460122 652898
rect 457805 652840 457810 652896
rect 457866 652840 460122 652896
rect 457805 652838 460122 652840
rect 457805 652835 457871 652838
rect 457621 650178 457687 650181
rect 460062 650178 460122 650760
rect 457621 650176 460122 650178
rect 457621 650120 457626 650176
rect 457682 650120 460122 650176
rect 457621 650118 460122 650120
rect 457621 650115 457687 650118
rect 458950 647668 458956 647732
rect 459020 647730 459026 647732
rect 460062 647730 460122 648312
rect 459020 647670 460122 647730
rect 459020 647668 459026 647670
rect 361757 645962 361823 645965
rect 359812 645960 361823 645962
rect 359812 645904 361762 645960
rect 361818 645904 361823 645960
rect 359812 645902 361823 645904
rect 361757 645899 361823 645902
rect 457529 645962 457595 645965
rect 457529 645960 460092 645962
rect 457529 645904 457534 645960
rect 457590 645904 460092 645960
rect 457529 645902 460092 645904
rect 457529 645899 457595 645902
rect -960 644996 480 645236
rect 580533 644058 580599 644061
rect 583520 644058 584960 644148
rect 580533 644056 584960 644058
rect 580533 644000 580538 644056
rect 580594 644000 584960 644056
rect 580533 643998 584960 644000
rect 580533 643995 580599 643998
rect 583520 643908 584960 643998
rect 457437 643242 457503 643245
rect 460062 643242 460122 643416
rect 457437 643240 460122 643242
rect 457437 643184 457442 643240
rect 457498 643184 460122 643240
rect 457437 643182 460122 643184
rect 457437 643179 457503 643182
rect 457345 640386 457411 640389
rect 460062 640386 460122 640968
rect 457345 640384 460122 640386
rect 457345 640328 457350 640384
rect 457406 640328 460122 640384
rect 457345 640326 460122 640328
rect 457345 640323 457411 640326
rect 459093 637938 459159 637941
rect 460062 637938 460122 638520
rect 459093 637936 460122 637938
rect 459093 637880 459098 637936
rect 459154 637880 460122 637936
rect 459093 637878 460122 637880
rect 459093 637875 459159 637878
rect 457253 635490 457319 635493
rect 460062 635490 460122 636072
rect 457253 635488 460122 635490
rect 457253 635432 457258 635488
rect 457314 635432 460122 635488
rect 457253 635430 460122 635432
rect 457253 635427 457319 635430
rect 361573 634946 361639 634949
rect 359812 634944 361639 634946
rect 359812 634888 361578 634944
rect 361634 634888 361639 634944
rect 359812 634886 361639 634888
rect 361573 634883 361639 634886
rect 459001 633450 459067 633453
rect 460062 633450 460122 633624
rect 459001 633448 460122 633450
rect 459001 633392 459006 633448
rect 459062 633392 460122 633448
rect 459001 633390 460122 633392
rect 459001 633387 459067 633390
rect -960 632090 480 632180
rect 3601 632090 3667 632093
rect -960 632088 3667 632090
rect -960 632032 3606 632088
rect 3662 632032 3667 632088
rect -960 632030 3667 632032
rect -960 631940 480 632030
rect 3601 632027 3667 632030
rect 458817 630730 458883 630733
rect 460062 630730 460122 631176
rect 580441 630866 580507 630869
rect 583520 630866 584960 630956
rect 580441 630864 584960 630866
rect 580441 630808 580446 630864
rect 580502 630808 584960 630864
rect 580441 630806 584960 630808
rect 580441 630803 580507 630806
rect 458817 630728 460122 630730
rect 458817 630672 458822 630728
rect 458878 630672 460122 630728
rect 583520 630716 584960 630806
rect 458817 630670 460122 630672
rect 458817 630667 458883 630670
rect 459369 628146 459435 628149
rect 460062 628146 460122 628728
rect 459369 628144 460122 628146
rect 459369 628088 459374 628144
rect 459430 628088 460122 628144
rect 459369 628086 460122 628088
rect 459369 628083 459435 628086
rect 459277 625834 459343 625837
rect 460062 625834 460122 626280
rect 459277 625832 460122 625834
rect 459277 625776 459282 625832
rect 459338 625776 460122 625832
rect 459277 625774 460122 625776
rect 459277 625771 459343 625774
rect 361573 623930 361639 623933
rect 359812 623928 361639 623930
rect 359812 623872 361578 623928
rect 361634 623872 361639 623928
rect 359812 623870 361639 623872
rect 361573 623867 361639 623870
rect 459185 623930 459251 623933
rect 459185 623928 460092 623930
rect 459185 623872 459190 623928
rect 459246 623872 460092 623928
rect 459185 623870 460092 623872
rect 459185 623867 459251 623870
rect 458909 621074 458975 621077
rect 460062 621074 460122 621384
rect 458909 621072 460122 621074
rect 458909 621016 458914 621072
rect 458970 621016 460122 621072
rect 458909 621014 460122 621016
rect 458909 621011 458975 621014
rect -960 619170 480 619260
rect 3550 619170 3556 619172
rect -960 619110 3556 619170
rect -960 619020 480 619110
rect 3550 619108 3556 619110
rect 3620 619108 3626 619172
rect 460062 618354 460122 618936
rect 460197 618354 460263 618357
rect 460062 618352 460263 618354
rect 460062 618296 460202 618352
rect 460258 618296 460263 618352
rect 460062 618294 460263 618296
rect 460197 618291 460263 618294
rect 579613 617538 579679 617541
rect 583520 617538 584960 617628
rect 579613 617536 584960 617538
rect 579613 617480 579618 617536
rect 579674 617480 584960 617536
rect 579613 617478 584960 617480
rect 579613 617475 579679 617478
rect 583520 617388 584960 617478
rect 459461 616042 459527 616045
rect 460062 616042 460122 616488
rect 459461 616040 460122 616042
rect 459461 615984 459466 616040
rect 459522 615984 460122 616040
rect 459461 615982 460122 615984
rect 459461 615979 459527 615982
rect 460062 613869 460122 614040
rect 460062 613864 460171 613869
rect 460062 613808 460110 613864
rect 460166 613808 460171 613864
rect 460062 613806 460171 613808
rect 460105 613803 460171 613806
rect 361573 612914 361639 612917
rect 359812 612912 361639 612914
rect 359812 612856 361578 612912
rect 361634 612856 361639 612912
rect 359812 612854 361639 612856
rect 361573 612851 361639 612854
rect 458633 611418 458699 611421
rect 460062 611418 460122 611592
rect 458633 611416 460122 611418
rect 458633 611360 458638 611416
rect 458694 611360 460122 611416
rect 458633 611358 460122 611360
rect 458633 611355 458699 611358
rect 460062 608701 460122 609144
rect 460013 608696 460122 608701
rect 460013 608640 460018 608696
rect 460074 608640 460122 608696
rect 460013 608638 460122 608640
rect 460013 608635 460079 608638
rect 459921 606386 459987 606389
rect 460062 606386 460122 606696
rect 459921 606384 460122 606386
rect 459921 606328 459926 606384
rect 459982 606328 460122 606384
rect 459921 606326 460122 606328
rect 459921 606323 459987 606326
rect -960 606114 480 606204
rect 3366 606114 3372 606116
rect -960 606054 3372 606114
rect -960 605964 480 606054
rect 3366 606052 3372 606054
rect 3436 606052 3442 606116
rect 459461 603666 459527 603669
rect 460062 603666 460122 604248
rect 583520 604060 584960 604300
rect 459461 603664 460122 603666
rect 459461 603608 459466 603664
rect 459522 603608 460122 603664
rect 459461 603606 460122 603608
rect 459461 603603 459527 603606
rect 460105 602034 460171 602037
rect 460062 602032 460171 602034
rect 460062 601976 460110 602032
rect 460166 601976 460171 602032
rect 460062 601971 460171 601976
rect 361757 601898 361823 601901
rect 359812 601896 361823 601898
rect 359812 601840 361762 601896
rect 361818 601840 361823 601896
rect 460062 601868 460122 601971
rect 359812 601838 361823 601840
rect 361757 601835 361823 601838
rect 458909 599586 458975 599589
rect 472014 599586 472020 599588
rect 458909 599584 472020 599586
rect 458909 599528 458914 599584
rect 458970 599528 472020 599584
rect 458909 599526 472020 599528
rect 458909 599523 458975 599526
rect 472014 599524 472020 599526
rect 472084 599524 472090 599588
rect 459134 596804 459140 596868
rect 459204 596866 459210 596868
rect 478822 596866 478828 596868
rect 459204 596806 478828 596866
rect 459204 596804 459210 596806
rect 478822 596804 478828 596806
rect 478892 596804 478898 596868
rect -960 592908 480 593148
rect 580165 591018 580231 591021
rect 583520 591018 584960 591108
rect 580165 591016 584960 591018
rect 580165 590960 580170 591016
rect 580226 590960 584960 591016
rect 580165 590958 584960 590960
rect 580165 590955 580231 590958
rect 361573 590882 361639 590885
rect 359812 590880 361639 590882
rect 359812 590824 361578 590880
rect 361634 590824 361639 590880
rect 583520 590868 584960 590958
rect 359812 590822 361639 590824
rect 361573 590819 361639 590822
rect -960 580002 480 580092
rect 3233 580002 3299 580005
rect -960 580000 3299 580002
rect -960 579944 3238 580000
rect 3294 579944 3299 580000
rect -960 579942 3299 579944
rect -960 579852 480 579942
rect 3233 579939 3299 579942
rect 361757 579866 361823 579869
rect 359812 579864 361823 579866
rect 359812 579808 361762 579864
rect 361818 579808 361823 579864
rect 359812 579806 361823 579808
rect 361757 579803 361823 579806
rect 579981 577690 580047 577693
rect 583520 577690 584960 577780
rect 579981 577688 584960 577690
rect 579981 577632 579986 577688
rect 580042 577632 584960 577688
rect 579981 577630 584960 577632
rect 579981 577627 580047 577630
rect 583520 577540 584960 577630
rect 361573 568850 361639 568853
rect 359812 568848 361639 568850
rect 359812 568792 361578 568848
rect 361634 568792 361639 568848
rect 359812 568790 361639 568792
rect 361573 568787 361639 568790
rect -960 566946 480 567036
rect 3325 566946 3391 566949
rect -960 566944 3391 566946
rect -960 566888 3330 566944
rect 3386 566888 3391 566944
rect -960 566886 3391 566888
rect -960 566796 480 566886
rect 3325 566883 3391 566886
rect 580165 564362 580231 564365
rect 583520 564362 584960 564452
rect 580165 564360 584960 564362
rect 580165 564304 580170 564360
rect 580226 564304 584960 564360
rect 580165 564302 584960 564304
rect 580165 564299 580231 564302
rect 583520 564212 584960 564302
rect 361665 557834 361731 557837
rect 359812 557832 361731 557834
rect 359812 557776 361670 557832
rect 361726 557776 361731 557832
rect 359812 557774 361731 557776
rect 361665 557771 361731 557774
rect -960 553890 480 553980
rect 4061 553890 4127 553893
rect -960 553888 4127 553890
rect -960 553832 4066 553888
rect 4122 553832 4127 553888
rect -960 553830 4127 553832
rect -960 553740 480 553830
rect 4061 553827 4127 553830
rect 583520 551020 584960 551260
rect 361757 546818 361823 546821
rect 359812 546816 361823 546818
rect 359812 546760 361762 546816
rect 361818 546760 361823 546816
rect 359812 546758 361823 546760
rect 361757 546755 361823 546758
rect 459093 543010 459159 543013
rect 474406 543010 474412 543012
rect 459093 543008 474412 543010
rect 459093 542952 459098 543008
rect 459154 542952 474412 543008
rect 459093 542950 474412 542952
rect 459093 542947 459159 542950
rect 474406 542948 474412 542950
rect 474476 542948 474482 543012
rect -960 540684 480 540924
rect 580165 537842 580231 537845
rect 583520 537842 584960 537932
rect 580165 537840 584960 537842
rect 580165 537784 580170 537840
rect 580226 537784 584960 537840
rect 580165 537782 584960 537784
rect 580165 537779 580231 537782
rect 583520 537692 584960 537782
rect 361757 535802 361823 535805
rect 359812 535800 361823 535802
rect 359812 535744 361762 535800
rect 361818 535744 361823 535800
rect 359812 535742 361823 535744
rect 361757 535739 361823 535742
rect -960 527914 480 528004
rect 3969 527914 4035 527917
rect -960 527912 4035 527914
rect -960 527856 3974 527912
rect 4030 527856 4035 527912
rect -960 527854 4035 527856
rect -960 527764 480 527854
rect 3969 527851 4035 527854
rect 361757 524786 361823 524789
rect 359812 524784 361823 524786
rect 359812 524728 361762 524784
rect 361818 524728 361823 524784
rect 359812 524726 361823 524728
rect 361757 524723 361823 524726
rect 580165 524514 580231 524517
rect 583520 524514 584960 524604
rect 580165 524512 584960 524514
rect 580165 524456 580170 524512
rect 580226 524456 584960 524512
rect 580165 524454 584960 524456
rect 580165 524451 580231 524454
rect 583520 524364 584960 524454
rect 458817 518258 458883 518261
rect 472198 518258 472204 518260
rect 458817 518256 472204 518258
rect 458817 518200 458822 518256
rect 458878 518200 472204 518256
rect 458817 518198 472204 518200
rect 458817 518195 458883 518198
rect 472198 518196 472204 518198
rect 472268 518196 472274 518260
rect 459502 518060 459508 518124
rect 459572 518122 459578 518124
rect 510613 518122 510679 518125
rect 459572 518120 510679 518122
rect 459572 518064 510618 518120
rect 510674 518064 510679 518120
rect 459572 518062 510679 518064
rect 459572 518060 459578 518062
rect 510613 518059 510679 518062
rect 458030 517516 458036 517580
rect 458100 517578 458106 517580
rect 463049 517578 463115 517581
rect 482737 517580 482803 517581
rect 458100 517576 463115 517578
rect 458100 517520 463054 517576
rect 463110 517520 463115 517576
rect 458100 517518 463115 517520
rect 458100 517516 458106 517518
rect 463049 517515 463115 517518
rect 482686 517516 482692 517580
rect 482756 517578 482803 517580
rect 482756 517576 482848 517578
rect 482798 517520 482848 517576
rect 482756 517518 482848 517520
rect 482756 517516 482803 517518
rect 482737 517515 482803 517516
rect 450445 516898 450511 516901
rect 500953 516898 501019 516901
rect 502241 516898 502307 516901
rect 450445 516896 502307 516898
rect 450445 516840 450450 516896
rect 450506 516840 500958 516896
rect 501014 516840 502246 516896
rect 502302 516840 502307 516896
rect 450445 516838 502307 516840
rect 450445 516835 450511 516838
rect 500953 516835 501019 516838
rect 502241 516835 502307 516838
rect 451038 516762 451044 516764
rect 450678 516702 451044 516762
rect 450678 516528 450738 516702
rect 451038 516700 451044 516702
rect 451108 516762 451114 516764
rect 507117 516762 507183 516765
rect 547873 516762 547939 516765
rect 451108 516760 547939 516762
rect 451108 516704 507122 516760
rect 507178 516704 547878 516760
rect 547934 516704 547939 516760
rect 451108 516702 547939 516704
rect 451108 516700 451114 516702
rect 507117 516699 507183 516702
rect 547873 516699 547939 516702
rect 491894 515946 491954 515984
rect 494329 515946 494395 515949
rect 491894 515944 494395 515946
rect 491894 515888 494334 515944
rect 494390 515888 494395 515944
rect 491894 515886 494395 515888
rect 494329 515883 494395 515886
rect -960 514858 480 514948
rect 3877 514858 3943 514861
rect -960 514856 3943 514858
rect -960 514800 3882 514856
rect 3938 514800 3943 514856
rect -960 514798 3943 514800
rect -960 514708 480 514798
rect 3877 514795 3943 514798
rect 450445 514722 450511 514725
rect 450445 514720 450554 514722
rect 450445 514664 450450 514720
rect 450506 514664 450554 514720
rect 450445 514659 450554 514664
rect 450494 514384 450554 514659
rect 450486 514320 450492 514384
rect 450556 514320 450562 514384
rect 361757 513770 361823 513773
rect 359812 513768 361823 513770
rect 359812 513712 361762 513768
rect 361818 513712 361823 513768
rect 359812 513710 361823 513712
rect 361757 513707 361823 513710
rect 492121 512478 492187 512481
rect 491924 512476 492187 512478
rect 491924 512420 492126 512476
rect 492182 512420 492187 512476
rect 491924 512418 492187 512420
rect 492121 512415 492187 512418
rect 450537 512410 450603 512413
rect 450494 512408 450603 512410
rect 450494 512352 450542 512408
rect 450598 512352 450603 512408
rect 450494 512347 450603 512352
rect 450494 512176 450554 512347
rect 580165 511322 580231 511325
rect 583520 511322 584960 511412
rect 580165 511320 584960 511322
rect 580165 511264 580170 511320
rect 580226 511264 584960 511320
rect 580165 511262 584960 511264
rect 580165 511259 580231 511262
rect 583520 511172 584960 511262
rect 450353 510234 450419 510237
rect 450310 510232 450419 510234
rect 450310 510176 450358 510232
rect 450414 510176 450419 510232
rect 450310 510171 450419 510176
rect 450310 510000 450370 510171
rect 491894 508874 491954 508912
rect 494145 508874 494211 508877
rect 491894 508872 494211 508874
rect 491894 508816 494150 508872
rect 494206 508816 494211 508872
rect 491894 508814 494211 508816
rect 494145 508811 494211 508814
rect 449985 507650 450051 507653
rect 450126 507650 450186 507824
rect 449985 507648 450186 507650
rect 449985 507592 449990 507648
rect 450046 507592 450186 507648
rect 449985 507590 450186 507592
rect 449985 507587 450051 507590
rect 494237 505746 494303 505749
rect 495065 505746 495131 505749
rect 491894 505744 495131 505746
rect 491894 505688 494242 505744
rect 494298 505688 495070 505744
rect 495126 505688 495131 505744
rect 491894 505686 495131 505688
rect 450126 505477 450186 505648
rect 450077 505474 450186 505477
rect 450629 505474 450695 505477
rect 450077 505472 450695 505474
rect 450077 505416 450082 505472
rect 450138 505416 450634 505472
rect 450690 505416 450695 505472
rect 450077 505414 450695 505416
rect 450077 505411 450143 505414
rect 450629 505411 450695 505414
rect 491894 505376 491954 505686
rect 494237 505683 494303 505686
rect 495065 505683 495131 505686
rect 449709 503502 449775 503505
rect 449709 503500 450156 503502
rect 449709 503444 449714 503500
rect 449770 503472 450156 503500
rect 449770 503444 450186 503472
rect 449709 503442 450186 503444
rect 449709 503439 449775 503442
rect 450126 503301 450186 503442
rect 450126 503296 450235 503301
rect 450126 503240 450174 503296
rect 450230 503240 450235 503296
rect 450126 503238 450235 503240
rect 450169 503235 450235 503238
rect 361757 502754 361823 502757
rect 359812 502752 361823 502754
rect 359812 502696 361762 502752
rect 361818 502696 361823 502752
rect 359812 502694 361823 502696
rect 361757 502691 361823 502694
rect 519629 502346 519695 502349
rect 527214 502346 527220 502348
rect 519629 502344 527220 502346
rect 519629 502288 519634 502344
rect 519690 502288 527220 502344
rect 519629 502286 527220 502288
rect 519629 502283 519695 502286
rect 527214 502284 527220 502286
rect 527284 502284 527290 502348
rect -960 501802 480 501892
rect 3785 501802 3851 501805
rect -960 501800 3851 501802
rect -960 501744 3790 501800
rect 3846 501744 3851 501800
rect -960 501742 3851 501744
rect -960 501652 480 501742
rect 3785 501739 3851 501742
rect 491894 501666 491954 501840
rect 470550 501606 491954 501666
rect 450678 501122 450738 501296
rect 463141 501122 463207 501125
rect 470550 501122 470610 501606
rect 491894 501258 491954 501606
rect 494697 501258 494763 501261
rect 491894 501256 494763 501258
rect 491894 501200 494702 501256
rect 494758 501200 494763 501256
rect 491894 501198 494763 501200
rect 494697 501195 494763 501198
rect 450678 501120 470610 501122
rect 450678 501064 463146 501120
rect 463202 501064 470610 501120
rect 450678 501062 470610 501064
rect 463141 501059 463207 501062
rect 583520 497844 584960 498084
rect 489177 496906 489243 496909
rect 489310 496906 489316 496908
rect 489177 496904 489316 496906
rect 489177 496848 489182 496904
rect 489238 496848 489316 496904
rect 489177 496846 489316 496848
rect 489177 496843 489243 496846
rect 489310 496844 489316 496846
rect 489380 496844 489386 496908
rect 361757 491738 361823 491741
rect 359812 491736 361823 491738
rect 359812 491680 361762 491736
rect 361818 491680 361823 491736
rect 359812 491678 361823 491680
rect 361757 491675 361823 491678
rect -960 488596 480 488836
rect 580165 484666 580231 484669
rect 583520 484666 584960 484756
rect 580165 484664 584960 484666
rect 580165 484608 580170 484664
rect 580226 484608 584960 484664
rect 580165 484606 584960 484608
rect 580165 484603 580231 484606
rect 583520 484516 584960 484606
rect 361757 480722 361823 480725
rect 359812 480720 361823 480722
rect 359812 480664 361762 480720
rect 361818 480664 361823 480720
rect 359812 480662 361823 480664
rect 361757 480659 361823 480662
rect -960 475690 480 475780
rect 3693 475690 3759 475693
rect -960 475688 3759 475690
rect -960 475632 3698 475688
rect 3754 475632 3759 475688
rect -960 475630 3759 475632
rect -960 475540 480 475630
rect 3693 475627 3759 475630
rect 580533 471474 580599 471477
rect 583520 471474 584960 471564
rect 580533 471472 584960 471474
rect 580533 471416 580538 471472
rect 580594 471416 584960 471472
rect 580533 471414 584960 471416
rect 580533 471411 580599 471414
rect 583520 471324 584960 471414
rect 361757 469706 361823 469709
rect 359812 469704 361823 469706
rect 359812 469648 361762 469704
rect 361818 469648 361823 469704
rect 359812 469646 361823 469648
rect 361757 469643 361823 469646
rect 473721 462906 473787 462909
rect 482686 462906 482692 462908
rect 473721 462904 482692 462906
rect 473721 462848 473726 462904
rect 473782 462848 482692 462904
rect 473721 462846 482692 462848
rect 473721 462843 473787 462846
rect 482686 462844 482692 462846
rect 482756 462906 482762 462908
rect 521745 462906 521811 462909
rect 482756 462904 521811 462906
rect 482756 462848 521750 462904
rect 521806 462848 521811 462904
rect 482756 462846 521811 462848
rect 482756 462844 482762 462846
rect 521745 462843 521811 462846
rect -960 462634 480 462724
rect 3509 462634 3575 462637
rect -960 462632 3575 462634
rect -960 462576 3514 462632
rect 3570 462576 3575 462632
rect -960 462574 3575 462576
rect -960 462484 480 462574
rect 3509 462571 3575 462574
rect 361757 458690 361823 458693
rect 359812 458688 361823 458690
rect 359812 458632 361762 458688
rect 361818 458632 361823 458688
rect 359812 458630 361823 458632
rect 361757 458627 361823 458630
rect 580165 458146 580231 458149
rect 583520 458146 584960 458236
rect 580165 458144 584960 458146
rect 580165 458088 580170 458144
rect 580226 458088 584960 458144
rect 580165 458086 584960 458088
rect 580165 458083 580231 458086
rect 583520 457996 584960 458086
rect -960 449578 480 449668
rect 3417 449578 3483 449581
rect -960 449576 3483 449578
rect -960 449520 3422 449576
rect 3478 449520 3483 449576
rect -960 449518 3483 449520
rect -960 449428 480 449518
rect 3417 449515 3483 449518
rect 361757 447674 361823 447677
rect 359812 447672 361823 447674
rect 359812 447616 361762 447672
rect 361818 447616 361823 447672
rect 359812 447614 361823 447616
rect 361757 447611 361823 447614
rect 447409 447266 447475 447269
rect 448278 447266 448284 447268
rect 447409 447264 448284 447266
rect 447409 447208 447414 447264
rect 447470 447208 448284 447264
rect 447409 447206 448284 447208
rect 447409 447203 447475 447206
rect 448278 447204 448284 447206
rect 448348 447204 448354 447268
rect 583520 444668 584960 444908
rect 557533 442914 557599 442917
rect 555956 442912 557599 442914
rect 555956 442856 557538 442912
rect 557594 442856 557599 442912
rect 555956 442854 557599 442856
rect 557533 442851 557599 442854
rect -960 436508 480 436748
rect 361757 436658 361823 436661
rect 359812 436656 361823 436658
rect 359812 436600 361762 436656
rect 361818 436600 361823 436656
rect 359812 436598 361823 436600
rect 361757 436595 361823 436598
rect 580625 431626 580691 431629
rect 583520 431626 584960 431716
rect 580625 431624 584960 431626
rect 580625 431568 580630 431624
rect 580686 431568 584960 431624
rect 580625 431566 584960 431568
rect 580625 431563 580691 431566
rect 583520 431476 584960 431566
rect 458950 428436 458956 428500
rect 459020 428498 459026 428500
rect 476113 428498 476179 428501
rect 459020 428496 476179 428498
rect 459020 428440 476118 428496
rect 476174 428440 476179 428496
rect 459020 428438 476179 428440
rect 459020 428436 459026 428438
rect 476113 428435 476179 428438
rect 361757 425642 361823 425645
rect 359812 425640 361823 425642
rect 359812 425584 361762 425640
rect 361818 425584 361823 425640
rect 359812 425582 361823 425584
rect 361757 425579 361823 425582
rect -960 423602 480 423692
rect 3601 423602 3667 423605
rect -960 423600 3667 423602
rect -960 423544 3606 423600
rect 3662 423544 3667 423600
rect -960 423542 3667 423544
rect -960 423452 480 423542
rect 3601 423539 3667 423542
rect 447777 422378 447843 422381
rect 444330 422376 447843 422378
rect 444330 422320 447782 422376
rect 447838 422320 447843 422376
rect 444330 422318 447843 422320
rect 443494 421908 443500 421972
rect 443564 421970 443570 421972
rect 444189 421970 444255 421973
rect 443564 421968 444255 421970
rect 443564 421912 444194 421968
rect 444250 421912 444255 421968
rect 443564 421910 444255 421912
rect 443564 421908 443570 421910
rect 444189 421907 444255 421910
rect 444046 421772 444052 421836
rect 444116 421834 444122 421836
rect 444330 421834 444390 422318
rect 447777 422315 447843 422318
rect 444116 421774 444390 421834
rect 444116 421772 444122 421774
rect 580717 418298 580783 418301
rect 583520 418298 584960 418388
rect 580717 418296 584960 418298
rect 580717 418240 580722 418296
rect 580778 418240 584960 418296
rect 580717 418238 584960 418240
rect 580717 418235 580783 418238
rect 583520 418148 584960 418238
rect 361573 414626 361639 414629
rect 359812 414624 361639 414626
rect 359812 414568 361578 414624
rect 361634 414568 361639 414624
rect 359812 414566 361639 414568
rect 361573 414563 361639 414566
rect -960 410546 480 410636
rect 3969 410546 4035 410549
rect -960 410544 4035 410546
rect -960 410488 3974 410544
rect 4030 410488 4035 410544
rect -960 410486 4035 410488
rect -960 410396 480 410486
rect 3969 410483 4035 410486
rect 580165 404970 580231 404973
rect 583520 404970 584960 405060
rect 580165 404968 584960 404970
rect 580165 404912 580170 404968
rect 580226 404912 584960 404968
rect 580165 404910 584960 404912
rect 580165 404907 580231 404910
rect 583520 404820 584960 404910
rect 361573 403610 361639 403613
rect 359812 403608 361639 403610
rect 359812 403552 361578 403608
rect 361634 403552 361639 403608
rect 359812 403550 361639 403552
rect 361573 403547 361639 403550
rect -960 397490 480 397580
rect 3785 397490 3851 397493
rect -960 397488 3851 397490
rect -960 397432 3790 397488
rect 3846 397432 3851 397488
rect -960 397430 3851 397432
rect -960 397340 480 397430
rect 3785 397427 3851 397430
rect 361573 392594 361639 392597
rect 359812 392592 361639 392594
rect 359812 392536 361578 392592
rect 361634 392536 361639 392592
rect 359812 392534 361639 392536
rect 361573 392531 361639 392534
rect 448094 392532 448100 392596
rect 448164 392594 448170 392596
rect 493317 392594 493383 392597
rect 448164 392592 493383 392594
rect 448164 392536 493322 392592
rect 493378 392536 493383 392592
rect 448164 392534 493383 392536
rect 448164 392532 448170 392534
rect 493317 392531 493383 392534
rect 583520 391628 584960 391868
rect 472157 389060 472223 389061
rect 474365 389060 474431 389061
rect 472157 389058 472204 389060
rect 472112 389056 472204 389058
rect 472112 389000 472162 389056
rect 472112 388998 472204 389000
rect 472157 388996 472204 388998
rect 472268 388996 472274 389060
rect 474365 389058 474412 389060
rect 474320 389056 474412 389058
rect 474320 389000 474370 389056
rect 474320 388998 474412 389000
rect 474365 388996 474412 388998
rect 474476 388996 474482 389060
rect 478822 388996 478828 389060
rect 478892 389058 478898 389060
rect 479517 389058 479583 389061
rect 478892 389056 479583 389058
rect 478892 389000 479522 389056
rect 479578 389000 479583 389056
rect 478892 388998 479583 389000
rect 478892 388996 478898 388998
rect 472157 388995 472223 388996
rect 474365 388995 474431 388996
rect 479517 388995 479583 388998
rect 472014 388860 472020 388924
rect 472084 388922 472090 388924
rect 472893 388922 472959 388925
rect 472084 388920 472959 388922
rect 472084 388864 472898 388920
rect 472954 388864 472959 388920
rect 472084 388862 472959 388864
rect 472084 388860 472090 388862
rect 472893 388859 472959 388862
rect 449065 387018 449131 387021
rect 489310 387018 489316 387020
rect 449065 387016 489316 387018
rect 449065 386960 449070 387016
rect 449126 386960 489316 387016
rect 449065 386958 489316 386960
rect 449065 386955 449131 386958
rect 489310 386956 489316 386958
rect 489380 386956 489386 387020
rect 513189 384706 513255 384709
rect 509956 384704 513255 384706
rect 509956 384648 513194 384704
rect 513250 384648 513255 384704
rect 509956 384646 513255 384648
rect 513189 384643 513255 384646
rect -960 384284 480 384524
rect 513281 384162 513347 384165
rect 509956 384160 513347 384162
rect 509956 384104 513286 384160
rect 513342 384104 513347 384160
rect 509956 384102 513347 384104
rect 513281 384099 513347 384102
rect 447133 383618 447199 383621
rect 512637 383618 512703 383621
rect 447133 383616 450156 383618
rect 447133 383560 447138 383616
rect 447194 383560 450156 383616
rect 447133 383558 450156 383560
rect 509956 383616 512703 383618
rect 509956 383560 512642 383616
rect 512698 383560 512703 383616
rect 509956 383558 512703 383560
rect 447133 383555 447199 383558
rect 512637 383555 512703 383558
rect 513005 383074 513071 383077
rect 509956 383072 513071 383074
rect 509956 383016 513010 383072
rect 513066 383016 513071 383072
rect 509956 383014 513071 383016
rect 513005 383011 513071 383014
rect 447225 382938 447291 382941
rect 447225 382936 450156 382938
rect 447225 382880 447230 382936
rect 447286 382880 450156 382936
rect 447225 382878 450156 382880
rect 447225 382875 447291 382878
rect 512453 382530 512519 382533
rect 509956 382528 512519 382530
rect 509956 382472 512458 382528
rect 512514 382472 512519 382528
rect 509956 382470 512519 382472
rect 512453 382467 512519 382470
rect 447133 382258 447199 382261
rect 447133 382256 450156 382258
rect 447133 382200 447138 382256
rect 447194 382200 450156 382256
rect 447133 382198 450156 382200
rect 447133 382195 447199 382198
rect 513005 381986 513071 381989
rect 509956 381984 513071 381986
rect 509956 381928 513010 381984
rect 513066 381928 513071 381984
rect 509956 381926 513071 381928
rect 513005 381923 513071 381926
rect 361573 381578 361639 381581
rect 359812 381576 361639 381578
rect 359812 381520 361578 381576
rect 361634 381520 361639 381576
rect 359812 381518 361639 381520
rect 361573 381515 361639 381518
rect 447225 381578 447291 381581
rect 447225 381576 450156 381578
rect 447225 381520 447230 381576
rect 447286 381520 450156 381576
rect 447225 381518 450156 381520
rect 447225 381515 447291 381518
rect 512453 381442 512519 381445
rect 509956 381440 512519 381442
rect 509956 381384 512458 381440
rect 512514 381384 512519 381440
rect 509956 381382 512519 381384
rect 512453 381379 512519 381382
rect 447225 380898 447291 380901
rect 513189 380898 513255 380901
rect 447225 380896 450156 380898
rect 447225 380840 447230 380896
rect 447286 380840 450156 380896
rect 447225 380838 450156 380840
rect 509956 380896 513255 380898
rect 509956 380840 513194 380896
rect 513250 380840 513255 380896
rect 509956 380838 513255 380840
rect 447225 380835 447291 380838
rect 513189 380835 513255 380838
rect 513281 380354 513347 380357
rect 509956 380352 513347 380354
rect 509956 380296 513286 380352
rect 513342 380296 513347 380352
rect 509956 380294 513347 380296
rect 513281 380291 513347 380294
rect 447133 380218 447199 380221
rect 447133 380216 450156 380218
rect 447133 380160 447138 380216
rect 447194 380160 450156 380216
rect 447133 380158 450156 380160
rect 447133 380155 447199 380158
rect 512545 379810 512611 379813
rect 509956 379808 512611 379810
rect 509956 379752 512550 379808
rect 512606 379752 512611 379808
rect 509956 379750 512611 379752
rect 512545 379747 512611 379750
rect 447409 379538 447475 379541
rect 447409 379536 450156 379538
rect 447409 379480 447414 379536
rect 447470 379480 450156 379536
rect 447409 379478 450156 379480
rect 447409 379475 447475 379478
rect 512821 379266 512887 379269
rect 509956 379264 512887 379266
rect 509956 379208 512826 379264
rect 512882 379208 512887 379264
rect 509956 379206 512887 379208
rect 512821 379203 512887 379206
rect 447133 378858 447199 378861
rect 447133 378856 450156 378858
rect 447133 378800 447138 378856
rect 447194 378800 450156 378856
rect 447133 378798 450156 378800
rect 447133 378795 447199 378798
rect 513281 378722 513347 378725
rect 509956 378720 513347 378722
rect 509956 378664 513286 378720
rect 513342 378664 513347 378720
rect 509956 378662 513347 378664
rect 513281 378659 513347 378662
rect 580165 378450 580231 378453
rect 583520 378450 584960 378540
rect 580165 378448 584960 378450
rect 580165 378392 580170 378448
rect 580226 378392 584960 378448
rect 580165 378390 584960 378392
rect 580165 378387 580231 378390
rect 583520 378300 584960 378390
rect 447317 378178 447383 378181
rect 512269 378178 512335 378181
rect 447317 378176 450156 378178
rect 447317 378120 447322 378176
rect 447378 378120 450156 378176
rect 447317 378118 450156 378120
rect 509956 378176 512335 378178
rect 509956 378120 512274 378176
rect 512330 378120 512335 378176
rect 509956 378118 512335 378120
rect 447317 378115 447383 378118
rect 512269 378115 512335 378118
rect 512453 377634 512519 377637
rect 509956 377632 512519 377634
rect 509956 377576 512458 377632
rect 512514 377576 512519 377632
rect 509956 377574 512519 377576
rect 512453 377571 512519 377574
rect 447133 377498 447199 377501
rect 447133 377496 450156 377498
rect 447133 377440 447138 377496
rect 447194 377440 450156 377496
rect 447133 377438 450156 377440
rect 447133 377435 447199 377438
rect 513189 377090 513255 377093
rect 509956 377088 513255 377090
rect 509956 377032 513194 377088
rect 513250 377032 513255 377088
rect 509956 377030 513255 377032
rect 513189 377027 513255 377030
rect 447225 376818 447291 376821
rect 447225 376816 450156 376818
rect 447225 376760 447230 376816
rect 447286 376760 450156 376816
rect 447225 376758 450156 376760
rect 447225 376755 447291 376758
rect 512361 376546 512427 376549
rect 509956 376544 512427 376546
rect 509956 376488 512366 376544
rect 512422 376488 512427 376544
rect 509956 376486 512427 376488
rect 512361 376483 512427 376486
rect 447133 376138 447199 376141
rect 447133 376136 450156 376138
rect 447133 376080 447138 376136
rect 447194 376080 450156 376136
rect 447133 376078 450156 376080
rect 447133 376075 447199 376078
rect 512085 376002 512151 376005
rect 509956 376000 512151 376002
rect 509956 375944 512090 376000
rect 512146 375944 512151 376000
rect 509956 375942 512151 375944
rect 512085 375939 512151 375942
rect 509325 375594 509391 375597
rect 509325 375592 509434 375594
rect 509325 375536 509330 375592
rect 509386 375536 509434 375592
rect 509325 375531 509434 375536
rect 447225 375458 447291 375461
rect 447225 375456 450156 375458
rect 447225 375400 447230 375456
rect 447286 375400 450156 375456
rect 509374 375428 509434 375531
rect 447225 375398 450156 375400
rect 447225 375395 447291 375398
rect 511993 374914 512059 374917
rect 509956 374912 512059 374914
rect 509956 374856 511998 374912
rect 512054 374856 512059 374912
rect 509956 374854 512059 374856
rect 511993 374851 512059 374854
rect 447133 374778 447199 374781
rect 447133 374776 450156 374778
rect 447133 374720 447138 374776
rect 447194 374720 450156 374776
rect 447133 374718 450156 374720
rect 447133 374715 447199 374718
rect 513281 374370 513347 374373
rect 509956 374368 513347 374370
rect 509956 374312 513286 374368
rect 513342 374312 513347 374368
rect 509956 374310 513347 374312
rect 513281 374307 513347 374310
rect 447225 374098 447291 374101
rect 447225 374096 450156 374098
rect 447225 374040 447230 374096
rect 447286 374040 450156 374096
rect 447225 374038 450156 374040
rect 447225 374035 447291 374038
rect 510705 373826 510771 373829
rect 509956 373824 510771 373826
rect 509956 373768 510710 373824
rect 510766 373768 510771 373824
rect 509956 373766 510771 373768
rect 510705 373763 510771 373766
rect 447133 373418 447199 373421
rect 447133 373416 450156 373418
rect 447133 373360 447138 373416
rect 447194 373360 450156 373416
rect 447133 373358 450156 373360
rect 447133 373355 447199 373358
rect 512637 373282 512703 373285
rect 509956 373280 512703 373282
rect 509956 373224 512642 373280
rect 512698 373224 512703 373280
rect 509956 373222 512703 373224
rect 512637 373219 512703 373222
rect 447225 372738 447291 372741
rect 513281 372738 513347 372741
rect 447225 372736 450156 372738
rect 447225 372680 447230 372736
rect 447286 372680 450156 372736
rect 447225 372678 450156 372680
rect 509956 372736 513347 372738
rect 509956 372680 513286 372736
rect 513342 372680 513347 372736
rect 509956 372678 513347 372680
rect 447225 372675 447291 372678
rect 513281 372675 513347 372678
rect 511993 372194 512059 372197
rect 509956 372192 512059 372194
rect 509956 372136 511998 372192
rect 512054 372136 512059 372192
rect 509956 372134 512059 372136
rect 511993 372131 512059 372134
rect 447133 372058 447199 372061
rect 447133 372056 450156 372058
rect 447133 372000 447138 372056
rect 447194 372000 450156 372056
rect 447133 371998 450156 372000
rect 447133 371995 447199 371998
rect 511993 371650 512059 371653
rect 509956 371648 512059 371650
rect 509956 371592 511998 371648
rect 512054 371592 512059 371648
rect 509956 371590 512059 371592
rect 511993 371587 512059 371590
rect -960 371378 480 371468
rect 3877 371378 3943 371381
rect -960 371376 3943 371378
rect -960 371320 3882 371376
rect 3938 371320 3943 371376
rect -960 371318 3943 371320
rect -960 371228 480 371318
rect 3877 371315 3943 371318
rect 447225 371378 447291 371381
rect 447225 371376 450156 371378
rect 447225 371320 447230 371376
rect 447286 371320 450156 371376
rect 447225 371318 450156 371320
rect 447225 371315 447291 371318
rect 512085 371106 512151 371109
rect 509956 371104 512151 371106
rect 509956 371048 512090 371104
rect 512146 371048 512151 371104
rect 509956 371046 512151 371048
rect 512085 371043 512151 371046
rect 447133 370698 447199 370701
rect 447133 370696 450156 370698
rect 447133 370640 447138 370696
rect 447194 370640 450156 370696
rect 447133 370638 450156 370640
rect 447133 370635 447199 370638
rect 361573 370562 361639 370565
rect 513281 370562 513347 370565
rect 359812 370560 361639 370562
rect 359812 370504 361578 370560
rect 361634 370504 361639 370560
rect 359812 370502 361639 370504
rect 509956 370560 513347 370562
rect 509956 370504 513286 370560
rect 513342 370504 513347 370560
rect 509956 370502 513347 370504
rect 361573 370499 361639 370502
rect 513281 370499 513347 370502
rect 447225 370018 447291 370021
rect 513281 370018 513347 370021
rect 447225 370016 450156 370018
rect 447225 369960 447230 370016
rect 447286 369960 450156 370016
rect 447225 369958 450156 369960
rect 509956 370016 513347 370018
rect 509956 369960 513286 370016
rect 513342 369960 513347 370016
rect 509956 369958 513347 369960
rect 447225 369955 447291 369958
rect 513281 369955 513347 369958
rect 512085 369474 512151 369477
rect 509956 369472 512151 369474
rect 509956 369416 512090 369472
rect 512146 369416 512151 369472
rect 509956 369414 512151 369416
rect 512085 369411 512151 369414
rect 447133 369338 447199 369341
rect 447133 369336 450156 369338
rect 447133 369280 447138 369336
rect 447194 369280 450156 369336
rect 447133 369278 450156 369280
rect 447133 369275 447199 369278
rect 512269 368930 512335 368933
rect 509956 368928 512335 368930
rect 509956 368872 512274 368928
rect 512330 368872 512335 368928
rect 509956 368870 512335 368872
rect 512269 368867 512335 368870
rect 447225 368658 447291 368661
rect 447225 368656 450156 368658
rect 447225 368600 447230 368656
rect 447286 368600 450156 368656
rect 447225 368598 450156 368600
rect 447225 368595 447291 368598
rect 512177 368386 512243 368389
rect 509956 368384 512243 368386
rect 509956 368328 512182 368384
rect 512238 368328 512243 368384
rect 509956 368326 512243 368328
rect 512177 368323 512243 368326
rect 447133 367978 447199 367981
rect 447133 367976 450156 367978
rect 447133 367920 447138 367976
rect 447194 367920 450156 367976
rect 447133 367918 450156 367920
rect 447133 367915 447199 367918
rect 513281 367842 513347 367845
rect 509956 367840 513347 367842
rect 509956 367784 513286 367840
rect 513342 367784 513347 367840
rect 509956 367782 513347 367784
rect 513281 367779 513347 367782
rect 447225 367298 447291 367301
rect 447225 367296 450156 367298
rect 447225 367240 447230 367296
rect 447286 367240 450156 367296
rect 447225 367238 450156 367240
rect 447225 367235 447291 367238
rect 509558 367029 509618 367268
rect 509509 367024 509618 367029
rect 509509 366968 509514 367024
rect 509570 366968 509618 367024
rect 509509 366966 509618 366968
rect 509509 366963 509575 366966
rect 513281 366754 513347 366757
rect 509956 366752 513347 366754
rect 509956 366696 513286 366752
rect 513342 366696 513347 366752
rect 509956 366694 513347 366696
rect 513281 366691 513347 366694
rect 447133 366618 447199 366621
rect 447133 366616 450156 366618
rect 447133 366560 447138 366616
rect 447194 366560 450156 366616
rect 447133 366558 450156 366560
rect 447133 366555 447199 366558
rect 513373 366210 513439 366213
rect 509956 366208 513439 366210
rect 509956 366152 513378 366208
rect 513434 366152 513439 366208
rect 509956 366150 513439 366152
rect 513373 366147 513439 366150
rect 447225 365938 447291 365941
rect 447225 365936 450156 365938
rect 447225 365880 447230 365936
rect 447286 365880 450156 365936
rect 447225 365878 450156 365880
rect 447225 365875 447291 365878
rect 511993 365666 512059 365669
rect 509956 365664 512059 365666
rect 509956 365608 511998 365664
rect 512054 365608 512059 365664
rect 509956 365606 512059 365608
rect 511993 365603 512059 365606
rect 447225 365258 447291 365261
rect 447225 365256 450156 365258
rect 447225 365200 447230 365256
rect 447286 365200 450156 365256
rect 447225 365198 450156 365200
rect 447225 365195 447291 365198
rect 512821 365122 512887 365125
rect 509956 365120 512887 365122
rect 509956 365064 512826 365120
rect 512882 365064 512887 365120
rect 509956 365062 512887 365064
rect 512821 365059 512887 365062
rect 580165 365122 580231 365125
rect 583520 365122 584960 365212
rect 580165 365120 584960 365122
rect 580165 365064 580170 365120
rect 580226 365064 584960 365120
rect 580165 365062 584960 365064
rect 580165 365059 580231 365062
rect 583520 364972 584960 365062
rect 447133 364578 447199 364581
rect 513281 364578 513347 364581
rect 447133 364576 450156 364578
rect 447133 364520 447138 364576
rect 447194 364520 450156 364576
rect 447133 364518 450156 364520
rect 509956 364576 513347 364578
rect 509956 364520 513286 364576
rect 513342 364520 513347 364576
rect 509956 364518 513347 364520
rect 447133 364515 447199 364518
rect 513281 364515 513347 364518
rect 511993 364034 512059 364037
rect 509956 364032 512059 364034
rect 509956 363976 511998 364032
rect 512054 363976 512059 364032
rect 509956 363974 512059 363976
rect 511993 363971 512059 363974
rect 447225 363898 447291 363901
rect 447225 363896 450156 363898
rect 447225 363840 447230 363896
rect 447286 363840 450156 363896
rect 447225 363838 450156 363840
rect 447225 363835 447291 363838
rect 512269 363490 512335 363493
rect 509956 363488 512335 363490
rect 509956 363432 512274 363488
rect 512330 363432 512335 363488
rect 509956 363430 512335 363432
rect 512269 363427 512335 363430
rect 447133 363218 447199 363221
rect 447133 363216 450156 363218
rect 447133 363160 447138 363216
rect 447194 363160 450156 363216
rect 447133 363158 450156 363160
rect 447133 363155 447199 363158
rect 513005 362946 513071 362949
rect 509956 362944 513071 362946
rect 509956 362888 513010 362944
rect 513066 362888 513071 362944
rect 509956 362886 513071 362888
rect 513005 362883 513071 362886
rect 447133 362538 447199 362541
rect 447133 362536 450156 362538
rect 447133 362480 447138 362536
rect 447194 362480 450156 362536
rect 447133 362478 450156 362480
rect 447133 362475 447199 362478
rect 511993 362402 512059 362405
rect 509956 362400 512059 362402
rect 509956 362344 511998 362400
rect 512054 362344 512059 362400
rect 509956 362342 512059 362344
rect 511993 362339 512059 362342
rect 447225 361858 447291 361861
rect 513281 361858 513347 361861
rect 447225 361856 450156 361858
rect 447225 361800 447230 361856
rect 447286 361800 450156 361856
rect 447225 361798 450156 361800
rect 509956 361856 513347 361858
rect 509956 361800 513286 361856
rect 513342 361800 513347 361856
rect 509956 361798 513347 361800
rect 447225 361795 447291 361798
rect 513281 361795 513347 361798
rect 512637 361314 512703 361317
rect 509956 361312 512703 361314
rect 509956 361256 512642 361312
rect 512698 361256 512703 361312
rect 509956 361254 512703 361256
rect 512637 361251 512703 361254
rect 447225 361178 447291 361181
rect 447225 361176 450156 361178
rect 447225 361120 447230 361176
rect 447286 361120 450156 361176
rect 447225 361118 450156 361120
rect 447225 361115 447291 361118
rect 511993 360770 512059 360773
rect 509956 360768 512059 360770
rect 509956 360712 511998 360768
rect 512054 360712 512059 360768
rect 509956 360710 512059 360712
rect 511993 360707 512059 360710
rect 447133 360498 447199 360501
rect 447133 360496 450156 360498
rect 447133 360440 447138 360496
rect 447194 360440 450156 360496
rect 447133 360438 450156 360440
rect 447133 360435 447199 360438
rect 512361 360226 512427 360229
rect 509956 360224 512427 360226
rect 509956 360168 512366 360224
rect 512422 360168 512427 360224
rect 509956 360166 512427 360168
rect 512361 360163 512427 360166
rect 447133 359818 447199 359821
rect 447133 359816 450156 359818
rect 447133 359760 447138 359816
rect 447194 359760 450156 359816
rect 447133 359758 450156 359760
rect 447133 359755 447199 359758
rect 513005 359682 513071 359685
rect 509956 359680 513071 359682
rect 509956 359624 513010 359680
rect 513066 359624 513071 359680
rect 509956 359622 513071 359624
rect 513005 359619 513071 359622
rect 362217 359546 362283 359549
rect 359812 359544 362283 359546
rect 359812 359488 362222 359544
rect 362278 359488 362283 359544
rect 359812 359486 362283 359488
rect 362217 359483 362283 359486
rect 447225 359138 447291 359141
rect 510797 359138 510863 359141
rect 447225 359136 450156 359138
rect 447225 359080 447230 359136
rect 447286 359080 450156 359136
rect 447225 359078 450156 359080
rect 509956 359136 510863 359138
rect 509956 359080 510802 359136
rect 510858 359080 510863 359136
rect 509956 359078 510863 359080
rect 447225 359075 447291 359078
rect 510797 359075 510863 359078
rect 512545 358594 512611 358597
rect 509956 358592 512611 358594
rect -960 358458 480 358548
rect 509956 358536 512550 358592
rect 512606 358536 512611 358592
rect 509956 358534 512611 358536
rect 512545 358531 512611 358534
rect 3509 358458 3575 358461
rect -960 358456 3575 358458
rect -960 358400 3514 358456
rect 3570 358400 3575 358456
rect -960 358398 3575 358400
rect -960 358308 480 358398
rect 3509 358395 3575 358398
rect 448973 358458 449039 358461
rect 448973 358456 450156 358458
rect 448973 358400 448978 358456
rect 449034 358400 450156 358456
rect 448973 358398 450156 358400
rect 448973 358395 449039 358398
rect 513557 358050 513623 358053
rect 509956 358048 513623 358050
rect 509956 357992 513562 358048
rect 513618 357992 513623 358048
rect 509956 357990 513623 357992
rect 513557 357987 513623 357990
rect 449617 357778 449683 357781
rect 449617 357776 450156 357778
rect 449617 357720 449622 357776
rect 449678 357720 450156 357776
rect 449617 357718 450156 357720
rect 449617 357715 449683 357718
rect 509417 357642 509483 357645
rect 509374 357640 509483 357642
rect 509374 357584 509422 357640
rect 509478 357584 509483 357640
rect 509374 357579 509483 357584
rect 509374 357476 509434 357579
rect 449065 357098 449131 357101
rect 449065 357096 450156 357098
rect 449065 357040 449070 357096
rect 449126 357040 450156 357096
rect 449065 357038 450156 357040
rect 449065 357035 449131 357038
rect 513281 356962 513347 356965
rect 509956 356960 513347 356962
rect 509956 356904 513286 356960
rect 513342 356904 513347 356960
rect 509956 356902 513347 356904
rect 513281 356899 513347 356902
rect 449709 356418 449775 356421
rect 512821 356418 512887 356421
rect 449709 356416 450156 356418
rect 449709 356360 449714 356416
rect 449770 356360 450156 356416
rect 449709 356358 450156 356360
rect 509956 356416 512887 356418
rect 509956 356360 512826 356416
rect 512882 356360 512887 356416
rect 509956 356358 512887 356360
rect 449709 356355 449775 356358
rect 512821 356355 512887 356358
rect 510981 355874 511047 355877
rect 509956 355872 511047 355874
rect 509956 355816 510986 355872
rect 511042 355816 511047 355872
rect 509956 355814 511047 355816
rect 510981 355811 511047 355814
rect 448421 355738 448487 355741
rect 448421 355736 450156 355738
rect 448421 355680 448426 355736
rect 448482 355680 450156 355736
rect 448421 355678 450156 355680
rect 448421 355675 448487 355678
rect 513281 355330 513347 355333
rect 509956 355328 513347 355330
rect 509956 355272 513286 355328
rect 513342 355272 513347 355328
rect 509956 355270 513347 355272
rect 513281 355267 513347 355270
rect 447501 355058 447567 355061
rect 447501 355056 450156 355058
rect 447501 355000 447506 355056
rect 447562 355000 450156 355056
rect 447501 354998 450156 355000
rect 447501 354995 447567 354998
rect 513281 354786 513347 354789
rect 509956 354784 513347 354786
rect 509956 354728 513286 354784
rect 513342 354728 513347 354784
rect 509956 354726 513347 354728
rect 513281 354723 513347 354726
rect 447777 354378 447843 354381
rect 447777 354376 450156 354378
rect 447777 354320 447782 354376
rect 447838 354320 450156 354376
rect 447777 354318 450156 354320
rect 447777 354315 447843 354318
rect 512085 354242 512151 354245
rect 509956 354240 512151 354242
rect 509956 354184 512090 354240
rect 512146 354184 512151 354240
rect 509956 354182 512151 354184
rect 512085 354179 512151 354182
rect 447685 353698 447751 353701
rect 513281 353698 513347 353701
rect 447685 353696 450156 353698
rect 447685 353640 447690 353696
rect 447746 353640 450156 353696
rect 447685 353638 450156 353640
rect 509956 353696 513347 353698
rect 509956 353640 513286 353696
rect 513342 353640 513347 353696
rect 509956 353638 513347 353640
rect 447685 353635 447751 353638
rect 513281 353635 513347 353638
rect 510889 353154 510955 353157
rect 509956 353152 510955 353154
rect 509956 353096 510894 353152
rect 510950 353096 510955 353152
rect 509956 353094 510955 353096
rect 510889 353091 510955 353094
rect 447869 353018 447935 353021
rect 447869 353016 450156 353018
rect 447869 352960 447874 353016
rect 447930 352960 450156 353016
rect 447869 352958 450156 352960
rect 447869 352955 447935 352958
rect 512453 352610 512519 352613
rect 509956 352608 512519 352610
rect 509956 352552 512458 352608
rect 512514 352552 512519 352608
rect 509956 352550 512519 352552
rect 512453 352547 512519 352550
rect 448053 352338 448119 352341
rect 448053 352336 450156 352338
rect 448053 352280 448058 352336
rect 448114 352280 450156 352336
rect 448053 352278 450156 352280
rect 448053 352275 448119 352278
rect 509742 351797 509802 352036
rect 580809 351930 580875 351933
rect 583520 351930 584960 352020
rect 580809 351928 584960 351930
rect 580809 351872 580814 351928
rect 580870 351872 584960 351928
rect 580809 351870 584960 351872
rect 580809 351867 580875 351870
rect 509742 351792 509851 351797
rect 509742 351736 509790 351792
rect 509846 351736 509851 351792
rect 583520 351780 584960 351870
rect 509742 351734 509851 351736
rect 509785 351731 509851 351734
rect 447317 351658 447383 351661
rect 447317 351656 450156 351658
rect 447317 351600 447322 351656
rect 447378 351600 450156 351656
rect 447317 351598 450156 351600
rect 447317 351595 447383 351598
rect 512913 351522 512979 351525
rect 509956 351520 512979 351522
rect 509956 351464 512918 351520
rect 512974 351464 512979 351520
rect 509956 351462 512979 351464
rect 512913 351459 512979 351462
rect 447133 350978 447199 350981
rect 512453 350978 512519 350981
rect 447133 350976 450156 350978
rect 447133 350920 447138 350976
rect 447194 350920 450156 350976
rect 447133 350918 450156 350920
rect 509956 350976 512519 350978
rect 509956 350920 512458 350976
rect 512514 350920 512519 350976
rect 509956 350918 512519 350920
rect 447133 350915 447199 350918
rect 512453 350915 512519 350918
rect 513281 350434 513347 350437
rect 509956 350432 513347 350434
rect 509956 350376 513286 350432
rect 513342 350376 513347 350432
rect 509956 350374 513347 350376
rect 513281 350371 513347 350374
rect 449709 350298 449775 350301
rect 449709 350296 450156 350298
rect 449709 350240 449714 350296
rect 449770 350240 450156 350296
rect 449709 350238 450156 350240
rect 449709 350235 449775 350238
rect 512821 349890 512887 349893
rect 509956 349888 512887 349890
rect 509956 349832 512826 349888
rect 512882 349832 512887 349888
rect 509956 349830 512887 349832
rect 512821 349827 512887 349830
rect 449801 349618 449867 349621
rect 449801 349616 450156 349618
rect 449801 349560 449806 349616
rect 449862 349560 450156 349616
rect 449801 349558 450156 349560
rect 449801 349555 449867 349558
rect 512085 349346 512151 349349
rect 509956 349344 512151 349346
rect 509956 349288 512090 349344
rect 512146 349288 512151 349344
rect 509956 349286 512151 349288
rect 512085 349283 512151 349286
rect 448145 348938 448211 348941
rect 448145 348936 450156 348938
rect 448145 348880 448150 348936
rect 448206 348880 450156 348936
rect 448145 348878 450156 348880
rect 448145 348875 448211 348878
rect 513281 348802 513347 348805
rect 509956 348800 513347 348802
rect 509956 348744 513286 348800
rect 513342 348744 513347 348800
rect 509956 348742 513347 348744
rect 513281 348739 513347 348742
rect 361757 348530 361823 348533
rect 359812 348528 361823 348530
rect 359812 348472 361762 348528
rect 361818 348472 361823 348528
rect 359812 348470 361823 348472
rect 361757 348467 361823 348470
rect 449433 348258 449499 348261
rect 513281 348258 513347 348261
rect 449433 348256 450156 348258
rect 449433 348200 449438 348256
rect 449494 348200 450156 348256
rect 449433 348198 450156 348200
rect 509956 348256 513347 348258
rect 509956 348200 513286 348256
rect 513342 348200 513347 348256
rect 509956 348198 513347 348200
rect 449433 348195 449499 348198
rect 513281 348195 513347 348198
rect 511073 347714 511139 347717
rect 509956 347712 511139 347714
rect 509956 347656 511078 347712
rect 511134 347656 511139 347712
rect 509956 347654 511139 347656
rect 511073 347651 511139 347654
rect 447133 347578 447199 347581
rect 447133 347576 450156 347578
rect 447133 347520 447138 347576
rect 447194 347520 450156 347576
rect 447133 347518 450156 347520
rect 447133 347515 447199 347518
rect 512085 347170 512151 347173
rect 509956 347168 512151 347170
rect 509956 347112 512090 347168
rect 512146 347112 512151 347168
rect 509956 347110 512151 347112
rect 512085 347107 512151 347110
rect 448237 346898 448303 346901
rect 448237 346896 450156 346898
rect 448237 346840 448242 346896
rect 448298 346840 450156 346896
rect 448237 346838 450156 346840
rect 448237 346835 448303 346838
rect 512637 346626 512703 346629
rect 509956 346624 512703 346626
rect 509956 346568 512642 346624
rect 512698 346568 512703 346624
rect 509956 346566 512703 346568
rect 512637 346563 512703 346566
rect 448094 346156 448100 346220
rect 448164 346218 448170 346220
rect 448164 346158 450156 346218
rect 448164 346156 448170 346158
rect 511165 346082 511231 346085
rect 509956 346080 511231 346082
rect 509956 346024 511170 346080
rect 511226 346024 511231 346080
rect 509956 346022 511231 346024
rect 511165 346019 511231 346022
rect 447869 345538 447935 345541
rect 512453 345538 512519 345541
rect 447869 345536 450156 345538
rect -960 345402 480 345492
rect 447869 345480 447874 345536
rect 447930 345480 450156 345536
rect 447869 345478 450156 345480
rect 509956 345536 512519 345538
rect 509956 345480 512458 345536
rect 512514 345480 512519 345536
rect 509956 345478 512519 345480
rect 447869 345475 447935 345478
rect 512453 345475 512519 345478
rect 3417 345402 3483 345405
rect -960 345400 3483 345402
rect -960 345344 3422 345400
rect 3478 345344 3483 345400
rect -960 345342 3483 345344
rect -960 345252 480 345342
rect 3417 345339 3483 345342
rect 512085 344994 512151 344997
rect 509956 344992 512151 344994
rect 509956 344936 512090 344992
rect 512146 344936 512151 344992
rect 509956 344934 512151 344936
rect 512085 344931 512151 344934
rect 448421 344858 448487 344861
rect 448421 344856 450156 344858
rect 448421 344800 448426 344856
rect 448482 344800 450156 344856
rect 448421 344798 450156 344800
rect 448421 344795 448487 344798
rect 449709 344178 449775 344181
rect 449709 344176 450156 344178
rect 449709 344120 449714 344176
rect 449770 344120 450156 344176
rect 449709 344118 450156 344120
rect 449709 344115 449775 344118
rect 509558 344045 509618 344420
rect 509558 344040 509667 344045
rect 509558 343984 509606 344040
rect 509662 343984 509667 344040
rect 509558 343982 509667 343984
rect 509601 343979 509667 343982
rect 512913 343906 512979 343909
rect 509956 343904 512979 343906
rect 509956 343848 512918 343904
rect 512974 343848 512979 343904
rect 509956 343846 512979 343848
rect 512913 343843 512979 343846
rect 448421 343498 448487 343501
rect 448421 343496 450156 343498
rect 448421 343440 448426 343496
rect 448482 343440 450156 343496
rect 448421 343438 450156 343440
rect 448421 343435 448487 343438
rect 513189 343362 513255 343365
rect 509956 343360 513255 343362
rect 509956 343304 513194 343360
rect 513250 343304 513255 343360
rect 509956 343302 513255 343304
rect 513189 343299 513255 343302
rect 449525 342818 449591 342821
rect 510654 342818 510660 342820
rect 449525 342816 450156 342818
rect 449525 342760 449530 342816
rect 449586 342760 450156 342816
rect 449525 342758 450156 342760
rect 509956 342758 510660 342818
rect 449525 342755 449591 342758
rect 510654 342756 510660 342758
rect 510724 342756 510730 342820
rect 513281 342274 513347 342277
rect 509956 342272 513347 342274
rect 509956 342216 513286 342272
rect 513342 342216 513347 342272
rect 509956 342214 513347 342216
rect 513281 342211 513347 342214
rect 447133 342138 447199 342141
rect 447133 342136 450156 342138
rect 447133 342080 447138 342136
rect 447194 342080 450156 342136
rect 447133 342078 450156 342080
rect 447133 342075 447199 342078
rect 512637 341730 512703 341733
rect 509956 341728 512703 341730
rect 509956 341672 512642 341728
rect 512698 341672 512703 341728
rect 509956 341670 512703 341672
rect 512637 341667 512703 341670
rect 447225 341458 447291 341461
rect 447225 341456 450156 341458
rect 447225 341400 447230 341456
rect 447286 341400 450156 341456
rect 447225 341398 450156 341400
rect 447225 341395 447291 341398
rect 512821 341186 512887 341189
rect 509956 341184 512887 341186
rect 509956 341128 512826 341184
rect 512882 341128 512887 341184
rect 509956 341126 512887 341128
rect 512821 341123 512887 341126
rect 447225 340778 447291 340781
rect 447225 340776 450156 340778
rect 447225 340720 447230 340776
rect 447286 340720 450156 340776
rect 447225 340718 450156 340720
rect 447225 340715 447291 340718
rect 513189 340642 513255 340645
rect 509956 340640 513255 340642
rect 509956 340584 513194 340640
rect 513250 340584 513255 340640
rect 509956 340582 513255 340584
rect 513189 340579 513255 340582
rect 447133 340098 447199 340101
rect 513281 340098 513347 340101
rect 447133 340096 450156 340098
rect 447133 340040 447138 340096
rect 447194 340040 450156 340096
rect 447133 340038 450156 340040
rect 509956 340096 513347 340098
rect 509956 340040 513286 340096
rect 513342 340040 513347 340096
rect 509956 340038 513347 340040
rect 447133 340035 447199 340038
rect 513281 340035 513347 340038
rect 517830 339554 517836 339556
rect 509956 339494 517836 339554
rect 517830 339492 517836 339494
rect 517900 339492 517906 339556
rect 447225 339418 447291 339421
rect 447225 339416 450156 339418
rect 447225 339360 447230 339416
rect 447286 339360 450156 339416
rect 447225 339358 450156 339360
rect 447225 339355 447291 339358
rect 512729 339010 512795 339013
rect 509956 339008 512795 339010
rect 509956 338952 512734 339008
rect 512790 338952 512795 339008
rect 509956 338950 512795 338952
rect 512729 338947 512795 338950
rect 447133 338738 447199 338741
rect 447133 338736 450156 338738
rect 447133 338680 447138 338736
rect 447194 338680 450156 338736
rect 447133 338678 450156 338680
rect 447133 338675 447199 338678
rect 513281 338466 513347 338469
rect 509956 338464 513347 338466
rect 509956 338408 513286 338464
rect 513342 338408 513347 338464
rect 583520 338452 584960 338692
rect 509956 338406 513347 338408
rect 513281 338403 513347 338406
rect 447501 338058 447567 338061
rect 447501 338056 450156 338058
rect 447501 338000 447506 338056
rect 447562 338000 450156 338056
rect 447501 337998 450156 338000
rect 447501 337995 447567 337998
rect 513097 337922 513163 337925
rect 509956 337920 513163 337922
rect 509956 337864 513102 337920
rect 513158 337864 513163 337920
rect 509956 337862 513163 337864
rect 513097 337859 513163 337862
rect 450261 337786 450327 337789
rect 450537 337786 450603 337789
rect 450261 337784 450603 337786
rect 450261 337728 450266 337784
rect 450322 337728 450542 337784
rect 450598 337728 450603 337784
rect 450261 337726 450603 337728
rect 450261 337723 450327 337726
rect 450537 337723 450603 337726
rect 361757 337514 361823 337517
rect 359812 337512 361823 337514
rect 359812 337456 361762 337512
rect 361818 337456 361823 337512
rect 359812 337454 361823 337456
rect 361757 337451 361823 337454
rect 447133 337378 447199 337381
rect 513189 337378 513255 337381
rect 447133 337376 450156 337378
rect 447133 337320 447138 337376
rect 447194 337320 450156 337376
rect 447133 337318 450156 337320
rect 509956 337376 513255 337378
rect 509956 337320 513194 337376
rect 513250 337320 513255 337376
rect 509956 337318 513255 337320
rect 447133 337315 447199 337318
rect 513189 337315 513255 337318
rect 427813 337106 427879 337109
rect 450261 337106 450327 337109
rect 427813 337104 450327 337106
rect 427813 337048 427818 337104
rect 427874 337048 450266 337104
rect 450322 337048 450327 337104
rect 427813 337046 450327 337048
rect 427813 337043 427879 337046
rect 450261 337043 450327 337046
rect 513281 336834 513347 336837
rect 509956 336832 513347 336834
rect 509956 336776 513286 336832
rect 513342 336776 513347 336832
rect 509956 336774 513347 336776
rect 513281 336771 513347 336774
rect 447409 336698 447475 336701
rect 447409 336696 450156 336698
rect 447409 336640 447414 336696
rect 447470 336640 450156 336696
rect 447409 336638 450156 336640
rect 447409 336635 447475 336638
rect 512821 336290 512887 336293
rect 509956 336288 512887 336290
rect 509956 336232 512826 336288
rect 512882 336232 512887 336288
rect 509956 336230 512887 336232
rect 512821 336227 512887 336230
rect 447133 336018 447199 336021
rect 447133 336016 450156 336018
rect 447133 335960 447138 336016
rect 447194 335960 450156 336016
rect 447133 335958 450156 335960
rect 447133 335955 447199 335958
rect 513281 335746 513347 335749
rect 509956 335744 513347 335746
rect 509956 335688 513286 335744
rect 513342 335688 513347 335744
rect 509956 335686 513347 335688
rect 513281 335683 513347 335686
rect 447225 335338 447291 335341
rect 447225 335336 450156 335338
rect 447225 335280 447230 335336
rect 447286 335280 450156 335336
rect 447225 335278 450156 335280
rect 447225 335275 447291 335278
rect 420361 335202 420427 335205
rect 513281 335202 513347 335205
rect 420361 335200 422310 335202
rect 420361 335144 420366 335200
rect 420422 335144 422310 335200
rect 420361 335142 422310 335144
rect 509956 335200 513347 335202
rect 509956 335144 513286 335200
rect 513342 335144 513347 335200
rect 509956 335142 513347 335144
rect 420361 335139 420427 335142
rect 422250 334658 422310 335142
rect 513281 335139 513347 335142
rect 447133 334658 447199 334661
rect 518014 334658 518020 334660
rect 422250 334598 431970 334658
rect 428089 334522 428155 334525
rect 428406 334522 428412 334524
rect 428089 334520 428412 334522
rect 428089 334464 428094 334520
rect 428150 334464 428412 334520
rect 428089 334462 428412 334464
rect 428089 334459 428155 334462
rect 428406 334460 428412 334462
rect 428476 334460 428482 334524
rect 431910 334522 431970 334598
rect 447133 334656 450156 334658
rect 447133 334600 447138 334656
rect 447194 334600 450156 334656
rect 447133 334598 450156 334600
rect 509956 334598 518020 334658
rect 447133 334595 447199 334598
rect 518014 334596 518020 334598
rect 518084 334596 518090 334660
rect 447910 334522 447916 334524
rect 431910 334462 447916 334522
rect 447910 334460 447916 334462
rect 447980 334460 447986 334524
rect 420453 334386 420519 334389
rect 424133 334386 424199 334389
rect 425830 334386 425836 334388
rect 420453 334384 421482 334386
rect 420453 334328 420458 334384
rect 420514 334328 421482 334384
rect 420453 334326 421482 334328
rect 420453 334323 420519 334326
rect 421422 334116 421482 334326
rect 424133 334384 425836 334386
rect 424133 334328 424138 334384
rect 424194 334328 425836 334384
rect 424133 334326 425836 334328
rect 424133 334323 424199 334326
rect 425830 334324 425836 334326
rect 425900 334386 425906 334388
rect 425900 334326 431970 334386
rect 425900 334324 425906 334326
rect 431910 334250 431970 334326
rect 450537 334250 450603 334253
rect 431910 334248 450603 334250
rect 431910 334192 450542 334248
rect 450598 334192 450603 334248
rect 431910 334190 450603 334192
rect 450537 334187 450603 334190
rect 421414 334052 421420 334116
rect 421484 334114 421490 334116
rect 449985 334114 450051 334117
rect 513281 334114 513347 334117
rect 421484 334112 450051 334114
rect 421484 334056 449990 334112
rect 450046 334056 450051 334112
rect 421484 334054 450051 334056
rect 509956 334112 513347 334114
rect 509956 334056 513286 334112
rect 513342 334056 513347 334112
rect 509956 334054 513347 334056
rect 421484 334052 421490 334054
rect 449985 334051 450051 334054
rect 513281 334051 513347 334054
rect 447225 333978 447291 333981
rect 447225 333976 450156 333978
rect 447225 333920 447230 333976
rect 447286 333920 450156 333976
rect 447225 333918 450156 333920
rect 447225 333915 447291 333918
rect 513005 333570 513071 333573
rect 509956 333568 513071 333570
rect 509956 333512 513010 333568
rect 513066 333512 513071 333568
rect 509956 333510 513071 333512
rect 513005 333507 513071 333510
rect 447133 333298 447199 333301
rect 447133 333296 450156 333298
rect 447133 333240 447138 333296
rect 447194 333240 450156 333296
rect 447133 333238 450156 333240
rect 447133 333235 447199 333238
rect 512637 333026 512703 333029
rect 509956 333024 512703 333026
rect 509956 332968 512642 333024
rect 512698 332968 512703 333024
rect 509956 332966 512703 332968
rect 512637 332963 512703 332966
rect 432873 332890 432939 332893
rect 429916 332888 432939 332890
rect 429916 332832 432878 332888
rect 432934 332832 432939 332888
rect 429916 332830 432939 332832
rect 432873 332827 432939 332830
rect 448053 332618 448119 332621
rect 448053 332616 450156 332618
rect 448053 332560 448058 332616
rect 448114 332560 450156 332616
rect 448053 332558 450156 332560
rect 448053 332555 448119 332558
rect 512637 332482 512703 332485
rect 509956 332480 512703 332482
rect -960 332196 480 332436
rect 509956 332424 512642 332480
rect 512698 332424 512703 332480
rect 509956 332422 512703 332424
rect 512637 332419 512703 332422
rect 448237 331938 448303 331941
rect 510838 331938 510844 331940
rect 448237 331936 450156 331938
rect 448237 331880 448242 331936
rect 448298 331880 450156 331936
rect 448237 331878 450156 331880
rect 509956 331878 510844 331938
rect 448237 331875 448303 331878
rect 510838 331876 510844 331878
rect 510908 331876 510914 331940
rect 515254 331394 515260 331396
rect 509956 331334 515260 331394
rect 515254 331332 515260 331334
rect 515324 331332 515330 331396
rect 447777 331258 447843 331261
rect 448329 331258 448395 331261
rect 447777 331256 450156 331258
rect 447777 331200 447782 331256
rect 447838 331200 448334 331256
rect 448390 331200 450156 331256
rect 447777 331198 450156 331200
rect 447777 331195 447843 331198
rect 448329 331195 448395 331198
rect 447961 330578 448027 330581
rect 447961 330576 450156 330578
rect 447961 330520 447966 330576
rect 448022 330520 450156 330576
rect 447961 330518 450156 330520
rect 447961 330515 448027 330518
rect 509926 330442 509986 330820
rect 509926 330382 514770 330442
rect 510061 330306 510127 330309
rect 509956 330304 510127 330306
rect 509956 330248 510066 330304
rect 510122 330248 510127 330304
rect 509956 330246 510127 330248
rect 510061 330243 510127 330246
rect 447133 329898 447199 329901
rect 448278 329898 448284 329900
rect 447133 329896 448284 329898
rect 447133 329840 447138 329896
rect 447194 329840 448284 329896
rect 447133 329838 448284 329840
rect 447133 329835 447199 329838
rect 448278 329836 448284 329838
rect 448348 329898 448354 329900
rect 514710 329898 514770 330382
rect 518934 329898 518940 329900
rect 448348 329838 450156 329898
rect 514710 329838 518940 329898
rect 448348 329836 448354 329838
rect 518934 329836 518940 329838
rect 519004 329836 519010 329900
rect 515070 329762 515076 329764
rect 509956 329702 515076 329762
rect 515070 329700 515076 329702
rect 515140 329700 515146 329764
rect 432781 329218 432847 329221
rect 429916 329216 432847 329218
rect 429916 329160 432786 329216
rect 432842 329160 432847 329216
rect 429916 329158 432847 329160
rect 432781 329155 432847 329158
rect 450126 329082 450186 329188
rect 450670 329156 450676 329220
rect 450740 329156 450746 329220
rect 513465 329218 513531 329221
rect 509956 329216 513531 329218
rect 509956 329160 513470 329216
rect 513526 329160 513531 329216
rect 509956 329158 513531 329160
rect 450678 329082 450738 329156
rect 513465 329155 513531 329158
rect 450126 329022 450738 329082
rect 449893 328946 449959 328949
rect 450126 328946 450186 329022
rect 449893 328944 450186 328946
rect 449893 328888 449898 328944
rect 449954 328888 450186 328944
rect 449893 328886 450186 328888
rect 449893 328883 449959 328886
rect 450445 328676 450511 328677
rect 450445 328674 450492 328676
rect 450404 328672 450492 328674
rect 450404 328616 450450 328672
rect 450404 328614 450492 328616
rect 450445 328612 450492 328614
rect 450556 328612 450562 328676
rect 450445 328611 450554 328612
rect 450494 328508 450554 328611
rect 509742 328405 509802 328644
rect 509693 328400 509802 328405
rect 509693 328344 509698 328400
rect 509754 328344 509802 328400
rect 509693 328342 509802 328344
rect 509693 328339 509759 328342
rect 450261 327994 450327 327997
rect 450261 327992 450370 327994
rect 450261 327936 450266 327992
rect 450322 327936 450370 327992
rect 450261 327931 450370 327936
rect 450310 327828 450370 327931
rect 509926 327725 509986 328100
rect 509877 327720 509986 327725
rect 509877 327664 509882 327720
rect 509938 327664 509986 327720
rect 509877 327662 509986 327664
rect 509877 327659 509943 327662
rect 511206 327586 511212 327588
rect 509956 327526 511212 327586
rect 511206 327524 511212 327526
rect 511276 327524 511282 327588
rect 450537 327314 450603 327317
rect 450494 327312 450603 327314
rect 450494 327256 450542 327312
rect 450598 327256 450603 327312
rect 450494 327251 450603 327256
rect 450494 327148 450554 327251
rect 514150 327042 514156 327044
rect 509956 326982 514156 327042
rect 514150 326980 514156 326982
rect 514220 326980 514226 327044
rect 449985 326634 450051 326637
rect 449985 326632 450186 326634
rect 449985 326576 449990 326632
rect 450046 326576 450186 326632
rect 449985 326574 450186 326576
rect 449985 326571 450051 326574
rect 362217 326498 362283 326501
rect 359812 326496 362283 326498
rect 359812 326440 362222 326496
rect 362278 326440 362283 326496
rect 450126 326468 450186 326574
rect 359812 326438 362283 326440
rect 362217 326435 362283 326438
rect 509926 326093 509986 326468
rect 509926 326088 510035 326093
rect 509926 326032 509974 326088
rect 510030 326032 510035 326088
rect 509926 326030 510035 326032
rect 509969 326027 510035 326030
rect 510286 325954 510292 325956
rect 509956 325894 510292 325954
rect 510286 325892 510292 325894
rect 510356 325892 510362 325956
rect 450494 325549 450554 325788
rect 432689 325546 432755 325549
rect 429916 325544 432755 325546
rect 429916 325488 432694 325544
rect 432750 325488 432755 325544
rect 429916 325486 432755 325488
rect 432689 325483 432755 325486
rect 450445 325544 450554 325549
rect 450445 325488 450450 325544
rect 450506 325488 450554 325544
rect 450445 325486 450554 325488
rect 450445 325483 450511 325486
rect 512729 325410 512795 325413
rect 509956 325408 512795 325410
rect 509956 325352 512734 325408
rect 512790 325352 512795 325408
rect 509956 325350 512795 325352
rect 512729 325347 512795 325350
rect 580165 325274 580231 325277
rect 583520 325274 584960 325364
rect 580165 325272 584960 325274
rect 580165 325216 580170 325272
rect 580226 325216 584960 325272
rect 580165 325214 584960 325216
rect 580165 325211 580231 325214
rect 583520 325124 584960 325214
rect 450310 324869 450370 325108
rect 450310 324864 450419 324869
rect 514886 324866 514892 324868
rect 450310 324808 450358 324864
rect 450414 324808 450419 324864
rect 450310 324806 450419 324808
rect 509956 324806 514892 324866
rect 450353 324803 450419 324806
rect 514886 324804 514892 324806
rect 514956 324804 514962 324868
rect 450077 324594 450143 324597
rect 450077 324592 450738 324594
rect 450077 324536 450082 324592
rect 450138 324536 450738 324592
rect 450077 324534 450738 324536
rect 450077 324531 450143 324534
rect 450678 324189 450738 324534
rect 511022 324322 511028 324324
rect 509956 324262 511028 324322
rect 511022 324260 511028 324262
rect 511092 324260 511098 324324
rect 450629 324184 450738 324189
rect 450629 324128 450634 324184
rect 450690 324128 450738 324184
rect 450629 324126 450738 324128
rect 450629 324123 450695 324126
rect 510470 323778 510476 323780
rect 509956 323718 510476 323778
rect 510470 323716 510476 323718
rect 510540 323716 510546 323780
rect 509374 322965 509434 323204
rect 509325 322960 509434 322965
rect 509325 322904 509330 322960
rect 509386 322904 509434 322960
rect 509325 322902 509434 322904
rect 509325 322899 509391 322902
rect 445569 322826 445635 322829
rect 445569 322824 482938 322826
rect 445569 322768 445574 322824
rect 445630 322768 482938 322824
rect 445569 322766 482938 322768
rect 445569 322763 445635 322766
rect 445201 322690 445267 322693
rect 482645 322690 482711 322693
rect 445201 322688 482711 322690
rect 445201 322632 445206 322688
rect 445262 322632 482650 322688
rect 482706 322632 482711 322688
rect 445201 322630 482711 322632
rect 482878 322690 482938 322766
rect 483749 322690 483815 322693
rect 482878 322688 483815 322690
rect 482878 322632 483754 322688
rect 483810 322632 483815 322688
rect 482878 322630 483815 322632
rect 445201 322627 445267 322630
rect 482645 322627 482711 322630
rect 483749 322627 483815 322630
rect 507117 322690 507183 322693
rect 510286 322690 510292 322692
rect 507117 322688 510292 322690
rect 507117 322632 507122 322688
rect 507178 322632 510292 322688
rect 507117 322630 510292 322632
rect 507117 322627 507183 322630
rect 510286 322628 510292 322630
rect 510356 322628 510362 322692
rect 446305 322554 446371 322557
rect 473537 322554 473603 322557
rect 446305 322552 473603 322554
rect 446305 322496 446310 322552
rect 446366 322496 473542 322552
rect 473598 322496 473603 322552
rect 446305 322494 473603 322496
rect 446305 322491 446371 322494
rect 473537 322491 473603 322494
rect 468753 322418 468819 322421
rect 470133 322418 470199 322421
rect 468753 322416 470199 322418
rect 468753 322360 468758 322416
rect 468814 322360 470138 322416
rect 470194 322360 470199 322416
rect 468753 322358 470199 322360
rect 468753 322355 468819 322358
rect 470133 322355 470199 322358
rect 432873 321874 432939 321877
rect 429916 321872 432939 321874
rect 429916 321816 432878 321872
rect 432934 321816 432939 321872
rect 429916 321814 432939 321816
rect 432873 321811 432939 321814
rect 449157 321466 449223 321469
rect 462221 321466 462287 321469
rect 449157 321464 462287 321466
rect 449157 321408 449162 321464
rect 449218 321408 462226 321464
rect 462282 321408 462287 321464
rect 449157 321406 462287 321408
rect 449157 321403 449223 321406
rect 462221 321403 462287 321406
rect 507485 321466 507551 321469
rect 511206 321466 511212 321468
rect 507485 321464 511212 321466
rect 507485 321408 507490 321464
rect 507546 321408 511212 321464
rect 507485 321406 511212 321408
rect 507485 321403 507551 321406
rect 511206 321404 511212 321406
rect 511276 321404 511282 321468
rect 444230 321268 444236 321332
rect 444300 321330 444306 321332
rect 461117 321330 461183 321333
rect 444300 321328 461183 321330
rect 444300 321272 461122 321328
rect 461178 321272 461183 321328
rect 444300 321270 461183 321272
rect 444300 321268 444306 321270
rect 461117 321267 461183 321270
rect 470501 321330 470567 321333
rect 530526 321330 530532 321332
rect 470501 321328 530532 321330
rect 470501 321272 470506 321328
rect 470562 321272 530532 321328
rect 470501 321270 530532 321272
rect 470501 321267 470567 321270
rect 530526 321268 530532 321270
rect 530596 321268 530602 321332
rect 447726 321132 447732 321196
rect 447796 321194 447802 321196
rect 462497 321194 462563 321197
rect 447796 321192 462563 321194
rect 447796 321136 462502 321192
rect 462558 321136 462563 321192
rect 447796 321134 462563 321136
rect 447796 321132 447802 321134
rect 462497 321131 462563 321134
rect 443494 320996 443500 321060
rect 443564 321058 443570 321060
rect 461945 321058 462011 321061
rect 443564 321056 462011 321058
rect 443564 321000 461950 321056
rect 462006 321000 462011 321056
rect 443564 320998 462011 321000
rect 443564 320996 443570 320998
rect 461945 320995 462011 320998
rect 458766 320724 458772 320788
rect 458836 320786 458842 320788
rect 509325 320786 509391 320789
rect 458836 320784 509391 320786
rect 458836 320728 509330 320784
rect 509386 320728 509391 320784
rect 458836 320726 509391 320728
rect 458836 320724 458842 320726
rect 509325 320723 509391 320726
rect 460013 320650 460079 320653
rect 558126 320650 558132 320652
rect 460013 320648 558132 320650
rect 460013 320592 460018 320648
rect 460074 320592 558132 320648
rect 460013 320590 558132 320592
rect 460013 320587 460079 320590
rect 558126 320588 558132 320590
rect 558196 320588 558202 320652
rect 444046 320044 444052 320108
rect 444116 320106 444122 320108
rect 460289 320106 460355 320109
rect 444116 320104 460355 320106
rect 444116 320048 460294 320104
rect 460350 320048 460355 320104
rect 444116 320046 460355 320048
rect 444116 320044 444122 320046
rect 460289 320043 460355 320046
rect 446254 319908 446260 319972
rect 446324 319970 446330 319972
rect 472709 319970 472775 319973
rect 446324 319968 472775 319970
rect 446324 319912 472714 319968
rect 472770 319912 472775 319968
rect 446324 319910 472775 319912
rect 446324 319908 446330 319910
rect 472709 319907 472775 319910
rect 447910 319772 447916 319836
rect 447980 319834 447986 319836
rect 474089 319834 474155 319837
rect 447980 319832 474155 319834
rect 447980 319776 474094 319832
rect 474150 319776 474155 319832
rect 447980 319774 474155 319776
rect 447980 319772 447986 319774
rect 474089 319771 474155 319774
rect 446765 319698 446831 319701
rect 472985 319698 473051 319701
rect 446765 319696 473051 319698
rect 446765 319640 446770 319696
rect 446826 319640 472990 319696
rect 473046 319640 473051 319696
rect 446765 319638 473051 319640
rect 446765 319635 446831 319638
rect 472985 319635 473051 319638
rect 449341 319562 449407 319565
rect 482921 319562 482987 319565
rect 449341 319560 482987 319562
rect 449341 319504 449346 319560
rect 449402 319504 482926 319560
rect 482982 319504 482987 319560
rect 449341 319502 482987 319504
rect 449341 319499 449407 319502
rect 482921 319499 482987 319502
rect 456149 319426 456215 319429
rect 486233 319426 486299 319429
rect 456149 319424 486299 319426
rect -960 319290 480 319380
rect 456149 319368 456154 319424
rect 456210 319368 486238 319424
rect 486294 319368 486299 319424
rect 456149 319366 486299 319368
rect 456149 319363 456215 319366
rect 486233 319363 486299 319366
rect 3969 319290 4035 319293
rect -960 319288 4035 319290
rect -960 319232 3974 319288
rect 4030 319232 4035 319288
rect -960 319230 4035 319232
rect -960 319140 480 319230
rect 3969 319227 4035 319230
rect 432781 318202 432847 318205
rect 429916 318200 432847 318202
rect 429916 318144 432786 318200
rect 432842 318144 432847 318200
rect 429916 318142 432847 318144
rect 432781 318139 432847 318142
rect 454677 317250 454743 317253
rect 510153 317250 510219 317253
rect 454677 317248 510219 317250
rect 454677 317192 454682 317248
rect 454738 317192 510158 317248
rect 510214 317192 510219 317248
rect 454677 317190 510219 317192
rect 454677 317187 454743 317190
rect 510153 317187 510219 317190
rect 450537 317114 450603 317117
rect 512545 317114 512611 317117
rect 450537 317112 512611 317114
rect 450537 317056 450542 317112
rect 450598 317056 512550 317112
rect 512606 317056 512611 317112
rect 450537 317054 512611 317056
rect 450537 317051 450603 317054
rect 512545 317051 512611 317054
rect 450905 316978 450971 316981
rect 514109 316978 514175 316981
rect 450905 316976 514175 316978
rect 450905 316920 450910 316976
rect 450966 316920 514114 316976
rect 514170 316920 514175 316976
rect 450905 316918 514175 316920
rect 450905 316915 450971 316918
rect 514109 316915 514175 316918
rect 451089 316842 451155 316845
rect 515121 316842 515187 316845
rect 451089 316840 515187 316842
rect 451089 316784 451094 316840
rect 451150 316784 515126 316840
rect 515182 316784 515187 316840
rect 451089 316782 515187 316784
rect 451089 316779 451155 316782
rect 515121 316779 515187 316782
rect 450721 316706 450787 316709
rect 515070 316706 515076 316708
rect 450721 316704 515076 316706
rect 450721 316648 450726 316704
rect 450782 316648 515076 316704
rect 450721 316646 515076 316648
rect 450721 316643 450787 316646
rect 515070 316644 515076 316646
rect 515140 316644 515146 316708
rect 361757 315482 361823 315485
rect 359812 315480 361823 315482
rect 359812 315424 361762 315480
rect 361818 315424 361823 315480
rect 359812 315422 361823 315424
rect 361757 315419 361823 315422
rect 432689 314530 432755 314533
rect 429916 314528 432755 314530
rect 429916 314472 432694 314528
rect 432750 314472 432755 314528
rect 429916 314470 432755 314472
rect 432689 314467 432755 314470
rect 580165 312082 580231 312085
rect 583520 312082 584960 312172
rect 580165 312080 584960 312082
rect 580165 312024 580170 312080
rect 580226 312024 584960 312080
rect 580165 312022 584960 312024
rect 580165 312019 580231 312022
rect 583520 311932 584960 312022
rect 497181 311130 497247 311133
rect 542670 311130 542676 311132
rect 497181 311128 542676 311130
rect 497181 311072 497186 311128
rect 497242 311072 542676 311128
rect 497181 311070 542676 311072
rect 497181 311067 497247 311070
rect 542670 311068 542676 311070
rect 542740 311068 542746 311132
rect 432045 310858 432111 310861
rect 429916 310856 432111 310858
rect 429916 310800 432050 310856
rect 432106 310800 432111 310856
rect 429916 310798 432111 310800
rect 432045 310795 432111 310798
rect 433149 307186 433215 307189
rect 429916 307184 433215 307186
rect 429916 307128 433154 307184
rect 433210 307128 433215 307184
rect 429916 307126 433215 307128
rect 433149 307123 433215 307126
rect -960 306234 480 306324
rect 3693 306234 3759 306237
rect -960 306232 3759 306234
rect -960 306176 3698 306232
rect 3754 306176 3759 306232
rect -960 306174 3759 306176
rect -960 306084 480 306174
rect 3693 306171 3759 306174
rect 406377 305962 406443 305965
rect 510470 305962 510476 305964
rect 406377 305960 510476 305962
rect 406377 305904 406382 305960
rect 406438 305904 510476 305960
rect 406377 305902 510476 305904
rect 406377 305899 406443 305902
rect 510470 305900 510476 305902
rect 510540 305900 510546 305964
rect 406745 305826 406811 305829
rect 510654 305826 510660 305828
rect 406745 305824 510660 305826
rect 406745 305768 406750 305824
rect 406806 305768 510660 305824
rect 406745 305766 510660 305768
rect 406745 305763 406811 305766
rect 510654 305764 510660 305766
rect 510724 305764 510730 305828
rect 406561 305690 406627 305693
rect 511022 305690 511028 305692
rect 406561 305688 511028 305690
rect 406561 305632 406566 305688
rect 406622 305632 511028 305688
rect 406561 305630 511028 305632
rect 406561 305627 406627 305630
rect 511022 305628 511028 305630
rect 511092 305628 511098 305692
rect 361757 304466 361823 304469
rect 359812 304464 361823 304466
rect 359812 304408 361762 304464
rect 361818 304408 361823 304464
rect 359812 304406 361823 304408
rect 361757 304403 361823 304406
rect 401225 302834 401291 302837
rect 509877 302834 509943 302837
rect 401225 302832 509943 302834
rect 401225 302776 401230 302832
rect 401286 302776 509882 302832
rect 509938 302776 509943 302832
rect 401225 302774 509943 302776
rect 401225 302771 401291 302774
rect 509877 302771 509943 302774
rect 395521 300658 395587 300661
rect 515254 300658 515260 300660
rect 395521 300656 515260 300658
rect 395521 300600 395526 300656
rect 395582 300600 515260 300656
rect 395521 300598 515260 300600
rect 395521 300595 395587 300598
rect 515254 300596 515260 300598
rect 515324 300596 515330 300660
rect 392577 300522 392643 300525
rect 514150 300522 514156 300524
rect 392577 300520 514156 300522
rect 392577 300464 392582 300520
rect 392638 300464 514156 300520
rect 392577 300462 514156 300464
rect 392577 300459 392643 300462
rect 514150 300460 514156 300462
rect 514220 300460 514226 300524
rect 392761 300386 392827 300389
rect 514886 300386 514892 300388
rect 392761 300384 514892 300386
rect 392761 300328 392766 300384
rect 392822 300328 514892 300384
rect 392761 300326 514892 300328
rect 392761 300323 392827 300326
rect 514886 300324 514892 300326
rect 514956 300324 514962 300388
rect 395337 300250 395403 300253
rect 518014 300250 518020 300252
rect 395337 300248 518020 300250
rect 395337 300192 395342 300248
rect 395398 300192 518020 300248
rect 395337 300190 518020 300192
rect 395337 300187 395403 300190
rect 518014 300188 518020 300190
rect 518084 300188 518090 300252
rect 392945 300114 393011 300117
rect 517830 300114 517836 300116
rect 392945 300112 517836 300114
rect 392945 300056 392950 300112
rect 393006 300056 517836 300112
rect 392945 300054 517836 300056
rect 392945 300051 393011 300054
rect 517830 300052 517836 300054
rect 517900 300052 517906 300116
rect 580165 298754 580231 298757
rect 583520 298754 584960 298844
rect 580165 298752 584960 298754
rect 580165 298696 580170 298752
rect 580226 298696 584960 298752
rect 580165 298694 584960 298696
rect 580165 298691 580231 298694
rect 583520 298604 584960 298694
rect 378961 294538 379027 294541
rect 510838 294538 510844 294540
rect 378961 294536 510844 294538
rect 378961 294480 378966 294536
rect 379022 294480 510844 294536
rect 378961 294478 510844 294480
rect 378961 294475 379027 294478
rect 510838 294476 510844 294478
rect 510908 294476 510914 294540
rect 361757 293450 361823 293453
rect 359812 293448 361823 293450
rect 359812 293392 361762 293448
rect 361818 293392 361823 293448
rect 359812 293390 361823 293392
rect 361757 293387 361823 293390
rect -960 293178 480 293268
rect 3601 293178 3667 293181
rect -960 293176 3667 293178
rect -960 293120 3606 293176
rect 3662 293120 3667 293176
rect -960 293118 3667 293120
rect -960 293028 480 293118
rect 3601 293115 3667 293118
rect 368105 291818 368171 291821
rect 518934 291818 518940 291820
rect 368105 291816 518940 291818
rect 368105 291760 368110 291816
rect 368166 291760 518940 291816
rect 368105 291758 518940 291760
rect 368105 291755 368171 291758
rect 518934 291756 518940 291758
rect 519004 291756 519010 291820
rect 583520 285276 584960 285516
rect 361757 282434 361823 282437
rect 359812 282432 361823 282434
rect 359812 282376 361762 282432
rect 361818 282376 361823 282432
rect 359812 282374 361823 282376
rect 361757 282371 361823 282374
rect -960 279972 480 280212
rect 502241 278082 502307 278085
rect 538254 278082 538260 278084
rect 502241 278080 538260 278082
rect 502241 278024 502246 278080
rect 502302 278024 538260 278080
rect 502241 278022 538260 278024
rect 502241 278019 502307 278022
rect 538254 278020 538260 278022
rect 538324 278020 538330 278084
rect 579889 272234 579955 272237
rect 583520 272234 584960 272324
rect 579889 272232 584960 272234
rect 579889 272176 579894 272232
rect 579950 272176 584960 272232
rect 579889 272174 584960 272176
rect 579889 272171 579955 272174
rect 583520 272084 584960 272174
rect 361757 271418 361823 271421
rect 359812 271416 361823 271418
rect 359812 271360 361762 271416
rect 361818 271360 361823 271416
rect 359812 271358 361823 271360
rect 361757 271355 361823 271358
rect -960 267202 480 267292
rect 3509 267202 3575 267205
rect -960 267200 3575 267202
rect -960 267144 3514 267200
rect 3570 267144 3575 267200
rect -960 267142 3575 267144
rect -960 267052 480 267142
rect 3509 267139 3575 267142
rect 456793 262714 456859 262717
rect 456793 262712 460092 262714
rect 456793 262656 456798 262712
rect 456854 262656 460092 262712
rect 456793 262654 460092 262656
rect 456793 262651 456859 262654
rect 530117 261082 530183 261085
rect 529828 261080 530183 261082
rect 529828 261024 530122 261080
rect 530178 261024 530183 261080
rect 529828 261022 530183 261024
rect 530117 261019 530183 261022
rect 361757 260402 361823 260405
rect 359812 260400 361823 260402
rect 359812 260344 361762 260400
rect 361818 260344 361823 260400
rect 359812 260342 361823 260344
rect 361757 260339 361823 260342
rect 580349 258906 580415 258909
rect 583520 258906 584960 258996
rect 580349 258904 584960 258906
rect 580349 258848 580354 258904
rect 580410 258848 584960 258904
rect 580349 258846 584960 258848
rect 580349 258843 580415 258846
rect 583520 258756 584960 258846
rect -960 254146 480 254236
rect 3417 254146 3483 254149
rect -960 254144 3483 254146
rect -960 254088 3422 254144
rect 3478 254088 3483 254144
rect -960 254086 3483 254088
rect -960 253996 480 254086
rect 3417 254083 3483 254086
rect 361757 249386 361823 249389
rect 359812 249384 361823 249386
rect 359812 249328 361762 249384
rect 361818 249328 361823 249384
rect 359812 249326 361823 249328
rect 361757 249323 361823 249326
rect 457805 248842 457871 248845
rect 457805 248840 460092 248842
rect 457805 248784 457810 248840
rect 457866 248784 460092 248840
rect 457805 248782 460092 248784
rect 457805 248779 457871 248782
rect 580165 245578 580231 245581
rect 583520 245578 584960 245668
rect 580165 245576 584960 245578
rect 580165 245520 580170 245576
rect 580226 245520 584960 245576
rect 580165 245518 584960 245520
rect 580165 245515 580231 245518
rect 583520 245428 584960 245518
rect 531313 243674 531379 243677
rect 529828 243672 531379 243674
rect 529828 243616 531318 243672
rect 531374 243616 531379 243672
rect 529828 243614 531379 243616
rect 531313 243611 531379 243614
rect -960 241090 480 241180
rect 3785 241090 3851 241093
rect -960 241088 3851 241090
rect -960 241032 3790 241088
rect 3846 241032 3851 241088
rect -960 241030 3851 241032
rect -960 240940 480 241030
rect 3785 241027 3851 241030
rect 361757 238370 361823 238373
rect 359812 238368 361823 238370
rect 359812 238312 361762 238368
rect 361818 238312 361823 238368
rect 359812 238310 361823 238312
rect 361757 238307 361823 238310
rect 457989 234970 458055 234973
rect 457989 234968 460092 234970
rect 457989 234912 457994 234968
rect 458050 234912 460092 234968
rect 457989 234910 460092 234912
rect 457989 234907 458055 234910
rect 580165 232386 580231 232389
rect 583520 232386 584960 232476
rect 580165 232384 584960 232386
rect 580165 232328 580170 232384
rect 580226 232328 584960 232384
rect 580165 232326 584960 232328
rect 580165 232323 580231 232326
rect 583520 232236 584960 232326
rect -960 227884 480 228124
rect 361757 227354 361823 227357
rect 359812 227352 361823 227354
rect 359812 227296 361762 227352
rect 361818 227296 361823 227352
rect 359812 227294 361823 227296
rect 361757 227291 361823 227294
rect 530117 226266 530183 226269
rect 529828 226264 530183 226266
rect 529828 226208 530122 226264
rect 530178 226208 530183 226264
rect 529828 226206 530183 226208
rect 530117 226203 530183 226206
rect 457989 221098 458055 221101
rect 457989 221096 460092 221098
rect 457989 221040 457994 221096
rect 458050 221040 460092 221096
rect 457989 221038 460092 221040
rect 457989 221035 458055 221038
rect 580257 219058 580323 219061
rect 583520 219058 584960 219148
rect 580257 219056 584960 219058
rect 580257 219000 580262 219056
rect 580318 219000 584960 219056
rect 580257 218998 584960 219000
rect 580257 218995 580323 218998
rect 583520 218908 584960 218998
rect 361573 216338 361639 216341
rect 359812 216336 361639 216338
rect 359812 216280 361578 216336
rect 361634 216280 361639 216336
rect 359812 216278 361639 216280
rect 361573 216275 361639 216278
rect -960 214978 480 215068
rect 3877 214978 3943 214981
rect -960 214976 3943 214978
rect -960 214920 3882 214976
rect 3938 214920 3943 214976
rect -960 214918 3943 214920
rect -960 214828 480 214918
rect 3877 214915 3943 214918
rect 529933 209266 529999 209269
rect 529798 209264 529999 209266
rect 529798 209208 529938 209264
rect 529994 209208 529999 209264
rect 529798 209206 529999 209208
rect 529798 208828 529858 209206
rect 529933 209203 529999 209206
rect 457713 207226 457779 207229
rect 458081 207226 458147 207229
rect 457713 207224 460092 207226
rect 457713 207168 457718 207224
rect 457774 207168 458086 207224
rect 458142 207168 460092 207224
rect 457713 207166 460092 207168
rect 457713 207163 457779 207166
rect 458081 207163 458147 207166
rect 579797 205730 579863 205733
rect 583520 205730 584960 205820
rect 579797 205728 584960 205730
rect 579797 205672 579802 205728
rect 579858 205672 584960 205728
rect 579797 205670 584960 205672
rect 579797 205667 579863 205670
rect 583520 205580 584960 205670
rect 361757 205322 361823 205325
rect 359812 205320 361823 205322
rect 359812 205264 361762 205320
rect 361818 205264 361823 205320
rect 359812 205262 361823 205264
rect 361757 205259 361823 205262
rect -960 201922 480 202012
rect 3969 201922 4035 201925
rect -960 201920 4035 201922
rect -960 201864 3974 201920
rect 4030 201864 4035 201920
rect -960 201862 4035 201864
rect -960 201772 480 201862
rect 3969 201859 4035 201862
rect 361665 194306 361731 194309
rect 359812 194304 361731 194306
rect 359812 194248 361670 194304
rect 361726 194248 361731 194304
rect 359812 194246 361731 194248
rect 361665 194243 361731 194246
rect 580165 192538 580231 192541
rect 583520 192538 584960 192628
rect 580165 192536 584960 192538
rect 580165 192480 580170 192536
rect 580226 192480 584960 192536
rect 580165 192478 584960 192480
rect 580165 192475 580231 192478
rect 583520 192388 584960 192478
rect -960 188866 480 188956
rect 4061 188866 4127 188869
rect -960 188864 4127 188866
rect -960 188808 4066 188864
rect 4122 188808 4127 188864
rect -960 188806 4127 188808
rect -960 188716 480 188806
rect 4061 188803 4127 188806
rect 361665 183290 361731 183293
rect 359812 183288 361731 183290
rect 359812 183232 361670 183288
rect 361726 183232 361731 183288
rect 359812 183230 361731 183232
rect 361665 183227 361731 183230
rect 580165 179210 580231 179213
rect 583520 179210 584960 179300
rect 580165 179208 584960 179210
rect 580165 179152 580170 179208
rect 580226 179152 584960 179208
rect 580165 179150 584960 179152
rect 580165 179147 580231 179150
rect 583520 179060 584960 179150
rect -960 175796 480 176036
rect 361665 172274 361731 172277
rect 359812 172272 361731 172274
rect 359812 172216 361670 172272
rect 361726 172216 361731 172272
rect 359812 172214 361731 172216
rect 361665 172211 361731 172214
rect 580165 165882 580231 165885
rect 583520 165882 584960 165972
rect 580165 165880 584960 165882
rect 580165 165824 580170 165880
rect 580226 165824 584960 165880
rect 580165 165822 584960 165824
rect 580165 165819 580231 165822
rect 583520 165732 584960 165822
rect -960 162890 480 162980
rect 3325 162890 3391 162893
rect -960 162888 3391 162890
rect -960 162832 3330 162888
rect 3386 162832 3391 162888
rect -960 162830 3391 162832
rect -960 162740 480 162830
rect 3325 162827 3391 162830
rect 421414 162692 421420 162756
rect 421484 162754 421490 162756
rect 422017 162754 422083 162757
rect 421484 162752 422083 162754
rect 421484 162696 422022 162752
rect 422078 162696 422083 162752
rect 421484 162694 422083 162696
rect 421484 162692 421490 162694
rect 422017 162691 422083 162694
rect 425830 162692 425836 162756
rect 425900 162754 425906 162756
rect 426341 162754 426407 162757
rect 425900 162752 426407 162754
rect 425900 162696 426346 162752
rect 426402 162696 426407 162752
rect 425900 162694 426407 162696
rect 425900 162692 425906 162694
rect 426341 162691 426407 162694
rect 428406 162692 428412 162756
rect 428476 162754 428482 162756
rect 428641 162754 428707 162757
rect 428476 162752 428707 162754
rect 428476 162696 428646 162752
rect 428702 162696 428707 162752
rect 428476 162694 428707 162696
rect 428476 162692 428482 162694
rect 428641 162691 428707 162694
rect 361757 161258 361823 161261
rect 359812 161256 361823 161258
rect 359812 161200 361762 161256
rect 361818 161200 361823 161256
rect 359812 161198 361823 161200
rect 361757 161195 361823 161198
rect 452561 158266 452627 158269
rect 449788 158264 452627 158266
rect 449788 158208 452566 158264
rect 452622 158208 452627 158264
rect 449788 158206 452627 158208
rect 452561 158203 452627 158206
rect 451917 156906 451983 156909
rect 449788 156904 451983 156906
rect 449788 156848 451922 156904
rect 451978 156848 451983 156904
rect 449788 156846 451983 156848
rect 451917 156843 451983 156846
rect 452561 155546 452627 155549
rect 449788 155544 452627 155546
rect 449788 155488 452566 155544
rect 452622 155488 452627 155544
rect 449788 155486 452627 155488
rect 452561 155483 452627 155486
rect 452377 154186 452443 154189
rect 449788 154184 452443 154186
rect 449788 154128 452382 154184
rect 452438 154128 452443 154184
rect 449788 154126 452443 154128
rect 452377 154123 452443 154126
rect 452285 152826 452351 152829
rect 449788 152824 452351 152826
rect 449788 152768 452290 152824
rect 452346 152768 452351 152824
rect 449788 152766 452351 152768
rect 452285 152763 452351 152766
rect 580165 152690 580231 152693
rect 583520 152690 584960 152780
rect 580165 152688 584960 152690
rect 580165 152632 580170 152688
rect 580226 152632 584960 152688
rect 580165 152630 584960 152632
rect 580165 152627 580231 152630
rect 583520 152540 584960 152630
rect 452009 151466 452075 151469
rect 449788 151464 452075 151466
rect 449788 151408 452014 151464
rect 452070 151408 452075 151464
rect 449788 151406 452075 151408
rect 452009 151403 452075 151406
rect 361757 150242 361823 150245
rect 359812 150240 361823 150242
rect 359812 150184 361762 150240
rect 361818 150184 361823 150240
rect 359812 150182 361823 150184
rect 361757 150179 361823 150182
rect 451549 150106 451615 150109
rect 449788 150104 451615 150106
rect 449788 150048 451554 150104
rect 451610 150048 451615 150104
rect 449788 150046 451615 150048
rect 451549 150043 451615 150046
rect -960 149834 480 149924
rect 3233 149834 3299 149837
rect -960 149832 3299 149834
rect -960 149776 3238 149832
rect 3294 149776 3299 149832
rect -960 149774 3299 149776
rect -960 149684 480 149774
rect 3233 149771 3299 149774
rect 451733 148746 451799 148749
rect 449788 148744 451799 148746
rect 449788 148688 451738 148744
rect 451794 148688 451799 148744
rect 449788 148686 451799 148688
rect 451733 148683 451799 148686
rect 451733 147386 451799 147389
rect 449788 147384 451799 147386
rect 449788 147328 451738 147384
rect 451794 147328 451799 147384
rect 449788 147326 451799 147328
rect 451733 147323 451799 147326
rect 452561 146026 452627 146029
rect 449788 146024 452627 146026
rect 449788 145968 452566 146024
rect 452622 145968 452627 146024
rect 449788 145966 452627 145968
rect 452561 145963 452627 145966
rect 452561 144666 452627 144669
rect 449788 144664 452627 144666
rect 449788 144608 452566 144664
rect 452622 144608 452627 144664
rect 449788 144606 452627 144608
rect 452561 144603 452627 144606
rect 452561 143306 452627 143309
rect 449788 143304 452627 143306
rect 449788 143248 452566 143304
rect 452622 143248 452627 143304
rect 449788 143246 452627 143248
rect 452561 143243 452627 143246
rect 452561 141946 452627 141949
rect 449788 141944 452627 141946
rect 449788 141888 452566 141944
rect 452622 141888 452627 141944
rect 449788 141886 452627 141888
rect 452561 141883 452627 141886
rect 452561 140586 452627 140589
rect 449788 140584 452627 140586
rect 449788 140528 452566 140584
rect 452622 140528 452627 140584
rect 449788 140526 452627 140528
rect 452561 140523 452627 140526
rect 580165 139362 580231 139365
rect 583520 139362 584960 139452
rect 580165 139360 584960 139362
rect 580165 139304 580170 139360
rect 580226 139304 584960 139360
rect 580165 139302 584960 139304
rect 580165 139299 580231 139302
rect 361757 139226 361823 139229
rect 451549 139226 451615 139229
rect 359812 139224 361823 139226
rect 359812 139168 361762 139224
rect 361818 139168 361823 139224
rect 359812 139166 361823 139168
rect 449788 139224 451615 139226
rect 449788 139168 451554 139224
rect 451610 139168 451615 139224
rect 583520 139212 584960 139302
rect 449788 139166 451615 139168
rect 361757 139163 361823 139166
rect 451549 139163 451615 139166
rect 538949 138002 539015 138005
rect 538949 138000 539610 138002
rect 538949 137944 538954 138000
rect 539010 137944 539610 138000
rect 538949 137942 539610 137944
rect 538949 137939 539015 137942
rect 452561 137866 452627 137869
rect 449788 137864 452627 137866
rect 449788 137808 452566 137864
rect 452622 137808 452627 137864
rect 449788 137806 452627 137808
rect 452561 137803 452627 137806
rect 539550 137428 539610 137942
rect -960 136778 480 136868
rect 2814 136778 2820 136780
rect -960 136718 2820 136778
rect -960 136628 480 136718
rect 2814 136716 2820 136718
rect 2884 136716 2890 136780
rect 452561 136506 452627 136509
rect 449788 136504 452627 136506
rect 449788 136448 452566 136504
rect 452622 136448 452627 136504
rect 449788 136446 452627 136448
rect 452561 136443 452627 136446
rect 539317 135690 539383 135693
rect 539317 135688 539426 135690
rect 539317 135632 539322 135688
rect 539378 135632 539426 135688
rect 539317 135627 539426 135632
rect 539366 135388 539426 135627
rect 452561 135146 452627 135149
rect 449788 135144 452627 135146
rect 449788 135088 452566 135144
rect 452622 135088 452627 135144
rect 449788 135086 452627 135088
rect 452561 135083 452627 135086
rect 452561 133786 452627 133789
rect 449788 133784 452627 133786
rect 449788 133728 452566 133784
rect 452622 133728 452627 133784
rect 449788 133726 452627 133728
rect 452561 133723 452627 133726
rect 543181 133378 543247 133381
rect 539948 133376 543247 133378
rect 539948 133320 543186 133376
rect 543242 133320 543247 133376
rect 539948 133318 543247 133320
rect 543181 133315 543247 133318
rect 452469 132426 452535 132429
rect 449788 132424 452535 132426
rect 449788 132368 452474 132424
rect 452530 132368 452535 132424
rect 449788 132366 452535 132368
rect 452469 132363 452535 132366
rect 543089 131338 543155 131341
rect 539948 131336 543155 131338
rect 539948 131280 543094 131336
rect 543150 131280 543155 131336
rect 539948 131278 543155 131280
rect 543089 131275 543155 131278
rect 452561 131066 452627 131069
rect 449788 131064 452627 131066
rect 449788 131008 452566 131064
rect 452622 131008 452627 131064
rect 449788 131006 452627 131008
rect 452561 131003 452627 131006
rect 452193 129706 452259 129709
rect 449788 129704 452259 129706
rect 449788 129648 452198 129704
rect 452254 129648 452259 129704
rect 449788 129646 452259 129648
rect 452193 129643 452259 129646
rect 542629 129298 542695 129301
rect 539948 129296 542695 129298
rect 539948 129240 542634 129296
rect 542690 129240 542695 129296
rect 539948 129238 542695 129240
rect 542629 129235 542695 129238
rect 452101 128346 452167 128349
rect 449788 128344 452167 128346
rect 449788 128288 452106 128344
rect 452162 128288 452167 128344
rect 449788 128286 452167 128288
rect 452101 128283 452167 128286
rect 361573 128210 361639 128213
rect 359812 128208 361639 128210
rect 359812 128152 361578 128208
rect 361634 128152 361639 128208
rect 359812 128150 361639 128152
rect 361573 128147 361639 128150
rect 539358 127196 539364 127260
rect 539428 127196 539434 127260
rect 452561 126986 452627 126989
rect 449788 126984 452627 126986
rect 449788 126928 452566 126984
rect 452622 126928 452627 126984
rect 449788 126926 452627 126928
rect 452561 126923 452627 126926
rect 580165 126034 580231 126037
rect 583520 126034 584960 126124
rect 580165 126032 584960 126034
rect 580165 125976 580170 126032
rect 580226 125976 584960 126032
rect 580165 125974 584960 125976
rect 580165 125971 580231 125974
rect 583520 125884 584960 125974
rect 451917 125626 451983 125629
rect 449788 125624 451983 125626
rect 449788 125568 451922 125624
rect 451978 125568 451983 125624
rect 449788 125566 451983 125568
rect 451917 125563 451983 125566
rect 542537 125218 542603 125221
rect 539948 125216 542603 125218
rect 539948 125160 542542 125216
rect 542598 125160 542603 125216
rect 539948 125158 542603 125160
rect 542537 125155 542603 125158
rect 451917 124266 451983 124269
rect 449788 124264 451983 124266
rect 449788 124208 451922 124264
rect 451978 124208 451983 124264
rect 449788 124206 451983 124208
rect 451917 124203 451983 124206
rect -960 123572 480 123812
rect 542997 123178 543063 123181
rect 539948 123176 543063 123178
rect 539948 123120 543002 123176
rect 543058 123120 543063 123176
rect 539948 123118 543063 123120
rect 542997 123115 543063 123118
rect 451917 122906 451983 122909
rect 449788 122904 451983 122906
rect 449788 122848 451922 122904
rect 451978 122848 451983 122904
rect 449788 122846 451983 122848
rect 451917 122843 451983 122846
rect 451733 121546 451799 121549
rect 449788 121544 451799 121546
rect 449788 121488 451738 121544
rect 451794 121488 451799 121544
rect 449788 121486 451799 121488
rect 451733 121483 451799 121486
rect 541065 121138 541131 121141
rect 539948 121136 541131 121138
rect 539948 121080 541070 121136
rect 541126 121080 541131 121136
rect 539948 121078 541131 121080
rect 541065 121075 541131 121078
rect 539869 119642 539935 119645
rect 539869 119640 539978 119642
rect 539869 119584 539874 119640
rect 539930 119584 539978 119640
rect 539869 119579 539978 119584
rect 539918 119068 539978 119579
rect 361573 117194 361639 117197
rect 359812 117192 361639 117194
rect 359812 117136 361578 117192
rect 361634 117136 361639 117192
rect 359812 117134 361639 117136
rect 361573 117131 361639 117134
rect 541433 117058 541499 117061
rect 539948 117056 541499 117058
rect 539948 117000 541438 117056
rect 541494 117000 541499 117056
rect 539948 116998 541499 117000
rect 541433 116995 541499 116998
rect 540237 115018 540303 115021
rect 539948 115016 540303 115018
rect 539948 114960 540242 115016
rect 540298 114960 540303 115016
rect 539948 114958 540303 114960
rect 540237 114955 540303 114958
rect 539777 113250 539843 113253
rect 539734 113248 539843 113250
rect 539734 113192 539782 113248
rect 539838 113192 539843 113248
rect 539734 113187 539843 113192
rect 539734 112948 539794 113187
rect 579797 112842 579863 112845
rect 583520 112842 584960 112932
rect 579797 112840 584960 112842
rect 579797 112784 579802 112840
rect 579858 112784 584960 112840
rect 579797 112782 584960 112784
rect 579797 112779 579863 112782
rect 583520 112692 584960 112782
rect 541157 110938 541223 110941
rect 539948 110936 541223 110938
rect 539948 110880 541162 110936
rect 541218 110880 541223 110936
rect 539948 110878 541223 110880
rect 541157 110875 541223 110878
rect -960 110666 480 110756
rect 3366 110666 3372 110668
rect -960 110606 3372 110666
rect -960 110516 480 110606
rect 3366 110604 3372 110606
rect 3436 110604 3442 110668
rect 539918 108762 539978 108868
rect 540053 108762 540119 108765
rect 539918 108760 540119 108762
rect 539918 108704 540058 108760
rect 540114 108704 540119 108760
rect 539918 108702 540119 108704
rect 540053 108699 540119 108702
rect 541341 106858 541407 106861
rect 539948 106856 541407 106858
rect 539948 106800 541346 106856
rect 541402 106800 541407 106856
rect 539948 106798 541407 106800
rect 541341 106795 541407 106798
rect 361573 106178 361639 106181
rect 359812 106176 361639 106178
rect 359812 106120 361578 106176
rect 361634 106120 361639 106176
rect 359812 106118 361639 106120
rect 361573 106115 361639 106118
rect 540145 104818 540211 104821
rect 539948 104816 540211 104818
rect 539948 104760 540150 104816
rect 540206 104760 540211 104816
rect 539948 104758 540211 104760
rect 540145 104755 540211 104758
rect 541249 102778 541315 102781
rect 539948 102776 541315 102778
rect 539948 102720 541254 102776
rect 541310 102720 541315 102776
rect 539948 102718 541315 102720
rect 541249 102715 541315 102718
rect 542905 100738 542971 100741
rect 539948 100736 542971 100738
rect 539948 100680 542910 100736
rect 542966 100680 542971 100736
rect 539948 100678 542971 100680
rect 542905 100675 542971 100678
rect 580165 99514 580231 99517
rect 583520 99514 584960 99604
rect 580165 99512 584960 99514
rect 580165 99456 580170 99512
rect 580226 99456 584960 99512
rect 580165 99454 584960 99456
rect 580165 99451 580231 99454
rect 583520 99364 584960 99454
rect 539961 99242 540027 99245
rect 539918 99240 540027 99242
rect 539918 99184 539966 99240
rect 540022 99184 540027 99240
rect 539918 99179 540027 99184
rect 2814 98636 2820 98700
rect 2884 98698 2890 98700
rect 3141 98698 3207 98701
rect 2884 98696 3207 98698
rect 2884 98640 3146 98696
rect 3202 98640 3207 98696
rect 539918 98668 539978 99179
rect 2884 98638 3207 98640
rect 2884 98636 2890 98638
rect 3141 98635 3207 98638
rect -960 97610 480 97700
rect 3550 97610 3556 97612
rect -960 97550 3556 97610
rect -960 97460 480 97550
rect 3550 97548 3556 97550
rect 3620 97548 3626 97612
rect 542721 96658 542787 96661
rect 539948 96656 542787 96658
rect 539948 96600 542726 96656
rect 542782 96600 542787 96656
rect 539948 96598 542787 96600
rect 542721 96595 542787 96598
rect 361757 95162 361823 95165
rect 359812 95160 361823 95162
rect 359812 95104 361762 95160
rect 361818 95104 361823 95160
rect 359812 95102 361823 95104
rect 361757 95099 361823 95102
rect 542813 94618 542879 94621
rect 539948 94616 542879 94618
rect 539948 94560 542818 94616
rect 542874 94560 542879 94616
rect 539948 94558 542879 94560
rect 542813 94555 542879 94558
rect 542445 92578 542511 92581
rect 539948 92576 542511 92578
rect 539948 92520 542450 92576
rect 542506 92520 542511 92576
rect 539948 92518 542511 92520
rect 542445 92515 542511 92518
rect 543273 90538 543339 90541
rect 539948 90536 543339 90538
rect 539948 90480 543278 90536
rect 543334 90480 543339 90536
rect 539948 90478 543339 90480
rect 543273 90475 543339 90478
rect 542670 88498 542676 88500
rect 539948 88438 542676 88498
rect 542670 88436 542676 88438
rect 542740 88436 542746 88500
rect 540973 86458 541039 86461
rect 539948 86456 541039 86458
rect 539948 86400 540978 86456
rect 541034 86400 541039 86456
rect 539948 86398 541039 86400
rect 540973 86395 541039 86398
rect 580165 86186 580231 86189
rect 583520 86186 584960 86276
rect 580165 86184 584960 86186
rect 580165 86128 580170 86184
rect 580226 86128 584960 86184
rect 580165 86126 584960 86128
rect 580165 86123 580231 86126
rect 583520 86036 584960 86126
rect 539685 84962 539751 84965
rect 539685 84960 539794 84962
rect 539685 84904 539690 84960
rect 539746 84904 539794 84960
rect 539685 84899 539794 84904
rect -960 84690 480 84780
rect 3734 84690 3740 84692
rect -960 84630 3740 84690
rect -960 84540 480 84630
rect 3734 84628 3740 84630
rect 3804 84628 3810 84692
rect 539734 84388 539794 84899
rect 361757 84146 361823 84149
rect 359812 84144 361823 84146
rect 359812 84088 361762 84144
rect 361818 84088 361823 84144
rect 359812 84086 361823 84088
rect 361757 84083 361823 84086
rect 539593 82786 539659 82789
rect 539550 82784 539659 82786
rect 539550 82728 539598 82784
rect 539654 82728 539659 82784
rect 539550 82723 539659 82728
rect 539550 82348 539610 82723
rect 20897 77210 20963 77213
rect 21449 77210 21515 77213
rect 20897 77208 21515 77210
rect 20897 77152 20902 77208
rect 20958 77152 21454 77208
rect 21510 77152 21515 77208
rect 20897 77150 21515 77152
rect 20897 77147 20963 77150
rect 21449 77147 21515 77150
rect 361757 73130 361823 73133
rect 359812 73128 361823 73130
rect 359812 73072 361762 73128
rect 361818 73072 361823 73128
rect 359812 73070 361823 73072
rect 361757 73067 361823 73070
rect 580165 72994 580231 72997
rect 583520 72994 584960 73084
rect 580165 72992 584960 72994
rect 580165 72936 580170 72992
rect 580226 72936 584960 72992
rect 580165 72934 584960 72936
rect 580165 72931 580231 72934
rect 583520 72844 584960 72934
rect -960 71634 480 71724
rect 3601 71634 3667 71637
rect -960 71632 3667 71634
rect -960 71576 3606 71632
rect 3662 71576 3667 71632
rect -960 71574 3667 71576
rect -960 71484 480 71574
rect 3601 71571 3667 71574
rect 361757 62114 361823 62117
rect 359812 62112 361823 62114
rect 359812 62056 361762 62112
rect 361818 62056 361823 62112
rect 359812 62054 361823 62056
rect 361757 62051 361823 62054
rect 580165 59666 580231 59669
rect 583520 59666 584960 59756
rect 580165 59664 584960 59666
rect 580165 59608 580170 59664
rect 580226 59608 584960 59664
rect 580165 59606 584960 59608
rect 580165 59603 580231 59606
rect 583520 59516 584960 59606
rect -960 58578 480 58668
rect 3509 58578 3575 58581
rect -960 58576 3575 58578
rect -960 58520 3514 58576
rect 3570 58520 3575 58576
rect -960 58518 3575 58520
rect -960 58428 480 58518
rect 3509 58515 3575 58518
rect 361757 51098 361823 51101
rect 359812 51096 361823 51098
rect 359812 51040 361762 51096
rect 361818 51040 361823 51096
rect 359812 51038 361823 51040
rect 361757 51035 361823 51038
rect 18781 49330 18847 49333
rect 22318 49330 22324 49332
rect 18781 49328 22324 49330
rect 18781 49272 18786 49328
rect 18842 49272 22324 49328
rect 18781 49270 22324 49272
rect 18781 49267 18847 49270
rect 22318 49268 22324 49270
rect 22388 49268 22394 49332
rect 11697 48922 11763 48925
rect 22134 48922 22140 48924
rect 11697 48920 22140 48922
rect 11697 48864 11702 48920
rect 11758 48864 22140 48920
rect 11697 48862 22140 48864
rect 11697 48859 11763 48862
rect 22134 48860 22140 48862
rect 22204 48860 22210 48924
rect 540605 48922 540671 48925
rect 540605 48920 540714 48922
rect 540605 48864 540610 48920
rect 540666 48864 540714 48920
rect 540605 48859 540714 48864
rect 540654 48348 540714 48859
rect 3366 46820 3372 46884
rect 3436 46882 3442 46884
rect 459001 46882 459067 46885
rect 3436 46880 459067 46882
rect 3436 46824 459006 46880
rect 459062 46824 459067 46880
rect 3436 46822 459067 46824
rect 3436 46820 3442 46822
rect 459001 46819 459067 46822
rect 3734 46684 3740 46748
rect 3804 46746 3810 46748
rect 459185 46746 459251 46749
rect 3804 46744 459251 46746
rect 3804 46688 459190 46744
rect 459246 46688 459251 46744
rect 3804 46686 459251 46688
rect 3804 46684 3810 46686
rect 459185 46683 459251 46686
rect 3550 46548 3556 46612
rect 3620 46610 3626 46612
rect 458817 46610 458883 46613
rect 3620 46608 458883 46610
rect 3620 46552 458822 46608
rect 458878 46552 458883 46608
rect 3620 46550 458883 46552
rect 3620 46548 3626 46550
rect 458817 46547 458883 46550
rect 22134 46412 22140 46476
rect 22204 46474 22210 46476
rect 361481 46474 361547 46477
rect 22204 46472 361547 46474
rect 22204 46416 361486 46472
rect 361542 46416 361547 46472
rect 22204 46414 361547 46416
rect 22204 46412 22210 46414
rect 361481 46411 361547 46414
rect 22318 46276 22324 46340
rect 22388 46338 22394 46340
rect 359549 46338 359615 46341
rect 22388 46336 359615 46338
rect 22388 46280 359554 46336
rect 359610 46280 359615 46336
rect 22388 46278 359615 46280
rect 22388 46276 22394 46278
rect 359549 46275 359615 46278
rect 580165 46338 580231 46341
rect 583520 46338 584960 46428
rect 580165 46336 584960 46338
rect 580165 46280 580170 46336
rect 580226 46280 584960 46336
rect 580165 46278 584960 46280
rect 580165 46275 580231 46278
rect 583520 46188 584960 46278
rect -960 45522 480 45612
rect 3509 45522 3575 45525
rect -960 45520 3575 45522
rect -960 45464 3514 45520
rect 3570 45464 3575 45520
rect -960 45462 3575 45464
rect -960 45372 480 45462
rect 3509 45459 3575 45462
rect 7649 44842 7715 44845
rect 406653 44842 406719 44845
rect 7649 44840 406719 44842
rect 7649 44784 7654 44840
rect 7710 44784 406658 44840
rect 406714 44784 406719 44840
rect 7649 44782 406719 44784
rect 7649 44779 7715 44782
rect 406653 44779 406719 44782
rect 536833 41034 536899 41037
rect 536833 41032 540132 41034
rect 536833 40976 536838 41032
rect 536894 40976 540132 41032
rect 536833 40974 540132 40976
rect 536833 40971 536899 40974
rect 540329 34234 540395 34237
rect 540286 34232 540395 34234
rect 540286 34176 540334 34232
rect 540390 34176 540395 34232
rect 540286 34171 540395 34176
rect 540286 33660 540346 34171
rect 580165 33146 580231 33149
rect 583520 33146 584960 33236
rect 580165 33144 584960 33146
rect 580165 33088 580170 33144
rect 580226 33088 584960 33144
rect 580165 33086 584960 33088
rect 580165 33083 580231 33086
rect 583520 32996 584960 33086
rect -960 32466 480 32556
rect 2865 32466 2931 32469
rect -960 32464 2931 32466
rect -960 32408 2870 32464
rect 2926 32408 2931 32464
rect -960 32406 2931 32408
rect -960 32316 480 32406
rect 2865 32403 2931 32406
rect 579981 19818 580047 19821
rect 583520 19818 584960 19908
rect 579981 19816 584960 19818
rect 579981 19760 579986 19816
rect 580042 19760 584960 19816
rect 579981 19758 584960 19760
rect 579981 19755 580047 19758
rect 583520 19668 584960 19758
rect -960 19410 480 19500
rect 3417 19410 3483 19413
rect -960 19408 3483 19410
rect -960 19352 3422 19408
rect 3478 19352 3483 19408
rect -960 19350 3483 19352
rect -960 19260 480 19350
rect 3417 19347 3483 19350
rect 580165 6626 580231 6629
rect 583520 6626 584960 6716
rect 580165 6624 584960 6626
rect -960 6490 480 6580
rect 580165 6568 580170 6624
rect 580226 6568 584960 6624
rect 580165 6566 584960 6568
rect 580165 6563 580231 6566
rect 3417 6490 3483 6493
rect -960 6488 3483 6490
rect -960 6432 3422 6488
rect 3478 6432 3483 6488
rect 583520 6476 584960 6566
rect -960 6430 3483 6432
rect -960 6340 480 6430
rect 3417 6427 3483 6430
rect 9949 4042 10015 4045
rect 376017 4042 376083 4045
rect 9949 4040 376083 4042
rect 9949 3984 9954 4040
rect 10010 3984 376022 4040
rect 376078 3984 376083 4040
rect 9949 3982 376083 3984
rect 9949 3979 10015 3982
rect 376017 3979 376083 3982
rect 13537 3906 13603 3909
rect 387057 3906 387123 3909
rect 13537 3904 387123 3906
rect 13537 3848 13542 3904
rect 13598 3848 387062 3904
rect 387118 3848 387123 3904
rect 13537 3846 387123 3848
rect 13537 3843 13603 3846
rect 387057 3843 387123 3846
rect 8753 3770 8819 3773
rect 392577 3770 392643 3773
rect 8753 3768 392643 3770
rect 8753 3712 8758 3768
rect 8814 3712 392582 3768
rect 392638 3712 392643 3768
rect 8753 3710 392643 3712
rect 8753 3707 8819 3710
rect 392577 3707 392643 3710
rect 2865 3634 2931 3637
rect 406561 3634 406627 3637
rect 2865 3632 406627 3634
rect 2865 3576 2870 3632
rect 2926 3576 406566 3632
rect 406622 3576 406627 3632
rect 2865 3574 406627 3576
rect 2865 3571 2931 3574
rect 406561 3571 406627 3574
rect 1669 3498 1735 3501
rect 406377 3498 406443 3501
rect 1669 3496 406443 3498
rect 1669 3440 1674 3496
rect 1730 3440 406382 3496
rect 406438 3440 406443 3496
rect 1669 3438 406443 3440
rect 1669 3435 1735 3438
rect 406377 3435 406443 3438
rect 565 3362 631 3365
rect 458766 3362 458772 3364
rect 565 3360 458772 3362
rect 565 3304 570 3360
rect 626 3304 458772 3360
rect 565 3302 458772 3304
rect 565 3299 631 3302
rect 458766 3300 458772 3302
rect 458836 3300 458842 3364
rect 5257 3226 5323 3229
rect 363597 3226 363663 3229
rect 5257 3224 363663 3226
rect 5257 3168 5262 3224
rect 5318 3168 363602 3224
rect 363658 3168 363663 3224
rect 5257 3166 363663 3168
rect 5257 3163 5323 3166
rect 363597 3163 363663 3166
<< via3 >>
rect 444236 700300 444300 700364
rect 530532 700300 530596 700364
rect 527220 699816 527284 699820
rect 527220 699760 527234 699816
rect 527234 699760 527284 699816
rect 527220 699756 527284 699760
rect 558132 699756 558196 699820
rect 446260 686428 446324 686492
rect 447732 684252 447796 684316
rect 3740 683300 3804 683364
rect 3556 683164 3620 683228
rect 3372 682756 3436 682820
rect 3740 671196 3804 671260
rect 459508 670516 459572 670580
rect 458036 665212 458100 665276
rect 459140 655692 459204 655756
rect 458956 647668 459020 647732
rect 3556 619108 3620 619172
rect 3372 606052 3436 606116
rect 472020 599524 472084 599588
rect 459140 596804 459204 596868
rect 478828 596804 478892 596868
rect 474412 542948 474476 543012
rect 472204 518196 472268 518260
rect 459508 518060 459572 518124
rect 458036 517516 458100 517580
rect 482692 517576 482756 517580
rect 482692 517520 482742 517576
rect 482742 517520 482756 517576
rect 482692 517516 482756 517520
rect 451044 516700 451108 516764
rect 450492 514320 450556 514384
rect 527220 502284 527284 502348
rect 489316 496844 489380 496908
rect 482692 462844 482756 462908
rect 448284 447204 448348 447268
rect 458956 428436 459020 428500
rect 443500 421908 443564 421972
rect 444052 421772 444116 421836
rect 448100 392532 448164 392596
rect 472204 389056 472268 389060
rect 472204 389000 472218 389056
rect 472218 389000 472268 389056
rect 472204 388996 472268 389000
rect 474412 389056 474476 389060
rect 474412 389000 474426 389056
rect 474426 389000 474476 389056
rect 474412 388996 474476 389000
rect 478828 388996 478892 389060
rect 472020 388860 472084 388924
rect 489316 386956 489380 387020
rect 448100 346156 448164 346220
rect 510660 342756 510724 342820
rect 517836 339492 517900 339556
rect 428412 334460 428476 334524
rect 518020 334596 518084 334660
rect 447916 334460 447980 334524
rect 425836 334324 425900 334388
rect 421420 334052 421484 334116
rect 510844 331876 510908 331940
rect 515260 331332 515324 331396
rect 448284 329836 448348 329900
rect 518940 329836 519004 329900
rect 515076 329700 515140 329764
rect 450676 329156 450740 329220
rect 450492 328672 450556 328676
rect 450492 328616 450506 328672
rect 450506 328616 450556 328672
rect 450492 328612 450556 328616
rect 511212 327524 511276 327588
rect 514156 326980 514220 327044
rect 510292 325892 510356 325956
rect 514892 324804 514956 324868
rect 511028 324260 511092 324324
rect 510476 323716 510540 323780
rect 510292 322628 510356 322692
rect 511212 321404 511276 321468
rect 444236 321268 444300 321332
rect 530532 321268 530596 321332
rect 447732 321132 447796 321196
rect 443500 320996 443564 321060
rect 458772 320724 458836 320788
rect 558132 320588 558196 320652
rect 444052 320044 444116 320108
rect 446260 319908 446324 319972
rect 447916 319772 447980 319836
rect 515076 316644 515140 316708
rect 542676 311068 542740 311132
rect 510476 305900 510540 305964
rect 510660 305764 510724 305828
rect 511028 305628 511092 305692
rect 515260 300596 515324 300660
rect 514156 300460 514220 300524
rect 514892 300324 514956 300388
rect 518020 300188 518084 300252
rect 517836 300052 517900 300116
rect 510844 294476 510908 294540
rect 518940 291756 519004 291820
rect 538260 278020 538324 278084
rect 421420 162692 421484 162756
rect 425836 162692 425900 162756
rect 428412 162692 428476 162756
rect 2820 136716 2884 136780
rect 539364 127196 539428 127260
rect 3372 110604 3436 110668
rect 2820 98636 2884 98700
rect 3556 97548 3620 97612
rect 542676 88436 542740 88500
rect 3740 84628 3804 84692
rect 22324 49268 22388 49332
rect 22140 48860 22204 48924
rect 3372 46820 3436 46884
rect 3740 46684 3804 46748
rect 3556 46548 3620 46612
rect 22140 46412 22204 46476
rect 22324 46276 22388 46340
rect 458772 3300 458836 3364
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 677494 -8106 711002
rect -8726 677258 -8694 677494
rect -8458 677258 -8374 677494
rect -8138 677258 -8106 677494
rect -8726 677174 -8106 677258
rect -8726 676938 -8694 677174
rect -8458 676938 -8374 677174
rect -8138 676938 -8106 677174
rect -8726 641494 -8106 676938
rect -8726 641258 -8694 641494
rect -8458 641258 -8374 641494
rect -8138 641258 -8106 641494
rect -8726 641174 -8106 641258
rect -8726 640938 -8694 641174
rect -8458 640938 -8374 641174
rect -8138 640938 -8106 641174
rect -8726 605494 -8106 640938
rect -8726 605258 -8694 605494
rect -8458 605258 -8374 605494
rect -8138 605258 -8106 605494
rect -8726 605174 -8106 605258
rect -8726 604938 -8694 605174
rect -8458 604938 -8374 605174
rect -8138 604938 -8106 605174
rect -8726 569494 -8106 604938
rect -8726 569258 -8694 569494
rect -8458 569258 -8374 569494
rect -8138 569258 -8106 569494
rect -8726 569174 -8106 569258
rect -8726 568938 -8694 569174
rect -8458 568938 -8374 569174
rect -8138 568938 -8106 569174
rect -8726 533494 -8106 568938
rect -8726 533258 -8694 533494
rect -8458 533258 -8374 533494
rect -8138 533258 -8106 533494
rect -8726 533174 -8106 533258
rect -8726 532938 -8694 533174
rect -8458 532938 -8374 533174
rect -8138 532938 -8106 533174
rect -8726 497494 -8106 532938
rect -8726 497258 -8694 497494
rect -8458 497258 -8374 497494
rect -8138 497258 -8106 497494
rect -8726 497174 -8106 497258
rect -8726 496938 -8694 497174
rect -8458 496938 -8374 497174
rect -8138 496938 -8106 497174
rect -8726 461494 -8106 496938
rect -8726 461258 -8694 461494
rect -8458 461258 -8374 461494
rect -8138 461258 -8106 461494
rect -8726 461174 -8106 461258
rect -8726 460938 -8694 461174
rect -8458 460938 -8374 461174
rect -8138 460938 -8106 461174
rect -8726 425494 -8106 460938
rect -8726 425258 -8694 425494
rect -8458 425258 -8374 425494
rect -8138 425258 -8106 425494
rect -8726 425174 -8106 425258
rect -8726 424938 -8694 425174
rect -8458 424938 -8374 425174
rect -8138 424938 -8106 425174
rect -8726 389494 -8106 424938
rect -8726 389258 -8694 389494
rect -8458 389258 -8374 389494
rect -8138 389258 -8106 389494
rect -8726 389174 -8106 389258
rect -8726 388938 -8694 389174
rect -8458 388938 -8374 389174
rect -8138 388938 -8106 389174
rect -8726 353494 -8106 388938
rect -8726 353258 -8694 353494
rect -8458 353258 -8374 353494
rect -8138 353258 -8106 353494
rect -8726 353174 -8106 353258
rect -8726 352938 -8694 353174
rect -8458 352938 -8374 353174
rect -8138 352938 -8106 353174
rect -8726 317494 -8106 352938
rect -8726 317258 -8694 317494
rect -8458 317258 -8374 317494
rect -8138 317258 -8106 317494
rect -8726 317174 -8106 317258
rect -8726 316938 -8694 317174
rect -8458 316938 -8374 317174
rect -8138 316938 -8106 317174
rect -8726 281494 -8106 316938
rect -8726 281258 -8694 281494
rect -8458 281258 -8374 281494
rect -8138 281258 -8106 281494
rect -8726 281174 -8106 281258
rect -8726 280938 -8694 281174
rect -8458 280938 -8374 281174
rect -8138 280938 -8106 281174
rect -8726 245494 -8106 280938
rect -8726 245258 -8694 245494
rect -8458 245258 -8374 245494
rect -8138 245258 -8106 245494
rect -8726 245174 -8106 245258
rect -8726 244938 -8694 245174
rect -8458 244938 -8374 245174
rect -8138 244938 -8106 245174
rect -8726 209494 -8106 244938
rect -8726 209258 -8694 209494
rect -8458 209258 -8374 209494
rect -8138 209258 -8106 209494
rect -8726 209174 -8106 209258
rect -8726 208938 -8694 209174
rect -8458 208938 -8374 209174
rect -8138 208938 -8106 209174
rect -8726 173494 -8106 208938
rect -8726 173258 -8694 173494
rect -8458 173258 -8374 173494
rect -8138 173258 -8106 173494
rect -8726 173174 -8106 173258
rect -8726 172938 -8694 173174
rect -8458 172938 -8374 173174
rect -8138 172938 -8106 173174
rect -8726 137494 -8106 172938
rect -8726 137258 -8694 137494
rect -8458 137258 -8374 137494
rect -8138 137258 -8106 137494
rect -8726 137174 -8106 137258
rect -8726 136938 -8694 137174
rect -8458 136938 -8374 137174
rect -8138 136938 -8106 137174
rect -8726 101494 -8106 136938
rect -8726 101258 -8694 101494
rect -8458 101258 -8374 101494
rect -8138 101258 -8106 101494
rect -8726 101174 -8106 101258
rect -8726 100938 -8694 101174
rect -8458 100938 -8374 101174
rect -8138 100938 -8106 101174
rect -8726 65494 -8106 100938
rect -8726 65258 -8694 65494
rect -8458 65258 -8374 65494
rect -8138 65258 -8106 65494
rect -8726 65174 -8106 65258
rect -8726 64938 -8694 65174
rect -8458 64938 -8374 65174
rect -8138 64938 -8106 65174
rect -8726 29494 -8106 64938
rect -8726 29258 -8694 29494
rect -8458 29258 -8374 29494
rect -8138 29258 -8106 29494
rect -8726 29174 -8106 29258
rect -8726 28938 -8694 29174
rect -8458 28938 -8374 29174
rect -8138 28938 -8106 29174
rect -8726 -7066 -8106 28938
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 673774 -7146 710042
rect -7766 673538 -7734 673774
rect -7498 673538 -7414 673774
rect -7178 673538 -7146 673774
rect -7766 673454 -7146 673538
rect -7766 673218 -7734 673454
rect -7498 673218 -7414 673454
rect -7178 673218 -7146 673454
rect -7766 637774 -7146 673218
rect -7766 637538 -7734 637774
rect -7498 637538 -7414 637774
rect -7178 637538 -7146 637774
rect -7766 637454 -7146 637538
rect -7766 637218 -7734 637454
rect -7498 637218 -7414 637454
rect -7178 637218 -7146 637454
rect -7766 601774 -7146 637218
rect -7766 601538 -7734 601774
rect -7498 601538 -7414 601774
rect -7178 601538 -7146 601774
rect -7766 601454 -7146 601538
rect -7766 601218 -7734 601454
rect -7498 601218 -7414 601454
rect -7178 601218 -7146 601454
rect -7766 565774 -7146 601218
rect -7766 565538 -7734 565774
rect -7498 565538 -7414 565774
rect -7178 565538 -7146 565774
rect -7766 565454 -7146 565538
rect -7766 565218 -7734 565454
rect -7498 565218 -7414 565454
rect -7178 565218 -7146 565454
rect -7766 529774 -7146 565218
rect -7766 529538 -7734 529774
rect -7498 529538 -7414 529774
rect -7178 529538 -7146 529774
rect -7766 529454 -7146 529538
rect -7766 529218 -7734 529454
rect -7498 529218 -7414 529454
rect -7178 529218 -7146 529454
rect -7766 493774 -7146 529218
rect -7766 493538 -7734 493774
rect -7498 493538 -7414 493774
rect -7178 493538 -7146 493774
rect -7766 493454 -7146 493538
rect -7766 493218 -7734 493454
rect -7498 493218 -7414 493454
rect -7178 493218 -7146 493454
rect -7766 457774 -7146 493218
rect -7766 457538 -7734 457774
rect -7498 457538 -7414 457774
rect -7178 457538 -7146 457774
rect -7766 457454 -7146 457538
rect -7766 457218 -7734 457454
rect -7498 457218 -7414 457454
rect -7178 457218 -7146 457454
rect -7766 421774 -7146 457218
rect -7766 421538 -7734 421774
rect -7498 421538 -7414 421774
rect -7178 421538 -7146 421774
rect -7766 421454 -7146 421538
rect -7766 421218 -7734 421454
rect -7498 421218 -7414 421454
rect -7178 421218 -7146 421454
rect -7766 385774 -7146 421218
rect -7766 385538 -7734 385774
rect -7498 385538 -7414 385774
rect -7178 385538 -7146 385774
rect -7766 385454 -7146 385538
rect -7766 385218 -7734 385454
rect -7498 385218 -7414 385454
rect -7178 385218 -7146 385454
rect -7766 349774 -7146 385218
rect -7766 349538 -7734 349774
rect -7498 349538 -7414 349774
rect -7178 349538 -7146 349774
rect -7766 349454 -7146 349538
rect -7766 349218 -7734 349454
rect -7498 349218 -7414 349454
rect -7178 349218 -7146 349454
rect -7766 313774 -7146 349218
rect -7766 313538 -7734 313774
rect -7498 313538 -7414 313774
rect -7178 313538 -7146 313774
rect -7766 313454 -7146 313538
rect -7766 313218 -7734 313454
rect -7498 313218 -7414 313454
rect -7178 313218 -7146 313454
rect -7766 277774 -7146 313218
rect -7766 277538 -7734 277774
rect -7498 277538 -7414 277774
rect -7178 277538 -7146 277774
rect -7766 277454 -7146 277538
rect -7766 277218 -7734 277454
rect -7498 277218 -7414 277454
rect -7178 277218 -7146 277454
rect -7766 241774 -7146 277218
rect -7766 241538 -7734 241774
rect -7498 241538 -7414 241774
rect -7178 241538 -7146 241774
rect -7766 241454 -7146 241538
rect -7766 241218 -7734 241454
rect -7498 241218 -7414 241454
rect -7178 241218 -7146 241454
rect -7766 205774 -7146 241218
rect -7766 205538 -7734 205774
rect -7498 205538 -7414 205774
rect -7178 205538 -7146 205774
rect -7766 205454 -7146 205538
rect -7766 205218 -7734 205454
rect -7498 205218 -7414 205454
rect -7178 205218 -7146 205454
rect -7766 169774 -7146 205218
rect -7766 169538 -7734 169774
rect -7498 169538 -7414 169774
rect -7178 169538 -7146 169774
rect -7766 169454 -7146 169538
rect -7766 169218 -7734 169454
rect -7498 169218 -7414 169454
rect -7178 169218 -7146 169454
rect -7766 133774 -7146 169218
rect -7766 133538 -7734 133774
rect -7498 133538 -7414 133774
rect -7178 133538 -7146 133774
rect -7766 133454 -7146 133538
rect -7766 133218 -7734 133454
rect -7498 133218 -7414 133454
rect -7178 133218 -7146 133454
rect -7766 97774 -7146 133218
rect -7766 97538 -7734 97774
rect -7498 97538 -7414 97774
rect -7178 97538 -7146 97774
rect -7766 97454 -7146 97538
rect -7766 97218 -7734 97454
rect -7498 97218 -7414 97454
rect -7178 97218 -7146 97454
rect -7766 61774 -7146 97218
rect -7766 61538 -7734 61774
rect -7498 61538 -7414 61774
rect -7178 61538 -7146 61774
rect -7766 61454 -7146 61538
rect -7766 61218 -7734 61454
rect -7498 61218 -7414 61454
rect -7178 61218 -7146 61454
rect -7766 25774 -7146 61218
rect -7766 25538 -7734 25774
rect -7498 25538 -7414 25774
rect -7178 25538 -7146 25774
rect -7766 25454 -7146 25538
rect -7766 25218 -7734 25454
rect -7498 25218 -7414 25454
rect -7178 25218 -7146 25454
rect -7766 -6106 -7146 25218
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 670054 -6186 709082
rect -6806 669818 -6774 670054
rect -6538 669818 -6454 670054
rect -6218 669818 -6186 670054
rect -6806 669734 -6186 669818
rect -6806 669498 -6774 669734
rect -6538 669498 -6454 669734
rect -6218 669498 -6186 669734
rect -6806 634054 -6186 669498
rect -6806 633818 -6774 634054
rect -6538 633818 -6454 634054
rect -6218 633818 -6186 634054
rect -6806 633734 -6186 633818
rect -6806 633498 -6774 633734
rect -6538 633498 -6454 633734
rect -6218 633498 -6186 633734
rect -6806 598054 -6186 633498
rect -6806 597818 -6774 598054
rect -6538 597818 -6454 598054
rect -6218 597818 -6186 598054
rect -6806 597734 -6186 597818
rect -6806 597498 -6774 597734
rect -6538 597498 -6454 597734
rect -6218 597498 -6186 597734
rect -6806 562054 -6186 597498
rect -6806 561818 -6774 562054
rect -6538 561818 -6454 562054
rect -6218 561818 -6186 562054
rect -6806 561734 -6186 561818
rect -6806 561498 -6774 561734
rect -6538 561498 -6454 561734
rect -6218 561498 -6186 561734
rect -6806 526054 -6186 561498
rect -6806 525818 -6774 526054
rect -6538 525818 -6454 526054
rect -6218 525818 -6186 526054
rect -6806 525734 -6186 525818
rect -6806 525498 -6774 525734
rect -6538 525498 -6454 525734
rect -6218 525498 -6186 525734
rect -6806 490054 -6186 525498
rect -6806 489818 -6774 490054
rect -6538 489818 -6454 490054
rect -6218 489818 -6186 490054
rect -6806 489734 -6186 489818
rect -6806 489498 -6774 489734
rect -6538 489498 -6454 489734
rect -6218 489498 -6186 489734
rect -6806 454054 -6186 489498
rect -6806 453818 -6774 454054
rect -6538 453818 -6454 454054
rect -6218 453818 -6186 454054
rect -6806 453734 -6186 453818
rect -6806 453498 -6774 453734
rect -6538 453498 -6454 453734
rect -6218 453498 -6186 453734
rect -6806 418054 -6186 453498
rect -6806 417818 -6774 418054
rect -6538 417818 -6454 418054
rect -6218 417818 -6186 418054
rect -6806 417734 -6186 417818
rect -6806 417498 -6774 417734
rect -6538 417498 -6454 417734
rect -6218 417498 -6186 417734
rect -6806 382054 -6186 417498
rect -6806 381818 -6774 382054
rect -6538 381818 -6454 382054
rect -6218 381818 -6186 382054
rect -6806 381734 -6186 381818
rect -6806 381498 -6774 381734
rect -6538 381498 -6454 381734
rect -6218 381498 -6186 381734
rect -6806 346054 -6186 381498
rect -6806 345818 -6774 346054
rect -6538 345818 -6454 346054
rect -6218 345818 -6186 346054
rect -6806 345734 -6186 345818
rect -6806 345498 -6774 345734
rect -6538 345498 -6454 345734
rect -6218 345498 -6186 345734
rect -6806 310054 -6186 345498
rect -6806 309818 -6774 310054
rect -6538 309818 -6454 310054
rect -6218 309818 -6186 310054
rect -6806 309734 -6186 309818
rect -6806 309498 -6774 309734
rect -6538 309498 -6454 309734
rect -6218 309498 -6186 309734
rect -6806 274054 -6186 309498
rect -6806 273818 -6774 274054
rect -6538 273818 -6454 274054
rect -6218 273818 -6186 274054
rect -6806 273734 -6186 273818
rect -6806 273498 -6774 273734
rect -6538 273498 -6454 273734
rect -6218 273498 -6186 273734
rect -6806 238054 -6186 273498
rect -6806 237818 -6774 238054
rect -6538 237818 -6454 238054
rect -6218 237818 -6186 238054
rect -6806 237734 -6186 237818
rect -6806 237498 -6774 237734
rect -6538 237498 -6454 237734
rect -6218 237498 -6186 237734
rect -6806 202054 -6186 237498
rect -6806 201818 -6774 202054
rect -6538 201818 -6454 202054
rect -6218 201818 -6186 202054
rect -6806 201734 -6186 201818
rect -6806 201498 -6774 201734
rect -6538 201498 -6454 201734
rect -6218 201498 -6186 201734
rect -6806 166054 -6186 201498
rect -6806 165818 -6774 166054
rect -6538 165818 -6454 166054
rect -6218 165818 -6186 166054
rect -6806 165734 -6186 165818
rect -6806 165498 -6774 165734
rect -6538 165498 -6454 165734
rect -6218 165498 -6186 165734
rect -6806 130054 -6186 165498
rect -6806 129818 -6774 130054
rect -6538 129818 -6454 130054
rect -6218 129818 -6186 130054
rect -6806 129734 -6186 129818
rect -6806 129498 -6774 129734
rect -6538 129498 -6454 129734
rect -6218 129498 -6186 129734
rect -6806 94054 -6186 129498
rect -6806 93818 -6774 94054
rect -6538 93818 -6454 94054
rect -6218 93818 -6186 94054
rect -6806 93734 -6186 93818
rect -6806 93498 -6774 93734
rect -6538 93498 -6454 93734
rect -6218 93498 -6186 93734
rect -6806 58054 -6186 93498
rect -6806 57818 -6774 58054
rect -6538 57818 -6454 58054
rect -6218 57818 -6186 58054
rect -6806 57734 -6186 57818
rect -6806 57498 -6774 57734
rect -6538 57498 -6454 57734
rect -6218 57498 -6186 57734
rect -6806 22054 -6186 57498
rect -6806 21818 -6774 22054
rect -6538 21818 -6454 22054
rect -6218 21818 -6186 22054
rect -6806 21734 -6186 21818
rect -6806 21498 -6774 21734
rect -6538 21498 -6454 21734
rect -6218 21498 -6186 21734
rect -6806 -5146 -6186 21498
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 666334 -5226 708122
rect -5846 666098 -5814 666334
rect -5578 666098 -5494 666334
rect -5258 666098 -5226 666334
rect -5846 666014 -5226 666098
rect -5846 665778 -5814 666014
rect -5578 665778 -5494 666014
rect -5258 665778 -5226 666014
rect -5846 630334 -5226 665778
rect -5846 630098 -5814 630334
rect -5578 630098 -5494 630334
rect -5258 630098 -5226 630334
rect -5846 630014 -5226 630098
rect -5846 629778 -5814 630014
rect -5578 629778 -5494 630014
rect -5258 629778 -5226 630014
rect -5846 594334 -5226 629778
rect -5846 594098 -5814 594334
rect -5578 594098 -5494 594334
rect -5258 594098 -5226 594334
rect -5846 594014 -5226 594098
rect -5846 593778 -5814 594014
rect -5578 593778 -5494 594014
rect -5258 593778 -5226 594014
rect -5846 558334 -5226 593778
rect -5846 558098 -5814 558334
rect -5578 558098 -5494 558334
rect -5258 558098 -5226 558334
rect -5846 558014 -5226 558098
rect -5846 557778 -5814 558014
rect -5578 557778 -5494 558014
rect -5258 557778 -5226 558014
rect -5846 522334 -5226 557778
rect -5846 522098 -5814 522334
rect -5578 522098 -5494 522334
rect -5258 522098 -5226 522334
rect -5846 522014 -5226 522098
rect -5846 521778 -5814 522014
rect -5578 521778 -5494 522014
rect -5258 521778 -5226 522014
rect -5846 486334 -5226 521778
rect -5846 486098 -5814 486334
rect -5578 486098 -5494 486334
rect -5258 486098 -5226 486334
rect -5846 486014 -5226 486098
rect -5846 485778 -5814 486014
rect -5578 485778 -5494 486014
rect -5258 485778 -5226 486014
rect -5846 450334 -5226 485778
rect -5846 450098 -5814 450334
rect -5578 450098 -5494 450334
rect -5258 450098 -5226 450334
rect -5846 450014 -5226 450098
rect -5846 449778 -5814 450014
rect -5578 449778 -5494 450014
rect -5258 449778 -5226 450014
rect -5846 414334 -5226 449778
rect -5846 414098 -5814 414334
rect -5578 414098 -5494 414334
rect -5258 414098 -5226 414334
rect -5846 414014 -5226 414098
rect -5846 413778 -5814 414014
rect -5578 413778 -5494 414014
rect -5258 413778 -5226 414014
rect -5846 378334 -5226 413778
rect -5846 378098 -5814 378334
rect -5578 378098 -5494 378334
rect -5258 378098 -5226 378334
rect -5846 378014 -5226 378098
rect -5846 377778 -5814 378014
rect -5578 377778 -5494 378014
rect -5258 377778 -5226 378014
rect -5846 342334 -5226 377778
rect -5846 342098 -5814 342334
rect -5578 342098 -5494 342334
rect -5258 342098 -5226 342334
rect -5846 342014 -5226 342098
rect -5846 341778 -5814 342014
rect -5578 341778 -5494 342014
rect -5258 341778 -5226 342014
rect -5846 306334 -5226 341778
rect -5846 306098 -5814 306334
rect -5578 306098 -5494 306334
rect -5258 306098 -5226 306334
rect -5846 306014 -5226 306098
rect -5846 305778 -5814 306014
rect -5578 305778 -5494 306014
rect -5258 305778 -5226 306014
rect -5846 270334 -5226 305778
rect -5846 270098 -5814 270334
rect -5578 270098 -5494 270334
rect -5258 270098 -5226 270334
rect -5846 270014 -5226 270098
rect -5846 269778 -5814 270014
rect -5578 269778 -5494 270014
rect -5258 269778 -5226 270014
rect -5846 234334 -5226 269778
rect -5846 234098 -5814 234334
rect -5578 234098 -5494 234334
rect -5258 234098 -5226 234334
rect -5846 234014 -5226 234098
rect -5846 233778 -5814 234014
rect -5578 233778 -5494 234014
rect -5258 233778 -5226 234014
rect -5846 198334 -5226 233778
rect -5846 198098 -5814 198334
rect -5578 198098 -5494 198334
rect -5258 198098 -5226 198334
rect -5846 198014 -5226 198098
rect -5846 197778 -5814 198014
rect -5578 197778 -5494 198014
rect -5258 197778 -5226 198014
rect -5846 162334 -5226 197778
rect -5846 162098 -5814 162334
rect -5578 162098 -5494 162334
rect -5258 162098 -5226 162334
rect -5846 162014 -5226 162098
rect -5846 161778 -5814 162014
rect -5578 161778 -5494 162014
rect -5258 161778 -5226 162014
rect -5846 126334 -5226 161778
rect -5846 126098 -5814 126334
rect -5578 126098 -5494 126334
rect -5258 126098 -5226 126334
rect -5846 126014 -5226 126098
rect -5846 125778 -5814 126014
rect -5578 125778 -5494 126014
rect -5258 125778 -5226 126014
rect -5846 90334 -5226 125778
rect -5846 90098 -5814 90334
rect -5578 90098 -5494 90334
rect -5258 90098 -5226 90334
rect -5846 90014 -5226 90098
rect -5846 89778 -5814 90014
rect -5578 89778 -5494 90014
rect -5258 89778 -5226 90014
rect -5846 54334 -5226 89778
rect -5846 54098 -5814 54334
rect -5578 54098 -5494 54334
rect -5258 54098 -5226 54334
rect -5846 54014 -5226 54098
rect -5846 53778 -5814 54014
rect -5578 53778 -5494 54014
rect -5258 53778 -5226 54014
rect -5846 18334 -5226 53778
rect -5846 18098 -5814 18334
rect -5578 18098 -5494 18334
rect -5258 18098 -5226 18334
rect -5846 18014 -5226 18098
rect -5846 17778 -5814 18014
rect -5578 17778 -5494 18014
rect -5258 17778 -5226 18014
rect -5846 -4186 -5226 17778
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 698614 -4266 707162
rect -4886 698378 -4854 698614
rect -4618 698378 -4534 698614
rect -4298 698378 -4266 698614
rect -4886 698294 -4266 698378
rect -4886 698058 -4854 698294
rect -4618 698058 -4534 698294
rect -4298 698058 -4266 698294
rect -4886 662614 -4266 698058
rect -4886 662378 -4854 662614
rect -4618 662378 -4534 662614
rect -4298 662378 -4266 662614
rect -4886 662294 -4266 662378
rect -4886 662058 -4854 662294
rect -4618 662058 -4534 662294
rect -4298 662058 -4266 662294
rect -4886 626614 -4266 662058
rect -4886 626378 -4854 626614
rect -4618 626378 -4534 626614
rect -4298 626378 -4266 626614
rect -4886 626294 -4266 626378
rect -4886 626058 -4854 626294
rect -4618 626058 -4534 626294
rect -4298 626058 -4266 626294
rect -4886 590614 -4266 626058
rect -4886 590378 -4854 590614
rect -4618 590378 -4534 590614
rect -4298 590378 -4266 590614
rect -4886 590294 -4266 590378
rect -4886 590058 -4854 590294
rect -4618 590058 -4534 590294
rect -4298 590058 -4266 590294
rect -4886 554614 -4266 590058
rect -4886 554378 -4854 554614
rect -4618 554378 -4534 554614
rect -4298 554378 -4266 554614
rect -4886 554294 -4266 554378
rect -4886 554058 -4854 554294
rect -4618 554058 -4534 554294
rect -4298 554058 -4266 554294
rect -4886 518614 -4266 554058
rect -4886 518378 -4854 518614
rect -4618 518378 -4534 518614
rect -4298 518378 -4266 518614
rect -4886 518294 -4266 518378
rect -4886 518058 -4854 518294
rect -4618 518058 -4534 518294
rect -4298 518058 -4266 518294
rect -4886 482614 -4266 518058
rect -4886 482378 -4854 482614
rect -4618 482378 -4534 482614
rect -4298 482378 -4266 482614
rect -4886 482294 -4266 482378
rect -4886 482058 -4854 482294
rect -4618 482058 -4534 482294
rect -4298 482058 -4266 482294
rect -4886 446614 -4266 482058
rect -4886 446378 -4854 446614
rect -4618 446378 -4534 446614
rect -4298 446378 -4266 446614
rect -4886 446294 -4266 446378
rect -4886 446058 -4854 446294
rect -4618 446058 -4534 446294
rect -4298 446058 -4266 446294
rect -4886 410614 -4266 446058
rect -4886 410378 -4854 410614
rect -4618 410378 -4534 410614
rect -4298 410378 -4266 410614
rect -4886 410294 -4266 410378
rect -4886 410058 -4854 410294
rect -4618 410058 -4534 410294
rect -4298 410058 -4266 410294
rect -4886 374614 -4266 410058
rect -4886 374378 -4854 374614
rect -4618 374378 -4534 374614
rect -4298 374378 -4266 374614
rect -4886 374294 -4266 374378
rect -4886 374058 -4854 374294
rect -4618 374058 -4534 374294
rect -4298 374058 -4266 374294
rect -4886 338614 -4266 374058
rect -4886 338378 -4854 338614
rect -4618 338378 -4534 338614
rect -4298 338378 -4266 338614
rect -4886 338294 -4266 338378
rect -4886 338058 -4854 338294
rect -4618 338058 -4534 338294
rect -4298 338058 -4266 338294
rect -4886 302614 -4266 338058
rect -4886 302378 -4854 302614
rect -4618 302378 -4534 302614
rect -4298 302378 -4266 302614
rect -4886 302294 -4266 302378
rect -4886 302058 -4854 302294
rect -4618 302058 -4534 302294
rect -4298 302058 -4266 302294
rect -4886 266614 -4266 302058
rect -4886 266378 -4854 266614
rect -4618 266378 -4534 266614
rect -4298 266378 -4266 266614
rect -4886 266294 -4266 266378
rect -4886 266058 -4854 266294
rect -4618 266058 -4534 266294
rect -4298 266058 -4266 266294
rect -4886 230614 -4266 266058
rect -4886 230378 -4854 230614
rect -4618 230378 -4534 230614
rect -4298 230378 -4266 230614
rect -4886 230294 -4266 230378
rect -4886 230058 -4854 230294
rect -4618 230058 -4534 230294
rect -4298 230058 -4266 230294
rect -4886 194614 -4266 230058
rect -4886 194378 -4854 194614
rect -4618 194378 -4534 194614
rect -4298 194378 -4266 194614
rect -4886 194294 -4266 194378
rect -4886 194058 -4854 194294
rect -4618 194058 -4534 194294
rect -4298 194058 -4266 194294
rect -4886 158614 -4266 194058
rect -4886 158378 -4854 158614
rect -4618 158378 -4534 158614
rect -4298 158378 -4266 158614
rect -4886 158294 -4266 158378
rect -4886 158058 -4854 158294
rect -4618 158058 -4534 158294
rect -4298 158058 -4266 158294
rect -4886 122614 -4266 158058
rect -4886 122378 -4854 122614
rect -4618 122378 -4534 122614
rect -4298 122378 -4266 122614
rect -4886 122294 -4266 122378
rect -4886 122058 -4854 122294
rect -4618 122058 -4534 122294
rect -4298 122058 -4266 122294
rect -4886 86614 -4266 122058
rect -4886 86378 -4854 86614
rect -4618 86378 -4534 86614
rect -4298 86378 -4266 86614
rect -4886 86294 -4266 86378
rect -4886 86058 -4854 86294
rect -4618 86058 -4534 86294
rect -4298 86058 -4266 86294
rect -4886 50614 -4266 86058
rect -4886 50378 -4854 50614
rect -4618 50378 -4534 50614
rect -4298 50378 -4266 50614
rect -4886 50294 -4266 50378
rect -4886 50058 -4854 50294
rect -4618 50058 -4534 50294
rect -4298 50058 -4266 50294
rect -4886 14614 -4266 50058
rect -4886 14378 -4854 14614
rect -4618 14378 -4534 14614
rect -4298 14378 -4266 14614
rect -4886 14294 -4266 14378
rect -4886 14058 -4854 14294
rect -4618 14058 -4534 14294
rect -4298 14058 -4266 14294
rect -4886 -3226 -4266 14058
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 694894 -3306 706202
rect -3926 694658 -3894 694894
rect -3658 694658 -3574 694894
rect -3338 694658 -3306 694894
rect -3926 694574 -3306 694658
rect -3926 694338 -3894 694574
rect -3658 694338 -3574 694574
rect -3338 694338 -3306 694574
rect -3926 658894 -3306 694338
rect -3926 658658 -3894 658894
rect -3658 658658 -3574 658894
rect -3338 658658 -3306 658894
rect -3926 658574 -3306 658658
rect -3926 658338 -3894 658574
rect -3658 658338 -3574 658574
rect -3338 658338 -3306 658574
rect -3926 622894 -3306 658338
rect -3926 622658 -3894 622894
rect -3658 622658 -3574 622894
rect -3338 622658 -3306 622894
rect -3926 622574 -3306 622658
rect -3926 622338 -3894 622574
rect -3658 622338 -3574 622574
rect -3338 622338 -3306 622574
rect -3926 586894 -3306 622338
rect -3926 586658 -3894 586894
rect -3658 586658 -3574 586894
rect -3338 586658 -3306 586894
rect -3926 586574 -3306 586658
rect -3926 586338 -3894 586574
rect -3658 586338 -3574 586574
rect -3338 586338 -3306 586574
rect -3926 550894 -3306 586338
rect -3926 550658 -3894 550894
rect -3658 550658 -3574 550894
rect -3338 550658 -3306 550894
rect -3926 550574 -3306 550658
rect -3926 550338 -3894 550574
rect -3658 550338 -3574 550574
rect -3338 550338 -3306 550574
rect -3926 514894 -3306 550338
rect -3926 514658 -3894 514894
rect -3658 514658 -3574 514894
rect -3338 514658 -3306 514894
rect -3926 514574 -3306 514658
rect -3926 514338 -3894 514574
rect -3658 514338 -3574 514574
rect -3338 514338 -3306 514574
rect -3926 478894 -3306 514338
rect -3926 478658 -3894 478894
rect -3658 478658 -3574 478894
rect -3338 478658 -3306 478894
rect -3926 478574 -3306 478658
rect -3926 478338 -3894 478574
rect -3658 478338 -3574 478574
rect -3338 478338 -3306 478574
rect -3926 442894 -3306 478338
rect -3926 442658 -3894 442894
rect -3658 442658 -3574 442894
rect -3338 442658 -3306 442894
rect -3926 442574 -3306 442658
rect -3926 442338 -3894 442574
rect -3658 442338 -3574 442574
rect -3338 442338 -3306 442574
rect -3926 406894 -3306 442338
rect -3926 406658 -3894 406894
rect -3658 406658 -3574 406894
rect -3338 406658 -3306 406894
rect -3926 406574 -3306 406658
rect -3926 406338 -3894 406574
rect -3658 406338 -3574 406574
rect -3338 406338 -3306 406574
rect -3926 370894 -3306 406338
rect -3926 370658 -3894 370894
rect -3658 370658 -3574 370894
rect -3338 370658 -3306 370894
rect -3926 370574 -3306 370658
rect -3926 370338 -3894 370574
rect -3658 370338 -3574 370574
rect -3338 370338 -3306 370574
rect -3926 334894 -3306 370338
rect -3926 334658 -3894 334894
rect -3658 334658 -3574 334894
rect -3338 334658 -3306 334894
rect -3926 334574 -3306 334658
rect -3926 334338 -3894 334574
rect -3658 334338 -3574 334574
rect -3338 334338 -3306 334574
rect -3926 298894 -3306 334338
rect -3926 298658 -3894 298894
rect -3658 298658 -3574 298894
rect -3338 298658 -3306 298894
rect -3926 298574 -3306 298658
rect -3926 298338 -3894 298574
rect -3658 298338 -3574 298574
rect -3338 298338 -3306 298574
rect -3926 262894 -3306 298338
rect -3926 262658 -3894 262894
rect -3658 262658 -3574 262894
rect -3338 262658 -3306 262894
rect -3926 262574 -3306 262658
rect -3926 262338 -3894 262574
rect -3658 262338 -3574 262574
rect -3338 262338 -3306 262574
rect -3926 226894 -3306 262338
rect -3926 226658 -3894 226894
rect -3658 226658 -3574 226894
rect -3338 226658 -3306 226894
rect -3926 226574 -3306 226658
rect -3926 226338 -3894 226574
rect -3658 226338 -3574 226574
rect -3338 226338 -3306 226574
rect -3926 190894 -3306 226338
rect -3926 190658 -3894 190894
rect -3658 190658 -3574 190894
rect -3338 190658 -3306 190894
rect -3926 190574 -3306 190658
rect -3926 190338 -3894 190574
rect -3658 190338 -3574 190574
rect -3338 190338 -3306 190574
rect -3926 154894 -3306 190338
rect -3926 154658 -3894 154894
rect -3658 154658 -3574 154894
rect -3338 154658 -3306 154894
rect -3926 154574 -3306 154658
rect -3926 154338 -3894 154574
rect -3658 154338 -3574 154574
rect -3338 154338 -3306 154574
rect -3926 118894 -3306 154338
rect -3926 118658 -3894 118894
rect -3658 118658 -3574 118894
rect -3338 118658 -3306 118894
rect -3926 118574 -3306 118658
rect -3926 118338 -3894 118574
rect -3658 118338 -3574 118574
rect -3338 118338 -3306 118574
rect -3926 82894 -3306 118338
rect -3926 82658 -3894 82894
rect -3658 82658 -3574 82894
rect -3338 82658 -3306 82894
rect -3926 82574 -3306 82658
rect -3926 82338 -3894 82574
rect -3658 82338 -3574 82574
rect -3338 82338 -3306 82574
rect -3926 46894 -3306 82338
rect -3926 46658 -3894 46894
rect -3658 46658 -3574 46894
rect -3338 46658 -3306 46894
rect -3926 46574 -3306 46658
rect -3926 46338 -3894 46574
rect -3658 46338 -3574 46574
rect -3338 46338 -3306 46574
rect -3926 10894 -3306 46338
rect -3926 10658 -3894 10894
rect -3658 10658 -3574 10894
rect -3338 10658 -3306 10894
rect -3926 10574 -3306 10658
rect -3926 10338 -3894 10574
rect -3658 10338 -3574 10574
rect -3338 10338 -3306 10574
rect -3926 -2266 -3306 10338
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 691174 -2346 705242
rect -2966 690938 -2934 691174
rect -2698 690938 -2614 691174
rect -2378 690938 -2346 691174
rect -2966 690854 -2346 690938
rect -2966 690618 -2934 690854
rect -2698 690618 -2614 690854
rect -2378 690618 -2346 690854
rect -2966 655174 -2346 690618
rect -2966 654938 -2934 655174
rect -2698 654938 -2614 655174
rect -2378 654938 -2346 655174
rect -2966 654854 -2346 654938
rect -2966 654618 -2934 654854
rect -2698 654618 -2614 654854
rect -2378 654618 -2346 654854
rect -2966 619174 -2346 654618
rect -2966 618938 -2934 619174
rect -2698 618938 -2614 619174
rect -2378 618938 -2346 619174
rect -2966 618854 -2346 618938
rect -2966 618618 -2934 618854
rect -2698 618618 -2614 618854
rect -2378 618618 -2346 618854
rect -2966 583174 -2346 618618
rect -2966 582938 -2934 583174
rect -2698 582938 -2614 583174
rect -2378 582938 -2346 583174
rect -2966 582854 -2346 582938
rect -2966 582618 -2934 582854
rect -2698 582618 -2614 582854
rect -2378 582618 -2346 582854
rect -2966 547174 -2346 582618
rect -2966 546938 -2934 547174
rect -2698 546938 -2614 547174
rect -2378 546938 -2346 547174
rect -2966 546854 -2346 546938
rect -2966 546618 -2934 546854
rect -2698 546618 -2614 546854
rect -2378 546618 -2346 546854
rect -2966 511174 -2346 546618
rect -2966 510938 -2934 511174
rect -2698 510938 -2614 511174
rect -2378 510938 -2346 511174
rect -2966 510854 -2346 510938
rect -2966 510618 -2934 510854
rect -2698 510618 -2614 510854
rect -2378 510618 -2346 510854
rect -2966 475174 -2346 510618
rect -2966 474938 -2934 475174
rect -2698 474938 -2614 475174
rect -2378 474938 -2346 475174
rect -2966 474854 -2346 474938
rect -2966 474618 -2934 474854
rect -2698 474618 -2614 474854
rect -2378 474618 -2346 474854
rect -2966 439174 -2346 474618
rect -2966 438938 -2934 439174
rect -2698 438938 -2614 439174
rect -2378 438938 -2346 439174
rect -2966 438854 -2346 438938
rect -2966 438618 -2934 438854
rect -2698 438618 -2614 438854
rect -2378 438618 -2346 438854
rect -2966 403174 -2346 438618
rect -2966 402938 -2934 403174
rect -2698 402938 -2614 403174
rect -2378 402938 -2346 403174
rect -2966 402854 -2346 402938
rect -2966 402618 -2934 402854
rect -2698 402618 -2614 402854
rect -2378 402618 -2346 402854
rect -2966 367174 -2346 402618
rect -2966 366938 -2934 367174
rect -2698 366938 -2614 367174
rect -2378 366938 -2346 367174
rect -2966 366854 -2346 366938
rect -2966 366618 -2934 366854
rect -2698 366618 -2614 366854
rect -2378 366618 -2346 366854
rect -2966 331174 -2346 366618
rect -2966 330938 -2934 331174
rect -2698 330938 -2614 331174
rect -2378 330938 -2346 331174
rect -2966 330854 -2346 330938
rect -2966 330618 -2934 330854
rect -2698 330618 -2614 330854
rect -2378 330618 -2346 330854
rect -2966 295174 -2346 330618
rect -2966 294938 -2934 295174
rect -2698 294938 -2614 295174
rect -2378 294938 -2346 295174
rect -2966 294854 -2346 294938
rect -2966 294618 -2934 294854
rect -2698 294618 -2614 294854
rect -2378 294618 -2346 294854
rect -2966 259174 -2346 294618
rect -2966 258938 -2934 259174
rect -2698 258938 -2614 259174
rect -2378 258938 -2346 259174
rect -2966 258854 -2346 258938
rect -2966 258618 -2934 258854
rect -2698 258618 -2614 258854
rect -2378 258618 -2346 258854
rect -2966 223174 -2346 258618
rect -2966 222938 -2934 223174
rect -2698 222938 -2614 223174
rect -2378 222938 -2346 223174
rect -2966 222854 -2346 222938
rect -2966 222618 -2934 222854
rect -2698 222618 -2614 222854
rect -2378 222618 -2346 222854
rect -2966 187174 -2346 222618
rect -2966 186938 -2934 187174
rect -2698 186938 -2614 187174
rect -2378 186938 -2346 187174
rect -2966 186854 -2346 186938
rect -2966 186618 -2934 186854
rect -2698 186618 -2614 186854
rect -2378 186618 -2346 186854
rect -2966 151174 -2346 186618
rect -2966 150938 -2934 151174
rect -2698 150938 -2614 151174
rect -2378 150938 -2346 151174
rect -2966 150854 -2346 150938
rect -2966 150618 -2934 150854
rect -2698 150618 -2614 150854
rect -2378 150618 -2346 150854
rect -2966 115174 -2346 150618
rect -2966 114938 -2934 115174
rect -2698 114938 -2614 115174
rect -2378 114938 -2346 115174
rect -2966 114854 -2346 114938
rect -2966 114618 -2934 114854
rect -2698 114618 -2614 114854
rect -2378 114618 -2346 114854
rect -2966 79174 -2346 114618
rect -2966 78938 -2934 79174
rect -2698 78938 -2614 79174
rect -2378 78938 -2346 79174
rect -2966 78854 -2346 78938
rect -2966 78618 -2934 78854
rect -2698 78618 -2614 78854
rect -2378 78618 -2346 78854
rect -2966 43174 -2346 78618
rect -2966 42938 -2934 43174
rect -2698 42938 -2614 43174
rect -2378 42938 -2346 43174
rect -2966 42854 -2346 42938
rect -2966 42618 -2934 42854
rect -2698 42618 -2614 42854
rect -2378 42618 -2346 42854
rect -2966 7174 -2346 42618
rect -2966 6938 -2934 7174
rect -2698 6938 -2614 7174
rect -2378 6938 -2346 7174
rect -2966 6854 -2346 6938
rect -2966 6618 -2934 6854
rect -2698 6618 -2614 6854
rect -2378 6618 -2346 6854
rect -2966 -1306 -2346 6618
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 687454 -1386 704282
rect -2006 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 -1386 687454
rect -2006 687134 -1386 687218
rect -2006 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 -1386 687134
rect -2006 651454 -1386 686898
rect -2006 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 -1386 651454
rect -2006 651134 -1386 651218
rect -2006 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 -1386 651134
rect -2006 615454 -1386 650898
rect -2006 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 -1386 615454
rect -2006 615134 -1386 615218
rect -2006 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 -1386 615134
rect -2006 579454 -1386 614898
rect -2006 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 -1386 579454
rect -2006 579134 -1386 579218
rect -2006 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 -1386 579134
rect -2006 543454 -1386 578898
rect -2006 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 -1386 543454
rect -2006 543134 -1386 543218
rect -2006 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 -1386 543134
rect -2006 507454 -1386 542898
rect -2006 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 -1386 507454
rect -2006 507134 -1386 507218
rect -2006 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 -1386 507134
rect -2006 471454 -1386 506898
rect -2006 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 -1386 471454
rect -2006 471134 -1386 471218
rect -2006 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 -1386 471134
rect -2006 435454 -1386 470898
rect -2006 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 -1386 435454
rect -2006 435134 -1386 435218
rect -2006 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 -1386 435134
rect -2006 399454 -1386 434898
rect -2006 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 -1386 399454
rect -2006 399134 -1386 399218
rect -2006 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 -1386 399134
rect -2006 363454 -1386 398898
rect -2006 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 -1386 363454
rect -2006 363134 -1386 363218
rect -2006 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 -1386 363134
rect -2006 327454 -1386 362898
rect -2006 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 -1386 327454
rect -2006 327134 -1386 327218
rect -2006 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 -1386 327134
rect -2006 291454 -1386 326898
rect -2006 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 -1386 291454
rect -2006 291134 -1386 291218
rect -2006 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 -1386 291134
rect -2006 255454 -1386 290898
rect -2006 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 -1386 255454
rect -2006 255134 -1386 255218
rect -2006 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 -1386 255134
rect -2006 219454 -1386 254898
rect -2006 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 -1386 219454
rect -2006 219134 -1386 219218
rect -2006 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 -1386 219134
rect -2006 183454 -1386 218898
rect -2006 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 -1386 183454
rect -2006 183134 -1386 183218
rect -2006 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 -1386 183134
rect -2006 147454 -1386 182898
rect -2006 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 -1386 147454
rect -2006 147134 -1386 147218
rect -2006 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 -1386 147134
rect -2006 111454 -1386 146898
rect -2006 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 -1386 111454
rect -2006 111134 -1386 111218
rect -2006 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 -1386 111134
rect -2006 75454 -1386 110898
rect -2006 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 -1386 75454
rect -2006 75134 -1386 75218
rect -2006 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 -1386 75134
rect -2006 39454 -1386 74898
rect -2006 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 -1386 39454
rect -2006 39134 -1386 39218
rect -2006 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 -1386 39134
rect -2006 3454 -1386 38898
rect -2006 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 -1386 3454
rect -2006 3134 -1386 3218
rect -2006 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 -1386 3134
rect -2006 -346 -1386 2898
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect 1794 704838 2414 711590
rect 1794 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 2414 704838
rect 1794 704518 2414 704602
rect 1794 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 2414 704518
rect 1794 687454 2414 704282
rect 1794 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 2414 687454
rect 1794 687134 2414 687218
rect 1794 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 2414 687134
rect 1794 651454 2414 686898
rect 5514 705798 6134 711590
rect 5514 705562 5546 705798
rect 5782 705562 5866 705798
rect 6102 705562 6134 705798
rect 5514 705478 6134 705562
rect 5514 705242 5546 705478
rect 5782 705242 5866 705478
rect 6102 705242 6134 705478
rect 5514 691174 6134 705242
rect 5514 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 6134 691174
rect 5514 690854 6134 690938
rect 5514 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 6134 690854
rect 3739 683364 3805 683365
rect 3739 683300 3740 683364
rect 3804 683300 3805 683364
rect 3739 683299 3805 683300
rect 3555 683228 3621 683229
rect 3555 683164 3556 683228
rect 3620 683164 3621 683228
rect 3555 683163 3621 683164
rect 3371 682820 3437 682821
rect 3371 682756 3372 682820
rect 3436 682756 3437 682820
rect 3371 682755 3437 682756
rect 1794 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 2414 651454
rect 1794 651134 2414 651218
rect 1794 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 2414 651134
rect 1794 615454 2414 650898
rect 1794 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 2414 615454
rect 1794 615134 2414 615218
rect 1794 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 2414 615134
rect 1794 579454 2414 614898
rect 3374 606117 3434 682755
rect 3558 619173 3618 683163
rect 3742 671261 3802 683299
rect 3739 671260 3805 671261
rect 3739 671196 3740 671260
rect 3804 671196 3805 671260
rect 3739 671195 3805 671196
rect 5514 655174 6134 690618
rect 5514 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 6134 655174
rect 5514 654854 6134 654938
rect 5514 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 6134 654854
rect 5514 619174 6134 654618
rect 3555 619172 3621 619173
rect 3555 619108 3556 619172
rect 3620 619108 3621 619172
rect 3555 619107 3621 619108
rect 5514 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 6134 619174
rect 5514 618854 6134 618938
rect 5514 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 6134 618854
rect 3371 606116 3437 606117
rect 3371 606052 3372 606116
rect 3436 606052 3437 606116
rect 3371 606051 3437 606052
rect 1794 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 2414 579454
rect 1794 579134 2414 579218
rect 1794 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 2414 579134
rect 1794 543454 2414 578898
rect 1794 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 2414 543454
rect 1794 543134 2414 543218
rect 1794 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 2414 543134
rect 1794 507454 2414 542898
rect 1794 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 2414 507454
rect 1794 507134 2414 507218
rect 1794 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 2414 507134
rect 1794 471454 2414 506898
rect 1794 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 2414 471454
rect 1794 471134 2414 471218
rect 1794 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 2414 471134
rect 1794 435454 2414 470898
rect 1794 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 2414 435454
rect 1794 435134 2414 435218
rect 1794 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 2414 435134
rect 1794 399454 2414 434898
rect 1794 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 2414 399454
rect 1794 399134 2414 399218
rect 1794 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 2414 399134
rect 1794 363454 2414 398898
rect 1794 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 2414 363454
rect 1794 363134 2414 363218
rect 1794 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 2414 363134
rect 1794 327454 2414 362898
rect 1794 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 2414 327454
rect 1794 327134 2414 327218
rect 1794 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 2414 327134
rect 1794 291454 2414 326898
rect 1794 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 2414 291454
rect 1794 291134 2414 291218
rect 1794 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 2414 291134
rect 1794 255454 2414 290898
rect 1794 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 2414 255454
rect 1794 255134 2414 255218
rect 1794 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 2414 255134
rect 1794 219454 2414 254898
rect 1794 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 2414 219454
rect 1794 219134 2414 219218
rect 1794 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 2414 219134
rect 1794 183454 2414 218898
rect 1794 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 2414 183454
rect 1794 183134 2414 183218
rect 1794 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 2414 183134
rect 1794 147454 2414 182898
rect 1794 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 2414 147454
rect 1794 147134 2414 147218
rect 1794 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 2414 147134
rect 1794 111454 2414 146898
rect 5514 583174 6134 618618
rect 5514 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 6134 583174
rect 5514 582854 6134 582938
rect 5514 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 6134 582854
rect 5514 547174 6134 582618
rect 5514 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 6134 547174
rect 5514 546854 6134 546938
rect 5514 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 6134 546854
rect 5514 511174 6134 546618
rect 5514 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 6134 511174
rect 5514 510854 6134 510938
rect 5514 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 6134 510854
rect 5514 475174 6134 510618
rect 5514 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 6134 475174
rect 5514 474854 6134 474938
rect 5514 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 6134 474854
rect 5514 439174 6134 474618
rect 5514 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 6134 439174
rect 5514 438854 6134 438938
rect 5514 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 6134 438854
rect 5514 403174 6134 438618
rect 5514 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 6134 403174
rect 5514 402854 6134 402938
rect 5514 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 6134 402854
rect 5514 367174 6134 402618
rect 5514 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 6134 367174
rect 5514 366854 6134 366938
rect 5514 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 6134 366854
rect 5514 331174 6134 366618
rect 5514 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 6134 331174
rect 5514 330854 6134 330938
rect 5514 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 6134 330854
rect 5514 295174 6134 330618
rect 5514 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 6134 295174
rect 5514 294854 6134 294938
rect 5514 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 6134 294854
rect 5514 259174 6134 294618
rect 5514 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 6134 259174
rect 5514 258854 6134 258938
rect 5514 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 6134 258854
rect 5514 223174 6134 258618
rect 5514 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 6134 223174
rect 5514 222854 6134 222938
rect 5514 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 6134 222854
rect 5514 187174 6134 222618
rect 5514 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 6134 187174
rect 5514 186854 6134 186938
rect 5514 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 6134 186854
rect 5514 151174 6134 186618
rect 5514 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 6134 151174
rect 5514 150854 6134 150938
rect 5514 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 6134 150854
rect 2819 136780 2885 136781
rect 2819 136716 2820 136780
rect 2884 136716 2885 136780
rect 2819 136715 2885 136716
rect 1794 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 2414 111454
rect 1794 111134 2414 111218
rect 1794 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 2414 111134
rect 1794 75454 2414 110898
rect 2822 98701 2882 136715
rect 5514 115174 6134 150618
rect 5514 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 6134 115174
rect 5514 114854 6134 114938
rect 5514 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 6134 114854
rect 3371 110668 3437 110669
rect 3371 110604 3372 110668
rect 3436 110604 3437 110668
rect 3371 110603 3437 110604
rect 2819 98700 2885 98701
rect 2819 98636 2820 98700
rect 2884 98636 2885 98700
rect 2819 98635 2885 98636
rect 1794 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 2414 75454
rect 1794 75134 2414 75218
rect 1794 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 2414 75134
rect 1794 39454 2414 74898
rect 3374 46885 3434 110603
rect 3555 97612 3621 97613
rect 3555 97548 3556 97612
rect 3620 97548 3621 97612
rect 3555 97547 3621 97548
rect 3371 46884 3437 46885
rect 3371 46820 3372 46884
rect 3436 46820 3437 46884
rect 3371 46819 3437 46820
rect 3558 46613 3618 97547
rect 3739 84692 3805 84693
rect 3739 84628 3740 84692
rect 3804 84628 3805 84692
rect 3739 84627 3805 84628
rect 3742 46749 3802 84627
rect 5514 79174 6134 114618
rect 5514 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 6134 79174
rect 5514 78854 6134 78938
rect 5514 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 6134 78854
rect 3739 46748 3805 46749
rect 3739 46684 3740 46748
rect 3804 46684 3805 46748
rect 3739 46683 3805 46684
rect 3555 46612 3621 46613
rect 3555 46548 3556 46612
rect 3620 46548 3621 46612
rect 3555 46547 3621 46548
rect 1794 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 2414 39454
rect 1794 39134 2414 39218
rect 1794 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 2414 39134
rect 1794 3454 2414 38898
rect 1794 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 2414 3454
rect 1794 3134 2414 3218
rect 1794 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 2414 3134
rect 1794 -346 2414 2898
rect 1794 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 2414 -346
rect 1794 -666 2414 -582
rect 1794 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 2414 -666
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 1794 -7654 2414 -902
rect 5514 43174 6134 78618
rect 5514 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 6134 43174
rect 5514 42854 6134 42938
rect 5514 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 6134 42854
rect 5514 7174 6134 42618
rect 5514 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 6134 7174
rect 5514 6854 6134 6938
rect 5514 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 6134 6854
rect 5514 -1306 6134 6618
rect 5514 -1542 5546 -1306
rect 5782 -1542 5866 -1306
rect 6102 -1542 6134 -1306
rect 5514 -1626 6134 -1542
rect 5514 -1862 5546 -1626
rect 5782 -1862 5866 -1626
rect 6102 -1862 6134 -1626
rect 5514 -7654 6134 -1862
rect 9234 706758 9854 711590
rect 9234 706522 9266 706758
rect 9502 706522 9586 706758
rect 9822 706522 9854 706758
rect 9234 706438 9854 706522
rect 9234 706202 9266 706438
rect 9502 706202 9586 706438
rect 9822 706202 9854 706438
rect 9234 694894 9854 706202
rect 9234 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 9854 694894
rect 9234 694574 9854 694658
rect 9234 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 9854 694574
rect 9234 658894 9854 694338
rect 9234 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 9854 658894
rect 9234 658574 9854 658658
rect 9234 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 9854 658574
rect 9234 622894 9854 658338
rect 9234 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 9854 622894
rect 9234 622574 9854 622658
rect 9234 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 9854 622574
rect 9234 586894 9854 622338
rect 9234 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 9854 586894
rect 9234 586574 9854 586658
rect 9234 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 9854 586574
rect 9234 550894 9854 586338
rect 9234 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 9854 550894
rect 9234 550574 9854 550658
rect 9234 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 9854 550574
rect 9234 514894 9854 550338
rect 9234 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 9854 514894
rect 9234 514574 9854 514658
rect 9234 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 9854 514574
rect 9234 478894 9854 514338
rect 9234 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 9854 478894
rect 9234 478574 9854 478658
rect 9234 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 9854 478574
rect 9234 442894 9854 478338
rect 9234 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 9854 442894
rect 9234 442574 9854 442658
rect 9234 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 9854 442574
rect 9234 406894 9854 442338
rect 9234 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 9854 406894
rect 9234 406574 9854 406658
rect 9234 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 9854 406574
rect 9234 370894 9854 406338
rect 9234 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 9854 370894
rect 9234 370574 9854 370658
rect 9234 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 9854 370574
rect 9234 334894 9854 370338
rect 9234 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 9854 334894
rect 9234 334574 9854 334658
rect 9234 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 9854 334574
rect 9234 298894 9854 334338
rect 9234 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 9854 298894
rect 9234 298574 9854 298658
rect 9234 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 9854 298574
rect 9234 262894 9854 298338
rect 9234 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 9854 262894
rect 9234 262574 9854 262658
rect 9234 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 9854 262574
rect 9234 226894 9854 262338
rect 9234 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 9854 226894
rect 9234 226574 9854 226658
rect 9234 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 9854 226574
rect 9234 190894 9854 226338
rect 9234 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 9854 190894
rect 9234 190574 9854 190658
rect 9234 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 9854 190574
rect 9234 154894 9854 190338
rect 9234 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 9854 154894
rect 9234 154574 9854 154658
rect 9234 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 9854 154574
rect 9234 118894 9854 154338
rect 9234 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 9854 118894
rect 9234 118574 9854 118658
rect 9234 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 9854 118574
rect 9234 82894 9854 118338
rect 9234 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 9854 82894
rect 9234 82574 9854 82658
rect 9234 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 9854 82574
rect 9234 46894 9854 82338
rect 9234 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 9854 46894
rect 9234 46574 9854 46658
rect 9234 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 9854 46574
rect 9234 10894 9854 46338
rect 9234 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 9854 10894
rect 9234 10574 9854 10658
rect 9234 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 9854 10574
rect 9234 -2266 9854 10338
rect 9234 -2502 9266 -2266
rect 9502 -2502 9586 -2266
rect 9822 -2502 9854 -2266
rect 9234 -2586 9854 -2502
rect 9234 -2822 9266 -2586
rect 9502 -2822 9586 -2586
rect 9822 -2822 9854 -2586
rect 9234 -7654 9854 -2822
rect 12954 707718 13574 711590
rect 12954 707482 12986 707718
rect 13222 707482 13306 707718
rect 13542 707482 13574 707718
rect 12954 707398 13574 707482
rect 12954 707162 12986 707398
rect 13222 707162 13306 707398
rect 13542 707162 13574 707398
rect 12954 698614 13574 707162
rect 12954 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 13574 698614
rect 12954 698294 13574 698378
rect 12954 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 13574 698294
rect 12954 662614 13574 698058
rect 12954 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 13574 662614
rect 12954 662294 13574 662378
rect 12954 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 13574 662294
rect 12954 626614 13574 662058
rect 12954 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 13574 626614
rect 12954 626294 13574 626378
rect 12954 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 13574 626294
rect 12954 590614 13574 626058
rect 12954 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 13574 590614
rect 12954 590294 13574 590378
rect 12954 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 13574 590294
rect 12954 554614 13574 590058
rect 12954 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 13574 554614
rect 12954 554294 13574 554378
rect 12954 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 13574 554294
rect 12954 518614 13574 554058
rect 12954 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 13574 518614
rect 12954 518294 13574 518378
rect 12954 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 13574 518294
rect 12954 482614 13574 518058
rect 12954 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 13574 482614
rect 12954 482294 13574 482378
rect 12954 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 13574 482294
rect 12954 446614 13574 482058
rect 12954 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 13574 446614
rect 12954 446294 13574 446378
rect 12954 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 13574 446294
rect 12954 410614 13574 446058
rect 12954 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 13574 410614
rect 12954 410294 13574 410378
rect 12954 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 13574 410294
rect 12954 374614 13574 410058
rect 12954 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 13574 374614
rect 12954 374294 13574 374378
rect 12954 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 13574 374294
rect 12954 338614 13574 374058
rect 12954 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 13574 338614
rect 12954 338294 13574 338378
rect 12954 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 13574 338294
rect 12954 302614 13574 338058
rect 12954 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 13574 302614
rect 12954 302294 13574 302378
rect 12954 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 13574 302294
rect 12954 266614 13574 302058
rect 12954 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 13574 266614
rect 12954 266294 13574 266378
rect 12954 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 13574 266294
rect 12954 230614 13574 266058
rect 12954 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 13574 230614
rect 12954 230294 13574 230378
rect 12954 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 13574 230294
rect 12954 194614 13574 230058
rect 12954 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 13574 194614
rect 12954 194294 13574 194378
rect 12954 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 13574 194294
rect 12954 158614 13574 194058
rect 12954 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 13574 158614
rect 12954 158294 13574 158378
rect 12954 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 13574 158294
rect 12954 122614 13574 158058
rect 12954 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 13574 122614
rect 12954 122294 13574 122378
rect 12954 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 13574 122294
rect 12954 86614 13574 122058
rect 12954 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 13574 86614
rect 12954 86294 13574 86378
rect 12954 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 13574 86294
rect 12954 50614 13574 86058
rect 12954 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 13574 50614
rect 12954 50294 13574 50378
rect 12954 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 13574 50294
rect 12954 14614 13574 50058
rect 12954 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 13574 14614
rect 12954 14294 13574 14378
rect 12954 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 13574 14294
rect 12954 -3226 13574 14058
rect 12954 -3462 12986 -3226
rect 13222 -3462 13306 -3226
rect 13542 -3462 13574 -3226
rect 12954 -3546 13574 -3462
rect 12954 -3782 12986 -3546
rect 13222 -3782 13306 -3546
rect 13542 -3782 13574 -3546
rect 12954 -7654 13574 -3782
rect 16674 708678 17294 711590
rect 16674 708442 16706 708678
rect 16942 708442 17026 708678
rect 17262 708442 17294 708678
rect 16674 708358 17294 708442
rect 16674 708122 16706 708358
rect 16942 708122 17026 708358
rect 17262 708122 17294 708358
rect 16674 666334 17294 708122
rect 16674 666098 16706 666334
rect 16942 666098 17026 666334
rect 17262 666098 17294 666334
rect 16674 666014 17294 666098
rect 16674 665778 16706 666014
rect 16942 665778 17026 666014
rect 17262 665778 17294 666014
rect 16674 630334 17294 665778
rect 16674 630098 16706 630334
rect 16942 630098 17026 630334
rect 17262 630098 17294 630334
rect 16674 630014 17294 630098
rect 16674 629778 16706 630014
rect 16942 629778 17026 630014
rect 17262 629778 17294 630014
rect 16674 594334 17294 629778
rect 16674 594098 16706 594334
rect 16942 594098 17026 594334
rect 17262 594098 17294 594334
rect 16674 594014 17294 594098
rect 16674 593778 16706 594014
rect 16942 593778 17026 594014
rect 17262 593778 17294 594014
rect 16674 558334 17294 593778
rect 16674 558098 16706 558334
rect 16942 558098 17026 558334
rect 17262 558098 17294 558334
rect 16674 558014 17294 558098
rect 16674 557778 16706 558014
rect 16942 557778 17026 558014
rect 17262 557778 17294 558014
rect 16674 522334 17294 557778
rect 16674 522098 16706 522334
rect 16942 522098 17026 522334
rect 17262 522098 17294 522334
rect 16674 522014 17294 522098
rect 16674 521778 16706 522014
rect 16942 521778 17026 522014
rect 17262 521778 17294 522014
rect 16674 486334 17294 521778
rect 16674 486098 16706 486334
rect 16942 486098 17026 486334
rect 17262 486098 17294 486334
rect 16674 486014 17294 486098
rect 16674 485778 16706 486014
rect 16942 485778 17026 486014
rect 17262 485778 17294 486014
rect 16674 450334 17294 485778
rect 16674 450098 16706 450334
rect 16942 450098 17026 450334
rect 17262 450098 17294 450334
rect 16674 450014 17294 450098
rect 16674 449778 16706 450014
rect 16942 449778 17026 450014
rect 17262 449778 17294 450014
rect 16674 414334 17294 449778
rect 16674 414098 16706 414334
rect 16942 414098 17026 414334
rect 17262 414098 17294 414334
rect 16674 414014 17294 414098
rect 16674 413778 16706 414014
rect 16942 413778 17026 414014
rect 17262 413778 17294 414014
rect 16674 378334 17294 413778
rect 16674 378098 16706 378334
rect 16942 378098 17026 378334
rect 17262 378098 17294 378334
rect 16674 378014 17294 378098
rect 16674 377778 16706 378014
rect 16942 377778 17026 378014
rect 17262 377778 17294 378014
rect 16674 342334 17294 377778
rect 16674 342098 16706 342334
rect 16942 342098 17026 342334
rect 17262 342098 17294 342334
rect 16674 342014 17294 342098
rect 16674 341778 16706 342014
rect 16942 341778 17026 342014
rect 17262 341778 17294 342014
rect 16674 306334 17294 341778
rect 16674 306098 16706 306334
rect 16942 306098 17026 306334
rect 17262 306098 17294 306334
rect 16674 306014 17294 306098
rect 16674 305778 16706 306014
rect 16942 305778 17026 306014
rect 17262 305778 17294 306014
rect 16674 270334 17294 305778
rect 16674 270098 16706 270334
rect 16942 270098 17026 270334
rect 17262 270098 17294 270334
rect 16674 270014 17294 270098
rect 16674 269778 16706 270014
rect 16942 269778 17026 270014
rect 17262 269778 17294 270014
rect 16674 234334 17294 269778
rect 16674 234098 16706 234334
rect 16942 234098 17026 234334
rect 17262 234098 17294 234334
rect 16674 234014 17294 234098
rect 16674 233778 16706 234014
rect 16942 233778 17026 234014
rect 17262 233778 17294 234014
rect 16674 198334 17294 233778
rect 16674 198098 16706 198334
rect 16942 198098 17026 198334
rect 17262 198098 17294 198334
rect 16674 198014 17294 198098
rect 16674 197778 16706 198014
rect 16942 197778 17026 198014
rect 17262 197778 17294 198014
rect 16674 162334 17294 197778
rect 16674 162098 16706 162334
rect 16942 162098 17026 162334
rect 17262 162098 17294 162334
rect 16674 162014 17294 162098
rect 16674 161778 16706 162014
rect 16942 161778 17026 162014
rect 17262 161778 17294 162014
rect 16674 126334 17294 161778
rect 16674 126098 16706 126334
rect 16942 126098 17026 126334
rect 17262 126098 17294 126334
rect 16674 126014 17294 126098
rect 16674 125778 16706 126014
rect 16942 125778 17026 126014
rect 17262 125778 17294 126014
rect 16674 90334 17294 125778
rect 16674 90098 16706 90334
rect 16942 90098 17026 90334
rect 17262 90098 17294 90334
rect 16674 90014 17294 90098
rect 16674 89778 16706 90014
rect 16942 89778 17026 90014
rect 17262 89778 17294 90014
rect 16674 54334 17294 89778
rect 16674 54098 16706 54334
rect 16942 54098 17026 54334
rect 17262 54098 17294 54334
rect 16674 54014 17294 54098
rect 16674 53778 16706 54014
rect 16942 53778 17026 54014
rect 17262 53778 17294 54014
rect 16674 18334 17294 53778
rect 16674 18098 16706 18334
rect 16942 18098 17026 18334
rect 17262 18098 17294 18334
rect 16674 18014 17294 18098
rect 16674 17778 16706 18014
rect 16942 17778 17026 18014
rect 17262 17778 17294 18014
rect 16674 -4186 17294 17778
rect 16674 -4422 16706 -4186
rect 16942 -4422 17026 -4186
rect 17262 -4422 17294 -4186
rect 16674 -4506 17294 -4422
rect 16674 -4742 16706 -4506
rect 16942 -4742 17026 -4506
rect 17262 -4742 17294 -4506
rect 16674 -7654 17294 -4742
rect 20394 709638 21014 711590
rect 20394 709402 20426 709638
rect 20662 709402 20746 709638
rect 20982 709402 21014 709638
rect 20394 709318 21014 709402
rect 20394 709082 20426 709318
rect 20662 709082 20746 709318
rect 20982 709082 21014 709318
rect 20394 670054 21014 709082
rect 20394 669818 20426 670054
rect 20662 669818 20746 670054
rect 20982 669818 21014 670054
rect 20394 669734 21014 669818
rect 20394 669498 20426 669734
rect 20662 669498 20746 669734
rect 20982 669498 21014 669734
rect 20394 634054 21014 669498
rect 27834 711558 28454 711590
rect 27834 711322 27866 711558
rect 28102 711322 28186 711558
rect 28422 711322 28454 711558
rect 27834 711238 28454 711322
rect 27834 711002 27866 711238
rect 28102 711002 28186 711238
rect 28422 711002 28454 711238
rect 27834 677494 28454 711002
rect 27834 677258 27866 677494
rect 28102 677258 28186 677494
rect 28422 677258 28454 677494
rect 27834 677174 28454 677258
rect 27834 676938 27866 677174
rect 28102 676938 28186 677174
rect 28422 676938 28454 677174
rect 24208 651454 24528 651486
rect 24208 651218 24250 651454
rect 24486 651218 24528 651454
rect 24208 651134 24528 651218
rect 24208 650898 24250 651134
rect 24486 650898 24528 651134
rect 24208 650866 24528 650898
rect 20394 633818 20426 634054
rect 20662 633818 20746 634054
rect 20982 633818 21014 634054
rect 20394 633734 21014 633818
rect 20394 633498 20426 633734
rect 20662 633498 20746 633734
rect 20982 633498 21014 633734
rect 20394 598054 21014 633498
rect 27834 641494 28454 676938
rect 37794 704838 38414 711590
rect 37794 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 38414 704838
rect 37794 704518 38414 704602
rect 37794 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 38414 704518
rect 37794 687454 38414 704282
rect 37794 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 38414 687454
rect 37794 687134 38414 687218
rect 37794 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 38414 687134
rect 37794 674393 38414 686898
rect 41514 705798 42134 711590
rect 41514 705562 41546 705798
rect 41782 705562 41866 705798
rect 42102 705562 42134 705798
rect 41514 705478 42134 705562
rect 41514 705242 41546 705478
rect 41782 705242 41866 705478
rect 42102 705242 42134 705478
rect 41514 691174 42134 705242
rect 41514 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 42134 691174
rect 41514 690854 42134 690938
rect 41514 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 42134 690854
rect 41514 674393 42134 690618
rect 45234 706758 45854 711590
rect 45234 706522 45266 706758
rect 45502 706522 45586 706758
rect 45822 706522 45854 706758
rect 45234 706438 45854 706522
rect 45234 706202 45266 706438
rect 45502 706202 45586 706438
rect 45822 706202 45854 706438
rect 45234 694894 45854 706202
rect 45234 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 45854 694894
rect 45234 694574 45854 694658
rect 45234 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 45854 694574
rect 45234 674393 45854 694338
rect 48954 707718 49574 711590
rect 48954 707482 48986 707718
rect 49222 707482 49306 707718
rect 49542 707482 49574 707718
rect 48954 707398 49574 707482
rect 48954 707162 48986 707398
rect 49222 707162 49306 707398
rect 49542 707162 49574 707398
rect 48954 698614 49574 707162
rect 48954 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 49574 698614
rect 48954 698294 49574 698378
rect 48954 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 49574 698294
rect 48954 674393 49574 698058
rect 63834 711558 64454 711590
rect 63834 711322 63866 711558
rect 64102 711322 64186 711558
rect 64422 711322 64454 711558
rect 63834 711238 64454 711322
rect 63834 711002 63866 711238
rect 64102 711002 64186 711238
rect 64422 711002 64454 711238
rect 63834 677494 64454 711002
rect 63834 677258 63866 677494
rect 64102 677258 64186 677494
rect 64422 677258 64454 677494
rect 63834 677174 64454 677258
rect 63834 676938 63866 677174
rect 64102 676938 64186 677174
rect 64422 676938 64454 677174
rect 63834 674393 64454 676938
rect 73794 704838 74414 711590
rect 73794 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 74414 704838
rect 73794 704518 74414 704602
rect 73794 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 74414 704518
rect 73794 687454 74414 704282
rect 73794 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 74414 687454
rect 73794 687134 74414 687218
rect 73794 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 74414 687134
rect 73794 674393 74414 686898
rect 77514 705798 78134 711590
rect 77514 705562 77546 705798
rect 77782 705562 77866 705798
rect 78102 705562 78134 705798
rect 77514 705478 78134 705562
rect 77514 705242 77546 705478
rect 77782 705242 77866 705478
rect 78102 705242 78134 705478
rect 77514 691174 78134 705242
rect 77514 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 78134 691174
rect 77514 690854 78134 690938
rect 77514 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 78134 690854
rect 77514 674393 78134 690618
rect 81234 706758 81854 711590
rect 81234 706522 81266 706758
rect 81502 706522 81586 706758
rect 81822 706522 81854 706758
rect 81234 706438 81854 706522
rect 81234 706202 81266 706438
rect 81502 706202 81586 706438
rect 81822 706202 81854 706438
rect 81234 694894 81854 706202
rect 81234 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 81854 694894
rect 81234 694574 81854 694658
rect 81234 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 81854 694574
rect 81234 674393 81854 694338
rect 84954 707718 85574 711590
rect 84954 707482 84986 707718
rect 85222 707482 85306 707718
rect 85542 707482 85574 707718
rect 84954 707398 85574 707482
rect 84954 707162 84986 707398
rect 85222 707162 85306 707398
rect 85542 707162 85574 707398
rect 84954 698614 85574 707162
rect 84954 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 85574 698614
rect 84954 698294 85574 698378
rect 84954 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 85574 698294
rect 84954 674393 85574 698058
rect 99834 711558 100454 711590
rect 99834 711322 99866 711558
rect 100102 711322 100186 711558
rect 100422 711322 100454 711558
rect 99834 711238 100454 711322
rect 99834 711002 99866 711238
rect 100102 711002 100186 711238
rect 100422 711002 100454 711238
rect 99834 677494 100454 711002
rect 99834 677258 99866 677494
rect 100102 677258 100186 677494
rect 100422 677258 100454 677494
rect 99834 677174 100454 677258
rect 99834 676938 99866 677174
rect 100102 676938 100186 677174
rect 100422 676938 100454 677174
rect 99834 674393 100454 676938
rect 109794 704838 110414 711590
rect 109794 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 110414 704838
rect 109794 704518 110414 704602
rect 109794 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 110414 704518
rect 109794 687454 110414 704282
rect 109794 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 110414 687454
rect 109794 687134 110414 687218
rect 109794 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 110414 687134
rect 109794 674393 110414 686898
rect 113514 705798 114134 711590
rect 113514 705562 113546 705798
rect 113782 705562 113866 705798
rect 114102 705562 114134 705798
rect 113514 705478 114134 705562
rect 113514 705242 113546 705478
rect 113782 705242 113866 705478
rect 114102 705242 114134 705478
rect 113514 691174 114134 705242
rect 113514 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 114134 691174
rect 113514 690854 114134 690938
rect 113514 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 114134 690854
rect 113514 674393 114134 690618
rect 117234 706758 117854 711590
rect 117234 706522 117266 706758
rect 117502 706522 117586 706758
rect 117822 706522 117854 706758
rect 117234 706438 117854 706522
rect 117234 706202 117266 706438
rect 117502 706202 117586 706438
rect 117822 706202 117854 706438
rect 117234 694894 117854 706202
rect 117234 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 117854 694894
rect 117234 694574 117854 694658
rect 117234 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 117854 694574
rect 117234 674393 117854 694338
rect 120954 707718 121574 711590
rect 120954 707482 120986 707718
rect 121222 707482 121306 707718
rect 121542 707482 121574 707718
rect 120954 707398 121574 707482
rect 120954 707162 120986 707398
rect 121222 707162 121306 707398
rect 121542 707162 121574 707398
rect 120954 698614 121574 707162
rect 120954 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 121574 698614
rect 120954 698294 121574 698378
rect 120954 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 121574 698294
rect 120954 674393 121574 698058
rect 135834 711558 136454 711590
rect 135834 711322 135866 711558
rect 136102 711322 136186 711558
rect 136422 711322 136454 711558
rect 135834 711238 136454 711322
rect 135834 711002 135866 711238
rect 136102 711002 136186 711238
rect 136422 711002 136454 711238
rect 135834 677494 136454 711002
rect 135834 677258 135866 677494
rect 136102 677258 136186 677494
rect 136422 677258 136454 677494
rect 135834 677174 136454 677258
rect 135834 676938 135866 677174
rect 136102 676938 136186 677174
rect 136422 676938 136454 677174
rect 135834 674393 136454 676938
rect 145794 704838 146414 711590
rect 145794 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 146414 704838
rect 145794 704518 146414 704602
rect 145794 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 146414 704518
rect 145794 687454 146414 704282
rect 145794 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 146414 687454
rect 145794 687134 146414 687218
rect 145794 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 146414 687134
rect 145794 674393 146414 686898
rect 149514 705798 150134 711590
rect 149514 705562 149546 705798
rect 149782 705562 149866 705798
rect 150102 705562 150134 705798
rect 149514 705478 150134 705562
rect 149514 705242 149546 705478
rect 149782 705242 149866 705478
rect 150102 705242 150134 705478
rect 149514 691174 150134 705242
rect 149514 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 150134 691174
rect 149514 690854 150134 690938
rect 149514 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 150134 690854
rect 149514 674393 150134 690618
rect 153234 706758 153854 711590
rect 153234 706522 153266 706758
rect 153502 706522 153586 706758
rect 153822 706522 153854 706758
rect 153234 706438 153854 706522
rect 153234 706202 153266 706438
rect 153502 706202 153586 706438
rect 153822 706202 153854 706438
rect 153234 694894 153854 706202
rect 153234 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 153854 694894
rect 153234 694574 153854 694658
rect 153234 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 153854 694574
rect 153234 674393 153854 694338
rect 156954 707718 157574 711590
rect 156954 707482 156986 707718
rect 157222 707482 157306 707718
rect 157542 707482 157574 707718
rect 156954 707398 157574 707482
rect 156954 707162 156986 707398
rect 157222 707162 157306 707398
rect 157542 707162 157574 707398
rect 156954 698614 157574 707162
rect 156954 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 157574 698614
rect 156954 698294 157574 698378
rect 156954 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 157574 698294
rect 156954 674393 157574 698058
rect 171834 711558 172454 711590
rect 171834 711322 171866 711558
rect 172102 711322 172186 711558
rect 172422 711322 172454 711558
rect 171834 711238 172454 711322
rect 171834 711002 171866 711238
rect 172102 711002 172186 711238
rect 172422 711002 172454 711238
rect 171834 677494 172454 711002
rect 171834 677258 171866 677494
rect 172102 677258 172186 677494
rect 172422 677258 172454 677494
rect 171834 677174 172454 677258
rect 171834 676938 171866 677174
rect 172102 676938 172186 677174
rect 172422 676938 172454 677174
rect 171834 674393 172454 676938
rect 181794 704838 182414 711590
rect 181794 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 182414 704838
rect 181794 704518 182414 704602
rect 181794 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 182414 704518
rect 181794 687454 182414 704282
rect 181794 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 182414 687454
rect 181794 687134 182414 687218
rect 181794 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 182414 687134
rect 181794 674393 182414 686898
rect 185514 705798 186134 711590
rect 185514 705562 185546 705798
rect 185782 705562 185866 705798
rect 186102 705562 186134 705798
rect 185514 705478 186134 705562
rect 185514 705242 185546 705478
rect 185782 705242 185866 705478
rect 186102 705242 186134 705478
rect 185514 691174 186134 705242
rect 185514 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 186134 691174
rect 185514 690854 186134 690938
rect 185514 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 186134 690854
rect 185514 674393 186134 690618
rect 189234 706758 189854 711590
rect 189234 706522 189266 706758
rect 189502 706522 189586 706758
rect 189822 706522 189854 706758
rect 189234 706438 189854 706522
rect 189234 706202 189266 706438
rect 189502 706202 189586 706438
rect 189822 706202 189854 706438
rect 189234 694894 189854 706202
rect 189234 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 189854 694894
rect 189234 694574 189854 694658
rect 189234 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 189854 694574
rect 189234 674393 189854 694338
rect 192954 707718 193574 711590
rect 192954 707482 192986 707718
rect 193222 707482 193306 707718
rect 193542 707482 193574 707718
rect 192954 707398 193574 707482
rect 192954 707162 192986 707398
rect 193222 707162 193306 707398
rect 193542 707162 193574 707398
rect 192954 698614 193574 707162
rect 192954 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 193574 698614
rect 192954 698294 193574 698378
rect 192954 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 193574 698294
rect 192954 684676 193574 698058
rect 207834 711558 208454 711590
rect 207834 711322 207866 711558
rect 208102 711322 208186 711558
rect 208422 711322 208454 711558
rect 207834 711238 208454 711322
rect 207834 711002 207866 711238
rect 208102 711002 208186 711238
rect 208422 711002 208454 711238
rect 207834 677494 208454 711002
rect 207834 677258 207866 677494
rect 208102 677258 208186 677494
rect 208422 677258 208454 677494
rect 207834 677174 208454 677258
rect 207834 676938 207866 677174
rect 208102 676938 208186 677174
rect 208422 676938 208454 677174
rect 207834 674393 208454 676938
rect 217794 704838 218414 711590
rect 217794 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 218414 704838
rect 217794 704518 218414 704602
rect 217794 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 218414 704518
rect 217794 687454 218414 704282
rect 217794 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 218414 687454
rect 217794 687134 218414 687218
rect 217794 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 218414 687134
rect 217794 674393 218414 686898
rect 221514 705798 222134 711590
rect 221514 705562 221546 705798
rect 221782 705562 221866 705798
rect 222102 705562 222134 705798
rect 221514 705478 222134 705562
rect 221514 705242 221546 705478
rect 221782 705242 221866 705478
rect 222102 705242 222134 705478
rect 221514 691174 222134 705242
rect 221514 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 222134 691174
rect 221514 690854 222134 690938
rect 221514 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 222134 690854
rect 221514 674393 222134 690618
rect 225234 706758 225854 711590
rect 225234 706522 225266 706758
rect 225502 706522 225586 706758
rect 225822 706522 225854 706758
rect 225234 706438 225854 706522
rect 225234 706202 225266 706438
rect 225502 706202 225586 706438
rect 225822 706202 225854 706438
rect 225234 694894 225854 706202
rect 225234 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 225854 694894
rect 225234 694574 225854 694658
rect 225234 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 225854 694574
rect 225234 674393 225854 694338
rect 228954 707718 229574 711590
rect 228954 707482 228986 707718
rect 229222 707482 229306 707718
rect 229542 707482 229574 707718
rect 228954 707398 229574 707482
rect 228954 707162 228986 707398
rect 229222 707162 229306 707398
rect 229542 707162 229574 707398
rect 228954 698614 229574 707162
rect 228954 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 229574 698614
rect 228954 698294 229574 698378
rect 228954 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 229574 698294
rect 228954 674393 229574 698058
rect 243834 711558 244454 711590
rect 243834 711322 243866 711558
rect 244102 711322 244186 711558
rect 244422 711322 244454 711558
rect 243834 711238 244454 711322
rect 243834 711002 243866 711238
rect 244102 711002 244186 711238
rect 244422 711002 244454 711238
rect 243834 677494 244454 711002
rect 243834 677258 243866 677494
rect 244102 677258 244186 677494
rect 244422 677258 244454 677494
rect 243834 677174 244454 677258
rect 243834 676938 243866 677174
rect 244102 676938 244186 677174
rect 244422 676938 244454 677174
rect 243834 674393 244454 676938
rect 253794 704838 254414 711590
rect 253794 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 254414 704838
rect 253794 704518 254414 704602
rect 253794 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 254414 704518
rect 253794 687454 254414 704282
rect 253794 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 254414 687454
rect 253794 687134 254414 687218
rect 253794 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 254414 687134
rect 253794 674393 254414 686898
rect 257514 705798 258134 711590
rect 257514 705562 257546 705798
rect 257782 705562 257866 705798
rect 258102 705562 258134 705798
rect 257514 705478 258134 705562
rect 257514 705242 257546 705478
rect 257782 705242 257866 705478
rect 258102 705242 258134 705478
rect 257514 691174 258134 705242
rect 257514 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 258134 691174
rect 257514 690854 258134 690938
rect 257514 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 258134 690854
rect 257514 674393 258134 690618
rect 261234 706758 261854 711590
rect 261234 706522 261266 706758
rect 261502 706522 261586 706758
rect 261822 706522 261854 706758
rect 261234 706438 261854 706522
rect 261234 706202 261266 706438
rect 261502 706202 261586 706438
rect 261822 706202 261854 706438
rect 261234 694894 261854 706202
rect 261234 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 261854 694894
rect 261234 694574 261854 694658
rect 261234 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 261854 694574
rect 261234 674393 261854 694338
rect 264954 707718 265574 711590
rect 264954 707482 264986 707718
rect 265222 707482 265306 707718
rect 265542 707482 265574 707718
rect 264954 707398 265574 707482
rect 264954 707162 264986 707398
rect 265222 707162 265306 707398
rect 265542 707162 265574 707398
rect 264954 698614 265574 707162
rect 264954 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 265574 698614
rect 264954 698294 265574 698378
rect 264954 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 265574 698294
rect 264954 674393 265574 698058
rect 279834 711558 280454 711590
rect 279834 711322 279866 711558
rect 280102 711322 280186 711558
rect 280422 711322 280454 711558
rect 279834 711238 280454 711322
rect 279834 711002 279866 711238
rect 280102 711002 280186 711238
rect 280422 711002 280454 711238
rect 279834 677494 280454 711002
rect 279834 677258 279866 677494
rect 280102 677258 280186 677494
rect 280422 677258 280454 677494
rect 279834 677174 280454 677258
rect 279834 676938 279866 677174
rect 280102 676938 280186 677174
rect 280422 676938 280454 677174
rect 279834 674393 280454 676938
rect 289794 704838 290414 711590
rect 289794 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 290414 704838
rect 289794 704518 290414 704602
rect 289794 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 290414 704518
rect 289794 687454 290414 704282
rect 289794 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 290414 687454
rect 289794 687134 290414 687218
rect 289794 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 290414 687134
rect 289794 674393 290414 686898
rect 293514 705798 294134 711590
rect 293514 705562 293546 705798
rect 293782 705562 293866 705798
rect 294102 705562 294134 705798
rect 293514 705478 294134 705562
rect 293514 705242 293546 705478
rect 293782 705242 293866 705478
rect 294102 705242 294134 705478
rect 293514 691174 294134 705242
rect 293514 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 294134 691174
rect 293514 690854 294134 690938
rect 293514 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 294134 690854
rect 293514 674393 294134 690618
rect 297234 706758 297854 711590
rect 297234 706522 297266 706758
rect 297502 706522 297586 706758
rect 297822 706522 297854 706758
rect 297234 706438 297854 706522
rect 297234 706202 297266 706438
rect 297502 706202 297586 706438
rect 297822 706202 297854 706438
rect 297234 694894 297854 706202
rect 297234 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 297854 694894
rect 297234 694574 297854 694658
rect 297234 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 297854 694574
rect 297234 674393 297854 694338
rect 300954 707718 301574 711590
rect 300954 707482 300986 707718
rect 301222 707482 301306 707718
rect 301542 707482 301574 707718
rect 300954 707398 301574 707482
rect 300954 707162 300986 707398
rect 301222 707162 301306 707398
rect 301542 707162 301574 707398
rect 300954 698614 301574 707162
rect 300954 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 301574 698614
rect 300954 698294 301574 698378
rect 300954 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 301574 698294
rect 300954 684676 301574 698058
rect 325794 704838 326414 711590
rect 325794 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 326414 704838
rect 325794 704518 326414 704602
rect 325794 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 326414 704518
rect 325794 687454 326414 704282
rect 325794 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 326414 687454
rect 325794 687134 326414 687218
rect 325794 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 326414 687134
rect 325794 674393 326414 686898
rect 329514 705798 330134 711590
rect 329514 705562 329546 705798
rect 329782 705562 329866 705798
rect 330102 705562 330134 705798
rect 329514 705478 330134 705562
rect 329514 705242 329546 705478
rect 329782 705242 329866 705478
rect 330102 705242 330134 705478
rect 329514 691174 330134 705242
rect 329514 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 330134 691174
rect 329514 690854 330134 690938
rect 329514 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 330134 690854
rect 329514 674393 330134 690618
rect 333234 706758 333854 711590
rect 333234 706522 333266 706758
rect 333502 706522 333586 706758
rect 333822 706522 333854 706758
rect 333234 706438 333854 706522
rect 333234 706202 333266 706438
rect 333502 706202 333586 706438
rect 333822 706202 333854 706438
rect 333234 694894 333854 706202
rect 333234 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 333854 694894
rect 333234 694574 333854 694658
rect 333234 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 333854 694574
rect 333234 674393 333854 694338
rect 336954 707718 337574 711590
rect 336954 707482 336986 707718
rect 337222 707482 337306 707718
rect 337542 707482 337574 707718
rect 336954 707398 337574 707482
rect 336954 707162 336986 707398
rect 337222 707162 337306 707398
rect 337542 707162 337574 707398
rect 336954 698614 337574 707162
rect 336954 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 337574 698614
rect 336954 698294 337574 698378
rect 336954 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 337574 698294
rect 336954 674393 337574 698058
rect 351834 711558 352454 711590
rect 351834 711322 351866 711558
rect 352102 711322 352186 711558
rect 352422 711322 352454 711558
rect 351834 711238 352454 711322
rect 351834 711002 351866 711238
rect 352102 711002 352186 711238
rect 352422 711002 352454 711238
rect 351834 677494 352454 711002
rect 351834 677258 351866 677494
rect 352102 677258 352186 677494
rect 352422 677258 352454 677494
rect 351834 677174 352454 677258
rect 351834 676938 351866 677174
rect 352102 676938 352186 677174
rect 352422 676938 352454 677174
rect 351834 674393 352454 676938
rect 361794 704838 362414 711590
rect 361794 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 362414 704838
rect 361794 704518 362414 704602
rect 361794 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 362414 704518
rect 361794 687454 362414 704282
rect 361794 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 362414 687454
rect 361794 687134 362414 687218
rect 361794 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 362414 687134
rect 39568 655174 39888 655206
rect 39568 654938 39610 655174
rect 39846 654938 39888 655174
rect 39568 654854 39888 654938
rect 39568 654618 39610 654854
rect 39846 654618 39888 654854
rect 39568 654586 39888 654618
rect 70288 655174 70608 655206
rect 70288 654938 70330 655174
rect 70566 654938 70608 655174
rect 70288 654854 70608 654938
rect 70288 654618 70330 654854
rect 70566 654618 70608 654854
rect 70288 654586 70608 654618
rect 101008 655174 101328 655206
rect 101008 654938 101050 655174
rect 101286 654938 101328 655174
rect 101008 654854 101328 654938
rect 101008 654618 101050 654854
rect 101286 654618 101328 654854
rect 101008 654586 101328 654618
rect 131728 655174 132048 655206
rect 131728 654938 131770 655174
rect 132006 654938 132048 655174
rect 131728 654854 132048 654938
rect 131728 654618 131770 654854
rect 132006 654618 132048 654854
rect 131728 654586 132048 654618
rect 162448 655174 162768 655206
rect 162448 654938 162490 655174
rect 162726 654938 162768 655174
rect 162448 654854 162768 654938
rect 162448 654618 162490 654854
rect 162726 654618 162768 654854
rect 162448 654586 162768 654618
rect 193168 655174 193488 655206
rect 193168 654938 193210 655174
rect 193446 654938 193488 655174
rect 193168 654854 193488 654938
rect 193168 654618 193210 654854
rect 193446 654618 193488 654854
rect 193168 654586 193488 654618
rect 223888 655174 224208 655206
rect 223888 654938 223930 655174
rect 224166 654938 224208 655174
rect 223888 654854 224208 654938
rect 223888 654618 223930 654854
rect 224166 654618 224208 654854
rect 223888 654586 224208 654618
rect 254608 655174 254928 655206
rect 254608 654938 254650 655174
rect 254886 654938 254928 655174
rect 254608 654854 254928 654938
rect 254608 654618 254650 654854
rect 254886 654618 254928 654854
rect 254608 654586 254928 654618
rect 285328 655174 285648 655206
rect 285328 654938 285370 655174
rect 285606 654938 285648 655174
rect 285328 654854 285648 654938
rect 285328 654618 285370 654854
rect 285606 654618 285648 654854
rect 285328 654586 285648 654618
rect 316048 655174 316368 655206
rect 316048 654938 316090 655174
rect 316326 654938 316368 655174
rect 316048 654854 316368 654938
rect 316048 654618 316090 654854
rect 316326 654618 316368 654854
rect 316048 654586 316368 654618
rect 346768 655174 347088 655206
rect 346768 654938 346810 655174
rect 347046 654938 347088 655174
rect 346768 654854 347088 654938
rect 346768 654618 346810 654854
rect 347046 654618 347088 654854
rect 346768 654586 347088 654618
rect 54928 651454 55248 651486
rect 54928 651218 54970 651454
rect 55206 651218 55248 651454
rect 54928 651134 55248 651218
rect 54928 650898 54970 651134
rect 55206 650898 55248 651134
rect 54928 650866 55248 650898
rect 85648 651454 85968 651486
rect 85648 651218 85690 651454
rect 85926 651218 85968 651454
rect 85648 651134 85968 651218
rect 85648 650898 85690 651134
rect 85926 650898 85968 651134
rect 85648 650866 85968 650898
rect 116368 651454 116688 651486
rect 116368 651218 116410 651454
rect 116646 651218 116688 651454
rect 116368 651134 116688 651218
rect 116368 650898 116410 651134
rect 116646 650898 116688 651134
rect 116368 650866 116688 650898
rect 147088 651454 147408 651486
rect 147088 651218 147130 651454
rect 147366 651218 147408 651454
rect 147088 651134 147408 651218
rect 147088 650898 147130 651134
rect 147366 650898 147408 651134
rect 147088 650866 147408 650898
rect 177808 651454 178128 651486
rect 177808 651218 177850 651454
rect 178086 651218 178128 651454
rect 177808 651134 178128 651218
rect 177808 650898 177850 651134
rect 178086 650898 178128 651134
rect 177808 650866 178128 650898
rect 208528 651454 208848 651486
rect 208528 651218 208570 651454
rect 208806 651218 208848 651454
rect 208528 651134 208848 651218
rect 208528 650898 208570 651134
rect 208806 650898 208848 651134
rect 208528 650866 208848 650898
rect 239248 651454 239568 651486
rect 239248 651218 239290 651454
rect 239526 651218 239568 651454
rect 239248 651134 239568 651218
rect 239248 650898 239290 651134
rect 239526 650898 239568 651134
rect 239248 650866 239568 650898
rect 269968 651454 270288 651486
rect 269968 651218 270010 651454
rect 270246 651218 270288 651454
rect 269968 651134 270288 651218
rect 269968 650898 270010 651134
rect 270246 650898 270288 651134
rect 269968 650866 270288 650898
rect 300688 651454 301008 651486
rect 300688 651218 300730 651454
rect 300966 651218 301008 651454
rect 300688 651134 301008 651218
rect 300688 650898 300730 651134
rect 300966 650898 301008 651134
rect 300688 650866 301008 650898
rect 331408 651454 331728 651486
rect 331408 651218 331450 651454
rect 331686 651218 331728 651454
rect 331408 651134 331728 651218
rect 331408 650898 331450 651134
rect 331686 650898 331728 651134
rect 331408 650866 331728 650898
rect 361794 651454 362414 686898
rect 361794 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 362414 651454
rect 361794 651134 362414 651218
rect 361794 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 362414 651134
rect 27834 641258 27866 641494
rect 28102 641258 28186 641494
rect 28422 641258 28454 641494
rect 27834 641174 28454 641258
rect 27834 640938 27866 641174
rect 28102 640938 28186 641174
rect 28422 640938 28454 641174
rect 24208 615454 24528 615486
rect 24208 615218 24250 615454
rect 24486 615218 24528 615454
rect 24208 615134 24528 615218
rect 24208 614898 24250 615134
rect 24486 614898 24528 615134
rect 24208 614866 24528 614898
rect 20394 597818 20426 598054
rect 20662 597818 20746 598054
rect 20982 597818 21014 598054
rect 20394 597734 21014 597818
rect 20394 597498 20426 597734
rect 20662 597498 20746 597734
rect 20982 597498 21014 597734
rect 20394 562054 21014 597498
rect 27834 605494 28454 640938
rect 39568 619174 39888 619206
rect 39568 618938 39610 619174
rect 39846 618938 39888 619174
rect 39568 618854 39888 618938
rect 39568 618618 39610 618854
rect 39846 618618 39888 618854
rect 39568 618586 39888 618618
rect 70288 619174 70608 619206
rect 70288 618938 70330 619174
rect 70566 618938 70608 619174
rect 70288 618854 70608 618938
rect 70288 618618 70330 618854
rect 70566 618618 70608 618854
rect 70288 618586 70608 618618
rect 101008 619174 101328 619206
rect 101008 618938 101050 619174
rect 101286 618938 101328 619174
rect 101008 618854 101328 618938
rect 101008 618618 101050 618854
rect 101286 618618 101328 618854
rect 101008 618586 101328 618618
rect 131728 619174 132048 619206
rect 131728 618938 131770 619174
rect 132006 618938 132048 619174
rect 131728 618854 132048 618938
rect 131728 618618 131770 618854
rect 132006 618618 132048 618854
rect 131728 618586 132048 618618
rect 162448 619174 162768 619206
rect 162448 618938 162490 619174
rect 162726 618938 162768 619174
rect 162448 618854 162768 618938
rect 162448 618618 162490 618854
rect 162726 618618 162768 618854
rect 162448 618586 162768 618618
rect 193168 619174 193488 619206
rect 193168 618938 193210 619174
rect 193446 618938 193488 619174
rect 193168 618854 193488 618938
rect 193168 618618 193210 618854
rect 193446 618618 193488 618854
rect 193168 618586 193488 618618
rect 223888 619174 224208 619206
rect 223888 618938 223930 619174
rect 224166 618938 224208 619174
rect 223888 618854 224208 618938
rect 223888 618618 223930 618854
rect 224166 618618 224208 618854
rect 223888 618586 224208 618618
rect 254608 619174 254928 619206
rect 254608 618938 254650 619174
rect 254886 618938 254928 619174
rect 254608 618854 254928 618938
rect 254608 618618 254650 618854
rect 254886 618618 254928 618854
rect 254608 618586 254928 618618
rect 285328 619174 285648 619206
rect 285328 618938 285370 619174
rect 285606 618938 285648 619174
rect 285328 618854 285648 618938
rect 285328 618618 285370 618854
rect 285606 618618 285648 618854
rect 285328 618586 285648 618618
rect 316048 619174 316368 619206
rect 316048 618938 316090 619174
rect 316326 618938 316368 619174
rect 316048 618854 316368 618938
rect 316048 618618 316090 618854
rect 316326 618618 316368 618854
rect 316048 618586 316368 618618
rect 346768 619174 347088 619206
rect 346768 618938 346810 619174
rect 347046 618938 347088 619174
rect 346768 618854 347088 618938
rect 346768 618618 346810 618854
rect 347046 618618 347088 618854
rect 346768 618586 347088 618618
rect 54928 615454 55248 615486
rect 54928 615218 54970 615454
rect 55206 615218 55248 615454
rect 54928 615134 55248 615218
rect 54928 614898 54970 615134
rect 55206 614898 55248 615134
rect 54928 614866 55248 614898
rect 85648 615454 85968 615486
rect 85648 615218 85690 615454
rect 85926 615218 85968 615454
rect 85648 615134 85968 615218
rect 85648 614898 85690 615134
rect 85926 614898 85968 615134
rect 85648 614866 85968 614898
rect 116368 615454 116688 615486
rect 116368 615218 116410 615454
rect 116646 615218 116688 615454
rect 116368 615134 116688 615218
rect 116368 614898 116410 615134
rect 116646 614898 116688 615134
rect 116368 614866 116688 614898
rect 147088 615454 147408 615486
rect 147088 615218 147130 615454
rect 147366 615218 147408 615454
rect 147088 615134 147408 615218
rect 147088 614898 147130 615134
rect 147366 614898 147408 615134
rect 147088 614866 147408 614898
rect 177808 615454 178128 615486
rect 177808 615218 177850 615454
rect 178086 615218 178128 615454
rect 177808 615134 178128 615218
rect 177808 614898 177850 615134
rect 178086 614898 178128 615134
rect 177808 614866 178128 614898
rect 208528 615454 208848 615486
rect 208528 615218 208570 615454
rect 208806 615218 208848 615454
rect 208528 615134 208848 615218
rect 208528 614898 208570 615134
rect 208806 614898 208848 615134
rect 208528 614866 208848 614898
rect 239248 615454 239568 615486
rect 239248 615218 239290 615454
rect 239526 615218 239568 615454
rect 239248 615134 239568 615218
rect 239248 614898 239290 615134
rect 239526 614898 239568 615134
rect 239248 614866 239568 614898
rect 269968 615454 270288 615486
rect 269968 615218 270010 615454
rect 270246 615218 270288 615454
rect 269968 615134 270288 615218
rect 269968 614898 270010 615134
rect 270246 614898 270288 615134
rect 269968 614866 270288 614898
rect 300688 615454 301008 615486
rect 300688 615218 300730 615454
rect 300966 615218 301008 615454
rect 300688 615134 301008 615218
rect 300688 614898 300730 615134
rect 300966 614898 301008 615134
rect 300688 614866 301008 614898
rect 331408 615454 331728 615486
rect 331408 615218 331450 615454
rect 331686 615218 331728 615454
rect 331408 615134 331728 615218
rect 331408 614898 331450 615134
rect 331686 614898 331728 615134
rect 331408 614866 331728 614898
rect 361794 615454 362414 650898
rect 361794 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 362414 615454
rect 361794 615134 362414 615218
rect 361794 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 362414 615134
rect 27834 605258 27866 605494
rect 28102 605258 28186 605494
rect 28422 605258 28454 605494
rect 27834 605174 28454 605258
rect 27834 604938 27866 605174
rect 28102 604938 28186 605174
rect 28422 604938 28454 605174
rect 24208 579454 24528 579486
rect 24208 579218 24250 579454
rect 24486 579218 24528 579454
rect 24208 579134 24528 579218
rect 24208 578898 24250 579134
rect 24486 578898 24528 579134
rect 24208 578866 24528 578898
rect 20394 561818 20426 562054
rect 20662 561818 20746 562054
rect 20982 561818 21014 562054
rect 20394 561734 21014 561818
rect 20394 561498 20426 561734
rect 20662 561498 20746 561734
rect 20982 561498 21014 561734
rect 20394 526054 21014 561498
rect 27834 569494 28454 604938
rect 39568 583174 39888 583206
rect 39568 582938 39610 583174
rect 39846 582938 39888 583174
rect 39568 582854 39888 582938
rect 39568 582618 39610 582854
rect 39846 582618 39888 582854
rect 39568 582586 39888 582618
rect 70288 583174 70608 583206
rect 70288 582938 70330 583174
rect 70566 582938 70608 583174
rect 70288 582854 70608 582938
rect 70288 582618 70330 582854
rect 70566 582618 70608 582854
rect 70288 582586 70608 582618
rect 101008 583174 101328 583206
rect 101008 582938 101050 583174
rect 101286 582938 101328 583174
rect 101008 582854 101328 582938
rect 101008 582618 101050 582854
rect 101286 582618 101328 582854
rect 101008 582586 101328 582618
rect 131728 583174 132048 583206
rect 131728 582938 131770 583174
rect 132006 582938 132048 583174
rect 131728 582854 132048 582938
rect 131728 582618 131770 582854
rect 132006 582618 132048 582854
rect 131728 582586 132048 582618
rect 162448 583174 162768 583206
rect 162448 582938 162490 583174
rect 162726 582938 162768 583174
rect 162448 582854 162768 582938
rect 162448 582618 162490 582854
rect 162726 582618 162768 582854
rect 162448 582586 162768 582618
rect 193168 583174 193488 583206
rect 193168 582938 193210 583174
rect 193446 582938 193488 583174
rect 193168 582854 193488 582938
rect 193168 582618 193210 582854
rect 193446 582618 193488 582854
rect 193168 582586 193488 582618
rect 223888 583174 224208 583206
rect 223888 582938 223930 583174
rect 224166 582938 224208 583174
rect 223888 582854 224208 582938
rect 223888 582618 223930 582854
rect 224166 582618 224208 582854
rect 223888 582586 224208 582618
rect 254608 583174 254928 583206
rect 254608 582938 254650 583174
rect 254886 582938 254928 583174
rect 254608 582854 254928 582938
rect 254608 582618 254650 582854
rect 254886 582618 254928 582854
rect 254608 582586 254928 582618
rect 285328 583174 285648 583206
rect 285328 582938 285370 583174
rect 285606 582938 285648 583174
rect 285328 582854 285648 582938
rect 285328 582618 285370 582854
rect 285606 582618 285648 582854
rect 285328 582586 285648 582618
rect 316048 583174 316368 583206
rect 316048 582938 316090 583174
rect 316326 582938 316368 583174
rect 316048 582854 316368 582938
rect 316048 582618 316090 582854
rect 316326 582618 316368 582854
rect 316048 582586 316368 582618
rect 346768 583174 347088 583206
rect 346768 582938 346810 583174
rect 347046 582938 347088 583174
rect 346768 582854 347088 582938
rect 346768 582618 346810 582854
rect 347046 582618 347088 582854
rect 346768 582586 347088 582618
rect 54928 579454 55248 579486
rect 54928 579218 54970 579454
rect 55206 579218 55248 579454
rect 54928 579134 55248 579218
rect 54928 578898 54970 579134
rect 55206 578898 55248 579134
rect 54928 578866 55248 578898
rect 85648 579454 85968 579486
rect 85648 579218 85690 579454
rect 85926 579218 85968 579454
rect 85648 579134 85968 579218
rect 85648 578898 85690 579134
rect 85926 578898 85968 579134
rect 85648 578866 85968 578898
rect 116368 579454 116688 579486
rect 116368 579218 116410 579454
rect 116646 579218 116688 579454
rect 116368 579134 116688 579218
rect 116368 578898 116410 579134
rect 116646 578898 116688 579134
rect 116368 578866 116688 578898
rect 147088 579454 147408 579486
rect 147088 579218 147130 579454
rect 147366 579218 147408 579454
rect 147088 579134 147408 579218
rect 147088 578898 147130 579134
rect 147366 578898 147408 579134
rect 147088 578866 147408 578898
rect 177808 579454 178128 579486
rect 177808 579218 177850 579454
rect 178086 579218 178128 579454
rect 177808 579134 178128 579218
rect 177808 578898 177850 579134
rect 178086 578898 178128 579134
rect 177808 578866 178128 578898
rect 208528 579454 208848 579486
rect 208528 579218 208570 579454
rect 208806 579218 208848 579454
rect 208528 579134 208848 579218
rect 208528 578898 208570 579134
rect 208806 578898 208848 579134
rect 208528 578866 208848 578898
rect 239248 579454 239568 579486
rect 239248 579218 239290 579454
rect 239526 579218 239568 579454
rect 239248 579134 239568 579218
rect 239248 578898 239290 579134
rect 239526 578898 239568 579134
rect 239248 578866 239568 578898
rect 269968 579454 270288 579486
rect 269968 579218 270010 579454
rect 270246 579218 270288 579454
rect 269968 579134 270288 579218
rect 269968 578898 270010 579134
rect 270246 578898 270288 579134
rect 269968 578866 270288 578898
rect 300688 579454 301008 579486
rect 300688 579218 300730 579454
rect 300966 579218 301008 579454
rect 300688 579134 301008 579218
rect 300688 578898 300730 579134
rect 300966 578898 301008 579134
rect 300688 578866 301008 578898
rect 331408 579454 331728 579486
rect 331408 579218 331450 579454
rect 331686 579218 331728 579454
rect 331408 579134 331728 579218
rect 331408 578898 331450 579134
rect 331686 578898 331728 579134
rect 331408 578866 331728 578898
rect 361794 579454 362414 614898
rect 361794 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 362414 579454
rect 361794 579134 362414 579218
rect 361794 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 362414 579134
rect 27834 569258 27866 569494
rect 28102 569258 28186 569494
rect 28422 569258 28454 569494
rect 27834 569174 28454 569258
rect 27834 568938 27866 569174
rect 28102 568938 28186 569174
rect 28422 568938 28454 569174
rect 24208 543454 24528 543486
rect 24208 543218 24250 543454
rect 24486 543218 24528 543454
rect 24208 543134 24528 543218
rect 24208 542898 24250 543134
rect 24486 542898 24528 543134
rect 24208 542866 24528 542898
rect 20394 525818 20426 526054
rect 20662 525818 20746 526054
rect 20982 525818 21014 526054
rect 20394 525734 21014 525818
rect 20394 525498 20426 525734
rect 20662 525498 20746 525734
rect 20982 525498 21014 525734
rect 20394 490054 21014 525498
rect 27834 533494 28454 568938
rect 39568 547174 39888 547206
rect 39568 546938 39610 547174
rect 39846 546938 39888 547174
rect 39568 546854 39888 546938
rect 39568 546618 39610 546854
rect 39846 546618 39888 546854
rect 39568 546586 39888 546618
rect 70288 547174 70608 547206
rect 70288 546938 70330 547174
rect 70566 546938 70608 547174
rect 70288 546854 70608 546938
rect 70288 546618 70330 546854
rect 70566 546618 70608 546854
rect 70288 546586 70608 546618
rect 101008 547174 101328 547206
rect 101008 546938 101050 547174
rect 101286 546938 101328 547174
rect 101008 546854 101328 546938
rect 101008 546618 101050 546854
rect 101286 546618 101328 546854
rect 101008 546586 101328 546618
rect 131728 547174 132048 547206
rect 131728 546938 131770 547174
rect 132006 546938 132048 547174
rect 131728 546854 132048 546938
rect 131728 546618 131770 546854
rect 132006 546618 132048 546854
rect 131728 546586 132048 546618
rect 162448 547174 162768 547206
rect 162448 546938 162490 547174
rect 162726 546938 162768 547174
rect 162448 546854 162768 546938
rect 162448 546618 162490 546854
rect 162726 546618 162768 546854
rect 162448 546586 162768 546618
rect 193168 547174 193488 547206
rect 193168 546938 193210 547174
rect 193446 546938 193488 547174
rect 193168 546854 193488 546938
rect 193168 546618 193210 546854
rect 193446 546618 193488 546854
rect 193168 546586 193488 546618
rect 223888 547174 224208 547206
rect 223888 546938 223930 547174
rect 224166 546938 224208 547174
rect 223888 546854 224208 546938
rect 223888 546618 223930 546854
rect 224166 546618 224208 546854
rect 223888 546586 224208 546618
rect 254608 547174 254928 547206
rect 254608 546938 254650 547174
rect 254886 546938 254928 547174
rect 254608 546854 254928 546938
rect 254608 546618 254650 546854
rect 254886 546618 254928 546854
rect 254608 546586 254928 546618
rect 285328 547174 285648 547206
rect 285328 546938 285370 547174
rect 285606 546938 285648 547174
rect 285328 546854 285648 546938
rect 285328 546618 285370 546854
rect 285606 546618 285648 546854
rect 285328 546586 285648 546618
rect 316048 547174 316368 547206
rect 316048 546938 316090 547174
rect 316326 546938 316368 547174
rect 316048 546854 316368 546938
rect 316048 546618 316090 546854
rect 316326 546618 316368 546854
rect 316048 546586 316368 546618
rect 346768 547174 347088 547206
rect 346768 546938 346810 547174
rect 347046 546938 347088 547174
rect 346768 546854 347088 546938
rect 346768 546618 346810 546854
rect 347046 546618 347088 546854
rect 346768 546586 347088 546618
rect 54928 543454 55248 543486
rect 54928 543218 54970 543454
rect 55206 543218 55248 543454
rect 54928 543134 55248 543218
rect 54928 542898 54970 543134
rect 55206 542898 55248 543134
rect 54928 542866 55248 542898
rect 85648 543454 85968 543486
rect 85648 543218 85690 543454
rect 85926 543218 85968 543454
rect 85648 543134 85968 543218
rect 85648 542898 85690 543134
rect 85926 542898 85968 543134
rect 85648 542866 85968 542898
rect 116368 543454 116688 543486
rect 116368 543218 116410 543454
rect 116646 543218 116688 543454
rect 116368 543134 116688 543218
rect 116368 542898 116410 543134
rect 116646 542898 116688 543134
rect 116368 542866 116688 542898
rect 147088 543454 147408 543486
rect 147088 543218 147130 543454
rect 147366 543218 147408 543454
rect 147088 543134 147408 543218
rect 147088 542898 147130 543134
rect 147366 542898 147408 543134
rect 147088 542866 147408 542898
rect 177808 543454 178128 543486
rect 177808 543218 177850 543454
rect 178086 543218 178128 543454
rect 177808 543134 178128 543218
rect 177808 542898 177850 543134
rect 178086 542898 178128 543134
rect 177808 542866 178128 542898
rect 208528 543454 208848 543486
rect 208528 543218 208570 543454
rect 208806 543218 208848 543454
rect 208528 543134 208848 543218
rect 208528 542898 208570 543134
rect 208806 542898 208848 543134
rect 208528 542866 208848 542898
rect 239248 543454 239568 543486
rect 239248 543218 239290 543454
rect 239526 543218 239568 543454
rect 239248 543134 239568 543218
rect 239248 542898 239290 543134
rect 239526 542898 239568 543134
rect 239248 542866 239568 542898
rect 269968 543454 270288 543486
rect 269968 543218 270010 543454
rect 270246 543218 270288 543454
rect 269968 543134 270288 543218
rect 269968 542898 270010 543134
rect 270246 542898 270288 543134
rect 269968 542866 270288 542898
rect 300688 543454 301008 543486
rect 300688 543218 300730 543454
rect 300966 543218 301008 543454
rect 300688 543134 301008 543218
rect 300688 542898 300730 543134
rect 300966 542898 301008 543134
rect 300688 542866 301008 542898
rect 331408 543454 331728 543486
rect 331408 543218 331450 543454
rect 331686 543218 331728 543454
rect 331408 543134 331728 543218
rect 331408 542898 331450 543134
rect 331686 542898 331728 543134
rect 331408 542866 331728 542898
rect 361794 543454 362414 578898
rect 361794 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 362414 543454
rect 361794 543134 362414 543218
rect 361794 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 362414 543134
rect 27834 533258 27866 533494
rect 28102 533258 28186 533494
rect 28422 533258 28454 533494
rect 27834 533174 28454 533258
rect 27834 532938 27866 533174
rect 28102 532938 28186 533174
rect 28422 532938 28454 533174
rect 24208 507454 24528 507486
rect 24208 507218 24250 507454
rect 24486 507218 24528 507454
rect 24208 507134 24528 507218
rect 24208 506898 24250 507134
rect 24486 506898 24528 507134
rect 24208 506866 24528 506898
rect 20394 489818 20426 490054
rect 20662 489818 20746 490054
rect 20982 489818 21014 490054
rect 20394 489734 21014 489818
rect 20394 489498 20426 489734
rect 20662 489498 20746 489734
rect 20982 489498 21014 489734
rect 20394 454054 21014 489498
rect 27834 497494 28454 532938
rect 39568 511174 39888 511206
rect 39568 510938 39610 511174
rect 39846 510938 39888 511174
rect 39568 510854 39888 510938
rect 39568 510618 39610 510854
rect 39846 510618 39888 510854
rect 39568 510586 39888 510618
rect 70288 511174 70608 511206
rect 70288 510938 70330 511174
rect 70566 510938 70608 511174
rect 70288 510854 70608 510938
rect 70288 510618 70330 510854
rect 70566 510618 70608 510854
rect 70288 510586 70608 510618
rect 101008 511174 101328 511206
rect 101008 510938 101050 511174
rect 101286 510938 101328 511174
rect 101008 510854 101328 510938
rect 101008 510618 101050 510854
rect 101286 510618 101328 510854
rect 101008 510586 101328 510618
rect 131728 511174 132048 511206
rect 131728 510938 131770 511174
rect 132006 510938 132048 511174
rect 131728 510854 132048 510938
rect 131728 510618 131770 510854
rect 132006 510618 132048 510854
rect 131728 510586 132048 510618
rect 162448 511174 162768 511206
rect 162448 510938 162490 511174
rect 162726 510938 162768 511174
rect 162448 510854 162768 510938
rect 162448 510618 162490 510854
rect 162726 510618 162768 510854
rect 162448 510586 162768 510618
rect 193168 511174 193488 511206
rect 193168 510938 193210 511174
rect 193446 510938 193488 511174
rect 193168 510854 193488 510938
rect 193168 510618 193210 510854
rect 193446 510618 193488 510854
rect 193168 510586 193488 510618
rect 223888 511174 224208 511206
rect 223888 510938 223930 511174
rect 224166 510938 224208 511174
rect 223888 510854 224208 510938
rect 223888 510618 223930 510854
rect 224166 510618 224208 510854
rect 223888 510586 224208 510618
rect 254608 511174 254928 511206
rect 254608 510938 254650 511174
rect 254886 510938 254928 511174
rect 254608 510854 254928 510938
rect 254608 510618 254650 510854
rect 254886 510618 254928 510854
rect 254608 510586 254928 510618
rect 285328 511174 285648 511206
rect 285328 510938 285370 511174
rect 285606 510938 285648 511174
rect 285328 510854 285648 510938
rect 285328 510618 285370 510854
rect 285606 510618 285648 510854
rect 285328 510586 285648 510618
rect 316048 511174 316368 511206
rect 316048 510938 316090 511174
rect 316326 510938 316368 511174
rect 316048 510854 316368 510938
rect 316048 510618 316090 510854
rect 316326 510618 316368 510854
rect 316048 510586 316368 510618
rect 346768 511174 347088 511206
rect 346768 510938 346810 511174
rect 347046 510938 347088 511174
rect 346768 510854 347088 510938
rect 346768 510618 346810 510854
rect 347046 510618 347088 510854
rect 346768 510586 347088 510618
rect 54928 507454 55248 507486
rect 54928 507218 54970 507454
rect 55206 507218 55248 507454
rect 54928 507134 55248 507218
rect 54928 506898 54970 507134
rect 55206 506898 55248 507134
rect 54928 506866 55248 506898
rect 85648 507454 85968 507486
rect 85648 507218 85690 507454
rect 85926 507218 85968 507454
rect 85648 507134 85968 507218
rect 85648 506898 85690 507134
rect 85926 506898 85968 507134
rect 85648 506866 85968 506898
rect 116368 507454 116688 507486
rect 116368 507218 116410 507454
rect 116646 507218 116688 507454
rect 116368 507134 116688 507218
rect 116368 506898 116410 507134
rect 116646 506898 116688 507134
rect 116368 506866 116688 506898
rect 147088 507454 147408 507486
rect 147088 507218 147130 507454
rect 147366 507218 147408 507454
rect 147088 507134 147408 507218
rect 147088 506898 147130 507134
rect 147366 506898 147408 507134
rect 147088 506866 147408 506898
rect 177808 507454 178128 507486
rect 177808 507218 177850 507454
rect 178086 507218 178128 507454
rect 177808 507134 178128 507218
rect 177808 506898 177850 507134
rect 178086 506898 178128 507134
rect 177808 506866 178128 506898
rect 208528 507454 208848 507486
rect 208528 507218 208570 507454
rect 208806 507218 208848 507454
rect 208528 507134 208848 507218
rect 208528 506898 208570 507134
rect 208806 506898 208848 507134
rect 208528 506866 208848 506898
rect 239248 507454 239568 507486
rect 239248 507218 239290 507454
rect 239526 507218 239568 507454
rect 239248 507134 239568 507218
rect 239248 506898 239290 507134
rect 239526 506898 239568 507134
rect 239248 506866 239568 506898
rect 269968 507454 270288 507486
rect 269968 507218 270010 507454
rect 270246 507218 270288 507454
rect 269968 507134 270288 507218
rect 269968 506898 270010 507134
rect 270246 506898 270288 507134
rect 269968 506866 270288 506898
rect 300688 507454 301008 507486
rect 300688 507218 300730 507454
rect 300966 507218 301008 507454
rect 300688 507134 301008 507218
rect 300688 506898 300730 507134
rect 300966 506898 301008 507134
rect 300688 506866 301008 506898
rect 331408 507454 331728 507486
rect 331408 507218 331450 507454
rect 331686 507218 331728 507454
rect 331408 507134 331728 507218
rect 331408 506898 331450 507134
rect 331686 506898 331728 507134
rect 331408 506866 331728 506898
rect 361794 507454 362414 542898
rect 361794 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 362414 507454
rect 361794 507134 362414 507218
rect 361794 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 362414 507134
rect 27834 497258 27866 497494
rect 28102 497258 28186 497494
rect 28422 497258 28454 497494
rect 27834 497174 28454 497258
rect 27834 496938 27866 497174
rect 28102 496938 28186 497174
rect 28422 496938 28454 497174
rect 24208 471454 24528 471486
rect 24208 471218 24250 471454
rect 24486 471218 24528 471454
rect 24208 471134 24528 471218
rect 24208 470898 24250 471134
rect 24486 470898 24528 471134
rect 24208 470866 24528 470898
rect 20394 453818 20426 454054
rect 20662 453818 20746 454054
rect 20982 453818 21014 454054
rect 20394 453734 21014 453818
rect 20394 453498 20426 453734
rect 20662 453498 20746 453734
rect 20982 453498 21014 453734
rect 20394 418054 21014 453498
rect 27834 461494 28454 496938
rect 39568 475174 39888 475206
rect 39568 474938 39610 475174
rect 39846 474938 39888 475174
rect 39568 474854 39888 474938
rect 39568 474618 39610 474854
rect 39846 474618 39888 474854
rect 39568 474586 39888 474618
rect 70288 475174 70608 475206
rect 70288 474938 70330 475174
rect 70566 474938 70608 475174
rect 70288 474854 70608 474938
rect 70288 474618 70330 474854
rect 70566 474618 70608 474854
rect 70288 474586 70608 474618
rect 101008 475174 101328 475206
rect 101008 474938 101050 475174
rect 101286 474938 101328 475174
rect 101008 474854 101328 474938
rect 101008 474618 101050 474854
rect 101286 474618 101328 474854
rect 101008 474586 101328 474618
rect 131728 475174 132048 475206
rect 131728 474938 131770 475174
rect 132006 474938 132048 475174
rect 131728 474854 132048 474938
rect 131728 474618 131770 474854
rect 132006 474618 132048 474854
rect 131728 474586 132048 474618
rect 162448 475174 162768 475206
rect 162448 474938 162490 475174
rect 162726 474938 162768 475174
rect 162448 474854 162768 474938
rect 162448 474618 162490 474854
rect 162726 474618 162768 474854
rect 162448 474586 162768 474618
rect 193168 475174 193488 475206
rect 193168 474938 193210 475174
rect 193446 474938 193488 475174
rect 193168 474854 193488 474938
rect 193168 474618 193210 474854
rect 193446 474618 193488 474854
rect 193168 474586 193488 474618
rect 223888 475174 224208 475206
rect 223888 474938 223930 475174
rect 224166 474938 224208 475174
rect 223888 474854 224208 474938
rect 223888 474618 223930 474854
rect 224166 474618 224208 474854
rect 223888 474586 224208 474618
rect 254608 475174 254928 475206
rect 254608 474938 254650 475174
rect 254886 474938 254928 475174
rect 254608 474854 254928 474938
rect 254608 474618 254650 474854
rect 254886 474618 254928 474854
rect 254608 474586 254928 474618
rect 285328 475174 285648 475206
rect 285328 474938 285370 475174
rect 285606 474938 285648 475174
rect 285328 474854 285648 474938
rect 285328 474618 285370 474854
rect 285606 474618 285648 474854
rect 285328 474586 285648 474618
rect 316048 475174 316368 475206
rect 316048 474938 316090 475174
rect 316326 474938 316368 475174
rect 316048 474854 316368 474938
rect 316048 474618 316090 474854
rect 316326 474618 316368 474854
rect 316048 474586 316368 474618
rect 346768 475174 347088 475206
rect 346768 474938 346810 475174
rect 347046 474938 347088 475174
rect 346768 474854 347088 474938
rect 346768 474618 346810 474854
rect 347046 474618 347088 474854
rect 346768 474586 347088 474618
rect 54928 471454 55248 471486
rect 54928 471218 54970 471454
rect 55206 471218 55248 471454
rect 54928 471134 55248 471218
rect 54928 470898 54970 471134
rect 55206 470898 55248 471134
rect 54928 470866 55248 470898
rect 85648 471454 85968 471486
rect 85648 471218 85690 471454
rect 85926 471218 85968 471454
rect 85648 471134 85968 471218
rect 85648 470898 85690 471134
rect 85926 470898 85968 471134
rect 85648 470866 85968 470898
rect 116368 471454 116688 471486
rect 116368 471218 116410 471454
rect 116646 471218 116688 471454
rect 116368 471134 116688 471218
rect 116368 470898 116410 471134
rect 116646 470898 116688 471134
rect 116368 470866 116688 470898
rect 147088 471454 147408 471486
rect 147088 471218 147130 471454
rect 147366 471218 147408 471454
rect 147088 471134 147408 471218
rect 147088 470898 147130 471134
rect 147366 470898 147408 471134
rect 147088 470866 147408 470898
rect 177808 471454 178128 471486
rect 177808 471218 177850 471454
rect 178086 471218 178128 471454
rect 177808 471134 178128 471218
rect 177808 470898 177850 471134
rect 178086 470898 178128 471134
rect 177808 470866 178128 470898
rect 208528 471454 208848 471486
rect 208528 471218 208570 471454
rect 208806 471218 208848 471454
rect 208528 471134 208848 471218
rect 208528 470898 208570 471134
rect 208806 470898 208848 471134
rect 208528 470866 208848 470898
rect 239248 471454 239568 471486
rect 239248 471218 239290 471454
rect 239526 471218 239568 471454
rect 239248 471134 239568 471218
rect 239248 470898 239290 471134
rect 239526 470898 239568 471134
rect 239248 470866 239568 470898
rect 269968 471454 270288 471486
rect 269968 471218 270010 471454
rect 270246 471218 270288 471454
rect 269968 471134 270288 471218
rect 269968 470898 270010 471134
rect 270246 470898 270288 471134
rect 269968 470866 270288 470898
rect 300688 471454 301008 471486
rect 300688 471218 300730 471454
rect 300966 471218 301008 471454
rect 300688 471134 301008 471218
rect 300688 470898 300730 471134
rect 300966 470898 301008 471134
rect 300688 470866 301008 470898
rect 331408 471454 331728 471486
rect 331408 471218 331450 471454
rect 331686 471218 331728 471454
rect 331408 471134 331728 471218
rect 331408 470898 331450 471134
rect 331686 470898 331728 471134
rect 331408 470866 331728 470898
rect 361794 471454 362414 506898
rect 361794 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 362414 471454
rect 361794 471134 362414 471218
rect 361794 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 362414 471134
rect 27834 461258 27866 461494
rect 28102 461258 28186 461494
rect 28422 461258 28454 461494
rect 27834 461174 28454 461258
rect 27834 460938 27866 461174
rect 28102 460938 28186 461174
rect 28422 460938 28454 461174
rect 24208 435454 24528 435486
rect 24208 435218 24250 435454
rect 24486 435218 24528 435454
rect 24208 435134 24528 435218
rect 24208 434898 24250 435134
rect 24486 434898 24528 435134
rect 24208 434866 24528 434898
rect 20394 417818 20426 418054
rect 20662 417818 20746 418054
rect 20982 417818 21014 418054
rect 20394 417734 21014 417818
rect 20394 417498 20426 417734
rect 20662 417498 20746 417734
rect 20982 417498 21014 417734
rect 20394 382054 21014 417498
rect 27834 425494 28454 460938
rect 39568 439174 39888 439206
rect 39568 438938 39610 439174
rect 39846 438938 39888 439174
rect 39568 438854 39888 438938
rect 39568 438618 39610 438854
rect 39846 438618 39888 438854
rect 39568 438586 39888 438618
rect 70288 439174 70608 439206
rect 70288 438938 70330 439174
rect 70566 438938 70608 439174
rect 70288 438854 70608 438938
rect 70288 438618 70330 438854
rect 70566 438618 70608 438854
rect 70288 438586 70608 438618
rect 101008 439174 101328 439206
rect 101008 438938 101050 439174
rect 101286 438938 101328 439174
rect 101008 438854 101328 438938
rect 101008 438618 101050 438854
rect 101286 438618 101328 438854
rect 101008 438586 101328 438618
rect 131728 439174 132048 439206
rect 131728 438938 131770 439174
rect 132006 438938 132048 439174
rect 131728 438854 132048 438938
rect 131728 438618 131770 438854
rect 132006 438618 132048 438854
rect 131728 438586 132048 438618
rect 162448 439174 162768 439206
rect 162448 438938 162490 439174
rect 162726 438938 162768 439174
rect 162448 438854 162768 438938
rect 162448 438618 162490 438854
rect 162726 438618 162768 438854
rect 162448 438586 162768 438618
rect 193168 439174 193488 439206
rect 193168 438938 193210 439174
rect 193446 438938 193488 439174
rect 193168 438854 193488 438938
rect 193168 438618 193210 438854
rect 193446 438618 193488 438854
rect 193168 438586 193488 438618
rect 223888 439174 224208 439206
rect 223888 438938 223930 439174
rect 224166 438938 224208 439174
rect 223888 438854 224208 438938
rect 223888 438618 223930 438854
rect 224166 438618 224208 438854
rect 223888 438586 224208 438618
rect 254608 439174 254928 439206
rect 254608 438938 254650 439174
rect 254886 438938 254928 439174
rect 254608 438854 254928 438938
rect 254608 438618 254650 438854
rect 254886 438618 254928 438854
rect 254608 438586 254928 438618
rect 285328 439174 285648 439206
rect 285328 438938 285370 439174
rect 285606 438938 285648 439174
rect 285328 438854 285648 438938
rect 285328 438618 285370 438854
rect 285606 438618 285648 438854
rect 285328 438586 285648 438618
rect 316048 439174 316368 439206
rect 316048 438938 316090 439174
rect 316326 438938 316368 439174
rect 316048 438854 316368 438938
rect 316048 438618 316090 438854
rect 316326 438618 316368 438854
rect 316048 438586 316368 438618
rect 346768 439174 347088 439206
rect 346768 438938 346810 439174
rect 347046 438938 347088 439174
rect 346768 438854 347088 438938
rect 346768 438618 346810 438854
rect 347046 438618 347088 438854
rect 346768 438586 347088 438618
rect 54928 435454 55248 435486
rect 54928 435218 54970 435454
rect 55206 435218 55248 435454
rect 54928 435134 55248 435218
rect 54928 434898 54970 435134
rect 55206 434898 55248 435134
rect 54928 434866 55248 434898
rect 85648 435454 85968 435486
rect 85648 435218 85690 435454
rect 85926 435218 85968 435454
rect 85648 435134 85968 435218
rect 85648 434898 85690 435134
rect 85926 434898 85968 435134
rect 85648 434866 85968 434898
rect 116368 435454 116688 435486
rect 116368 435218 116410 435454
rect 116646 435218 116688 435454
rect 116368 435134 116688 435218
rect 116368 434898 116410 435134
rect 116646 434898 116688 435134
rect 116368 434866 116688 434898
rect 147088 435454 147408 435486
rect 147088 435218 147130 435454
rect 147366 435218 147408 435454
rect 147088 435134 147408 435218
rect 147088 434898 147130 435134
rect 147366 434898 147408 435134
rect 147088 434866 147408 434898
rect 177808 435454 178128 435486
rect 177808 435218 177850 435454
rect 178086 435218 178128 435454
rect 177808 435134 178128 435218
rect 177808 434898 177850 435134
rect 178086 434898 178128 435134
rect 177808 434866 178128 434898
rect 208528 435454 208848 435486
rect 208528 435218 208570 435454
rect 208806 435218 208848 435454
rect 208528 435134 208848 435218
rect 208528 434898 208570 435134
rect 208806 434898 208848 435134
rect 208528 434866 208848 434898
rect 239248 435454 239568 435486
rect 239248 435218 239290 435454
rect 239526 435218 239568 435454
rect 239248 435134 239568 435218
rect 239248 434898 239290 435134
rect 239526 434898 239568 435134
rect 239248 434866 239568 434898
rect 269968 435454 270288 435486
rect 269968 435218 270010 435454
rect 270246 435218 270288 435454
rect 269968 435134 270288 435218
rect 269968 434898 270010 435134
rect 270246 434898 270288 435134
rect 269968 434866 270288 434898
rect 300688 435454 301008 435486
rect 300688 435218 300730 435454
rect 300966 435218 301008 435454
rect 300688 435134 301008 435218
rect 300688 434898 300730 435134
rect 300966 434898 301008 435134
rect 300688 434866 301008 434898
rect 331408 435454 331728 435486
rect 331408 435218 331450 435454
rect 331686 435218 331728 435454
rect 331408 435134 331728 435218
rect 331408 434898 331450 435134
rect 331686 434898 331728 435134
rect 331408 434866 331728 434898
rect 361794 435454 362414 470898
rect 361794 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 362414 435454
rect 361794 435134 362414 435218
rect 361794 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 362414 435134
rect 27834 425258 27866 425494
rect 28102 425258 28186 425494
rect 28422 425258 28454 425494
rect 27834 425174 28454 425258
rect 27834 424938 27866 425174
rect 28102 424938 28186 425174
rect 28422 424938 28454 425174
rect 24208 399454 24528 399486
rect 24208 399218 24250 399454
rect 24486 399218 24528 399454
rect 24208 399134 24528 399218
rect 24208 398898 24250 399134
rect 24486 398898 24528 399134
rect 24208 398866 24528 398898
rect 20394 381818 20426 382054
rect 20662 381818 20746 382054
rect 20982 381818 21014 382054
rect 20394 381734 21014 381818
rect 20394 381498 20426 381734
rect 20662 381498 20746 381734
rect 20982 381498 21014 381734
rect 20394 346054 21014 381498
rect 27834 389494 28454 424938
rect 39568 403174 39888 403206
rect 39568 402938 39610 403174
rect 39846 402938 39888 403174
rect 39568 402854 39888 402938
rect 39568 402618 39610 402854
rect 39846 402618 39888 402854
rect 39568 402586 39888 402618
rect 70288 403174 70608 403206
rect 70288 402938 70330 403174
rect 70566 402938 70608 403174
rect 70288 402854 70608 402938
rect 70288 402618 70330 402854
rect 70566 402618 70608 402854
rect 70288 402586 70608 402618
rect 101008 403174 101328 403206
rect 101008 402938 101050 403174
rect 101286 402938 101328 403174
rect 101008 402854 101328 402938
rect 101008 402618 101050 402854
rect 101286 402618 101328 402854
rect 101008 402586 101328 402618
rect 131728 403174 132048 403206
rect 131728 402938 131770 403174
rect 132006 402938 132048 403174
rect 131728 402854 132048 402938
rect 131728 402618 131770 402854
rect 132006 402618 132048 402854
rect 131728 402586 132048 402618
rect 162448 403174 162768 403206
rect 162448 402938 162490 403174
rect 162726 402938 162768 403174
rect 162448 402854 162768 402938
rect 162448 402618 162490 402854
rect 162726 402618 162768 402854
rect 162448 402586 162768 402618
rect 193168 403174 193488 403206
rect 193168 402938 193210 403174
rect 193446 402938 193488 403174
rect 193168 402854 193488 402938
rect 193168 402618 193210 402854
rect 193446 402618 193488 402854
rect 193168 402586 193488 402618
rect 223888 403174 224208 403206
rect 223888 402938 223930 403174
rect 224166 402938 224208 403174
rect 223888 402854 224208 402938
rect 223888 402618 223930 402854
rect 224166 402618 224208 402854
rect 223888 402586 224208 402618
rect 254608 403174 254928 403206
rect 254608 402938 254650 403174
rect 254886 402938 254928 403174
rect 254608 402854 254928 402938
rect 254608 402618 254650 402854
rect 254886 402618 254928 402854
rect 254608 402586 254928 402618
rect 285328 403174 285648 403206
rect 285328 402938 285370 403174
rect 285606 402938 285648 403174
rect 285328 402854 285648 402938
rect 285328 402618 285370 402854
rect 285606 402618 285648 402854
rect 285328 402586 285648 402618
rect 316048 403174 316368 403206
rect 316048 402938 316090 403174
rect 316326 402938 316368 403174
rect 316048 402854 316368 402938
rect 316048 402618 316090 402854
rect 316326 402618 316368 402854
rect 316048 402586 316368 402618
rect 346768 403174 347088 403206
rect 346768 402938 346810 403174
rect 347046 402938 347088 403174
rect 346768 402854 347088 402938
rect 346768 402618 346810 402854
rect 347046 402618 347088 402854
rect 346768 402586 347088 402618
rect 54928 399454 55248 399486
rect 54928 399218 54970 399454
rect 55206 399218 55248 399454
rect 54928 399134 55248 399218
rect 54928 398898 54970 399134
rect 55206 398898 55248 399134
rect 54928 398866 55248 398898
rect 85648 399454 85968 399486
rect 85648 399218 85690 399454
rect 85926 399218 85968 399454
rect 85648 399134 85968 399218
rect 85648 398898 85690 399134
rect 85926 398898 85968 399134
rect 85648 398866 85968 398898
rect 116368 399454 116688 399486
rect 116368 399218 116410 399454
rect 116646 399218 116688 399454
rect 116368 399134 116688 399218
rect 116368 398898 116410 399134
rect 116646 398898 116688 399134
rect 116368 398866 116688 398898
rect 147088 399454 147408 399486
rect 147088 399218 147130 399454
rect 147366 399218 147408 399454
rect 147088 399134 147408 399218
rect 147088 398898 147130 399134
rect 147366 398898 147408 399134
rect 147088 398866 147408 398898
rect 177808 399454 178128 399486
rect 177808 399218 177850 399454
rect 178086 399218 178128 399454
rect 177808 399134 178128 399218
rect 177808 398898 177850 399134
rect 178086 398898 178128 399134
rect 177808 398866 178128 398898
rect 208528 399454 208848 399486
rect 208528 399218 208570 399454
rect 208806 399218 208848 399454
rect 208528 399134 208848 399218
rect 208528 398898 208570 399134
rect 208806 398898 208848 399134
rect 208528 398866 208848 398898
rect 239248 399454 239568 399486
rect 239248 399218 239290 399454
rect 239526 399218 239568 399454
rect 239248 399134 239568 399218
rect 239248 398898 239290 399134
rect 239526 398898 239568 399134
rect 239248 398866 239568 398898
rect 269968 399454 270288 399486
rect 269968 399218 270010 399454
rect 270246 399218 270288 399454
rect 269968 399134 270288 399218
rect 269968 398898 270010 399134
rect 270246 398898 270288 399134
rect 269968 398866 270288 398898
rect 300688 399454 301008 399486
rect 300688 399218 300730 399454
rect 300966 399218 301008 399454
rect 300688 399134 301008 399218
rect 300688 398898 300730 399134
rect 300966 398898 301008 399134
rect 300688 398866 301008 398898
rect 331408 399454 331728 399486
rect 331408 399218 331450 399454
rect 331686 399218 331728 399454
rect 331408 399134 331728 399218
rect 331408 398898 331450 399134
rect 331686 398898 331728 399134
rect 331408 398866 331728 398898
rect 361794 399454 362414 434898
rect 361794 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 362414 399454
rect 361794 399134 362414 399218
rect 361794 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 362414 399134
rect 27834 389258 27866 389494
rect 28102 389258 28186 389494
rect 28422 389258 28454 389494
rect 27834 389174 28454 389258
rect 27834 388938 27866 389174
rect 28102 388938 28186 389174
rect 28422 388938 28454 389174
rect 24208 363454 24528 363486
rect 24208 363218 24250 363454
rect 24486 363218 24528 363454
rect 24208 363134 24528 363218
rect 24208 362898 24250 363134
rect 24486 362898 24528 363134
rect 24208 362866 24528 362898
rect 20394 345818 20426 346054
rect 20662 345818 20746 346054
rect 20982 345818 21014 346054
rect 20394 345734 21014 345818
rect 20394 345498 20426 345734
rect 20662 345498 20746 345734
rect 20982 345498 21014 345734
rect 20394 310054 21014 345498
rect 27834 353494 28454 388938
rect 39568 367174 39888 367206
rect 39568 366938 39610 367174
rect 39846 366938 39888 367174
rect 39568 366854 39888 366938
rect 39568 366618 39610 366854
rect 39846 366618 39888 366854
rect 39568 366586 39888 366618
rect 70288 367174 70608 367206
rect 70288 366938 70330 367174
rect 70566 366938 70608 367174
rect 70288 366854 70608 366938
rect 70288 366618 70330 366854
rect 70566 366618 70608 366854
rect 70288 366586 70608 366618
rect 101008 367174 101328 367206
rect 101008 366938 101050 367174
rect 101286 366938 101328 367174
rect 101008 366854 101328 366938
rect 101008 366618 101050 366854
rect 101286 366618 101328 366854
rect 101008 366586 101328 366618
rect 131728 367174 132048 367206
rect 131728 366938 131770 367174
rect 132006 366938 132048 367174
rect 131728 366854 132048 366938
rect 131728 366618 131770 366854
rect 132006 366618 132048 366854
rect 131728 366586 132048 366618
rect 162448 367174 162768 367206
rect 162448 366938 162490 367174
rect 162726 366938 162768 367174
rect 162448 366854 162768 366938
rect 162448 366618 162490 366854
rect 162726 366618 162768 366854
rect 162448 366586 162768 366618
rect 193168 367174 193488 367206
rect 193168 366938 193210 367174
rect 193446 366938 193488 367174
rect 193168 366854 193488 366938
rect 193168 366618 193210 366854
rect 193446 366618 193488 366854
rect 193168 366586 193488 366618
rect 223888 367174 224208 367206
rect 223888 366938 223930 367174
rect 224166 366938 224208 367174
rect 223888 366854 224208 366938
rect 223888 366618 223930 366854
rect 224166 366618 224208 366854
rect 223888 366586 224208 366618
rect 254608 367174 254928 367206
rect 254608 366938 254650 367174
rect 254886 366938 254928 367174
rect 254608 366854 254928 366938
rect 254608 366618 254650 366854
rect 254886 366618 254928 366854
rect 254608 366586 254928 366618
rect 285328 367174 285648 367206
rect 285328 366938 285370 367174
rect 285606 366938 285648 367174
rect 285328 366854 285648 366938
rect 285328 366618 285370 366854
rect 285606 366618 285648 366854
rect 285328 366586 285648 366618
rect 316048 367174 316368 367206
rect 316048 366938 316090 367174
rect 316326 366938 316368 367174
rect 316048 366854 316368 366938
rect 316048 366618 316090 366854
rect 316326 366618 316368 366854
rect 316048 366586 316368 366618
rect 346768 367174 347088 367206
rect 346768 366938 346810 367174
rect 347046 366938 347088 367174
rect 346768 366854 347088 366938
rect 346768 366618 346810 366854
rect 347046 366618 347088 366854
rect 346768 366586 347088 366618
rect 54928 363454 55248 363486
rect 54928 363218 54970 363454
rect 55206 363218 55248 363454
rect 54928 363134 55248 363218
rect 54928 362898 54970 363134
rect 55206 362898 55248 363134
rect 54928 362866 55248 362898
rect 85648 363454 85968 363486
rect 85648 363218 85690 363454
rect 85926 363218 85968 363454
rect 85648 363134 85968 363218
rect 85648 362898 85690 363134
rect 85926 362898 85968 363134
rect 85648 362866 85968 362898
rect 116368 363454 116688 363486
rect 116368 363218 116410 363454
rect 116646 363218 116688 363454
rect 116368 363134 116688 363218
rect 116368 362898 116410 363134
rect 116646 362898 116688 363134
rect 116368 362866 116688 362898
rect 147088 363454 147408 363486
rect 147088 363218 147130 363454
rect 147366 363218 147408 363454
rect 147088 363134 147408 363218
rect 147088 362898 147130 363134
rect 147366 362898 147408 363134
rect 147088 362866 147408 362898
rect 177808 363454 178128 363486
rect 177808 363218 177850 363454
rect 178086 363218 178128 363454
rect 177808 363134 178128 363218
rect 177808 362898 177850 363134
rect 178086 362898 178128 363134
rect 177808 362866 178128 362898
rect 208528 363454 208848 363486
rect 208528 363218 208570 363454
rect 208806 363218 208848 363454
rect 208528 363134 208848 363218
rect 208528 362898 208570 363134
rect 208806 362898 208848 363134
rect 208528 362866 208848 362898
rect 239248 363454 239568 363486
rect 239248 363218 239290 363454
rect 239526 363218 239568 363454
rect 239248 363134 239568 363218
rect 239248 362898 239290 363134
rect 239526 362898 239568 363134
rect 239248 362866 239568 362898
rect 269968 363454 270288 363486
rect 269968 363218 270010 363454
rect 270246 363218 270288 363454
rect 269968 363134 270288 363218
rect 269968 362898 270010 363134
rect 270246 362898 270288 363134
rect 269968 362866 270288 362898
rect 300688 363454 301008 363486
rect 300688 363218 300730 363454
rect 300966 363218 301008 363454
rect 300688 363134 301008 363218
rect 300688 362898 300730 363134
rect 300966 362898 301008 363134
rect 300688 362866 301008 362898
rect 331408 363454 331728 363486
rect 331408 363218 331450 363454
rect 331686 363218 331728 363454
rect 331408 363134 331728 363218
rect 331408 362898 331450 363134
rect 331686 362898 331728 363134
rect 331408 362866 331728 362898
rect 361794 363454 362414 398898
rect 361794 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 362414 363454
rect 361794 363134 362414 363218
rect 361794 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 362414 363134
rect 27834 353258 27866 353494
rect 28102 353258 28186 353494
rect 28422 353258 28454 353494
rect 27834 353174 28454 353258
rect 27834 352938 27866 353174
rect 28102 352938 28186 353174
rect 28422 352938 28454 353174
rect 24208 327454 24528 327486
rect 24208 327218 24250 327454
rect 24486 327218 24528 327454
rect 24208 327134 24528 327218
rect 24208 326898 24250 327134
rect 24486 326898 24528 327134
rect 24208 326866 24528 326898
rect 20394 309818 20426 310054
rect 20662 309818 20746 310054
rect 20982 309818 21014 310054
rect 20394 309734 21014 309818
rect 20394 309498 20426 309734
rect 20662 309498 20746 309734
rect 20982 309498 21014 309734
rect 20394 274054 21014 309498
rect 27834 317494 28454 352938
rect 39568 331174 39888 331206
rect 39568 330938 39610 331174
rect 39846 330938 39888 331174
rect 39568 330854 39888 330938
rect 39568 330618 39610 330854
rect 39846 330618 39888 330854
rect 39568 330586 39888 330618
rect 70288 331174 70608 331206
rect 70288 330938 70330 331174
rect 70566 330938 70608 331174
rect 70288 330854 70608 330938
rect 70288 330618 70330 330854
rect 70566 330618 70608 330854
rect 70288 330586 70608 330618
rect 101008 331174 101328 331206
rect 101008 330938 101050 331174
rect 101286 330938 101328 331174
rect 101008 330854 101328 330938
rect 101008 330618 101050 330854
rect 101286 330618 101328 330854
rect 101008 330586 101328 330618
rect 131728 331174 132048 331206
rect 131728 330938 131770 331174
rect 132006 330938 132048 331174
rect 131728 330854 132048 330938
rect 131728 330618 131770 330854
rect 132006 330618 132048 330854
rect 131728 330586 132048 330618
rect 162448 331174 162768 331206
rect 162448 330938 162490 331174
rect 162726 330938 162768 331174
rect 162448 330854 162768 330938
rect 162448 330618 162490 330854
rect 162726 330618 162768 330854
rect 162448 330586 162768 330618
rect 193168 331174 193488 331206
rect 193168 330938 193210 331174
rect 193446 330938 193488 331174
rect 193168 330854 193488 330938
rect 193168 330618 193210 330854
rect 193446 330618 193488 330854
rect 193168 330586 193488 330618
rect 223888 331174 224208 331206
rect 223888 330938 223930 331174
rect 224166 330938 224208 331174
rect 223888 330854 224208 330938
rect 223888 330618 223930 330854
rect 224166 330618 224208 330854
rect 223888 330586 224208 330618
rect 254608 331174 254928 331206
rect 254608 330938 254650 331174
rect 254886 330938 254928 331174
rect 254608 330854 254928 330938
rect 254608 330618 254650 330854
rect 254886 330618 254928 330854
rect 254608 330586 254928 330618
rect 285328 331174 285648 331206
rect 285328 330938 285370 331174
rect 285606 330938 285648 331174
rect 285328 330854 285648 330938
rect 285328 330618 285370 330854
rect 285606 330618 285648 330854
rect 285328 330586 285648 330618
rect 316048 331174 316368 331206
rect 316048 330938 316090 331174
rect 316326 330938 316368 331174
rect 316048 330854 316368 330938
rect 316048 330618 316090 330854
rect 316326 330618 316368 330854
rect 316048 330586 316368 330618
rect 346768 331174 347088 331206
rect 346768 330938 346810 331174
rect 347046 330938 347088 331174
rect 346768 330854 347088 330938
rect 346768 330618 346810 330854
rect 347046 330618 347088 330854
rect 346768 330586 347088 330618
rect 54928 327454 55248 327486
rect 54928 327218 54970 327454
rect 55206 327218 55248 327454
rect 54928 327134 55248 327218
rect 54928 326898 54970 327134
rect 55206 326898 55248 327134
rect 54928 326866 55248 326898
rect 85648 327454 85968 327486
rect 85648 327218 85690 327454
rect 85926 327218 85968 327454
rect 85648 327134 85968 327218
rect 85648 326898 85690 327134
rect 85926 326898 85968 327134
rect 85648 326866 85968 326898
rect 116368 327454 116688 327486
rect 116368 327218 116410 327454
rect 116646 327218 116688 327454
rect 116368 327134 116688 327218
rect 116368 326898 116410 327134
rect 116646 326898 116688 327134
rect 116368 326866 116688 326898
rect 147088 327454 147408 327486
rect 147088 327218 147130 327454
rect 147366 327218 147408 327454
rect 147088 327134 147408 327218
rect 147088 326898 147130 327134
rect 147366 326898 147408 327134
rect 147088 326866 147408 326898
rect 177808 327454 178128 327486
rect 177808 327218 177850 327454
rect 178086 327218 178128 327454
rect 177808 327134 178128 327218
rect 177808 326898 177850 327134
rect 178086 326898 178128 327134
rect 177808 326866 178128 326898
rect 208528 327454 208848 327486
rect 208528 327218 208570 327454
rect 208806 327218 208848 327454
rect 208528 327134 208848 327218
rect 208528 326898 208570 327134
rect 208806 326898 208848 327134
rect 208528 326866 208848 326898
rect 239248 327454 239568 327486
rect 239248 327218 239290 327454
rect 239526 327218 239568 327454
rect 239248 327134 239568 327218
rect 239248 326898 239290 327134
rect 239526 326898 239568 327134
rect 239248 326866 239568 326898
rect 269968 327454 270288 327486
rect 269968 327218 270010 327454
rect 270246 327218 270288 327454
rect 269968 327134 270288 327218
rect 269968 326898 270010 327134
rect 270246 326898 270288 327134
rect 269968 326866 270288 326898
rect 300688 327454 301008 327486
rect 300688 327218 300730 327454
rect 300966 327218 301008 327454
rect 300688 327134 301008 327218
rect 300688 326898 300730 327134
rect 300966 326898 301008 327134
rect 300688 326866 301008 326898
rect 331408 327454 331728 327486
rect 331408 327218 331450 327454
rect 331686 327218 331728 327454
rect 331408 327134 331728 327218
rect 331408 326898 331450 327134
rect 331686 326898 331728 327134
rect 331408 326866 331728 326898
rect 361794 327454 362414 362898
rect 361794 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 362414 327454
rect 361794 327134 362414 327218
rect 361794 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 362414 327134
rect 27834 317258 27866 317494
rect 28102 317258 28186 317494
rect 28422 317258 28454 317494
rect 27834 317174 28454 317258
rect 27834 316938 27866 317174
rect 28102 316938 28186 317174
rect 28422 316938 28454 317174
rect 24208 291454 24528 291486
rect 24208 291218 24250 291454
rect 24486 291218 24528 291454
rect 24208 291134 24528 291218
rect 24208 290898 24250 291134
rect 24486 290898 24528 291134
rect 24208 290866 24528 290898
rect 20394 273818 20426 274054
rect 20662 273818 20746 274054
rect 20982 273818 21014 274054
rect 20394 273734 21014 273818
rect 20394 273498 20426 273734
rect 20662 273498 20746 273734
rect 20982 273498 21014 273734
rect 20394 238054 21014 273498
rect 27834 281494 28454 316938
rect 39568 295174 39888 295206
rect 39568 294938 39610 295174
rect 39846 294938 39888 295174
rect 39568 294854 39888 294938
rect 39568 294618 39610 294854
rect 39846 294618 39888 294854
rect 39568 294586 39888 294618
rect 70288 295174 70608 295206
rect 70288 294938 70330 295174
rect 70566 294938 70608 295174
rect 70288 294854 70608 294938
rect 70288 294618 70330 294854
rect 70566 294618 70608 294854
rect 70288 294586 70608 294618
rect 101008 295174 101328 295206
rect 101008 294938 101050 295174
rect 101286 294938 101328 295174
rect 101008 294854 101328 294938
rect 101008 294618 101050 294854
rect 101286 294618 101328 294854
rect 101008 294586 101328 294618
rect 131728 295174 132048 295206
rect 131728 294938 131770 295174
rect 132006 294938 132048 295174
rect 131728 294854 132048 294938
rect 131728 294618 131770 294854
rect 132006 294618 132048 294854
rect 131728 294586 132048 294618
rect 162448 295174 162768 295206
rect 162448 294938 162490 295174
rect 162726 294938 162768 295174
rect 162448 294854 162768 294938
rect 162448 294618 162490 294854
rect 162726 294618 162768 294854
rect 162448 294586 162768 294618
rect 193168 295174 193488 295206
rect 193168 294938 193210 295174
rect 193446 294938 193488 295174
rect 193168 294854 193488 294938
rect 193168 294618 193210 294854
rect 193446 294618 193488 294854
rect 193168 294586 193488 294618
rect 223888 295174 224208 295206
rect 223888 294938 223930 295174
rect 224166 294938 224208 295174
rect 223888 294854 224208 294938
rect 223888 294618 223930 294854
rect 224166 294618 224208 294854
rect 223888 294586 224208 294618
rect 254608 295174 254928 295206
rect 254608 294938 254650 295174
rect 254886 294938 254928 295174
rect 254608 294854 254928 294938
rect 254608 294618 254650 294854
rect 254886 294618 254928 294854
rect 254608 294586 254928 294618
rect 285328 295174 285648 295206
rect 285328 294938 285370 295174
rect 285606 294938 285648 295174
rect 285328 294854 285648 294938
rect 285328 294618 285370 294854
rect 285606 294618 285648 294854
rect 285328 294586 285648 294618
rect 316048 295174 316368 295206
rect 316048 294938 316090 295174
rect 316326 294938 316368 295174
rect 316048 294854 316368 294938
rect 316048 294618 316090 294854
rect 316326 294618 316368 294854
rect 316048 294586 316368 294618
rect 346768 295174 347088 295206
rect 346768 294938 346810 295174
rect 347046 294938 347088 295174
rect 346768 294854 347088 294938
rect 346768 294618 346810 294854
rect 347046 294618 347088 294854
rect 346768 294586 347088 294618
rect 54928 291454 55248 291486
rect 54928 291218 54970 291454
rect 55206 291218 55248 291454
rect 54928 291134 55248 291218
rect 54928 290898 54970 291134
rect 55206 290898 55248 291134
rect 54928 290866 55248 290898
rect 85648 291454 85968 291486
rect 85648 291218 85690 291454
rect 85926 291218 85968 291454
rect 85648 291134 85968 291218
rect 85648 290898 85690 291134
rect 85926 290898 85968 291134
rect 85648 290866 85968 290898
rect 116368 291454 116688 291486
rect 116368 291218 116410 291454
rect 116646 291218 116688 291454
rect 116368 291134 116688 291218
rect 116368 290898 116410 291134
rect 116646 290898 116688 291134
rect 116368 290866 116688 290898
rect 147088 291454 147408 291486
rect 147088 291218 147130 291454
rect 147366 291218 147408 291454
rect 147088 291134 147408 291218
rect 147088 290898 147130 291134
rect 147366 290898 147408 291134
rect 147088 290866 147408 290898
rect 177808 291454 178128 291486
rect 177808 291218 177850 291454
rect 178086 291218 178128 291454
rect 177808 291134 178128 291218
rect 177808 290898 177850 291134
rect 178086 290898 178128 291134
rect 177808 290866 178128 290898
rect 208528 291454 208848 291486
rect 208528 291218 208570 291454
rect 208806 291218 208848 291454
rect 208528 291134 208848 291218
rect 208528 290898 208570 291134
rect 208806 290898 208848 291134
rect 208528 290866 208848 290898
rect 239248 291454 239568 291486
rect 239248 291218 239290 291454
rect 239526 291218 239568 291454
rect 239248 291134 239568 291218
rect 239248 290898 239290 291134
rect 239526 290898 239568 291134
rect 239248 290866 239568 290898
rect 269968 291454 270288 291486
rect 269968 291218 270010 291454
rect 270246 291218 270288 291454
rect 269968 291134 270288 291218
rect 269968 290898 270010 291134
rect 270246 290898 270288 291134
rect 269968 290866 270288 290898
rect 300688 291454 301008 291486
rect 300688 291218 300730 291454
rect 300966 291218 301008 291454
rect 300688 291134 301008 291218
rect 300688 290898 300730 291134
rect 300966 290898 301008 291134
rect 300688 290866 301008 290898
rect 331408 291454 331728 291486
rect 331408 291218 331450 291454
rect 331686 291218 331728 291454
rect 331408 291134 331728 291218
rect 331408 290898 331450 291134
rect 331686 290898 331728 291134
rect 331408 290866 331728 290898
rect 361794 291454 362414 326898
rect 361794 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 362414 291454
rect 361794 291134 362414 291218
rect 361794 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 362414 291134
rect 27834 281258 27866 281494
rect 28102 281258 28186 281494
rect 28422 281258 28454 281494
rect 27834 281174 28454 281258
rect 27834 280938 27866 281174
rect 28102 280938 28186 281174
rect 28422 280938 28454 281174
rect 24208 255454 24528 255486
rect 24208 255218 24250 255454
rect 24486 255218 24528 255454
rect 24208 255134 24528 255218
rect 24208 254898 24250 255134
rect 24486 254898 24528 255134
rect 24208 254866 24528 254898
rect 20394 237818 20426 238054
rect 20662 237818 20746 238054
rect 20982 237818 21014 238054
rect 20394 237734 21014 237818
rect 20394 237498 20426 237734
rect 20662 237498 20746 237734
rect 20982 237498 21014 237734
rect 20394 202054 21014 237498
rect 27834 245494 28454 280938
rect 39568 259174 39888 259206
rect 39568 258938 39610 259174
rect 39846 258938 39888 259174
rect 39568 258854 39888 258938
rect 39568 258618 39610 258854
rect 39846 258618 39888 258854
rect 39568 258586 39888 258618
rect 70288 259174 70608 259206
rect 70288 258938 70330 259174
rect 70566 258938 70608 259174
rect 70288 258854 70608 258938
rect 70288 258618 70330 258854
rect 70566 258618 70608 258854
rect 70288 258586 70608 258618
rect 101008 259174 101328 259206
rect 101008 258938 101050 259174
rect 101286 258938 101328 259174
rect 101008 258854 101328 258938
rect 101008 258618 101050 258854
rect 101286 258618 101328 258854
rect 101008 258586 101328 258618
rect 131728 259174 132048 259206
rect 131728 258938 131770 259174
rect 132006 258938 132048 259174
rect 131728 258854 132048 258938
rect 131728 258618 131770 258854
rect 132006 258618 132048 258854
rect 131728 258586 132048 258618
rect 162448 259174 162768 259206
rect 162448 258938 162490 259174
rect 162726 258938 162768 259174
rect 162448 258854 162768 258938
rect 162448 258618 162490 258854
rect 162726 258618 162768 258854
rect 162448 258586 162768 258618
rect 193168 259174 193488 259206
rect 193168 258938 193210 259174
rect 193446 258938 193488 259174
rect 193168 258854 193488 258938
rect 193168 258618 193210 258854
rect 193446 258618 193488 258854
rect 193168 258586 193488 258618
rect 223888 259174 224208 259206
rect 223888 258938 223930 259174
rect 224166 258938 224208 259174
rect 223888 258854 224208 258938
rect 223888 258618 223930 258854
rect 224166 258618 224208 258854
rect 223888 258586 224208 258618
rect 254608 259174 254928 259206
rect 254608 258938 254650 259174
rect 254886 258938 254928 259174
rect 254608 258854 254928 258938
rect 254608 258618 254650 258854
rect 254886 258618 254928 258854
rect 254608 258586 254928 258618
rect 285328 259174 285648 259206
rect 285328 258938 285370 259174
rect 285606 258938 285648 259174
rect 285328 258854 285648 258938
rect 285328 258618 285370 258854
rect 285606 258618 285648 258854
rect 285328 258586 285648 258618
rect 316048 259174 316368 259206
rect 316048 258938 316090 259174
rect 316326 258938 316368 259174
rect 316048 258854 316368 258938
rect 316048 258618 316090 258854
rect 316326 258618 316368 258854
rect 316048 258586 316368 258618
rect 346768 259174 347088 259206
rect 346768 258938 346810 259174
rect 347046 258938 347088 259174
rect 346768 258854 347088 258938
rect 346768 258618 346810 258854
rect 347046 258618 347088 258854
rect 346768 258586 347088 258618
rect 54928 255454 55248 255486
rect 54928 255218 54970 255454
rect 55206 255218 55248 255454
rect 54928 255134 55248 255218
rect 54928 254898 54970 255134
rect 55206 254898 55248 255134
rect 54928 254866 55248 254898
rect 85648 255454 85968 255486
rect 85648 255218 85690 255454
rect 85926 255218 85968 255454
rect 85648 255134 85968 255218
rect 85648 254898 85690 255134
rect 85926 254898 85968 255134
rect 85648 254866 85968 254898
rect 116368 255454 116688 255486
rect 116368 255218 116410 255454
rect 116646 255218 116688 255454
rect 116368 255134 116688 255218
rect 116368 254898 116410 255134
rect 116646 254898 116688 255134
rect 116368 254866 116688 254898
rect 147088 255454 147408 255486
rect 147088 255218 147130 255454
rect 147366 255218 147408 255454
rect 147088 255134 147408 255218
rect 147088 254898 147130 255134
rect 147366 254898 147408 255134
rect 147088 254866 147408 254898
rect 177808 255454 178128 255486
rect 177808 255218 177850 255454
rect 178086 255218 178128 255454
rect 177808 255134 178128 255218
rect 177808 254898 177850 255134
rect 178086 254898 178128 255134
rect 177808 254866 178128 254898
rect 208528 255454 208848 255486
rect 208528 255218 208570 255454
rect 208806 255218 208848 255454
rect 208528 255134 208848 255218
rect 208528 254898 208570 255134
rect 208806 254898 208848 255134
rect 208528 254866 208848 254898
rect 239248 255454 239568 255486
rect 239248 255218 239290 255454
rect 239526 255218 239568 255454
rect 239248 255134 239568 255218
rect 239248 254898 239290 255134
rect 239526 254898 239568 255134
rect 239248 254866 239568 254898
rect 269968 255454 270288 255486
rect 269968 255218 270010 255454
rect 270246 255218 270288 255454
rect 269968 255134 270288 255218
rect 269968 254898 270010 255134
rect 270246 254898 270288 255134
rect 269968 254866 270288 254898
rect 300688 255454 301008 255486
rect 300688 255218 300730 255454
rect 300966 255218 301008 255454
rect 300688 255134 301008 255218
rect 300688 254898 300730 255134
rect 300966 254898 301008 255134
rect 300688 254866 301008 254898
rect 331408 255454 331728 255486
rect 331408 255218 331450 255454
rect 331686 255218 331728 255454
rect 331408 255134 331728 255218
rect 331408 254898 331450 255134
rect 331686 254898 331728 255134
rect 331408 254866 331728 254898
rect 361794 255454 362414 290898
rect 361794 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 362414 255454
rect 361794 255134 362414 255218
rect 361794 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 362414 255134
rect 27834 245258 27866 245494
rect 28102 245258 28186 245494
rect 28422 245258 28454 245494
rect 27834 245174 28454 245258
rect 27834 244938 27866 245174
rect 28102 244938 28186 245174
rect 28422 244938 28454 245174
rect 24208 219454 24528 219486
rect 24208 219218 24250 219454
rect 24486 219218 24528 219454
rect 24208 219134 24528 219218
rect 24208 218898 24250 219134
rect 24486 218898 24528 219134
rect 24208 218866 24528 218898
rect 20394 201818 20426 202054
rect 20662 201818 20746 202054
rect 20982 201818 21014 202054
rect 20394 201734 21014 201818
rect 20394 201498 20426 201734
rect 20662 201498 20746 201734
rect 20982 201498 21014 201734
rect 20394 166054 21014 201498
rect 27834 209494 28454 244938
rect 39568 223174 39888 223206
rect 39568 222938 39610 223174
rect 39846 222938 39888 223174
rect 39568 222854 39888 222938
rect 39568 222618 39610 222854
rect 39846 222618 39888 222854
rect 39568 222586 39888 222618
rect 70288 223174 70608 223206
rect 70288 222938 70330 223174
rect 70566 222938 70608 223174
rect 70288 222854 70608 222938
rect 70288 222618 70330 222854
rect 70566 222618 70608 222854
rect 70288 222586 70608 222618
rect 101008 223174 101328 223206
rect 101008 222938 101050 223174
rect 101286 222938 101328 223174
rect 101008 222854 101328 222938
rect 101008 222618 101050 222854
rect 101286 222618 101328 222854
rect 101008 222586 101328 222618
rect 131728 223174 132048 223206
rect 131728 222938 131770 223174
rect 132006 222938 132048 223174
rect 131728 222854 132048 222938
rect 131728 222618 131770 222854
rect 132006 222618 132048 222854
rect 131728 222586 132048 222618
rect 162448 223174 162768 223206
rect 162448 222938 162490 223174
rect 162726 222938 162768 223174
rect 162448 222854 162768 222938
rect 162448 222618 162490 222854
rect 162726 222618 162768 222854
rect 162448 222586 162768 222618
rect 193168 223174 193488 223206
rect 193168 222938 193210 223174
rect 193446 222938 193488 223174
rect 193168 222854 193488 222938
rect 193168 222618 193210 222854
rect 193446 222618 193488 222854
rect 193168 222586 193488 222618
rect 223888 223174 224208 223206
rect 223888 222938 223930 223174
rect 224166 222938 224208 223174
rect 223888 222854 224208 222938
rect 223888 222618 223930 222854
rect 224166 222618 224208 222854
rect 223888 222586 224208 222618
rect 254608 223174 254928 223206
rect 254608 222938 254650 223174
rect 254886 222938 254928 223174
rect 254608 222854 254928 222938
rect 254608 222618 254650 222854
rect 254886 222618 254928 222854
rect 254608 222586 254928 222618
rect 285328 223174 285648 223206
rect 285328 222938 285370 223174
rect 285606 222938 285648 223174
rect 285328 222854 285648 222938
rect 285328 222618 285370 222854
rect 285606 222618 285648 222854
rect 285328 222586 285648 222618
rect 316048 223174 316368 223206
rect 316048 222938 316090 223174
rect 316326 222938 316368 223174
rect 316048 222854 316368 222938
rect 316048 222618 316090 222854
rect 316326 222618 316368 222854
rect 316048 222586 316368 222618
rect 346768 223174 347088 223206
rect 346768 222938 346810 223174
rect 347046 222938 347088 223174
rect 346768 222854 347088 222938
rect 346768 222618 346810 222854
rect 347046 222618 347088 222854
rect 346768 222586 347088 222618
rect 54928 219454 55248 219486
rect 54928 219218 54970 219454
rect 55206 219218 55248 219454
rect 54928 219134 55248 219218
rect 54928 218898 54970 219134
rect 55206 218898 55248 219134
rect 54928 218866 55248 218898
rect 85648 219454 85968 219486
rect 85648 219218 85690 219454
rect 85926 219218 85968 219454
rect 85648 219134 85968 219218
rect 85648 218898 85690 219134
rect 85926 218898 85968 219134
rect 85648 218866 85968 218898
rect 116368 219454 116688 219486
rect 116368 219218 116410 219454
rect 116646 219218 116688 219454
rect 116368 219134 116688 219218
rect 116368 218898 116410 219134
rect 116646 218898 116688 219134
rect 116368 218866 116688 218898
rect 147088 219454 147408 219486
rect 147088 219218 147130 219454
rect 147366 219218 147408 219454
rect 147088 219134 147408 219218
rect 147088 218898 147130 219134
rect 147366 218898 147408 219134
rect 147088 218866 147408 218898
rect 177808 219454 178128 219486
rect 177808 219218 177850 219454
rect 178086 219218 178128 219454
rect 177808 219134 178128 219218
rect 177808 218898 177850 219134
rect 178086 218898 178128 219134
rect 177808 218866 178128 218898
rect 208528 219454 208848 219486
rect 208528 219218 208570 219454
rect 208806 219218 208848 219454
rect 208528 219134 208848 219218
rect 208528 218898 208570 219134
rect 208806 218898 208848 219134
rect 208528 218866 208848 218898
rect 239248 219454 239568 219486
rect 239248 219218 239290 219454
rect 239526 219218 239568 219454
rect 239248 219134 239568 219218
rect 239248 218898 239290 219134
rect 239526 218898 239568 219134
rect 239248 218866 239568 218898
rect 269968 219454 270288 219486
rect 269968 219218 270010 219454
rect 270246 219218 270288 219454
rect 269968 219134 270288 219218
rect 269968 218898 270010 219134
rect 270246 218898 270288 219134
rect 269968 218866 270288 218898
rect 300688 219454 301008 219486
rect 300688 219218 300730 219454
rect 300966 219218 301008 219454
rect 300688 219134 301008 219218
rect 300688 218898 300730 219134
rect 300966 218898 301008 219134
rect 300688 218866 301008 218898
rect 331408 219454 331728 219486
rect 331408 219218 331450 219454
rect 331686 219218 331728 219454
rect 331408 219134 331728 219218
rect 331408 218898 331450 219134
rect 331686 218898 331728 219134
rect 331408 218866 331728 218898
rect 361794 219454 362414 254898
rect 361794 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 362414 219454
rect 361794 219134 362414 219218
rect 361794 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 362414 219134
rect 27834 209258 27866 209494
rect 28102 209258 28186 209494
rect 28422 209258 28454 209494
rect 27834 209174 28454 209258
rect 27834 208938 27866 209174
rect 28102 208938 28186 209174
rect 28422 208938 28454 209174
rect 24208 183454 24528 183486
rect 24208 183218 24250 183454
rect 24486 183218 24528 183454
rect 24208 183134 24528 183218
rect 24208 182898 24250 183134
rect 24486 182898 24528 183134
rect 24208 182866 24528 182898
rect 20394 165818 20426 166054
rect 20662 165818 20746 166054
rect 20982 165818 21014 166054
rect 20394 165734 21014 165818
rect 20394 165498 20426 165734
rect 20662 165498 20746 165734
rect 20982 165498 21014 165734
rect 20394 130054 21014 165498
rect 27834 173494 28454 208938
rect 39568 187174 39888 187206
rect 39568 186938 39610 187174
rect 39846 186938 39888 187174
rect 39568 186854 39888 186938
rect 39568 186618 39610 186854
rect 39846 186618 39888 186854
rect 39568 186586 39888 186618
rect 70288 187174 70608 187206
rect 70288 186938 70330 187174
rect 70566 186938 70608 187174
rect 70288 186854 70608 186938
rect 70288 186618 70330 186854
rect 70566 186618 70608 186854
rect 70288 186586 70608 186618
rect 101008 187174 101328 187206
rect 101008 186938 101050 187174
rect 101286 186938 101328 187174
rect 101008 186854 101328 186938
rect 101008 186618 101050 186854
rect 101286 186618 101328 186854
rect 101008 186586 101328 186618
rect 131728 187174 132048 187206
rect 131728 186938 131770 187174
rect 132006 186938 132048 187174
rect 131728 186854 132048 186938
rect 131728 186618 131770 186854
rect 132006 186618 132048 186854
rect 131728 186586 132048 186618
rect 162448 187174 162768 187206
rect 162448 186938 162490 187174
rect 162726 186938 162768 187174
rect 162448 186854 162768 186938
rect 162448 186618 162490 186854
rect 162726 186618 162768 186854
rect 162448 186586 162768 186618
rect 193168 187174 193488 187206
rect 193168 186938 193210 187174
rect 193446 186938 193488 187174
rect 193168 186854 193488 186938
rect 193168 186618 193210 186854
rect 193446 186618 193488 186854
rect 193168 186586 193488 186618
rect 223888 187174 224208 187206
rect 223888 186938 223930 187174
rect 224166 186938 224208 187174
rect 223888 186854 224208 186938
rect 223888 186618 223930 186854
rect 224166 186618 224208 186854
rect 223888 186586 224208 186618
rect 254608 187174 254928 187206
rect 254608 186938 254650 187174
rect 254886 186938 254928 187174
rect 254608 186854 254928 186938
rect 254608 186618 254650 186854
rect 254886 186618 254928 186854
rect 254608 186586 254928 186618
rect 285328 187174 285648 187206
rect 285328 186938 285370 187174
rect 285606 186938 285648 187174
rect 285328 186854 285648 186938
rect 285328 186618 285370 186854
rect 285606 186618 285648 186854
rect 285328 186586 285648 186618
rect 316048 187174 316368 187206
rect 316048 186938 316090 187174
rect 316326 186938 316368 187174
rect 316048 186854 316368 186938
rect 316048 186618 316090 186854
rect 316326 186618 316368 186854
rect 316048 186586 316368 186618
rect 346768 187174 347088 187206
rect 346768 186938 346810 187174
rect 347046 186938 347088 187174
rect 346768 186854 347088 186938
rect 346768 186618 346810 186854
rect 347046 186618 347088 186854
rect 346768 186586 347088 186618
rect 54928 183454 55248 183486
rect 54928 183218 54970 183454
rect 55206 183218 55248 183454
rect 54928 183134 55248 183218
rect 54928 182898 54970 183134
rect 55206 182898 55248 183134
rect 54928 182866 55248 182898
rect 85648 183454 85968 183486
rect 85648 183218 85690 183454
rect 85926 183218 85968 183454
rect 85648 183134 85968 183218
rect 85648 182898 85690 183134
rect 85926 182898 85968 183134
rect 85648 182866 85968 182898
rect 116368 183454 116688 183486
rect 116368 183218 116410 183454
rect 116646 183218 116688 183454
rect 116368 183134 116688 183218
rect 116368 182898 116410 183134
rect 116646 182898 116688 183134
rect 116368 182866 116688 182898
rect 147088 183454 147408 183486
rect 147088 183218 147130 183454
rect 147366 183218 147408 183454
rect 147088 183134 147408 183218
rect 147088 182898 147130 183134
rect 147366 182898 147408 183134
rect 147088 182866 147408 182898
rect 177808 183454 178128 183486
rect 177808 183218 177850 183454
rect 178086 183218 178128 183454
rect 177808 183134 178128 183218
rect 177808 182898 177850 183134
rect 178086 182898 178128 183134
rect 177808 182866 178128 182898
rect 208528 183454 208848 183486
rect 208528 183218 208570 183454
rect 208806 183218 208848 183454
rect 208528 183134 208848 183218
rect 208528 182898 208570 183134
rect 208806 182898 208848 183134
rect 208528 182866 208848 182898
rect 239248 183454 239568 183486
rect 239248 183218 239290 183454
rect 239526 183218 239568 183454
rect 239248 183134 239568 183218
rect 239248 182898 239290 183134
rect 239526 182898 239568 183134
rect 239248 182866 239568 182898
rect 269968 183454 270288 183486
rect 269968 183218 270010 183454
rect 270246 183218 270288 183454
rect 269968 183134 270288 183218
rect 269968 182898 270010 183134
rect 270246 182898 270288 183134
rect 269968 182866 270288 182898
rect 300688 183454 301008 183486
rect 300688 183218 300730 183454
rect 300966 183218 301008 183454
rect 300688 183134 301008 183218
rect 300688 182898 300730 183134
rect 300966 182898 301008 183134
rect 300688 182866 301008 182898
rect 331408 183454 331728 183486
rect 331408 183218 331450 183454
rect 331686 183218 331728 183454
rect 331408 183134 331728 183218
rect 331408 182898 331450 183134
rect 331686 182898 331728 183134
rect 331408 182866 331728 182898
rect 361794 183454 362414 218898
rect 361794 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 362414 183454
rect 361794 183134 362414 183218
rect 361794 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 362414 183134
rect 27834 173258 27866 173494
rect 28102 173258 28186 173494
rect 28422 173258 28454 173494
rect 27834 173174 28454 173258
rect 27834 172938 27866 173174
rect 28102 172938 28186 173174
rect 28422 172938 28454 173174
rect 24208 147454 24528 147486
rect 24208 147218 24250 147454
rect 24486 147218 24528 147454
rect 24208 147134 24528 147218
rect 24208 146898 24250 147134
rect 24486 146898 24528 147134
rect 24208 146866 24528 146898
rect 20394 129818 20426 130054
rect 20662 129818 20746 130054
rect 20982 129818 21014 130054
rect 20394 129734 21014 129818
rect 20394 129498 20426 129734
rect 20662 129498 20746 129734
rect 20982 129498 21014 129734
rect 20394 94054 21014 129498
rect 27834 137494 28454 172938
rect 39568 151174 39888 151206
rect 39568 150938 39610 151174
rect 39846 150938 39888 151174
rect 39568 150854 39888 150938
rect 39568 150618 39610 150854
rect 39846 150618 39888 150854
rect 39568 150586 39888 150618
rect 70288 151174 70608 151206
rect 70288 150938 70330 151174
rect 70566 150938 70608 151174
rect 70288 150854 70608 150938
rect 70288 150618 70330 150854
rect 70566 150618 70608 150854
rect 70288 150586 70608 150618
rect 101008 151174 101328 151206
rect 101008 150938 101050 151174
rect 101286 150938 101328 151174
rect 101008 150854 101328 150938
rect 101008 150618 101050 150854
rect 101286 150618 101328 150854
rect 101008 150586 101328 150618
rect 131728 151174 132048 151206
rect 131728 150938 131770 151174
rect 132006 150938 132048 151174
rect 131728 150854 132048 150938
rect 131728 150618 131770 150854
rect 132006 150618 132048 150854
rect 131728 150586 132048 150618
rect 162448 151174 162768 151206
rect 162448 150938 162490 151174
rect 162726 150938 162768 151174
rect 162448 150854 162768 150938
rect 162448 150618 162490 150854
rect 162726 150618 162768 150854
rect 162448 150586 162768 150618
rect 193168 151174 193488 151206
rect 193168 150938 193210 151174
rect 193446 150938 193488 151174
rect 193168 150854 193488 150938
rect 193168 150618 193210 150854
rect 193446 150618 193488 150854
rect 193168 150586 193488 150618
rect 223888 151174 224208 151206
rect 223888 150938 223930 151174
rect 224166 150938 224208 151174
rect 223888 150854 224208 150938
rect 223888 150618 223930 150854
rect 224166 150618 224208 150854
rect 223888 150586 224208 150618
rect 254608 151174 254928 151206
rect 254608 150938 254650 151174
rect 254886 150938 254928 151174
rect 254608 150854 254928 150938
rect 254608 150618 254650 150854
rect 254886 150618 254928 150854
rect 254608 150586 254928 150618
rect 285328 151174 285648 151206
rect 285328 150938 285370 151174
rect 285606 150938 285648 151174
rect 285328 150854 285648 150938
rect 285328 150618 285370 150854
rect 285606 150618 285648 150854
rect 285328 150586 285648 150618
rect 316048 151174 316368 151206
rect 316048 150938 316090 151174
rect 316326 150938 316368 151174
rect 316048 150854 316368 150938
rect 316048 150618 316090 150854
rect 316326 150618 316368 150854
rect 316048 150586 316368 150618
rect 346768 151174 347088 151206
rect 346768 150938 346810 151174
rect 347046 150938 347088 151174
rect 346768 150854 347088 150938
rect 346768 150618 346810 150854
rect 347046 150618 347088 150854
rect 346768 150586 347088 150618
rect 54928 147454 55248 147486
rect 54928 147218 54970 147454
rect 55206 147218 55248 147454
rect 54928 147134 55248 147218
rect 54928 146898 54970 147134
rect 55206 146898 55248 147134
rect 54928 146866 55248 146898
rect 85648 147454 85968 147486
rect 85648 147218 85690 147454
rect 85926 147218 85968 147454
rect 85648 147134 85968 147218
rect 85648 146898 85690 147134
rect 85926 146898 85968 147134
rect 85648 146866 85968 146898
rect 116368 147454 116688 147486
rect 116368 147218 116410 147454
rect 116646 147218 116688 147454
rect 116368 147134 116688 147218
rect 116368 146898 116410 147134
rect 116646 146898 116688 147134
rect 116368 146866 116688 146898
rect 147088 147454 147408 147486
rect 147088 147218 147130 147454
rect 147366 147218 147408 147454
rect 147088 147134 147408 147218
rect 147088 146898 147130 147134
rect 147366 146898 147408 147134
rect 147088 146866 147408 146898
rect 177808 147454 178128 147486
rect 177808 147218 177850 147454
rect 178086 147218 178128 147454
rect 177808 147134 178128 147218
rect 177808 146898 177850 147134
rect 178086 146898 178128 147134
rect 177808 146866 178128 146898
rect 208528 147454 208848 147486
rect 208528 147218 208570 147454
rect 208806 147218 208848 147454
rect 208528 147134 208848 147218
rect 208528 146898 208570 147134
rect 208806 146898 208848 147134
rect 208528 146866 208848 146898
rect 239248 147454 239568 147486
rect 239248 147218 239290 147454
rect 239526 147218 239568 147454
rect 239248 147134 239568 147218
rect 239248 146898 239290 147134
rect 239526 146898 239568 147134
rect 239248 146866 239568 146898
rect 269968 147454 270288 147486
rect 269968 147218 270010 147454
rect 270246 147218 270288 147454
rect 269968 147134 270288 147218
rect 269968 146898 270010 147134
rect 270246 146898 270288 147134
rect 269968 146866 270288 146898
rect 300688 147454 301008 147486
rect 300688 147218 300730 147454
rect 300966 147218 301008 147454
rect 300688 147134 301008 147218
rect 300688 146898 300730 147134
rect 300966 146898 301008 147134
rect 300688 146866 301008 146898
rect 331408 147454 331728 147486
rect 331408 147218 331450 147454
rect 331686 147218 331728 147454
rect 331408 147134 331728 147218
rect 331408 146898 331450 147134
rect 331686 146898 331728 147134
rect 331408 146866 331728 146898
rect 361794 147454 362414 182898
rect 361794 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 362414 147454
rect 361794 147134 362414 147218
rect 361794 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 362414 147134
rect 27834 137258 27866 137494
rect 28102 137258 28186 137494
rect 28422 137258 28454 137494
rect 27834 137174 28454 137258
rect 27834 136938 27866 137174
rect 28102 136938 28186 137174
rect 28422 136938 28454 137174
rect 24208 111454 24528 111486
rect 24208 111218 24250 111454
rect 24486 111218 24528 111454
rect 24208 111134 24528 111218
rect 24208 110898 24250 111134
rect 24486 110898 24528 111134
rect 24208 110866 24528 110898
rect 20394 93818 20426 94054
rect 20662 93818 20746 94054
rect 20982 93818 21014 94054
rect 20394 93734 21014 93818
rect 20394 93498 20426 93734
rect 20662 93498 20746 93734
rect 20982 93498 21014 93734
rect 20394 58054 21014 93498
rect 27834 101494 28454 136938
rect 39568 115174 39888 115206
rect 39568 114938 39610 115174
rect 39846 114938 39888 115174
rect 39568 114854 39888 114938
rect 39568 114618 39610 114854
rect 39846 114618 39888 114854
rect 39568 114586 39888 114618
rect 70288 115174 70608 115206
rect 70288 114938 70330 115174
rect 70566 114938 70608 115174
rect 70288 114854 70608 114938
rect 70288 114618 70330 114854
rect 70566 114618 70608 114854
rect 70288 114586 70608 114618
rect 101008 115174 101328 115206
rect 101008 114938 101050 115174
rect 101286 114938 101328 115174
rect 101008 114854 101328 114938
rect 101008 114618 101050 114854
rect 101286 114618 101328 114854
rect 101008 114586 101328 114618
rect 131728 115174 132048 115206
rect 131728 114938 131770 115174
rect 132006 114938 132048 115174
rect 131728 114854 132048 114938
rect 131728 114618 131770 114854
rect 132006 114618 132048 114854
rect 131728 114586 132048 114618
rect 162448 115174 162768 115206
rect 162448 114938 162490 115174
rect 162726 114938 162768 115174
rect 162448 114854 162768 114938
rect 162448 114618 162490 114854
rect 162726 114618 162768 114854
rect 162448 114586 162768 114618
rect 193168 115174 193488 115206
rect 193168 114938 193210 115174
rect 193446 114938 193488 115174
rect 193168 114854 193488 114938
rect 193168 114618 193210 114854
rect 193446 114618 193488 114854
rect 193168 114586 193488 114618
rect 223888 115174 224208 115206
rect 223888 114938 223930 115174
rect 224166 114938 224208 115174
rect 223888 114854 224208 114938
rect 223888 114618 223930 114854
rect 224166 114618 224208 114854
rect 223888 114586 224208 114618
rect 254608 115174 254928 115206
rect 254608 114938 254650 115174
rect 254886 114938 254928 115174
rect 254608 114854 254928 114938
rect 254608 114618 254650 114854
rect 254886 114618 254928 114854
rect 254608 114586 254928 114618
rect 285328 115174 285648 115206
rect 285328 114938 285370 115174
rect 285606 114938 285648 115174
rect 285328 114854 285648 114938
rect 285328 114618 285370 114854
rect 285606 114618 285648 114854
rect 285328 114586 285648 114618
rect 316048 115174 316368 115206
rect 316048 114938 316090 115174
rect 316326 114938 316368 115174
rect 316048 114854 316368 114938
rect 316048 114618 316090 114854
rect 316326 114618 316368 114854
rect 316048 114586 316368 114618
rect 346768 115174 347088 115206
rect 346768 114938 346810 115174
rect 347046 114938 347088 115174
rect 346768 114854 347088 114938
rect 346768 114618 346810 114854
rect 347046 114618 347088 114854
rect 346768 114586 347088 114618
rect 54928 111454 55248 111486
rect 54928 111218 54970 111454
rect 55206 111218 55248 111454
rect 54928 111134 55248 111218
rect 54928 110898 54970 111134
rect 55206 110898 55248 111134
rect 54928 110866 55248 110898
rect 85648 111454 85968 111486
rect 85648 111218 85690 111454
rect 85926 111218 85968 111454
rect 85648 111134 85968 111218
rect 85648 110898 85690 111134
rect 85926 110898 85968 111134
rect 85648 110866 85968 110898
rect 116368 111454 116688 111486
rect 116368 111218 116410 111454
rect 116646 111218 116688 111454
rect 116368 111134 116688 111218
rect 116368 110898 116410 111134
rect 116646 110898 116688 111134
rect 116368 110866 116688 110898
rect 147088 111454 147408 111486
rect 147088 111218 147130 111454
rect 147366 111218 147408 111454
rect 147088 111134 147408 111218
rect 147088 110898 147130 111134
rect 147366 110898 147408 111134
rect 147088 110866 147408 110898
rect 177808 111454 178128 111486
rect 177808 111218 177850 111454
rect 178086 111218 178128 111454
rect 177808 111134 178128 111218
rect 177808 110898 177850 111134
rect 178086 110898 178128 111134
rect 177808 110866 178128 110898
rect 208528 111454 208848 111486
rect 208528 111218 208570 111454
rect 208806 111218 208848 111454
rect 208528 111134 208848 111218
rect 208528 110898 208570 111134
rect 208806 110898 208848 111134
rect 208528 110866 208848 110898
rect 239248 111454 239568 111486
rect 239248 111218 239290 111454
rect 239526 111218 239568 111454
rect 239248 111134 239568 111218
rect 239248 110898 239290 111134
rect 239526 110898 239568 111134
rect 239248 110866 239568 110898
rect 269968 111454 270288 111486
rect 269968 111218 270010 111454
rect 270246 111218 270288 111454
rect 269968 111134 270288 111218
rect 269968 110898 270010 111134
rect 270246 110898 270288 111134
rect 269968 110866 270288 110898
rect 300688 111454 301008 111486
rect 300688 111218 300730 111454
rect 300966 111218 301008 111454
rect 300688 111134 301008 111218
rect 300688 110898 300730 111134
rect 300966 110898 301008 111134
rect 300688 110866 301008 110898
rect 331408 111454 331728 111486
rect 331408 111218 331450 111454
rect 331686 111218 331728 111454
rect 331408 111134 331728 111218
rect 331408 110898 331450 111134
rect 331686 110898 331728 111134
rect 331408 110866 331728 110898
rect 361794 111454 362414 146898
rect 361794 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 362414 111454
rect 361794 111134 362414 111218
rect 361794 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 362414 111134
rect 27834 101258 27866 101494
rect 28102 101258 28186 101494
rect 28422 101258 28454 101494
rect 27834 101174 28454 101258
rect 27834 100938 27866 101174
rect 28102 100938 28186 101174
rect 28422 100938 28454 101174
rect 24208 75454 24528 75486
rect 24208 75218 24250 75454
rect 24486 75218 24528 75454
rect 24208 75134 24528 75218
rect 24208 74898 24250 75134
rect 24486 74898 24528 75134
rect 24208 74866 24528 74898
rect 20394 57818 20426 58054
rect 20662 57818 20746 58054
rect 20982 57818 21014 58054
rect 20394 57734 21014 57818
rect 20394 57498 20426 57734
rect 20662 57498 20746 57734
rect 20982 57498 21014 57734
rect 20394 22054 21014 57498
rect 27834 65494 28454 100938
rect 39568 79174 39888 79206
rect 39568 78938 39610 79174
rect 39846 78938 39888 79174
rect 39568 78854 39888 78938
rect 39568 78618 39610 78854
rect 39846 78618 39888 78854
rect 39568 78586 39888 78618
rect 70288 79174 70608 79206
rect 70288 78938 70330 79174
rect 70566 78938 70608 79174
rect 70288 78854 70608 78938
rect 70288 78618 70330 78854
rect 70566 78618 70608 78854
rect 70288 78586 70608 78618
rect 101008 79174 101328 79206
rect 101008 78938 101050 79174
rect 101286 78938 101328 79174
rect 101008 78854 101328 78938
rect 101008 78618 101050 78854
rect 101286 78618 101328 78854
rect 101008 78586 101328 78618
rect 131728 79174 132048 79206
rect 131728 78938 131770 79174
rect 132006 78938 132048 79174
rect 131728 78854 132048 78938
rect 131728 78618 131770 78854
rect 132006 78618 132048 78854
rect 131728 78586 132048 78618
rect 162448 79174 162768 79206
rect 162448 78938 162490 79174
rect 162726 78938 162768 79174
rect 162448 78854 162768 78938
rect 162448 78618 162490 78854
rect 162726 78618 162768 78854
rect 162448 78586 162768 78618
rect 193168 79174 193488 79206
rect 193168 78938 193210 79174
rect 193446 78938 193488 79174
rect 193168 78854 193488 78938
rect 193168 78618 193210 78854
rect 193446 78618 193488 78854
rect 193168 78586 193488 78618
rect 223888 79174 224208 79206
rect 223888 78938 223930 79174
rect 224166 78938 224208 79174
rect 223888 78854 224208 78938
rect 223888 78618 223930 78854
rect 224166 78618 224208 78854
rect 223888 78586 224208 78618
rect 254608 79174 254928 79206
rect 254608 78938 254650 79174
rect 254886 78938 254928 79174
rect 254608 78854 254928 78938
rect 254608 78618 254650 78854
rect 254886 78618 254928 78854
rect 254608 78586 254928 78618
rect 285328 79174 285648 79206
rect 285328 78938 285370 79174
rect 285606 78938 285648 79174
rect 285328 78854 285648 78938
rect 285328 78618 285370 78854
rect 285606 78618 285648 78854
rect 285328 78586 285648 78618
rect 316048 79174 316368 79206
rect 316048 78938 316090 79174
rect 316326 78938 316368 79174
rect 316048 78854 316368 78938
rect 316048 78618 316090 78854
rect 316326 78618 316368 78854
rect 316048 78586 316368 78618
rect 346768 79174 347088 79206
rect 346768 78938 346810 79174
rect 347046 78938 347088 79174
rect 346768 78854 347088 78938
rect 346768 78618 346810 78854
rect 347046 78618 347088 78854
rect 346768 78586 347088 78618
rect 54928 75454 55248 75486
rect 54928 75218 54970 75454
rect 55206 75218 55248 75454
rect 54928 75134 55248 75218
rect 54928 74898 54970 75134
rect 55206 74898 55248 75134
rect 54928 74866 55248 74898
rect 85648 75454 85968 75486
rect 85648 75218 85690 75454
rect 85926 75218 85968 75454
rect 85648 75134 85968 75218
rect 85648 74898 85690 75134
rect 85926 74898 85968 75134
rect 85648 74866 85968 74898
rect 116368 75454 116688 75486
rect 116368 75218 116410 75454
rect 116646 75218 116688 75454
rect 116368 75134 116688 75218
rect 116368 74898 116410 75134
rect 116646 74898 116688 75134
rect 116368 74866 116688 74898
rect 147088 75454 147408 75486
rect 147088 75218 147130 75454
rect 147366 75218 147408 75454
rect 147088 75134 147408 75218
rect 147088 74898 147130 75134
rect 147366 74898 147408 75134
rect 147088 74866 147408 74898
rect 177808 75454 178128 75486
rect 177808 75218 177850 75454
rect 178086 75218 178128 75454
rect 177808 75134 178128 75218
rect 177808 74898 177850 75134
rect 178086 74898 178128 75134
rect 177808 74866 178128 74898
rect 208528 75454 208848 75486
rect 208528 75218 208570 75454
rect 208806 75218 208848 75454
rect 208528 75134 208848 75218
rect 208528 74898 208570 75134
rect 208806 74898 208848 75134
rect 208528 74866 208848 74898
rect 239248 75454 239568 75486
rect 239248 75218 239290 75454
rect 239526 75218 239568 75454
rect 239248 75134 239568 75218
rect 239248 74898 239290 75134
rect 239526 74898 239568 75134
rect 239248 74866 239568 74898
rect 269968 75454 270288 75486
rect 269968 75218 270010 75454
rect 270246 75218 270288 75454
rect 269968 75134 270288 75218
rect 269968 74898 270010 75134
rect 270246 74898 270288 75134
rect 269968 74866 270288 74898
rect 300688 75454 301008 75486
rect 300688 75218 300730 75454
rect 300966 75218 301008 75454
rect 300688 75134 301008 75218
rect 300688 74898 300730 75134
rect 300966 74898 301008 75134
rect 300688 74866 301008 74898
rect 331408 75454 331728 75486
rect 331408 75218 331450 75454
rect 331686 75218 331728 75454
rect 331408 75134 331728 75218
rect 331408 74898 331450 75134
rect 331686 74898 331728 75134
rect 331408 74866 331728 74898
rect 361794 75454 362414 110898
rect 361794 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 362414 75454
rect 361794 75134 362414 75218
rect 361794 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 362414 75134
rect 27834 65258 27866 65494
rect 28102 65258 28186 65494
rect 28422 65258 28454 65494
rect 27834 65174 28454 65258
rect 27834 64938 27866 65174
rect 28102 64938 28186 65174
rect 28422 64938 28454 65174
rect 22323 49332 22389 49333
rect 22323 49268 22324 49332
rect 22388 49268 22389 49332
rect 22323 49267 22389 49268
rect 22139 48924 22205 48925
rect 22139 48860 22140 48924
rect 22204 48860 22205 48924
rect 22139 48859 22205 48860
rect 22142 46477 22202 48859
rect 22139 46476 22205 46477
rect 22139 46412 22140 46476
rect 22204 46412 22205 46476
rect 22139 46411 22205 46412
rect 22326 46341 22386 49267
rect 22323 46340 22389 46341
rect 22323 46276 22324 46340
rect 22388 46276 22389 46340
rect 22323 46275 22389 46276
rect 20394 21818 20426 22054
rect 20662 21818 20746 22054
rect 20982 21818 21014 22054
rect 20394 21734 21014 21818
rect 20394 21498 20426 21734
rect 20662 21498 20746 21734
rect 20982 21498 21014 21734
rect 20394 -5146 21014 21498
rect 20394 -5382 20426 -5146
rect 20662 -5382 20746 -5146
rect 20982 -5382 21014 -5146
rect 20394 -5466 21014 -5382
rect 20394 -5702 20426 -5466
rect 20662 -5702 20746 -5466
rect 20982 -5702 21014 -5466
rect 20394 -7654 21014 -5702
rect 24114 25774 24734 45068
rect 24114 25538 24146 25774
rect 24382 25538 24466 25774
rect 24702 25538 24734 25774
rect 24114 25454 24734 25538
rect 24114 25218 24146 25454
rect 24382 25218 24466 25454
rect 24702 25218 24734 25454
rect 24114 -6106 24734 25218
rect 24114 -6342 24146 -6106
rect 24382 -6342 24466 -6106
rect 24702 -6342 24734 -6106
rect 24114 -6426 24734 -6342
rect 24114 -6662 24146 -6426
rect 24382 -6662 24466 -6426
rect 24702 -6662 24734 -6426
rect 24114 -7654 24734 -6662
rect 27834 29494 28454 64938
rect 27834 29258 27866 29494
rect 28102 29258 28186 29494
rect 28422 29258 28454 29494
rect 27834 29174 28454 29258
rect 27834 28938 27866 29174
rect 28102 28938 28186 29174
rect 28422 28938 28454 29174
rect 27834 -7066 28454 28938
rect 27834 -7302 27866 -7066
rect 28102 -7302 28186 -7066
rect 28422 -7302 28454 -7066
rect 27834 -7386 28454 -7302
rect 27834 -7622 27866 -7386
rect 28102 -7622 28186 -7386
rect 28422 -7622 28454 -7386
rect 27834 -7654 28454 -7622
rect 37794 39454 38414 49367
rect 37794 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 38414 39454
rect 37794 39134 38414 39218
rect 37794 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 38414 39134
rect 37794 3454 38414 38898
rect 37794 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 38414 3454
rect 37794 3134 38414 3218
rect 37794 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 38414 3134
rect 37794 -346 38414 2898
rect 37794 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 38414 -346
rect 37794 -666 38414 -582
rect 37794 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 38414 -666
rect 37794 -7654 38414 -902
rect 41514 43174 42134 49367
rect 41514 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 42134 43174
rect 41514 42854 42134 42938
rect 41514 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 42134 42854
rect 41514 7174 42134 42618
rect 41514 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 42134 7174
rect 41514 6854 42134 6938
rect 41514 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 42134 6854
rect 41514 -1306 42134 6618
rect 41514 -1542 41546 -1306
rect 41782 -1542 41866 -1306
rect 42102 -1542 42134 -1306
rect 41514 -1626 42134 -1542
rect 41514 -1862 41546 -1626
rect 41782 -1862 41866 -1626
rect 42102 -1862 42134 -1626
rect 41514 -7654 42134 -1862
rect 45234 46894 45854 49367
rect 45234 46658 45266 46894
rect 45502 46658 45586 46894
rect 45822 46658 45854 46894
rect 45234 46574 45854 46658
rect 45234 46338 45266 46574
rect 45502 46338 45586 46574
rect 45822 46338 45854 46574
rect 45234 10894 45854 46338
rect 45234 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 45854 10894
rect 45234 10574 45854 10658
rect 45234 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 45854 10574
rect 45234 -2266 45854 10338
rect 45234 -2502 45266 -2266
rect 45502 -2502 45586 -2266
rect 45822 -2502 45854 -2266
rect 45234 -2586 45854 -2502
rect 45234 -2822 45266 -2586
rect 45502 -2822 45586 -2586
rect 45822 -2822 45854 -2586
rect 45234 -7654 45854 -2822
rect 48954 14614 49574 49367
rect 48954 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 49574 14614
rect 48954 14294 49574 14378
rect 48954 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 49574 14294
rect 48954 -3226 49574 14058
rect 48954 -3462 48986 -3226
rect 49222 -3462 49306 -3226
rect 49542 -3462 49574 -3226
rect 48954 -3546 49574 -3462
rect 48954 -3782 48986 -3546
rect 49222 -3782 49306 -3546
rect 49542 -3782 49574 -3546
rect 48954 -7654 49574 -3782
rect 52674 18334 53294 49367
rect 52674 18098 52706 18334
rect 52942 18098 53026 18334
rect 53262 18098 53294 18334
rect 52674 18014 53294 18098
rect 52674 17778 52706 18014
rect 52942 17778 53026 18014
rect 53262 17778 53294 18014
rect 52674 -4186 53294 17778
rect 52674 -4422 52706 -4186
rect 52942 -4422 53026 -4186
rect 53262 -4422 53294 -4186
rect 52674 -4506 53294 -4422
rect 52674 -4742 52706 -4506
rect 52942 -4742 53026 -4506
rect 53262 -4742 53294 -4506
rect 52674 -7654 53294 -4742
rect 56394 22054 57014 49367
rect 56394 21818 56426 22054
rect 56662 21818 56746 22054
rect 56982 21818 57014 22054
rect 56394 21734 57014 21818
rect 56394 21498 56426 21734
rect 56662 21498 56746 21734
rect 56982 21498 57014 21734
rect 56394 -5146 57014 21498
rect 56394 -5382 56426 -5146
rect 56662 -5382 56746 -5146
rect 56982 -5382 57014 -5146
rect 56394 -5466 57014 -5382
rect 56394 -5702 56426 -5466
rect 56662 -5702 56746 -5466
rect 56982 -5702 57014 -5466
rect 56394 -7654 57014 -5702
rect 60114 25774 60734 49367
rect 60114 25538 60146 25774
rect 60382 25538 60466 25774
rect 60702 25538 60734 25774
rect 60114 25454 60734 25538
rect 60114 25218 60146 25454
rect 60382 25218 60466 25454
rect 60702 25218 60734 25454
rect 60114 -6106 60734 25218
rect 60114 -6342 60146 -6106
rect 60382 -6342 60466 -6106
rect 60702 -6342 60734 -6106
rect 60114 -6426 60734 -6342
rect 60114 -6662 60146 -6426
rect 60382 -6662 60466 -6426
rect 60702 -6662 60734 -6426
rect 60114 -7654 60734 -6662
rect 63834 29494 64454 49367
rect 63834 29258 63866 29494
rect 64102 29258 64186 29494
rect 64422 29258 64454 29494
rect 63834 29174 64454 29258
rect 63834 28938 63866 29174
rect 64102 28938 64186 29174
rect 64422 28938 64454 29174
rect 63834 -7066 64454 28938
rect 63834 -7302 63866 -7066
rect 64102 -7302 64186 -7066
rect 64422 -7302 64454 -7066
rect 63834 -7386 64454 -7302
rect 63834 -7622 63866 -7386
rect 64102 -7622 64186 -7386
rect 64422 -7622 64454 -7386
rect 63834 -7654 64454 -7622
rect 73794 39454 74414 49367
rect 73794 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 74414 39454
rect 73794 39134 74414 39218
rect 73794 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 74414 39134
rect 73794 3454 74414 38898
rect 73794 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 74414 3454
rect 73794 3134 74414 3218
rect 73794 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 74414 3134
rect 73794 -346 74414 2898
rect 73794 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 74414 -346
rect 73794 -666 74414 -582
rect 73794 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 74414 -666
rect 73794 -7654 74414 -902
rect 77514 43174 78134 49367
rect 77514 42938 77546 43174
rect 77782 42938 77866 43174
rect 78102 42938 78134 43174
rect 77514 42854 78134 42938
rect 77514 42618 77546 42854
rect 77782 42618 77866 42854
rect 78102 42618 78134 42854
rect 77514 7174 78134 42618
rect 77514 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 78134 7174
rect 77514 6854 78134 6938
rect 77514 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 78134 6854
rect 77514 -1306 78134 6618
rect 77514 -1542 77546 -1306
rect 77782 -1542 77866 -1306
rect 78102 -1542 78134 -1306
rect 77514 -1626 78134 -1542
rect 77514 -1862 77546 -1626
rect 77782 -1862 77866 -1626
rect 78102 -1862 78134 -1626
rect 77514 -7654 78134 -1862
rect 81234 46894 81854 49367
rect 81234 46658 81266 46894
rect 81502 46658 81586 46894
rect 81822 46658 81854 46894
rect 81234 46574 81854 46658
rect 81234 46338 81266 46574
rect 81502 46338 81586 46574
rect 81822 46338 81854 46574
rect 81234 10894 81854 46338
rect 81234 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 81854 10894
rect 81234 10574 81854 10658
rect 81234 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 81854 10574
rect 81234 -2266 81854 10338
rect 81234 -2502 81266 -2266
rect 81502 -2502 81586 -2266
rect 81822 -2502 81854 -2266
rect 81234 -2586 81854 -2502
rect 81234 -2822 81266 -2586
rect 81502 -2822 81586 -2586
rect 81822 -2822 81854 -2586
rect 81234 -7654 81854 -2822
rect 84954 14614 85574 49367
rect 84954 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 85574 14614
rect 84954 14294 85574 14378
rect 84954 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 85574 14294
rect 84954 -3226 85574 14058
rect 84954 -3462 84986 -3226
rect 85222 -3462 85306 -3226
rect 85542 -3462 85574 -3226
rect 84954 -3546 85574 -3462
rect 84954 -3782 84986 -3546
rect 85222 -3782 85306 -3546
rect 85542 -3782 85574 -3546
rect 84954 -7654 85574 -3782
rect 88674 18334 89294 49367
rect 88674 18098 88706 18334
rect 88942 18098 89026 18334
rect 89262 18098 89294 18334
rect 88674 18014 89294 18098
rect 88674 17778 88706 18014
rect 88942 17778 89026 18014
rect 89262 17778 89294 18014
rect 88674 -4186 89294 17778
rect 88674 -4422 88706 -4186
rect 88942 -4422 89026 -4186
rect 89262 -4422 89294 -4186
rect 88674 -4506 89294 -4422
rect 88674 -4742 88706 -4506
rect 88942 -4742 89026 -4506
rect 89262 -4742 89294 -4506
rect 88674 -7654 89294 -4742
rect 92394 22054 93014 49367
rect 92394 21818 92426 22054
rect 92662 21818 92746 22054
rect 92982 21818 93014 22054
rect 92394 21734 93014 21818
rect 92394 21498 92426 21734
rect 92662 21498 92746 21734
rect 92982 21498 93014 21734
rect 92394 -5146 93014 21498
rect 92394 -5382 92426 -5146
rect 92662 -5382 92746 -5146
rect 92982 -5382 93014 -5146
rect 92394 -5466 93014 -5382
rect 92394 -5702 92426 -5466
rect 92662 -5702 92746 -5466
rect 92982 -5702 93014 -5466
rect 92394 -7654 93014 -5702
rect 96114 25774 96734 49367
rect 96114 25538 96146 25774
rect 96382 25538 96466 25774
rect 96702 25538 96734 25774
rect 96114 25454 96734 25538
rect 96114 25218 96146 25454
rect 96382 25218 96466 25454
rect 96702 25218 96734 25454
rect 96114 -6106 96734 25218
rect 96114 -6342 96146 -6106
rect 96382 -6342 96466 -6106
rect 96702 -6342 96734 -6106
rect 96114 -6426 96734 -6342
rect 96114 -6662 96146 -6426
rect 96382 -6662 96466 -6426
rect 96702 -6662 96734 -6426
rect 96114 -7654 96734 -6662
rect 99834 29494 100454 49367
rect 99834 29258 99866 29494
rect 100102 29258 100186 29494
rect 100422 29258 100454 29494
rect 99834 29174 100454 29258
rect 99834 28938 99866 29174
rect 100102 28938 100186 29174
rect 100422 28938 100454 29174
rect 99834 -7066 100454 28938
rect 99834 -7302 99866 -7066
rect 100102 -7302 100186 -7066
rect 100422 -7302 100454 -7066
rect 99834 -7386 100454 -7302
rect 99834 -7622 99866 -7386
rect 100102 -7622 100186 -7386
rect 100422 -7622 100454 -7386
rect 99834 -7654 100454 -7622
rect 109794 39454 110414 49367
rect 109794 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 110414 39454
rect 109794 39134 110414 39218
rect 109794 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 110414 39134
rect 109794 3454 110414 38898
rect 109794 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 110414 3454
rect 109794 3134 110414 3218
rect 109794 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 110414 3134
rect 109794 -346 110414 2898
rect 109794 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 110414 -346
rect 109794 -666 110414 -582
rect 109794 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 110414 -666
rect 109794 -7654 110414 -902
rect 113514 43174 114134 49367
rect 113514 42938 113546 43174
rect 113782 42938 113866 43174
rect 114102 42938 114134 43174
rect 113514 42854 114134 42938
rect 113514 42618 113546 42854
rect 113782 42618 113866 42854
rect 114102 42618 114134 42854
rect 113514 7174 114134 42618
rect 113514 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 114134 7174
rect 113514 6854 114134 6938
rect 113514 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 114134 6854
rect 113514 -1306 114134 6618
rect 113514 -1542 113546 -1306
rect 113782 -1542 113866 -1306
rect 114102 -1542 114134 -1306
rect 113514 -1626 114134 -1542
rect 113514 -1862 113546 -1626
rect 113782 -1862 113866 -1626
rect 114102 -1862 114134 -1626
rect 113514 -7654 114134 -1862
rect 117234 46894 117854 49367
rect 117234 46658 117266 46894
rect 117502 46658 117586 46894
rect 117822 46658 117854 46894
rect 117234 46574 117854 46658
rect 117234 46338 117266 46574
rect 117502 46338 117586 46574
rect 117822 46338 117854 46574
rect 117234 10894 117854 46338
rect 117234 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 117854 10894
rect 117234 10574 117854 10658
rect 117234 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 117854 10574
rect 117234 -2266 117854 10338
rect 117234 -2502 117266 -2266
rect 117502 -2502 117586 -2266
rect 117822 -2502 117854 -2266
rect 117234 -2586 117854 -2502
rect 117234 -2822 117266 -2586
rect 117502 -2822 117586 -2586
rect 117822 -2822 117854 -2586
rect 117234 -7654 117854 -2822
rect 120954 14614 121574 49367
rect 120954 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 121574 14614
rect 120954 14294 121574 14378
rect 120954 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 121574 14294
rect 120954 -3226 121574 14058
rect 120954 -3462 120986 -3226
rect 121222 -3462 121306 -3226
rect 121542 -3462 121574 -3226
rect 120954 -3546 121574 -3462
rect 120954 -3782 120986 -3546
rect 121222 -3782 121306 -3546
rect 121542 -3782 121574 -3546
rect 120954 -7654 121574 -3782
rect 124674 18334 125294 49367
rect 124674 18098 124706 18334
rect 124942 18098 125026 18334
rect 125262 18098 125294 18334
rect 124674 18014 125294 18098
rect 124674 17778 124706 18014
rect 124942 17778 125026 18014
rect 125262 17778 125294 18014
rect 124674 -4186 125294 17778
rect 124674 -4422 124706 -4186
rect 124942 -4422 125026 -4186
rect 125262 -4422 125294 -4186
rect 124674 -4506 125294 -4422
rect 124674 -4742 124706 -4506
rect 124942 -4742 125026 -4506
rect 125262 -4742 125294 -4506
rect 124674 -7654 125294 -4742
rect 128394 22054 129014 49367
rect 128394 21818 128426 22054
rect 128662 21818 128746 22054
rect 128982 21818 129014 22054
rect 128394 21734 129014 21818
rect 128394 21498 128426 21734
rect 128662 21498 128746 21734
rect 128982 21498 129014 21734
rect 128394 -5146 129014 21498
rect 128394 -5382 128426 -5146
rect 128662 -5382 128746 -5146
rect 128982 -5382 129014 -5146
rect 128394 -5466 129014 -5382
rect 128394 -5702 128426 -5466
rect 128662 -5702 128746 -5466
rect 128982 -5702 129014 -5466
rect 128394 -7654 129014 -5702
rect 132114 25774 132734 49367
rect 132114 25538 132146 25774
rect 132382 25538 132466 25774
rect 132702 25538 132734 25774
rect 132114 25454 132734 25538
rect 132114 25218 132146 25454
rect 132382 25218 132466 25454
rect 132702 25218 132734 25454
rect 132114 -6106 132734 25218
rect 132114 -6342 132146 -6106
rect 132382 -6342 132466 -6106
rect 132702 -6342 132734 -6106
rect 132114 -6426 132734 -6342
rect 132114 -6662 132146 -6426
rect 132382 -6662 132466 -6426
rect 132702 -6662 132734 -6426
rect 132114 -7654 132734 -6662
rect 135834 29494 136454 49367
rect 135834 29258 135866 29494
rect 136102 29258 136186 29494
rect 136422 29258 136454 29494
rect 135834 29174 136454 29258
rect 135834 28938 135866 29174
rect 136102 28938 136186 29174
rect 136422 28938 136454 29174
rect 135834 -7066 136454 28938
rect 135834 -7302 135866 -7066
rect 136102 -7302 136186 -7066
rect 136422 -7302 136454 -7066
rect 135834 -7386 136454 -7302
rect 135834 -7622 135866 -7386
rect 136102 -7622 136186 -7386
rect 136422 -7622 136454 -7386
rect 135834 -7654 136454 -7622
rect 145794 39454 146414 49367
rect 145794 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 146414 39454
rect 145794 39134 146414 39218
rect 145794 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 146414 39134
rect 145794 3454 146414 38898
rect 145794 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 146414 3454
rect 145794 3134 146414 3218
rect 145794 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 146414 3134
rect 145794 -346 146414 2898
rect 145794 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 146414 -346
rect 145794 -666 146414 -582
rect 145794 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 146414 -666
rect 145794 -7654 146414 -902
rect 149514 43174 150134 49367
rect 149514 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 150134 43174
rect 149514 42854 150134 42938
rect 149514 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 150134 42854
rect 149514 7174 150134 42618
rect 149514 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 150134 7174
rect 149514 6854 150134 6938
rect 149514 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 150134 6854
rect 149514 -1306 150134 6618
rect 149514 -1542 149546 -1306
rect 149782 -1542 149866 -1306
rect 150102 -1542 150134 -1306
rect 149514 -1626 150134 -1542
rect 149514 -1862 149546 -1626
rect 149782 -1862 149866 -1626
rect 150102 -1862 150134 -1626
rect 149514 -7654 150134 -1862
rect 153234 46894 153854 49367
rect 153234 46658 153266 46894
rect 153502 46658 153586 46894
rect 153822 46658 153854 46894
rect 153234 46574 153854 46658
rect 153234 46338 153266 46574
rect 153502 46338 153586 46574
rect 153822 46338 153854 46574
rect 153234 10894 153854 46338
rect 153234 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 153854 10894
rect 153234 10574 153854 10658
rect 153234 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 153854 10574
rect 153234 -2266 153854 10338
rect 153234 -2502 153266 -2266
rect 153502 -2502 153586 -2266
rect 153822 -2502 153854 -2266
rect 153234 -2586 153854 -2502
rect 153234 -2822 153266 -2586
rect 153502 -2822 153586 -2586
rect 153822 -2822 153854 -2586
rect 153234 -7654 153854 -2822
rect 156954 14614 157574 49367
rect 156954 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 157574 14614
rect 156954 14294 157574 14378
rect 156954 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 157574 14294
rect 156954 -3226 157574 14058
rect 156954 -3462 156986 -3226
rect 157222 -3462 157306 -3226
rect 157542 -3462 157574 -3226
rect 156954 -3546 157574 -3462
rect 156954 -3782 156986 -3546
rect 157222 -3782 157306 -3546
rect 157542 -3782 157574 -3546
rect 156954 -7654 157574 -3782
rect 160674 18334 161294 49367
rect 160674 18098 160706 18334
rect 160942 18098 161026 18334
rect 161262 18098 161294 18334
rect 160674 18014 161294 18098
rect 160674 17778 160706 18014
rect 160942 17778 161026 18014
rect 161262 17778 161294 18014
rect 160674 -4186 161294 17778
rect 160674 -4422 160706 -4186
rect 160942 -4422 161026 -4186
rect 161262 -4422 161294 -4186
rect 160674 -4506 161294 -4422
rect 160674 -4742 160706 -4506
rect 160942 -4742 161026 -4506
rect 161262 -4742 161294 -4506
rect 160674 -7654 161294 -4742
rect 164394 22054 165014 49367
rect 164394 21818 164426 22054
rect 164662 21818 164746 22054
rect 164982 21818 165014 22054
rect 164394 21734 165014 21818
rect 164394 21498 164426 21734
rect 164662 21498 164746 21734
rect 164982 21498 165014 21734
rect 164394 -5146 165014 21498
rect 164394 -5382 164426 -5146
rect 164662 -5382 164746 -5146
rect 164982 -5382 165014 -5146
rect 164394 -5466 165014 -5382
rect 164394 -5702 164426 -5466
rect 164662 -5702 164746 -5466
rect 164982 -5702 165014 -5466
rect 164394 -7654 165014 -5702
rect 168114 25774 168734 49367
rect 168114 25538 168146 25774
rect 168382 25538 168466 25774
rect 168702 25538 168734 25774
rect 168114 25454 168734 25538
rect 168114 25218 168146 25454
rect 168382 25218 168466 25454
rect 168702 25218 168734 25454
rect 168114 -6106 168734 25218
rect 168114 -6342 168146 -6106
rect 168382 -6342 168466 -6106
rect 168702 -6342 168734 -6106
rect 168114 -6426 168734 -6342
rect 168114 -6662 168146 -6426
rect 168382 -6662 168466 -6426
rect 168702 -6662 168734 -6426
rect 168114 -7654 168734 -6662
rect 171834 29494 172454 49367
rect 171834 29258 171866 29494
rect 172102 29258 172186 29494
rect 172422 29258 172454 29494
rect 171834 29174 172454 29258
rect 171834 28938 171866 29174
rect 172102 28938 172186 29174
rect 172422 28938 172454 29174
rect 171834 -7066 172454 28938
rect 171834 -7302 171866 -7066
rect 172102 -7302 172186 -7066
rect 172422 -7302 172454 -7066
rect 171834 -7386 172454 -7302
rect 171834 -7622 171866 -7386
rect 172102 -7622 172186 -7386
rect 172422 -7622 172454 -7386
rect 171834 -7654 172454 -7622
rect 181794 39454 182414 49367
rect 181794 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 182414 39454
rect 181794 39134 182414 39218
rect 181794 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 182414 39134
rect 181794 3454 182414 38898
rect 181794 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 182414 3454
rect 181794 3134 182414 3218
rect 181794 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 182414 3134
rect 181794 -346 182414 2898
rect 181794 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 182414 -346
rect 181794 -666 182414 -582
rect 181794 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 182414 -666
rect 181794 -7654 182414 -902
rect 185514 43174 186134 49367
rect 185514 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 186134 43174
rect 185514 42854 186134 42938
rect 185514 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 186134 42854
rect 185514 7174 186134 42618
rect 185514 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 186134 7174
rect 185514 6854 186134 6938
rect 185514 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 186134 6854
rect 185514 -1306 186134 6618
rect 185514 -1542 185546 -1306
rect 185782 -1542 185866 -1306
rect 186102 -1542 186134 -1306
rect 185514 -1626 186134 -1542
rect 185514 -1862 185546 -1626
rect 185782 -1862 185866 -1626
rect 186102 -1862 186134 -1626
rect 185514 -7654 186134 -1862
rect 189234 46894 189854 49367
rect 189234 46658 189266 46894
rect 189502 46658 189586 46894
rect 189822 46658 189854 46894
rect 189234 46574 189854 46658
rect 189234 46338 189266 46574
rect 189502 46338 189586 46574
rect 189822 46338 189854 46574
rect 189234 10894 189854 46338
rect 189234 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 189854 10894
rect 189234 10574 189854 10658
rect 189234 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 189854 10574
rect 189234 -2266 189854 10338
rect 189234 -2502 189266 -2266
rect 189502 -2502 189586 -2266
rect 189822 -2502 189854 -2266
rect 189234 -2586 189854 -2502
rect 189234 -2822 189266 -2586
rect 189502 -2822 189586 -2586
rect 189822 -2822 189854 -2586
rect 189234 -7654 189854 -2822
rect 192954 14614 193574 45068
rect 192954 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 193574 14614
rect 192954 14294 193574 14378
rect 192954 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 193574 14294
rect 192954 -3226 193574 14058
rect 192954 -3462 192986 -3226
rect 193222 -3462 193306 -3226
rect 193542 -3462 193574 -3226
rect 192954 -3546 193574 -3462
rect 192954 -3782 192986 -3546
rect 193222 -3782 193306 -3546
rect 193542 -3782 193574 -3546
rect 192954 -7654 193574 -3782
rect 196674 18334 197294 49367
rect 196674 18098 196706 18334
rect 196942 18098 197026 18334
rect 197262 18098 197294 18334
rect 196674 18014 197294 18098
rect 196674 17778 196706 18014
rect 196942 17778 197026 18014
rect 197262 17778 197294 18014
rect 196674 -4186 197294 17778
rect 196674 -4422 196706 -4186
rect 196942 -4422 197026 -4186
rect 197262 -4422 197294 -4186
rect 196674 -4506 197294 -4422
rect 196674 -4742 196706 -4506
rect 196942 -4742 197026 -4506
rect 197262 -4742 197294 -4506
rect 196674 -7654 197294 -4742
rect 200394 22054 201014 49367
rect 200394 21818 200426 22054
rect 200662 21818 200746 22054
rect 200982 21818 201014 22054
rect 200394 21734 201014 21818
rect 200394 21498 200426 21734
rect 200662 21498 200746 21734
rect 200982 21498 201014 21734
rect 200394 -5146 201014 21498
rect 200394 -5382 200426 -5146
rect 200662 -5382 200746 -5146
rect 200982 -5382 201014 -5146
rect 200394 -5466 201014 -5382
rect 200394 -5702 200426 -5466
rect 200662 -5702 200746 -5466
rect 200982 -5702 201014 -5466
rect 200394 -7654 201014 -5702
rect 204114 25774 204734 49367
rect 204114 25538 204146 25774
rect 204382 25538 204466 25774
rect 204702 25538 204734 25774
rect 204114 25454 204734 25538
rect 204114 25218 204146 25454
rect 204382 25218 204466 25454
rect 204702 25218 204734 25454
rect 204114 -6106 204734 25218
rect 204114 -6342 204146 -6106
rect 204382 -6342 204466 -6106
rect 204702 -6342 204734 -6106
rect 204114 -6426 204734 -6342
rect 204114 -6662 204146 -6426
rect 204382 -6662 204466 -6426
rect 204702 -6662 204734 -6426
rect 204114 -7654 204734 -6662
rect 207834 29494 208454 49367
rect 207834 29258 207866 29494
rect 208102 29258 208186 29494
rect 208422 29258 208454 29494
rect 207834 29174 208454 29258
rect 207834 28938 207866 29174
rect 208102 28938 208186 29174
rect 208422 28938 208454 29174
rect 207834 -7066 208454 28938
rect 207834 -7302 207866 -7066
rect 208102 -7302 208186 -7066
rect 208422 -7302 208454 -7066
rect 207834 -7386 208454 -7302
rect 207834 -7622 207866 -7386
rect 208102 -7622 208186 -7386
rect 208422 -7622 208454 -7386
rect 207834 -7654 208454 -7622
rect 217794 39454 218414 49367
rect 217794 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 218414 39454
rect 217794 39134 218414 39218
rect 217794 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 218414 39134
rect 217794 3454 218414 38898
rect 217794 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 218414 3454
rect 217794 3134 218414 3218
rect 217794 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 218414 3134
rect 217794 -346 218414 2898
rect 217794 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 218414 -346
rect 217794 -666 218414 -582
rect 217794 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 218414 -666
rect 217794 -7654 218414 -902
rect 221514 43174 222134 49367
rect 221514 42938 221546 43174
rect 221782 42938 221866 43174
rect 222102 42938 222134 43174
rect 221514 42854 222134 42938
rect 221514 42618 221546 42854
rect 221782 42618 221866 42854
rect 222102 42618 222134 42854
rect 221514 7174 222134 42618
rect 221514 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 222134 7174
rect 221514 6854 222134 6938
rect 221514 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 222134 6854
rect 221514 -1306 222134 6618
rect 221514 -1542 221546 -1306
rect 221782 -1542 221866 -1306
rect 222102 -1542 222134 -1306
rect 221514 -1626 222134 -1542
rect 221514 -1862 221546 -1626
rect 221782 -1862 221866 -1626
rect 222102 -1862 222134 -1626
rect 221514 -7654 222134 -1862
rect 225234 46894 225854 49367
rect 225234 46658 225266 46894
rect 225502 46658 225586 46894
rect 225822 46658 225854 46894
rect 225234 46574 225854 46658
rect 225234 46338 225266 46574
rect 225502 46338 225586 46574
rect 225822 46338 225854 46574
rect 225234 10894 225854 46338
rect 225234 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 225854 10894
rect 225234 10574 225854 10658
rect 225234 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 225854 10574
rect 225234 -2266 225854 10338
rect 225234 -2502 225266 -2266
rect 225502 -2502 225586 -2266
rect 225822 -2502 225854 -2266
rect 225234 -2586 225854 -2502
rect 225234 -2822 225266 -2586
rect 225502 -2822 225586 -2586
rect 225822 -2822 225854 -2586
rect 225234 -7654 225854 -2822
rect 228954 14614 229574 49367
rect 228954 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 229574 14614
rect 228954 14294 229574 14378
rect 228954 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 229574 14294
rect 228954 -3226 229574 14058
rect 228954 -3462 228986 -3226
rect 229222 -3462 229306 -3226
rect 229542 -3462 229574 -3226
rect 228954 -3546 229574 -3462
rect 228954 -3782 228986 -3546
rect 229222 -3782 229306 -3546
rect 229542 -3782 229574 -3546
rect 228954 -7654 229574 -3782
rect 232674 18334 233294 49367
rect 232674 18098 232706 18334
rect 232942 18098 233026 18334
rect 233262 18098 233294 18334
rect 232674 18014 233294 18098
rect 232674 17778 232706 18014
rect 232942 17778 233026 18014
rect 233262 17778 233294 18014
rect 232674 -4186 233294 17778
rect 232674 -4422 232706 -4186
rect 232942 -4422 233026 -4186
rect 233262 -4422 233294 -4186
rect 232674 -4506 233294 -4422
rect 232674 -4742 232706 -4506
rect 232942 -4742 233026 -4506
rect 233262 -4742 233294 -4506
rect 232674 -7654 233294 -4742
rect 236394 22054 237014 49367
rect 236394 21818 236426 22054
rect 236662 21818 236746 22054
rect 236982 21818 237014 22054
rect 236394 21734 237014 21818
rect 236394 21498 236426 21734
rect 236662 21498 236746 21734
rect 236982 21498 237014 21734
rect 236394 -5146 237014 21498
rect 236394 -5382 236426 -5146
rect 236662 -5382 236746 -5146
rect 236982 -5382 237014 -5146
rect 236394 -5466 237014 -5382
rect 236394 -5702 236426 -5466
rect 236662 -5702 236746 -5466
rect 236982 -5702 237014 -5466
rect 236394 -7654 237014 -5702
rect 240114 25774 240734 49367
rect 240114 25538 240146 25774
rect 240382 25538 240466 25774
rect 240702 25538 240734 25774
rect 240114 25454 240734 25538
rect 240114 25218 240146 25454
rect 240382 25218 240466 25454
rect 240702 25218 240734 25454
rect 240114 -6106 240734 25218
rect 240114 -6342 240146 -6106
rect 240382 -6342 240466 -6106
rect 240702 -6342 240734 -6106
rect 240114 -6426 240734 -6342
rect 240114 -6662 240146 -6426
rect 240382 -6662 240466 -6426
rect 240702 -6662 240734 -6426
rect 240114 -7654 240734 -6662
rect 243834 29494 244454 49367
rect 243834 29258 243866 29494
rect 244102 29258 244186 29494
rect 244422 29258 244454 29494
rect 243834 29174 244454 29258
rect 243834 28938 243866 29174
rect 244102 28938 244186 29174
rect 244422 28938 244454 29174
rect 243834 -7066 244454 28938
rect 243834 -7302 243866 -7066
rect 244102 -7302 244186 -7066
rect 244422 -7302 244454 -7066
rect 243834 -7386 244454 -7302
rect 243834 -7622 243866 -7386
rect 244102 -7622 244186 -7386
rect 244422 -7622 244454 -7386
rect 243834 -7654 244454 -7622
rect 253794 39454 254414 49367
rect 253794 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 254414 39454
rect 253794 39134 254414 39218
rect 253794 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 254414 39134
rect 253794 3454 254414 38898
rect 253794 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 254414 3454
rect 253794 3134 254414 3218
rect 253794 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 254414 3134
rect 253794 -346 254414 2898
rect 253794 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 254414 -346
rect 253794 -666 254414 -582
rect 253794 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 254414 -666
rect 253794 -7654 254414 -902
rect 257514 43174 258134 49367
rect 257514 42938 257546 43174
rect 257782 42938 257866 43174
rect 258102 42938 258134 43174
rect 257514 42854 258134 42938
rect 257514 42618 257546 42854
rect 257782 42618 257866 42854
rect 258102 42618 258134 42854
rect 257514 7174 258134 42618
rect 257514 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 258134 7174
rect 257514 6854 258134 6938
rect 257514 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 258134 6854
rect 257514 -1306 258134 6618
rect 257514 -1542 257546 -1306
rect 257782 -1542 257866 -1306
rect 258102 -1542 258134 -1306
rect 257514 -1626 258134 -1542
rect 257514 -1862 257546 -1626
rect 257782 -1862 257866 -1626
rect 258102 -1862 258134 -1626
rect 257514 -7654 258134 -1862
rect 261234 46894 261854 49367
rect 261234 46658 261266 46894
rect 261502 46658 261586 46894
rect 261822 46658 261854 46894
rect 261234 46574 261854 46658
rect 261234 46338 261266 46574
rect 261502 46338 261586 46574
rect 261822 46338 261854 46574
rect 261234 10894 261854 46338
rect 261234 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 261854 10894
rect 261234 10574 261854 10658
rect 261234 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 261854 10574
rect 261234 -2266 261854 10338
rect 261234 -2502 261266 -2266
rect 261502 -2502 261586 -2266
rect 261822 -2502 261854 -2266
rect 261234 -2586 261854 -2502
rect 261234 -2822 261266 -2586
rect 261502 -2822 261586 -2586
rect 261822 -2822 261854 -2586
rect 261234 -7654 261854 -2822
rect 264954 14614 265574 49367
rect 264954 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 265574 14614
rect 264954 14294 265574 14378
rect 264954 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 265574 14294
rect 264954 -3226 265574 14058
rect 264954 -3462 264986 -3226
rect 265222 -3462 265306 -3226
rect 265542 -3462 265574 -3226
rect 264954 -3546 265574 -3462
rect 264954 -3782 264986 -3546
rect 265222 -3782 265306 -3546
rect 265542 -3782 265574 -3546
rect 264954 -7654 265574 -3782
rect 268674 18334 269294 49367
rect 268674 18098 268706 18334
rect 268942 18098 269026 18334
rect 269262 18098 269294 18334
rect 268674 18014 269294 18098
rect 268674 17778 268706 18014
rect 268942 17778 269026 18014
rect 269262 17778 269294 18014
rect 268674 -4186 269294 17778
rect 268674 -4422 268706 -4186
rect 268942 -4422 269026 -4186
rect 269262 -4422 269294 -4186
rect 268674 -4506 269294 -4422
rect 268674 -4742 268706 -4506
rect 268942 -4742 269026 -4506
rect 269262 -4742 269294 -4506
rect 268674 -7654 269294 -4742
rect 272394 22054 273014 49367
rect 272394 21818 272426 22054
rect 272662 21818 272746 22054
rect 272982 21818 273014 22054
rect 272394 21734 273014 21818
rect 272394 21498 272426 21734
rect 272662 21498 272746 21734
rect 272982 21498 273014 21734
rect 272394 -5146 273014 21498
rect 272394 -5382 272426 -5146
rect 272662 -5382 272746 -5146
rect 272982 -5382 273014 -5146
rect 272394 -5466 273014 -5382
rect 272394 -5702 272426 -5466
rect 272662 -5702 272746 -5466
rect 272982 -5702 273014 -5466
rect 272394 -7654 273014 -5702
rect 276114 25774 276734 49367
rect 276114 25538 276146 25774
rect 276382 25538 276466 25774
rect 276702 25538 276734 25774
rect 276114 25454 276734 25538
rect 276114 25218 276146 25454
rect 276382 25218 276466 25454
rect 276702 25218 276734 25454
rect 276114 -6106 276734 25218
rect 276114 -6342 276146 -6106
rect 276382 -6342 276466 -6106
rect 276702 -6342 276734 -6106
rect 276114 -6426 276734 -6342
rect 276114 -6662 276146 -6426
rect 276382 -6662 276466 -6426
rect 276702 -6662 276734 -6426
rect 276114 -7654 276734 -6662
rect 279834 29494 280454 49367
rect 279834 29258 279866 29494
rect 280102 29258 280186 29494
rect 280422 29258 280454 29494
rect 279834 29174 280454 29258
rect 279834 28938 279866 29174
rect 280102 28938 280186 29174
rect 280422 28938 280454 29174
rect 279834 -7066 280454 28938
rect 279834 -7302 279866 -7066
rect 280102 -7302 280186 -7066
rect 280422 -7302 280454 -7066
rect 279834 -7386 280454 -7302
rect 279834 -7622 279866 -7386
rect 280102 -7622 280186 -7386
rect 280422 -7622 280454 -7386
rect 279834 -7654 280454 -7622
rect 289794 39454 290414 49367
rect 289794 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 290414 39454
rect 289794 39134 290414 39218
rect 289794 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 290414 39134
rect 289794 3454 290414 38898
rect 289794 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 290414 3454
rect 289794 3134 290414 3218
rect 289794 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 290414 3134
rect 289794 -346 290414 2898
rect 289794 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 290414 -346
rect 289794 -666 290414 -582
rect 289794 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 290414 -666
rect 289794 -7654 290414 -902
rect 293514 43174 294134 49367
rect 293514 42938 293546 43174
rect 293782 42938 293866 43174
rect 294102 42938 294134 43174
rect 293514 42854 294134 42938
rect 293514 42618 293546 42854
rect 293782 42618 293866 42854
rect 294102 42618 294134 42854
rect 293514 7174 294134 42618
rect 293514 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 294134 7174
rect 293514 6854 294134 6938
rect 293514 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 294134 6854
rect 293514 -1306 294134 6618
rect 293514 -1542 293546 -1306
rect 293782 -1542 293866 -1306
rect 294102 -1542 294134 -1306
rect 293514 -1626 294134 -1542
rect 293514 -1862 293546 -1626
rect 293782 -1862 293866 -1626
rect 294102 -1862 294134 -1626
rect 293514 -7654 294134 -1862
rect 297234 46894 297854 49367
rect 297234 46658 297266 46894
rect 297502 46658 297586 46894
rect 297822 46658 297854 46894
rect 297234 46574 297854 46658
rect 297234 46338 297266 46574
rect 297502 46338 297586 46574
rect 297822 46338 297854 46574
rect 297234 10894 297854 46338
rect 297234 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 297854 10894
rect 297234 10574 297854 10658
rect 297234 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 297854 10574
rect 297234 -2266 297854 10338
rect 297234 -2502 297266 -2266
rect 297502 -2502 297586 -2266
rect 297822 -2502 297854 -2266
rect 297234 -2586 297854 -2502
rect 297234 -2822 297266 -2586
rect 297502 -2822 297586 -2586
rect 297822 -2822 297854 -2586
rect 297234 -7654 297854 -2822
rect 300954 14614 301574 45068
rect 300954 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 301574 14614
rect 300954 14294 301574 14378
rect 300954 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 301574 14294
rect 300954 -3226 301574 14058
rect 300954 -3462 300986 -3226
rect 301222 -3462 301306 -3226
rect 301542 -3462 301574 -3226
rect 300954 -3546 301574 -3462
rect 300954 -3782 300986 -3546
rect 301222 -3782 301306 -3546
rect 301542 -3782 301574 -3546
rect 300954 -7654 301574 -3782
rect 304674 18334 305294 49367
rect 304674 18098 304706 18334
rect 304942 18098 305026 18334
rect 305262 18098 305294 18334
rect 304674 18014 305294 18098
rect 304674 17778 304706 18014
rect 304942 17778 305026 18014
rect 305262 17778 305294 18014
rect 304674 -4186 305294 17778
rect 304674 -4422 304706 -4186
rect 304942 -4422 305026 -4186
rect 305262 -4422 305294 -4186
rect 304674 -4506 305294 -4422
rect 304674 -4742 304706 -4506
rect 304942 -4742 305026 -4506
rect 305262 -4742 305294 -4506
rect 304674 -7654 305294 -4742
rect 308394 22054 309014 49367
rect 308394 21818 308426 22054
rect 308662 21818 308746 22054
rect 308982 21818 309014 22054
rect 308394 21734 309014 21818
rect 308394 21498 308426 21734
rect 308662 21498 308746 21734
rect 308982 21498 309014 21734
rect 308394 -5146 309014 21498
rect 308394 -5382 308426 -5146
rect 308662 -5382 308746 -5146
rect 308982 -5382 309014 -5146
rect 308394 -5466 309014 -5382
rect 308394 -5702 308426 -5466
rect 308662 -5702 308746 -5466
rect 308982 -5702 309014 -5466
rect 308394 -7654 309014 -5702
rect 312114 25774 312734 49367
rect 312114 25538 312146 25774
rect 312382 25538 312466 25774
rect 312702 25538 312734 25774
rect 312114 25454 312734 25538
rect 312114 25218 312146 25454
rect 312382 25218 312466 25454
rect 312702 25218 312734 25454
rect 312114 -6106 312734 25218
rect 312114 -6342 312146 -6106
rect 312382 -6342 312466 -6106
rect 312702 -6342 312734 -6106
rect 312114 -6426 312734 -6342
rect 312114 -6662 312146 -6426
rect 312382 -6662 312466 -6426
rect 312702 -6662 312734 -6426
rect 312114 -7654 312734 -6662
rect 315834 29494 316454 45068
rect 315834 29258 315866 29494
rect 316102 29258 316186 29494
rect 316422 29258 316454 29494
rect 315834 29174 316454 29258
rect 315834 28938 315866 29174
rect 316102 28938 316186 29174
rect 316422 28938 316454 29174
rect 315834 -7066 316454 28938
rect 315834 -7302 315866 -7066
rect 316102 -7302 316186 -7066
rect 316422 -7302 316454 -7066
rect 315834 -7386 316454 -7302
rect 315834 -7622 315866 -7386
rect 316102 -7622 316186 -7386
rect 316422 -7622 316454 -7386
rect 315834 -7654 316454 -7622
rect 325794 39454 326414 49367
rect 325794 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 326414 39454
rect 325794 39134 326414 39218
rect 325794 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 326414 39134
rect 325794 3454 326414 38898
rect 325794 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 326414 3454
rect 325794 3134 326414 3218
rect 325794 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 326414 3134
rect 325794 -346 326414 2898
rect 325794 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 326414 -346
rect 325794 -666 326414 -582
rect 325794 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 326414 -666
rect 325794 -7654 326414 -902
rect 329514 43174 330134 49367
rect 329514 42938 329546 43174
rect 329782 42938 329866 43174
rect 330102 42938 330134 43174
rect 329514 42854 330134 42938
rect 329514 42618 329546 42854
rect 329782 42618 329866 42854
rect 330102 42618 330134 42854
rect 329514 7174 330134 42618
rect 329514 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 330134 7174
rect 329514 6854 330134 6938
rect 329514 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 330134 6854
rect 329514 -1306 330134 6618
rect 329514 -1542 329546 -1306
rect 329782 -1542 329866 -1306
rect 330102 -1542 330134 -1306
rect 329514 -1626 330134 -1542
rect 329514 -1862 329546 -1626
rect 329782 -1862 329866 -1626
rect 330102 -1862 330134 -1626
rect 329514 -7654 330134 -1862
rect 333234 46894 333854 49367
rect 333234 46658 333266 46894
rect 333502 46658 333586 46894
rect 333822 46658 333854 46894
rect 333234 46574 333854 46658
rect 333234 46338 333266 46574
rect 333502 46338 333586 46574
rect 333822 46338 333854 46574
rect 333234 10894 333854 46338
rect 333234 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 333854 10894
rect 333234 10574 333854 10658
rect 333234 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 333854 10574
rect 333234 -2266 333854 10338
rect 333234 -2502 333266 -2266
rect 333502 -2502 333586 -2266
rect 333822 -2502 333854 -2266
rect 333234 -2586 333854 -2502
rect 333234 -2822 333266 -2586
rect 333502 -2822 333586 -2586
rect 333822 -2822 333854 -2586
rect 333234 -7654 333854 -2822
rect 336954 14614 337574 49367
rect 336954 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 337574 14614
rect 336954 14294 337574 14378
rect 336954 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 337574 14294
rect 336954 -3226 337574 14058
rect 336954 -3462 336986 -3226
rect 337222 -3462 337306 -3226
rect 337542 -3462 337574 -3226
rect 336954 -3546 337574 -3462
rect 336954 -3782 336986 -3546
rect 337222 -3782 337306 -3546
rect 337542 -3782 337574 -3546
rect 336954 -7654 337574 -3782
rect 340674 18334 341294 49367
rect 340674 18098 340706 18334
rect 340942 18098 341026 18334
rect 341262 18098 341294 18334
rect 340674 18014 341294 18098
rect 340674 17778 340706 18014
rect 340942 17778 341026 18014
rect 341262 17778 341294 18014
rect 340674 -4186 341294 17778
rect 340674 -4422 340706 -4186
rect 340942 -4422 341026 -4186
rect 341262 -4422 341294 -4186
rect 340674 -4506 341294 -4422
rect 340674 -4742 340706 -4506
rect 340942 -4742 341026 -4506
rect 341262 -4742 341294 -4506
rect 340674 -7654 341294 -4742
rect 344394 22054 345014 49367
rect 344394 21818 344426 22054
rect 344662 21818 344746 22054
rect 344982 21818 345014 22054
rect 344394 21734 345014 21818
rect 344394 21498 344426 21734
rect 344662 21498 344746 21734
rect 344982 21498 345014 21734
rect 344394 -5146 345014 21498
rect 344394 -5382 344426 -5146
rect 344662 -5382 344746 -5146
rect 344982 -5382 345014 -5146
rect 344394 -5466 345014 -5382
rect 344394 -5702 344426 -5466
rect 344662 -5702 344746 -5466
rect 344982 -5702 345014 -5466
rect 344394 -7654 345014 -5702
rect 348114 25774 348734 49367
rect 348114 25538 348146 25774
rect 348382 25538 348466 25774
rect 348702 25538 348734 25774
rect 348114 25454 348734 25538
rect 348114 25218 348146 25454
rect 348382 25218 348466 25454
rect 348702 25218 348734 25454
rect 348114 -6106 348734 25218
rect 348114 -6342 348146 -6106
rect 348382 -6342 348466 -6106
rect 348702 -6342 348734 -6106
rect 348114 -6426 348734 -6342
rect 348114 -6662 348146 -6426
rect 348382 -6662 348466 -6426
rect 348702 -6662 348734 -6426
rect 348114 -7654 348734 -6662
rect 351834 29494 352454 49367
rect 351834 29258 351866 29494
rect 352102 29258 352186 29494
rect 352422 29258 352454 29494
rect 351834 29174 352454 29258
rect 351834 28938 351866 29174
rect 352102 28938 352186 29174
rect 352422 28938 352454 29174
rect 351834 -7066 352454 28938
rect 351834 -7302 351866 -7066
rect 352102 -7302 352186 -7066
rect 352422 -7302 352454 -7066
rect 351834 -7386 352454 -7302
rect 351834 -7622 351866 -7386
rect 352102 -7622 352186 -7386
rect 352422 -7622 352454 -7386
rect 351834 -7654 352454 -7622
rect 361794 39454 362414 74898
rect 361794 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 362414 39454
rect 361794 39134 362414 39218
rect 361794 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 362414 39134
rect 361794 3454 362414 38898
rect 361794 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 362414 3454
rect 361794 3134 362414 3218
rect 361794 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 362414 3134
rect 361794 -346 362414 2898
rect 361794 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 362414 -346
rect 361794 -666 362414 -582
rect 361794 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 362414 -666
rect 361794 -7654 362414 -902
rect 365514 705798 366134 711590
rect 365514 705562 365546 705798
rect 365782 705562 365866 705798
rect 366102 705562 366134 705798
rect 365514 705478 366134 705562
rect 365514 705242 365546 705478
rect 365782 705242 365866 705478
rect 366102 705242 366134 705478
rect 365514 691174 366134 705242
rect 365514 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 366134 691174
rect 365514 690854 366134 690938
rect 365514 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 366134 690854
rect 365514 655174 366134 690618
rect 365514 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 366134 655174
rect 365514 654854 366134 654938
rect 365514 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 366134 654854
rect 365514 619174 366134 654618
rect 365514 618938 365546 619174
rect 365782 618938 365866 619174
rect 366102 618938 366134 619174
rect 365514 618854 366134 618938
rect 365514 618618 365546 618854
rect 365782 618618 365866 618854
rect 366102 618618 366134 618854
rect 365514 583174 366134 618618
rect 365514 582938 365546 583174
rect 365782 582938 365866 583174
rect 366102 582938 366134 583174
rect 365514 582854 366134 582938
rect 365514 582618 365546 582854
rect 365782 582618 365866 582854
rect 366102 582618 366134 582854
rect 365514 547174 366134 582618
rect 365514 546938 365546 547174
rect 365782 546938 365866 547174
rect 366102 546938 366134 547174
rect 365514 546854 366134 546938
rect 365514 546618 365546 546854
rect 365782 546618 365866 546854
rect 366102 546618 366134 546854
rect 365514 511174 366134 546618
rect 365514 510938 365546 511174
rect 365782 510938 365866 511174
rect 366102 510938 366134 511174
rect 365514 510854 366134 510938
rect 365514 510618 365546 510854
rect 365782 510618 365866 510854
rect 366102 510618 366134 510854
rect 365514 475174 366134 510618
rect 365514 474938 365546 475174
rect 365782 474938 365866 475174
rect 366102 474938 366134 475174
rect 365514 474854 366134 474938
rect 365514 474618 365546 474854
rect 365782 474618 365866 474854
rect 366102 474618 366134 474854
rect 365514 439174 366134 474618
rect 365514 438938 365546 439174
rect 365782 438938 365866 439174
rect 366102 438938 366134 439174
rect 365514 438854 366134 438938
rect 365514 438618 365546 438854
rect 365782 438618 365866 438854
rect 366102 438618 366134 438854
rect 365514 403174 366134 438618
rect 365514 402938 365546 403174
rect 365782 402938 365866 403174
rect 366102 402938 366134 403174
rect 365514 402854 366134 402938
rect 365514 402618 365546 402854
rect 365782 402618 365866 402854
rect 366102 402618 366134 402854
rect 365514 367174 366134 402618
rect 365514 366938 365546 367174
rect 365782 366938 365866 367174
rect 366102 366938 366134 367174
rect 365514 366854 366134 366938
rect 365514 366618 365546 366854
rect 365782 366618 365866 366854
rect 366102 366618 366134 366854
rect 365514 331174 366134 366618
rect 365514 330938 365546 331174
rect 365782 330938 365866 331174
rect 366102 330938 366134 331174
rect 365514 330854 366134 330938
rect 365514 330618 365546 330854
rect 365782 330618 365866 330854
rect 366102 330618 366134 330854
rect 365514 295174 366134 330618
rect 365514 294938 365546 295174
rect 365782 294938 365866 295174
rect 366102 294938 366134 295174
rect 365514 294854 366134 294938
rect 365514 294618 365546 294854
rect 365782 294618 365866 294854
rect 366102 294618 366134 294854
rect 365514 259174 366134 294618
rect 365514 258938 365546 259174
rect 365782 258938 365866 259174
rect 366102 258938 366134 259174
rect 365514 258854 366134 258938
rect 365514 258618 365546 258854
rect 365782 258618 365866 258854
rect 366102 258618 366134 258854
rect 365514 223174 366134 258618
rect 365514 222938 365546 223174
rect 365782 222938 365866 223174
rect 366102 222938 366134 223174
rect 365514 222854 366134 222938
rect 365514 222618 365546 222854
rect 365782 222618 365866 222854
rect 366102 222618 366134 222854
rect 365514 187174 366134 222618
rect 365514 186938 365546 187174
rect 365782 186938 365866 187174
rect 366102 186938 366134 187174
rect 365514 186854 366134 186938
rect 365514 186618 365546 186854
rect 365782 186618 365866 186854
rect 366102 186618 366134 186854
rect 365514 151174 366134 186618
rect 365514 150938 365546 151174
rect 365782 150938 365866 151174
rect 366102 150938 366134 151174
rect 365514 150854 366134 150938
rect 365514 150618 365546 150854
rect 365782 150618 365866 150854
rect 366102 150618 366134 150854
rect 365514 115174 366134 150618
rect 365514 114938 365546 115174
rect 365782 114938 365866 115174
rect 366102 114938 366134 115174
rect 365514 114854 366134 114938
rect 365514 114618 365546 114854
rect 365782 114618 365866 114854
rect 366102 114618 366134 114854
rect 365514 79174 366134 114618
rect 365514 78938 365546 79174
rect 365782 78938 365866 79174
rect 366102 78938 366134 79174
rect 365514 78854 366134 78938
rect 365514 78618 365546 78854
rect 365782 78618 365866 78854
rect 366102 78618 366134 78854
rect 365514 43174 366134 78618
rect 365514 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 366134 43174
rect 365514 42854 366134 42938
rect 365514 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 366134 42854
rect 365514 7174 366134 42618
rect 365514 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 366134 7174
rect 365514 6854 366134 6938
rect 365514 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 366134 6854
rect 365514 -1306 366134 6618
rect 365514 -1542 365546 -1306
rect 365782 -1542 365866 -1306
rect 366102 -1542 366134 -1306
rect 365514 -1626 366134 -1542
rect 365514 -1862 365546 -1626
rect 365782 -1862 365866 -1626
rect 366102 -1862 366134 -1626
rect 365514 -7654 366134 -1862
rect 369234 706758 369854 711590
rect 369234 706522 369266 706758
rect 369502 706522 369586 706758
rect 369822 706522 369854 706758
rect 369234 706438 369854 706522
rect 369234 706202 369266 706438
rect 369502 706202 369586 706438
rect 369822 706202 369854 706438
rect 369234 694894 369854 706202
rect 369234 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 369854 694894
rect 369234 694574 369854 694658
rect 369234 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 369854 694574
rect 369234 658894 369854 694338
rect 369234 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 369854 658894
rect 369234 658574 369854 658658
rect 369234 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 369854 658574
rect 369234 622894 369854 658338
rect 369234 622658 369266 622894
rect 369502 622658 369586 622894
rect 369822 622658 369854 622894
rect 369234 622574 369854 622658
rect 369234 622338 369266 622574
rect 369502 622338 369586 622574
rect 369822 622338 369854 622574
rect 369234 586894 369854 622338
rect 369234 586658 369266 586894
rect 369502 586658 369586 586894
rect 369822 586658 369854 586894
rect 369234 586574 369854 586658
rect 369234 586338 369266 586574
rect 369502 586338 369586 586574
rect 369822 586338 369854 586574
rect 369234 550894 369854 586338
rect 369234 550658 369266 550894
rect 369502 550658 369586 550894
rect 369822 550658 369854 550894
rect 369234 550574 369854 550658
rect 369234 550338 369266 550574
rect 369502 550338 369586 550574
rect 369822 550338 369854 550574
rect 369234 514894 369854 550338
rect 369234 514658 369266 514894
rect 369502 514658 369586 514894
rect 369822 514658 369854 514894
rect 369234 514574 369854 514658
rect 369234 514338 369266 514574
rect 369502 514338 369586 514574
rect 369822 514338 369854 514574
rect 369234 478894 369854 514338
rect 369234 478658 369266 478894
rect 369502 478658 369586 478894
rect 369822 478658 369854 478894
rect 369234 478574 369854 478658
rect 369234 478338 369266 478574
rect 369502 478338 369586 478574
rect 369822 478338 369854 478574
rect 369234 442894 369854 478338
rect 369234 442658 369266 442894
rect 369502 442658 369586 442894
rect 369822 442658 369854 442894
rect 369234 442574 369854 442658
rect 369234 442338 369266 442574
rect 369502 442338 369586 442574
rect 369822 442338 369854 442574
rect 369234 406894 369854 442338
rect 369234 406658 369266 406894
rect 369502 406658 369586 406894
rect 369822 406658 369854 406894
rect 369234 406574 369854 406658
rect 369234 406338 369266 406574
rect 369502 406338 369586 406574
rect 369822 406338 369854 406574
rect 369234 370894 369854 406338
rect 369234 370658 369266 370894
rect 369502 370658 369586 370894
rect 369822 370658 369854 370894
rect 369234 370574 369854 370658
rect 369234 370338 369266 370574
rect 369502 370338 369586 370574
rect 369822 370338 369854 370574
rect 369234 334894 369854 370338
rect 369234 334658 369266 334894
rect 369502 334658 369586 334894
rect 369822 334658 369854 334894
rect 369234 334574 369854 334658
rect 369234 334338 369266 334574
rect 369502 334338 369586 334574
rect 369822 334338 369854 334574
rect 369234 298894 369854 334338
rect 369234 298658 369266 298894
rect 369502 298658 369586 298894
rect 369822 298658 369854 298894
rect 369234 298574 369854 298658
rect 369234 298338 369266 298574
rect 369502 298338 369586 298574
rect 369822 298338 369854 298574
rect 369234 262894 369854 298338
rect 369234 262658 369266 262894
rect 369502 262658 369586 262894
rect 369822 262658 369854 262894
rect 369234 262574 369854 262658
rect 369234 262338 369266 262574
rect 369502 262338 369586 262574
rect 369822 262338 369854 262574
rect 369234 226894 369854 262338
rect 369234 226658 369266 226894
rect 369502 226658 369586 226894
rect 369822 226658 369854 226894
rect 369234 226574 369854 226658
rect 369234 226338 369266 226574
rect 369502 226338 369586 226574
rect 369822 226338 369854 226574
rect 369234 190894 369854 226338
rect 369234 190658 369266 190894
rect 369502 190658 369586 190894
rect 369822 190658 369854 190894
rect 369234 190574 369854 190658
rect 369234 190338 369266 190574
rect 369502 190338 369586 190574
rect 369822 190338 369854 190574
rect 369234 154894 369854 190338
rect 369234 154658 369266 154894
rect 369502 154658 369586 154894
rect 369822 154658 369854 154894
rect 369234 154574 369854 154658
rect 369234 154338 369266 154574
rect 369502 154338 369586 154574
rect 369822 154338 369854 154574
rect 369234 118894 369854 154338
rect 369234 118658 369266 118894
rect 369502 118658 369586 118894
rect 369822 118658 369854 118894
rect 369234 118574 369854 118658
rect 369234 118338 369266 118574
rect 369502 118338 369586 118574
rect 369822 118338 369854 118574
rect 369234 82894 369854 118338
rect 369234 82658 369266 82894
rect 369502 82658 369586 82894
rect 369822 82658 369854 82894
rect 369234 82574 369854 82658
rect 369234 82338 369266 82574
rect 369502 82338 369586 82574
rect 369822 82338 369854 82574
rect 369234 46894 369854 82338
rect 369234 46658 369266 46894
rect 369502 46658 369586 46894
rect 369822 46658 369854 46894
rect 369234 46574 369854 46658
rect 369234 46338 369266 46574
rect 369502 46338 369586 46574
rect 369822 46338 369854 46574
rect 369234 10894 369854 46338
rect 369234 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 369854 10894
rect 369234 10574 369854 10658
rect 369234 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 369854 10574
rect 369234 -2266 369854 10338
rect 369234 -2502 369266 -2266
rect 369502 -2502 369586 -2266
rect 369822 -2502 369854 -2266
rect 369234 -2586 369854 -2502
rect 369234 -2822 369266 -2586
rect 369502 -2822 369586 -2586
rect 369822 -2822 369854 -2586
rect 369234 -7654 369854 -2822
rect 372954 707718 373574 711590
rect 372954 707482 372986 707718
rect 373222 707482 373306 707718
rect 373542 707482 373574 707718
rect 372954 707398 373574 707482
rect 372954 707162 372986 707398
rect 373222 707162 373306 707398
rect 373542 707162 373574 707398
rect 372954 698614 373574 707162
rect 372954 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 373574 698614
rect 372954 698294 373574 698378
rect 372954 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 373574 698294
rect 372954 662614 373574 698058
rect 372954 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 373574 662614
rect 372954 662294 373574 662378
rect 372954 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 373574 662294
rect 372954 626614 373574 662058
rect 372954 626378 372986 626614
rect 373222 626378 373306 626614
rect 373542 626378 373574 626614
rect 372954 626294 373574 626378
rect 372954 626058 372986 626294
rect 373222 626058 373306 626294
rect 373542 626058 373574 626294
rect 372954 590614 373574 626058
rect 372954 590378 372986 590614
rect 373222 590378 373306 590614
rect 373542 590378 373574 590614
rect 372954 590294 373574 590378
rect 372954 590058 372986 590294
rect 373222 590058 373306 590294
rect 373542 590058 373574 590294
rect 372954 554614 373574 590058
rect 372954 554378 372986 554614
rect 373222 554378 373306 554614
rect 373542 554378 373574 554614
rect 372954 554294 373574 554378
rect 372954 554058 372986 554294
rect 373222 554058 373306 554294
rect 373542 554058 373574 554294
rect 372954 518614 373574 554058
rect 372954 518378 372986 518614
rect 373222 518378 373306 518614
rect 373542 518378 373574 518614
rect 372954 518294 373574 518378
rect 372954 518058 372986 518294
rect 373222 518058 373306 518294
rect 373542 518058 373574 518294
rect 372954 482614 373574 518058
rect 372954 482378 372986 482614
rect 373222 482378 373306 482614
rect 373542 482378 373574 482614
rect 372954 482294 373574 482378
rect 372954 482058 372986 482294
rect 373222 482058 373306 482294
rect 373542 482058 373574 482294
rect 372954 446614 373574 482058
rect 372954 446378 372986 446614
rect 373222 446378 373306 446614
rect 373542 446378 373574 446614
rect 372954 446294 373574 446378
rect 372954 446058 372986 446294
rect 373222 446058 373306 446294
rect 373542 446058 373574 446294
rect 372954 410614 373574 446058
rect 372954 410378 372986 410614
rect 373222 410378 373306 410614
rect 373542 410378 373574 410614
rect 372954 410294 373574 410378
rect 372954 410058 372986 410294
rect 373222 410058 373306 410294
rect 373542 410058 373574 410294
rect 372954 374614 373574 410058
rect 372954 374378 372986 374614
rect 373222 374378 373306 374614
rect 373542 374378 373574 374614
rect 372954 374294 373574 374378
rect 372954 374058 372986 374294
rect 373222 374058 373306 374294
rect 373542 374058 373574 374294
rect 372954 338614 373574 374058
rect 372954 338378 372986 338614
rect 373222 338378 373306 338614
rect 373542 338378 373574 338614
rect 372954 338294 373574 338378
rect 372954 338058 372986 338294
rect 373222 338058 373306 338294
rect 373542 338058 373574 338294
rect 372954 302614 373574 338058
rect 372954 302378 372986 302614
rect 373222 302378 373306 302614
rect 373542 302378 373574 302614
rect 372954 302294 373574 302378
rect 372954 302058 372986 302294
rect 373222 302058 373306 302294
rect 373542 302058 373574 302294
rect 372954 266614 373574 302058
rect 372954 266378 372986 266614
rect 373222 266378 373306 266614
rect 373542 266378 373574 266614
rect 372954 266294 373574 266378
rect 372954 266058 372986 266294
rect 373222 266058 373306 266294
rect 373542 266058 373574 266294
rect 372954 230614 373574 266058
rect 372954 230378 372986 230614
rect 373222 230378 373306 230614
rect 373542 230378 373574 230614
rect 372954 230294 373574 230378
rect 372954 230058 372986 230294
rect 373222 230058 373306 230294
rect 373542 230058 373574 230294
rect 372954 194614 373574 230058
rect 372954 194378 372986 194614
rect 373222 194378 373306 194614
rect 373542 194378 373574 194614
rect 372954 194294 373574 194378
rect 372954 194058 372986 194294
rect 373222 194058 373306 194294
rect 373542 194058 373574 194294
rect 372954 158614 373574 194058
rect 372954 158378 372986 158614
rect 373222 158378 373306 158614
rect 373542 158378 373574 158614
rect 372954 158294 373574 158378
rect 372954 158058 372986 158294
rect 373222 158058 373306 158294
rect 373542 158058 373574 158294
rect 372954 122614 373574 158058
rect 372954 122378 372986 122614
rect 373222 122378 373306 122614
rect 373542 122378 373574 122614
rect 372954 122294 373574 122378
rect 372954 122058 372986 122294
rect 373222 122058 373306 122294
rect 373542 122058 373574 122294
rect 372954 86614 373574 122058
rect 372954 86378 372986 86614
rect 373222 86378 373306 86614
rect 373542 86378 373574 86614
rect 372954 86294 373574 86378
rect 372954 86058 372986 86294
rect 373222 86058 373306 86294
rect 373542 86058 373574 86294
rect 372954 50614 373574 86058
rect 372954 50378 372986 50614
rect 373222 50378 373306 50614
rect 373542 50378 373574 50614
rect 372954 50294 373574 50378
rect 372954 50058 372986 50294
rect 373222 50058 373306 50294
rect 373542 50058 373574 50294
rect 372954 14614 373574 50058
rect 372954 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 373574 14614
rect 372954 14294 373574 14378
rect 372954 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 373574 14294
rect 372954 -3226 373574 14058
rect 372954 -3462 372986 -3226
rect 373222 -3462 373306 -3226
rect 373542 -3462 373574 -3226
rect 372954 -3546 373574 -3462
rect 372954 -3782 372986 -3546
rect 373222 -3782 373306 -3546
rect 373542 -3782 373574 -3546
rect 372954 -7654 373574 -3782
rect 376674 708678 377294 711590
rect 376674 708442 376706 708678
rect 376942 708442 377026 708678
rect 377262 708442 377294 708678
rect 376674 708358 377294 708442
rect 376674 708122 376706 708358
rect 376942 708122 377026 708358
rect 377262 708122 377294 708358
rect 376674 666334 377294 708122
rect 376674 666098 376706 666334
rect 376942 666098 377026 666334
rect 377262 666098 377294 666334
rect 376674 666014 377294 666098
rect 376674 665778 376706 666014
rect 376942 665778 377026 666014
rect 377262 665778 377294 666014
rect 376674 630334 377294 665778
rect 376674 630098 376706 630334
rect 376942 630098 377026 630334
rect 377262 630098 377294 630334
rect 376674 630014 377294 630098
rect 376674 629778 376706 630014
rect 376942 629778 377026 630014
rect 377262 629778 377294 630014
rect 376674 594334 377294 629778
rect 376674 594098 376706 594334
rect 376942 594098 377026 594334
rect 377262 594098 377294 594334
rect 376674 594014 377294 594098
rect 376674 593778 376706 594014
rect 376942 593778 377026 594014
rect 377262 593778 377294 594014
rect 376674 558334 377294 593778
rect 376674 558098 376706 558334
rect 376942 558098 377026 558334
rect 377262 558098 377294 558334
rect 376674 558014 377294 558098
rect 376674 557778 376706 558014
rect 376942 557778 377026 558014
rect 377262 557778 377294 558014
rect 376674 522334 377294 557778
rect 376674 522098 376706 522334
rect 376942 522098 377026 522334
rect 377262 522098 377294 522334
rect 376674 522014 377294 522098
rect 376674 521778 376706 522014
rect 376942 521778 377026 522014
rect 377262 521778 377294 522014
rect 376674 486334 377294 521778
rect 376674 486098 376706 486334
rect 376942 486098 377026 486334
rect 377262 486098 377294 486334
rect 376674 486014 377294 486098
rect 376674 485778 376706 486014
rect 376942 485778 377026 486014
rect 377262 485778 377294 486014
rect 376674 450334 377294 485778
rect 376674 450098 376706 450334
rect 376942 450098 377026 450334
rect 377262 450098 377294 450334
rect 376674 450014 377294 450098
rect 376674 449778 376706 450014
rect 376942 449778 377026 450014
rect 377262 449778 377294 450014
rect 376674 414334 377294 449778
rect 376674 414098 376706 414334
rect 376942 414098 377026 414334
rect 377262 414098 377294 414334
rect 376674 414014 377294 414098
rect 376674 413778 376706 414014
rect 376942 413778 377026 414014
rect 377262 413778 377294 414014
rect 376674 378334 377294 413778
rect 376674 378098 376706 378334
rect 376942 378098 377026 378334
rect 377262 378098 377294 378334
rect 376674 378014 377294 378098
rect 376674 377778 376706 378014
rect 376942 377778 377026 378014
rect 377262 377778 377294 378014
rect 376674 342334 377294 377778
rect 376674 342098 376706 342334
rect 376942 342098 377026 342334
rect 377262 342098 377294 342334
rect 376674 342014 377294 342098
rect 376674 341778 376706 342014
rect 376942 341778 377026 342014
rect 377262 341778 377294 342014
rect 376674 306334 377294 341778
rect 376674 306098 376706 306334
rect 376942 306098 377026 306334
rect 377262 306098 377294 306334
rect 376674 306014 377294 306098
rect 376674 305778 376706 306014
rect 376942 305778 377026 306014
rect 377262 305778 377294 306014
rect 376674 270334 377294 305778
rect 376674 270098 376706 270334
rect 376942 270098 377026 270334
rect 377262 270098 377294 270334
rect 376674 270014 377294 270098
rect 376674 269778 376706 270014
rect 376942 269778 377026 270014
rect 377262 269778 377294 270014
rect 376674 234334 377294 269778
rect 376674 234098 376706 234334
rect 376942 234098 377026 234334
rect 377262 234098 377294 234334
rect 376674 234014 377294 234098
rect 376674 233778 376706 234014
rect 376942 233778 377026 234014
rect 377262 233778 377294 234014
rect 376674 198334 377294 233778
rect 376674 198098 376706 198334
rect 376942 198098 377026 198334
rect 377262 198098 377294 198334
rect 376674 198014 377294 198098
rect 376674 197778 376706 198014
rect 376942 197778 377026 198014
rect 377262 197778 377294 198014
rect 376674 162334 377294 197778
rect 376674 162098 376706 162334
rect 376942 162098 377026 162334
rect 377262 162098 377294 162334
rect 376674 162014 377294 162098
rect 376674 161778 376706 162014
rect 376942 161778 377026 162014
rect 377262 161778 377294 162014
rect 376674 126334 377294 161778
rect 376674 126098 376706 126334
rect 376942 126098 377026 126334
rect 377262 126098 377294 126334
rect 376674 126014 377294 126098
rect 376674 125778 376706 126014
rect 376942 125778 377026 126014
rect 377262 125778 377294 126014
rect 376674 90334 377294 125778
rect 376674 90098 376706 90334
rect 376942 90098 377026 90334
rect 377262 90098 377294 90334
rect 376674 90014 377294 90098
rect 376674 89778 376706 90014
rect 376942 89778 377026 90014
rect 377262 89778 377294 90014
rect 376674 54334 377294 89778
rect 376674 54098 376706 54334
rect 376942 54098 377026 54334
rect 377262 54098 377294 54334
rect 376674 54014 377294 54098
rect 376674 53778 376706 54014
rect 376942 53778 377026 54014
rect 377262 53778 377294 54014
rect 376674 18334 377294 53778
rect 376674 18098 376706 18334
rect 376942 18098 377026 18334
rect 377262 18098 377294 18334
rect 376674 18014 377294 18098
rect 376674 17778 376706 18014
rect 376942 17778 377026 18014
rect 377262 17778 377294 18014
rect 376674 -4186 377294 17778
rect 376674 -4422 376706 -4186
rect 376942 -4422 377026 -4186
rect 377262 -4422 377294 -4186
rect 376674 -4506 377294 -4422
rect 376674 -4742 376706 -4506
rect 376942 -4742 377026 -4506
rect 377262 -4742 377294 -4506
rect 376674 -7654 377294 -4742
rect 380394 709638 381014 711590
rect 380394 709402 380426 709638
rect 380662 709402 380746 709638
rect 380982 709402 381014 709638
rect 380394 709318 381014 709402
rect 380394 709082 380426 709318
rect 380662 709082 380746 709318
rect 380982 709082 381014 709318
rect 380394 670054 381014 709082
rect 380394 669818 380426 670054
rect 380662 669818 380746 670054
rect 380982 669818 381014 670054
rect 380394 669734 381014 669818
rect 380394 669498 380426 669734
rect 380662 669498 380746 669734
rect 380982 669498 381014 669734
rect 380394 634054 381014 669498
rect 380394 633818 380426 634054
rect 380662 633818 380746 634054
rect 380982 633818 381014 634054
rect 380394 633734 381014 633818
rect 380394 633498 380426 633734
rect 380662 633498 380746 633734
rect 380982 633498 381014 633734
rect 380394 598054 381014 633498
rect 380394 597818 380426 598054
rect 380662 597818 380746 598054
rect 380982 597818 381014 598054
rect 380394 597734 381014 597818
rect 380394 597498 380426 597734
rect 380662 597498 380746 597734
rect 380982 597498 381014 597734
rect 380394 562054 381014 597498
rect 380394 561818 380426 562054
rect 380662 561818 380746 562054
rect 380982 561818 381014 562054
rect 380394 561734 381014 561818
rect 380394 561498 380426 561734
rect 380662 561498 380746 561734
rect 380982 561498 381014 561734
rect 380394 526054 381014 561498
rect 380394 525818 380426 526054
rect 380662 525818 380746 526054
rect 380982 525818 381014 526054
rect 380394 525734 381014 525818
rect 380394 525498 380426 525734
rect 380662 525498 380746 525734
rect 380982 525498 381014 525734
rect 380394 490054 381014 525498
rect 380394 489818 380426 490054
rect 380662 489818 380746 490054
rect 380982 489818 381014 490054
rect 380394 489734 381014 489818
rect 380394 489498 380426 489734
rect 380662 489498 380746 489734
rect 380982 489498 381014 489734
rect 380394 454054 381014 489498
rect 380394 453818 380426 454054
rect 380662 453818 380746 454054
rect 380982 453818 381014 454054
rect 380394 453734 381014 453818
rect 380394 453498 380426 453734
rect 380662 453498 380746 453734
rect 380982 453498 381014 453734
rect 380394 418054 381014 453498
rect 380394 417818 380426 418054
rect 380662 417818 380746 418054
rect 380982 417818 381014 418054
rect 380394 417734 381014 417818
rect 380394 417498 380426 417734
rect 380662 417498 380746 417734
rect 380982 417498 381014 417734
rect 380394 382054 381014 417498
rect 380394 381818 380426 382054
rect 380662 381818 380746 382054
rect 380982 381818 381014 382054
rect 380394 381734 381014 381818
rect 380394 381498 380426 381734
rect 380662 381498 380746 381734
rect 380982 381498 381014 381734
rect 380394 346054 381014 381498
rect 380394 345818 380426 346054
rect 380662 345818 380746 346054
rect 380982 345818 381014 346054
rect 380394 345734 381014 345818
rect 380394 345498 380426 345734
rect 380662 345498 380746 345734
rect 380982 345498 381014 345734
rect 380394 310054 381014 345498
rect 380394 309818 380426 310054
rect 380662 309818 380746 310054
rect 380982 309818 381014 310054
rect 380394 309734 381014 309818
rect 380394 309498 380426 309734
rect 380662 309498 380746 309734
rect 380982 309498 381014 309734
rect 380394 274054 381014 309498
rect 380394 273818 380426 274054
rect 380662 273818 380746 274054
rect 380982 273818 381014 274054
rect 380394 273734 381014 273818
rect 380394 273498 380426 273734
rect 380662 273498 380746 273734
rect 380982 273498 381014 273734
rect 380394 238054 381014 273498
rect 380394 237818 380426 238054
rect 380662 237818 380746 238054
rect 380982 237818 381014 238054
rect 380394 237734 381014 237818
rect 380394 237498 380426 237734
rect 380662 237498 380746 237734
rect 380982 237498 381014 237734
rect 380394 202054 381014 237498
rect 380394 201818 380426 202054
rect 380662 201818 380746 202054
rect 380982 201818 381014 202054
rect 380394 201734 381014 201818
rect 380394 201498 380426 201734
rect 380662 201498 380746 201734
rect 380982 201498 381014 201734
rect 380394 166054 381014 201498
rect 380394 165818 380426 166054
rect 380662 165818 380746 166054
rect 380982 165818 381014 166054
rect 380394 165734 381014 165818
rect 380394 165498 380426 165734
rect 380662 165498 380746 165734
rect 380982 165498 381014 165734
rect 380394 130054 381014 165498
rect 380394 129818 380426 130054
rect 380662 129818 380746 130054
rect 380982 129818 381014 130054
rect 380394 129734 381014 129818
rect 380394 129498 380426 129734
rect 380662 129498 380746 129734
rect 380982 129498 381014 129734
rect 380394 94054 381014 129498
rect 380394 93818 380426 94054
rect 380662 93818 380746 94054
rect 380982 93818 381014 94054
rect 380394 93734 381014 93818
rect 380394 93498 380426 93734
rect 380662 93498 380746 93734
rect 380982 93498 381014 93734
rect 380394 58054 381014 93498
rect 380394 57818 380426 58054
rect 380662 57818 380746 58054
rect 380982 57818 381014 58054
rect 380394 57734 381014 57818
rect 380394 57498 380426 57734
rect 380662 57498 380746 57734
rect 380982 57498 381014 57734
rect 380394 22054 381014 57498
rect 380394 21818 380426 22054
rect 380662 21818 380746 22054
rect 380982 21818 381014 22054
rect 380394 21734 381014 21818
rect 380394 21498 380426 21734
rect 380662 21498 380746 21734
rect 380982 21498 381014 21734
rect 380394 -5146 381014 21498
rect 380394 -5382 380426 -5146
rect 380662 -5382 380746 -5146
rect 380982 -5382 381014 -5146
rect 380394 -5466 381014 -5382
rect 380394 -5702 380426 -5466
rect 380662 -5702 380746 -5466
rect 380982 -5702 381014 -5466
rect 380394 -7654 381014 -5702
rect 384114 710598 384734 711590
rect 384114 710362 384146 710598
rect 384382 710362 384466 710598
rect 384702 710362 384734 710598
rect 384114 710278 384734 710362
rect 384114 710042 384146 710278
rect 384382 710042 384466 710278
rect 384702 710042 384734 710278
rect 384114 673774 384734 710042
rect 384114 673538 384146 673774
rect 384382 673538 384466 673774
rect 384702 673538 384734 673774
rect 384114 673454 384734 673538
rect 384114 673218 384146 673454
rect 384382 673218 384466 673454
rect 384702 673218 384734 673454
rect 384114 637774 384734 673218
rect 384114 637538 384146 637774
rect 384382 637538 384466 637774
rect 384702 637538 384734 637774
rect 384114 637454 384734 637538
rect 384114 637218 384146 637454
rect 384382 637218 384466 637454
rect 384702 637218 384734 637454
rect 384114 601774 384734 637218
rect 384114 601538 384146 601774
rect 384382 601538 384466 601774
rect 384702 601538 384734 601774
rect 384114 601454 384734 601538
rect 384114 601218 384146 601454
rect 384382 601218 384466 601454
rect 384702 601218 384734 601454
rect 384114 565774 384734 601218
rect 384114 565538 384146 565774
rect 384382 565538 384466 565774
rect 384702 565538 384734 565774
rect 384114 565454 384734 565538
rect 384114 565218 384146 565454
rect 384382 565218 384466 565454
rect 384702 565218 384734 565454
rect 384114 529774 384734 565218
rect 384114 529538 384146 529774
rect 384382 529538 384466 529774
rect 384702 529538 384734 529774
rect 384114 529454 384734 529538
rect 384114 529218 384146 529454
rect 384382 529218 384466 529454
rect 384702 529218 384734 529454
rect 384114 493774 384734 529218
rect 384114 493538 384146 493774
rect 384382 493538 384466 493774
rect 384702 493538 384734 493774
rect 384114 493454 384734 493538
rect 384114 493218 384146 493454
rect 384382 493218 384466 493454
rect 384702 493218 384734 493454
rect 384114 457774 384734 493218
rect 384114 457538 384146 457774
rect 384382 457538 384466 457774
rect 384702 457538 384734 457774
rect 384114 457454 384734 457538
rect 384114 457218 384146 457454
rect 384382 457218 384466 457454
rect 384702 457218 384734 457454
rect 384114 421774 384734 457218
rect 384114 421538 384146 421774
rect 384382 421538 384466 421774
rect 384702 421538 384734 421774
rect 384114 421454 384734 421538
rect 384114 421218 384146 421454
rect 384382 421218 384466 421454
rect 384702 421218 384734 421454
rect 384114 385774 384734 421218
rect 384114 385538 384146 385774
rect 384382 385538 384466 385774
rect 384702 385538 384734 385774
rect 384114 385454 384734 385538
rect 384114 385218 384146 385454
rect 384382 385218 384466 385454
rect 384702 385218 384734 385454
rect 384114 349774 384734 385218
rect 384114 349538 384146 349774
rect 384382 349538 384466 349774
rect 384702 349538 384734 349774
rect 384114 349454 384734 349538
rect 384114 349218 384146 349454
rect 384382 349218 384466 349454
rect 384702 349218 384734 349454
rect 384114 313774 384734 349218
rect 384114 313538 384146 313774
rect 384382 313538 384466 313774
rect 384702 313538 384734 313774
rect 384114 313454 384734 313538
rect 384114 313218 384146 313454
rect 384382 313218 384466 313454
rect 384702 313218 384734 313454
rect 384114 277774 384734 313218
rect 384114 277538 384146 277774
rect 384382 277538 384466 277774
rect 384702 277538 384734 277774
rect 384114 277454 384734 277538
rect 384114 277218 384146 277454
rect 384382 277218 384466 277454
rect 384702 277218 384734 277454
rect 384114 241774 384734 277218
rect 384114 241538 384146 241774
rect 384382 241538 384466 241774
rect 384702 241538 384734 241774
rect 384114 241454 384734 241538
rect 384114 241218 384146 241454
rect 384382 241218 384466 241454
rect 384702 241218 384734 241454
rect 384114 205774 384734 241218
rect 384114 205538 384146 205774
rect 384382 205538 384466 205774
rect 384702 205538 384734 205774
rect 384114 205454 384734 205538
rect 384114 205218 384146 205454
rect 384382 205218 384466 205454
rect 384702 205218 384734 205454
rect 384114 169774 384734 205218
rect 384114 169538 384146 169774
rect 384382 169538 384466 169774
rect 384702 169538 384734 169774
rect 384114 169454 384734 169538
rect 384114 169218 384146 169454
rect 384382 169218 384466 169454
rect 384702 169218 384734 169454
rect 384114 133774 384734 169218
rect 384114 133538 384146 133774
rect 384382 133538 384466 133774
rect 384702 133538 384734 133774
rect 384114 133454 384734 133538
rect 384114 133218 384146 133454
rect 384382 133218 384466 133454
rect 384702 133218 384734 133454
rect 384114 97774 384734 133218
rect 384114 97538 384146 97774
rect 384382 97538 384466 97774
rect 384702 97538 384734 97774
rect 384114 97454 384734 97538
rect 384114 97218 384146 97454
rect 384382 97218 384466 97454
rect 384702 97218 384734 97454
rect 384114 61774 384734 97218
rect 384114 61538 384146 61774
rect 384382 61538 384466 61774
rect 384702 61538 384734 61774
rect 384114 61454 384734 61538
rect 384114 61218 384146 61454
rect 384382 61218 384466 61454
rect 384702 61218 384734 61454
rect 384114 25774 384734 61218
rect 384114 25538 384146 25774
rect 384382 25538 384466 25774
rect 384702 25538 384734 25774
rect 384114 25454 384734 25538
rect 384114 25218 384146 25454
rect 384382 25218 384466 25454
rect 384702 25218 384734 25454
rect 384114 -6106 384734 25218
rect 384114 -6342 384146 -6106
rect 384382 -6342 384466 -6106
rect 384702 -6342 384734 -6106
rect 384114 -6426 384734 -6342
rect 384114 -6662 384146 -6426
rect 384382 -6662 384466 -6426
rect 384702 -6662 384734 -6426
rect 384114 -7654 384734 -6662
rect 387834 711558 388454 711590
rect 387834 711322 387866 711558
rect 388102 711322 388186 711558
rect 388422 711322 388454 711558
rect 387834 711238 388454 711322
rect 387834 711002 387866 711238
rect 388102 711002 388186 711238
rect 388422 711002 388454 711238
rect 387834 677494 388454 711002
rect 387834 677258 387866 677494
rect 388102 677258 388186 677494
rect 388422 677258 388454 677494
rect 387834 677174 388454 677258
rect 387834 676938 387866 677174
rect 388102 676938 388186 677174
rect 388422 676938 388454 677174
rect 387834 641494 388454 676938
rect 387834 641258 387866 641494
rect 388102 641258 388186 641494
rect 388422 641258 388454 641494
rect 387834 641174 388454 641258
rect 387834 640938 387866 641174
rect 388102 640938 388186 641174
rect 388422 640938 388454 641174
rect 387834 605494 388454 640938
rect 387834 605258 387866 605494
rect 388102 605258 388186 605494
rect 388422 605258 388454 605494
rect 387834 605174 388454 605258
rect 387834 604938 387866 605174
rect 388102 604938 388186 605174
rect 388422 604938 388454 605174
rect 387834 569494 388454 604938
rect 387834 569258 387866 569494
rect 388102 569258 388186 569494
rect 388422 569258 388454 569494
rect 387834 569174 388454 569258
rect 387834 568938 387866 569174
rect 388102 568938 388186 569174
rect 388422 568938 388454 569174
rect 387834 533494 388454 568938
rect 387834 533258 387866 533494
rect 388102 533258 388186 533494
rect 388422 533258 388454 533494
rect 387834 533174 388454 533258
rect 387834 532938 387866 533174
rect 388102 532938 388186 533174
rect 388422 532938 388454 533174
rect 387834 497494 388454 532938
rect 387834 497258 387866 497494
rect 388102 497258 388186 497494
rect 388422 497258 388454 497494
rect 387834 497174 388454 497258
rect 387834 496938 387866 497174
rect 388102 496938 388186 497174
rect 388422 496938 388454 497174
rect 387834 461494 388454 496938
rect 387834 461258 387866 461494
rect 388102 461258 388186 461494
rect 388422 461258 388454 461494
rect 387834 461174 388454 461258
rect 387834 460938 387866 461174
rect 388102 460938 388186 461174
rect 388422 460938 388454 461174
rect 387834 425494 388454 460938
rect 387834 425258 387866 425494
rect 388102 425258 388186 425494
rect 388422 425258 388454 425494
rect 387834 425174 388454 425258
rect 387834 424938 387866 425174
rect 388102 424938 388186 425174
rect 388422 424938 388454 425174
rect 387834 389494 388454 424938
rect 387834 389258 387866 389494
rect 388102 389258 388186 389494
rect 388422 389258 388454 389494
rect 387834 389174 388454 389258
rect 387834 388938 387866 389174
rect 388102 388938 388186 389174
rect 388422 388938 388454 389174
rect 387834 353494 388454 388938
rect 387834 353258 387866 353494
rect 388102 353258 388186 353494
rect 388422 353258 388454 353494
rect 387834 353174 388454 353258
rect 387834 352938 387866 353174
rect 388102 352938 388186 353174
rect 388422 352938 388454 353174
rect 387834 317494 388454 352938
rect 387834 317258 387866 317494
rect 388102 317258 388186 317494
rect 388422 317258 388454 317494
rect 387834 317174 388454 317258
rect 387834 316938 387866 317174
rect 388102 316938 388186 317174
rect 388422 316938 388454 317174
rect 387834 281494 388454 316938
rect 387834 281258 387866 281494
rect 388102 281258 388186 281494
rect 388422 281258 388454 281494
rect 387834 281174 388454 281258
rect 387834 280938 387866 281174
rect 388102 280938 388186 281174
rect 388422 280938 388454 281174
rect 387834 245494 388454 280938
rect 387834 245258 387866 245494
rect 388102 245258 388186 245494
rect 388422 245258 388454 245494
rect 387834 245174 388454 245258
rect 387834 244938 387866 245174
rect 388102 244938 388186 245174
rect 388422 244938 388454 245174
rect 387834 209494 388454 244938
rect 387834 209258 387866 209494
rect 388102 209258 388186 209494
rect 388422 209258 388454 209494
rect 387834 209174 388454 209258
rect 387834 208938 387866 209174
rect 388102 208938 388186 209174
rect 388422 208938 388454 209174
rect 387834 173494 388454 208938
rect 387834 173258 387866 173494
rect 388102 173258 388186 173494
rect 388422 173258 388454 173494
rect 387834 173174 388454 173258
rect 387834 172938 387866 173174
rect 388102 172938 388186 173174
rect 388422 172938 388454 173174
rect 387834 137494 388454 172938
rect 387834 137258 387866 137494
rect 388102 137258 388186 137494
rect 388422 137258 388454 137494
rect 387834 137174 388454 137258
rect 387834 136938 387866 137174
rect 388102 136938 388186 137174
rect 388422 136938 388454 137174
rect 387834 101494 388454 136938
rect 387834 101258 387866 101494
rect 388102 101258 388186 101494
rect 388422 101258 388454 101494
rect 387834 101174 388454 101258
rect 387834 100938 387866 101174
rect 388102 100938 388186 101174
rect 388422 100938 388454 101174
rect 387834 65494 388454 100938
rect 387834 65258 387866 65494
rect 388102 65258 388186 65494
rect 388422 65258 388454 65494
rect 387834 65174 388454 65258
rect 387834 64938 387866 65174
rect 388102 64938 388186 65174
rect 388422 64938 388454 65174
rect 387834 29494 388454 64938
rect 387834 29258 387866 29494
rect 388102 29258 388186 29494
rect 388422 29258 388454 29494
rect 387834 29174 388454 29258
rect 387834 28938 387866 29174
rect 388102 28938 388186 29174
rect 388422 28938 388454 29174
rect 387834 -7066 388454 28938
rect 387834 -7302 387866 -7066
rect 388102 -7302 388186 -7066
rect 388422 -7302 388454 -7066
rect 387834 -7386 388454 -7302
rect 387834 -7622 387866 -7386
rect 388102 -7622 388186 -7386
rect 388422 -7622 388454 -7386
rect 387834 -7654 388454 -7622
rect 397794 704838 398414 711590
rect 397794 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 398414 704838
rect 397794 704518 398414 704602
rect 397794 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 398414 704518
rect 397794 687454 398414 704282
rect 397794 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 398414 687454
rect 397794 687134 398414 687218
rect 397794 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 398414 687134
rect 397794 651454 398414 686898
rect 397794 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 398414 651454
rect 397794 651134 398414 651218
rect 397794 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 398414 651134
rect 397794 615454 398414 650898
rect 397794 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 398414 615454
rect 397794 615134 398414 615218
rect 397794 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 398414 615134
rect 397794 579454 398414 614898
rect 397794 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 398414 579454
rect 397794 579134 398414 579218
rect 397794 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 398414 579134
rect 397794 543454 398414 578898
rect 397794 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 398414 543454
rect 397794 543134 398414 543218
rect 397794 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 398414 543134
rect 397794 507454 398414 542898
rect 397794 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 398414 507454
rect 397794 507134 398414 507218
rect 397794 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 398414 507134
rect 397794 471454 398414 506898
rect 397794 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 398414 471454
rect 397794 471134 398414 471218
rect 397794 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 398414 471134
rect 397794 435454 398414 470898
rect 397794 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 398414 435454
rect 397794 435134 398414 435218
rect 397794 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 398414 435134
rect 397794 399454 398414 434898
rect 397794 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 398414 399454
rect 397794 399134 398414 399218
rect 397794 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 398414 399134
rect 397794 363454 398414 398898
rect 397794 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 398414 363454
rect 397794 363134 398414 363218
rect 397794 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 398414 363134
rect 397794 327454 398414 362898
rect 397794 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 398414 327454
rect 397794 327134 398414 327218
rect 397794 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 398414 327134
rect 397794 291454 398414 326898
rect 397794 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 398414 291454
rect 397794 291134 398414 291218
rect 397794 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 398414 291134
rect 397794 255454 398414 290898
rect 397794 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 398414 255454
rect 397794 255134 398414 255218
rect 397794 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 398414 255134
rect 397794 219454 398414 254898
rect 397794 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 398414 219454
rect 397794 219134 398414 219218
rect 397794 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 398414 219134
rect 397794 183454 398414 218898
rect 397794 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 398414 183454
rect 397794 183134 398414 183218
rect 397794 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 398414 183134
rect 397794 147454 398414 182898
rect 397794 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 398414 147454
rect 397794 147134 398414 147218
rect 397794 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 398414 147134
rect 397794 111454 398414 146898
rect 397794 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 398414 111454
rect 397794 111134 398414 111218
rect 397794 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 398414 111134
rect 397794 75454 398414 110898
rect 397794 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 398414 75454
rect 397794 75134 398414 75218
rect 397794 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 398414 75134
rect 397794 39454 398414 74898
rect 397794 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 398414 39454
rect 397794 39134 398414 39218
rect 397794 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 398414 39134
rect 397794 3454 398414 38898
rect 397794 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 398414 3454
rect 397794 3134 398414 3218
rect 397794 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 398414 3134
rect 397794 -346 398414 2898
rect 397794 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 398414 -346
rect 397794 -666 398414 -582
rect 397794 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 398414 -666
rect 397794 -7654 398414 -902
rect 401514 705798 402134 711590
rect 401514 705562 401546 705798
rect 401782 705562 401866 705798
rect 402102 705562 402134 705798
rect 401514 705478 402134 705562
rect 401514 705242 401546 705478
rect 401782 705242 401866 705478
rect 402102 705242 402134 705478
rect 401514 691174 402134 705242
rect 401514 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 402134 691174
rect 401514 690854 402134 690938
rect 401514 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 402134 690854
rect 401514 655174 402134 690618
rect 401514 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 402134 655174
rect 401514 654854 402134 654938
rect 401514 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 402134 654854
rect 401514 619174 402134 654618
rect 401514 618938 401546 619174
rect 401782 618938 401866 619174
rect 402102 618938 402134 619174
rect 401514 618854 402134 618938
rect 401514 618618 401546 618854
rect 401782 618618 401866 618854
rect 402102 618618 402134 618854
rect 401514 583174 402134 618618
rect 401514 582938 401546 583174
rect 401782 582938 401866 583174
rect 402102 582938 402134 583174
rect 401514 582854 402134 582938
rect 401514 582618 401546 582854
rect 401782 582618 401866 582854
rect 402102 582618 402134 582854
rect 401514 547174 402134 582618
rect 401514 546938 401546 547174
rect 401782 546938 401866 547174
rect 402102 546938 402134 547174
rect 401514 546854 402134 546938
rect 401514 546618 401546 546854
rect 401782 546618 401866 546854
rect 402102 546618 402134 546854
rect 401514 511174 402134 546618
rect 401514 510938 401546 511174
rect 401782 510938 401866 511174
rect 402102 510938 402134 511174
rect 401514 510854 402134 510938
rect 401514 510618 401546 510854
rect 401782 510618 401866 510854
rect 402102 510618 402134 510854
rect 401514 475174 402134 510618
rect 401514 474938 401546 475174
rect 401782 474938 401866 475174
rect 402102 474938 402134 475174
rect 401514 474854 402134 474938
rect 401514 474618 401546 474854
rect 401782 474618 401866 474854
rect 402102 474618 402134 474854
rect 401514 439174 402134 474618
rect 401514 438938 401546 439174
rect 401782 438938 401866 439174
rect 402102 438938 402134 439174
rect 401514 438854 402134 438938
rect 401514 438618 401546 438854
rect 401782 438618 401866 438854
rect 402102 438618 402134 438854
rect 401514 403174 402134 438618
rect 401514 402938 401546 403174
rect 401782 402938 401866 403174
rect 402102 402938 402134 403174
rect 401514 402854 402134 402938
rect 401514 402618 401546 402854
rect 401782 402618 401866 402854
rect 402102 402618 402134 402854
rect 401514 367174 402134 402618
rect 401514 366938 401546 367174
rect 401782 366938 401866 367174
rect 402102 366938 402134 367174
rect 401514 366854 402134 366938
rect 401514 366618 401546 366854
rect 401782 366618 401866 366854
rect 402102 366618 402134 366854
rect 401514 331174 402134 366618
rect 401514 330938 401546 331174
rect 401782 330938 401866 331174
rect 402102 330938 402134 331174
rect 401514 330854 402134 330938
rect 401514 330618 401546 330854
rect 401782 330618 401866 330854
rect 402102 330618 402134 330854
rect 401514 295174 402134 330618
rect 405234 706758 405854 711590
rect 405234 706522 405266 706758
rect 405502 706522 405586 706758
rect 405822 706522 405854 706758
rect 405234 706438 405854 706522
rect 405234 706202 405266 706438
rect 405502 706202 405586 706438
rect 405822 706202 405854 706438
rect 405234 694894 405854 706202
rect 405234 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 405854 694894
rect 405234 694574 405854 694658
rect 405234 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 405854 694574
rect 405234 658894 405854 694338
rect 405234 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 405854 658894
rect 405234 658574 405854 658658
rect 405234 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 405854 658574
rect 405234 622894 405854 658338
rect 405234 622658 405266 622894
rect 405502 622658 405586 622894
rect 405822 622658 405854 622894
rect 405234 622574 405854 622658
rect 405234 622338 405266 622574
rect 405502 622338 405586 622574
rect 405822 622338 405854 622574
rect 405234 586894 405854 622338
rect 405234 586658 405266 586894
rect 405502 586658 405586 586894
rect 405822 586658 405854 586894
rect 405234 586574 405854 586658
rect 405234 586338 405266 586574
rect 405502 586338 405586 586574
rect 405822 586338 405854 586574
rect 405234 550894 405854 586338
rect 405234 550658 405266 550894
rect 405502 550658 405586 550894
rect 405822 550658 405854 550894
rect 405234 550574 405854 550658
rect 405234 550338 405266 550574
rect 405502 550338 405586 550574
rect 405822 550338 405854 550574
rect 405234 514894 405854 550338
rect 405234 514658 405266 514894
rect 405502 514658 405586 514894
rect 405822 514658 405854 514894
rect 405234 514574 405854 514658
rect 405234 514338 405266 514574
rect 405502 514338 405586 514574
rect 405822 514338 405854 514574
rect 405234 478894 405854 514338
rect 405234 478658 405266 478894
rect 405502 478658 405586 478894
rect 405822 478658 405854 478894
rect 405234 478574 405854 478658
rect 405234 478338 405266 478574
rect 405502 478338 405586 478574
rect 405822 478338 405854 478574
rect 405234 442894 405854 478338
rect 405234 442658 405266 442894
rect 405502 442658 405586 442894
rect 405822 442658 405854 442894
rect 405234 442574 405854 442658
rect 405234 442338 405266 442574
rect 405502 442338 405586 442574
rect 405822 442338 405854 442574
rect 405234 406894 405854 442338
rect 405234 406658 405266 406894
rect 405502 406658 405586 406894
rect 405822 406658 405854 406894
rect 405234 406574 405854 406658
rect 405234 406338 405266 406574
rect 405502 406338 405586 406574
rect 405822 406338 405854 406574
rect 405234 370894 405854 406338
rect 405234 370658 405266 370894
rect 405502 370658 405586 370894
rect 405822 370658 405854 370894
rect 405234 370574 405854 370658
rect 405234 370338 405266 370574
rect 405502 370338 405586 370574
rect 405822 370338 405854 370574
rect 405234 334894 405854 370338
rect 405234 334658 405266 334894
rect 405502 334658 405586 334894
rect 405822 334658 405854 334894
rect 405234 334574 405854 334658
rect 405234 334338 405266 334574
rect 405502 334338 405586 334574
rect 405822 334338 405854 334574
rect 404417 327454 404737 327486
rect 404417 327218 404459 327454
rect 404695 327218 404737 327454
rect 404417 327134 404737 327218
rect 404417 326898 404459 327134
rect 404695 326898 404737 327134
rect 404417 326866 404737 326898
rect 401514 294938 401546 295174
rect 401782 294938 401866 295174
rect 402102 294938 402134 295174
rect 401514 294854 402134 294938
rect 401514 294618 401546 294854
rect 401782 294618 401866 294854
rect 402102 294618 402134 294854
rect 401514 259174 402134 294618
rect 401514 258938 401546 259174
rect 401782 258938 401866 259174
rect 402102 258938 402134 259174
rect 401514 258854 402134 258938
rect 401514 258618 401546 258854
rect 401782 258618 401866 258854
rect 402102 258618 402134 258854
rect 401514 223174 402134 258618
rect 401514 222938 401546 223174
rect 401782 222938 401866 223174
rect 402102 222938 402134 223174
rect 401514 222854 402134 222938
rect 401514 222618 401546 222854
rect 401782 222618 401866 222854
rect 402102 222618 402134 222854
rect 401514 187174 402134 222618
rect 401514 186938 401546 187174
rect 401782 186938 401866 187174
rect 402102 186938 402134 187174
rect 401514 186854 402134 186938
rect 401514 186618 401546 186854
rect 401782 186618 401866 186854
rect 402102 186618 402134 186854
rect 401514 151174 402134 186618
rect 401514 150938 401546 151174
rect 401782 150938 401866 151174
rect 402102 150938 402134 151174
rect 401514 150854 402134 150938
rect 401514 150618 401546 150854
rect 401782 150618 401866 150854
rect 402102 150618 402134 150854
rect 401514 115174 402134 150618
rect 401514 114938 401546 115174
rect 401782 114938 401866 115174
rect 402102 114938 402134 115174
rect 401514 114854 402134 114938
rect 401514 114618 401546 114854
rect 401782 114618 401866 114854
rect 402102 114618 402134 114854
rect 401514 79174 402134 114618
rect 401514 78938 401546 79174
rect 401782 78938 401866 79174
rect 402102 78938 402134 79174
rect 401514 78854 402134 78938
rect 401514 78618 401546 78854
rect 401782 78618 401866 78854
rect 402102 78618 402134 78854
rect 401514 43174 402134 78618
rect 401514 42938 401546 43174
rect 401782 42938 401866 43174
rect 402102 42938 402134 43174
rect 401514 42854 402134 42938
rect 401514 42618 401546 42854
rect 401782 42618 401866 42854
rect 402102 42618 402134 42854
rect 401514 7174 402134 42618
rect 401514 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 402134 7174
rect 401514 6854 402134 6938
rect 401514 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 402134 6854
rect 401514 -1306 402134 6618
rect 401514 -1542 401546 -1306
rect 401782 -1542 401866 -1306
rect 402102 -1542 402134 -1306
rect 401514 -1626 402134 -1542
rect 401514 -1862 401546 -1626
rect 401782 -1862 401866 -1626
rect 402102 -1862 402134 -1626
rect 401514 -7654 402134 -1862
rect 405234 298894 405854 334338
rect 408954 707718 409574 711590
rect 408954 707482 408986 707718
rect 409222 707482 409306 707718
rect 409542 707482 409574 707718
rect 408954 707398 409574 707482
rect 408954 707162 408986 707398
rect 409222 707162 409306 707398
rect 409542 707162 409574 707398
rect 408954 698614 409574 707162
rect 408954 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 409574 698614
rect 408954 698294 409574 698378
rect 408954 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 409574 698294
rect 408954 662614 409574 698058
rect 408954 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 409574 662614
rect 408954 662294 409574 662378
rect 408954 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 409574 662294
rect 408954 626614 409574 662058
rect 408954 626378 408986 626614
rect 409222 626378 409306 626614
rect 409542 626378 409574 626614
rect 408954 626294 409574 626378
rect 408954 626058 408986 626294
rect 409222 626058 409306 626294
rect 409542 626058 409574 626294
rect 408954 590614 409574 626058
rect 408954 590378 408986 590614
rect 409222 590378 409306 590614
rect 409542 590378 409574 590614
rect 408954 590294 409574 590378
rect 408954 590058 408986 590294
rect 409222 590058 409306 590294
rect 409542 590058 409574 590294
rect 408954 554614 409574 590058
rect 408954 554378 408986 554614
rect 409222 554378 409306 554614
rect 409542 554378 409574 554614
rect 408954 554294 409574 554378
rect 408954 554058 408986 554294
rect 409222 554058 409306 554294
rect 409542 554058 409574 554294
rect 408954 518614 409574 554058
rect 408954 518378 408986 518614
rect 409222 518378 409306 518614
rect 409542 518378 409574 518614
rect 408954 518294 409574 518378
rect 408954 518058 408986 518294
rect 409222 518058 409306 518294
rect 409542 518058 409574 518294
rect 408954 482614 409574 518058
rect 408954 482378 408986 482614
rect 409222 482378 409306 482614
rect 409542 482378 409574 482614
rect 408954 482294 409574 482378
rect 408954 482058 408986 482294
rect 409222 482058 409306 482294
rect 409542 482058 409574 482294
rect 408954 446614 409574 482058
rect 408954 446378 408986 446614
rect 409222 446378 409306 446614
rect 409542 446378 409574 446614
rect 408954 446294 409574 446378
rect 408954 446058 408986 446294
rect 409222 446058 409306 446294
rect 409542 446058 409574 446294
rect 408954 410614 409574 446058
rect 408954 410378 408986 410614
rect 409222 410378 409306 410614
rect 409542 410378 409574 410614
rect 408954 410294 409574 410378
rect 408954 410058 408986 410294
rect 409222 410058 409306 410294
rect 409542 410058 409574 410294
rect 408954 374614 409574 410058
rect 408954 374378 408986 374614
rect 409222 374378 409306 374614
rect 409542 374378 409574 374614
rect 408954 374294 409574 374378
rect 408954 374058 408986 374294
rect 409222 374058 409306 374294
rect 409542 374058 409574 374294
rect 408954 338614 409574 374058
rect 408954 338378 408986 338614
rect 409222 338378 409306 338614
rect 409542 338378 409574 338614
rect 408954 338294 409574 338378
rect 408954 338058 408986 338294
rect 409222 338058 409306 338294
rect 409542 338058 409574 338294
rect 407890 331174 408210 331206
rect 407890 330938 407932 331174
rect 408168 330938 408210 331174
rect 407890 330854 408210 330938
rect 407890 330618 407932 330854
rect 408168 330618 408210 330854
rect 407890 330586 408210 330618
rect 405234 298658 405266 298894
rect 405502 298658 405586 298894
rect 405822 298658 405854 298894
rect 405234 298574 405854 298658
rect 405234 298338 405266 298574
rect 405502 298338 405586 298574
rect 405822 298338 405854 298574
rect 405234 262894 405854 298338
rect 405234 262658 405266 262894
rect 405502 262658 405586 262894
rect 405822 262658 405854 262894
rect 405234 262574 405854 262658
rect 405234 262338 405266 262574
rect 405502 262338 405586 262574
rect 405822 262338 405854 262574
rect 405234 226894 405854 262338
rect 405234 226658 405266 226894
rect 405502 226658 405586 226894
rect 405822 226658 405854 226894
rect 405234 226574 405854 226658
rect 405234 226338 405266 226574
rect 405502 226338 405586 226574
rect 405822 226338 405854 226574
rect 405234 190894 405854 226338
rect 405234 190658 405266 190894
rect 405502 190658 405586 190894
rect 405822 190658 405854 190894
rect 405234 190574 405854 190658
rect 405234 190338 405266 190574
rect 405502 190338 405586 190574
rect 405822 190338 405854 190574
rect 405234 154894 405854 190338
rect 405234 154658 405266 154894
rect 405502 154658 405586 154894
rect 405822 154658 405854 154894
rect 405234 154574 405854 154658
rect 405234 154338 405266 154574
rect 405502 154338 405586 154574
rect 405822 154338 405854 154574
rect 405234 118894 405854 154338
rect 405234 118658 405266 118894
rect 405502 118658 405586 118894
rect 405822 118658 405854 118894
rect 405234 118574 405854 118658
rect 405234 118338 405266 118574
rect 405502 118338 405586 118574
rect 405822 118338 405854 118574
rect 405234 82894 405854 118338
rect 405234 82658 405266 82894
rect 405502 82658 405586 82894
rect 405822 82658 405854 82894
rect 405234 82574 405854 82658
rect 405234 82338 405266 82574
rect 405502 82338 405586 82574
rect 405822 82338 405854 82574
rect 405234 46894 405854 82338
rect 405234 46658 405266 46894
rect 405502 46658 405586 46894
rect 405822 46658 405854 46894
rect 405234 46574 405854 46658
rect 405234 46338 405266 46574
rect 405502 46338 405586 46574
rect 405822 46338 405854 46574
rect 405234 10894 405854 46338
rect 405234 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 405854 10894
rect 405234 10574 405854 10658
rect 405234 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 405854 10574
rect 405234 -2266 405854 10338
rect 405234 -2502 405266 -2266
rect 405502 -2502 405586 -2266
rect 405822 -2502 405854 -2266
rect 405234 -2586 405854 -2502
rect 405234 -2822 405266 -2586
rect 405502 -2822 405586 -2586
rect 405822 -2822 405854 -2586
rect 405234 -7654 405854 -2822
rect 408954 302614 409574 338058
rect 412674 708678 413294 711590
rect 412674 708442 412706 708678
rect 412942 708442 413026 708678
rect 413262 708442 413294 708678
rect 412674 708358 413294 708442
rect 412674 708122 412706 708358
rect 412942 708122 413026 708358
rect 413262 708122 413294 708358
rect 412674 666334 413294 708122
rect 412674 666098 412706 666334
rect 412942 666098 413026 666334
rect 413262 666098 413294 666334
rect 412674 666014 413294 666098
rect 412674 665778 412706 666014
rect 412942 665778 413026 666014
rect 413262 665778 413294 666014
rect 412674 630334 413294 665778
rect 412674 630098 412706 630334
rect 412942 630098 413026 630334
rect 413262 630098 413294 630334
rect 412674 630014 413294 630098
rect 412674 629778 412706 630014
rect 412942 629778 413026 630014
rect 413262 629778 413294 630014
rect 412674 594334 413294 629778
rect 412674 594098 412706 594334
rect 412942 594098 413026 594334
rect 413262 594098 413294 594334
rect 412674 594014 413294 594098
rect 412674 593778 412706 594014
rect 412942 593778 413026 594014
rect 413262 593778 413294 594014
rect 412674 558334 413294 593778
rect 412674 558098 412706 558334
rect 412942 558098 413026 558334
rect 413262 558098 413294 558334
rect 412674 558014 413294 558098
rect 412674 557778 412706 558014
rect 412942 557778 413026 558014
rect 413262 557778 413294 558014
rect 412674 522334 413294 557778
rect 412674 522098 412706 522334
rect 412942 522098 413026 522334
rect 413262 522098 413294 522334
rect 412674 522014 413294 522098
rect 412674 521778 412706 522014
rect 412942 521778 413026 522014
rect 413262 521778 413294 522014
rect 412674 486334 413294 521778
rect 412674 486098 412706 486334
rect 412942 486098 413026 486334
rect 413262 486098 413294 486334
rect 412674 486014 413294 486098
rect 412674 485778 412706 486014
rect 412942 485778 413026 486014
rect 413262 485778 413294 486014
rect 412674 450334 413294 485778
rect 412674 450098 412706 450334
rect 412942 450098 413026 450334
rect 413262 450098 413294 450334
rect 412674 450014 413294 450098
rect 412674 449778 412706 450014
rect 412942 449778 413026 450014
rect 413262 449778 413294 450014
rect 412674 414334 413294 449778
rect 412674 414098 412706 414334
rect 412942 414098 413026 414334
rect 413262 414098 413294 414334
rect 412674 414014 413294 414098
rect 412674 413778 412706 414014
rect 412942 413778 413026 414014
rect 413262 413778 413294 414014
rect 412674 378334 413294 413778
rect 412674 378098 412706 378334
rect 412942 378098 413026 378334
rect 413262 378098 413294 378334
rect 412674 378014 413294 378098
rect 412674 377778 412706 378014
rect 412942 377778 413026 378014
rect 413262 377778 413294 378014
rect 412674 342334 413294 377778
rect 412674 342098 412706 342334
rect 412942 342098 413026 342334
rect 413262 342098 413294 342334
rect 412674 342014 413294 342098
rect 412674 341778 412706 342014
rect 412942 341778 413026 342014
rect 413262 341778 413294 342014
rect 411363 327454 411683 327486
rect 411363 327218 411405 327454
rect 411641 327218 411683 327454
rect 411363 327134 411683 327218
rect 411363 326898 411405 327134
rect 411641 326898 411683 327134
rect 411363 326866 411683 326898
rect 408954 302378 408986 302614
rect 409222 302378 409306 302614
rect 409542 302378 409574 302614
rect 408954 302294 409574 302378
rect 408954 302058 408986 302294
rect 409222 302058 409306 302294
rect 409542 302058 409574 302294
rect 408954 266614 409574 302058
rect 408954 266378 408986 266614
rect 409222 266378 409306 266614
rect 409542 266378 409574 266614
rect 408954 266294 409574 266378
rect 408954 266058 408986 266294
rect 409222 266058 409306 266294
rect 409542 266058 409574 266294
rect 408954 230614 409574 266058
rect 408954 230378 408986 230614
rect 409222 230378 409306 230614
rect 409542 230378 409574 230614
rect 408954 230294 409574 230378
rect 408954 230058 408986 230294
rect 409222 230058 409306 230294
rect 409542 230058 409574 230294
rect 408954 194614 409574 230058
rect 408954 194378 408986 194614
rect 409222 194378 409306 194614
rect 409542 194378 409574 194614
rect 408954 194294 409574 194378
rect 408954 194058 408986 194294
rect 409222 194058 409306 194294
rect 409542 194058 409574 194294
rect 408954 158614 409574 194058
rect 408954 158378 408986 158614
rect 409222 158378 409306 158614
rect 409542 158378 409574 158614
rect 408954 158294 409574 158378
rect 408954 158058 408986 158294
rect 409222 158058 409306 158294
rect 409542 158058 409574 158294
rect 408954 122614 409574 158058
rect 408954 122378 408986 122614
rect 409222 122378 409306 122614
rect 409542 122378 409574 122614
rect 408954 122294 409574 122378
rect 408954 122058 408986 122294
rect 409222 122058 409306 122294
rect 409542 122058 409574 122294
rect 408954 86614 409574 122058
rect 408954 86378 408986 86614
rect 409222 86378 409306 86614
rect 409542 86378 409574 86614
rect 408954 86294 409574 86378
rect 408954 86058 408986 86294
rect 409222 86058 409306 86294
rect 409542 86058 409574 86294
rect 408954 50614 409574 86058
rect 408954 50378 408986 50614
rect 409222 50378 409306 50614
rect 409542 50378 409574 50614
rect 408954 50294 409574 50378
rect 408954 50058 408986 50294
rect 409222 50058 409306 50294
rect 409542 50058 409574 50294
rect 408954 14614 409574 50058
rect 408954 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 409574 14614
rect 408954 14294 409574 14378
rect 408954 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 409574 14294
rect 408954 -3226 409574 14058
rect 408954 -3462 408986 -3226
rect 409222 -3462 409306 -3226
rect 409542 -3462 409574 -3226
rect 408954 -3546 409574 -3462
rect 408954 -3782 408986 -3546
rect 409222 -3782 409306 -3546
rect 409542 -3782 409574 -3546
rect 408954 -7654 409574 -3782
rect 412674 306334 413294 341778
rect 416394 709638 417014 711590
rect 416394 709402 416426 709638
rect 416662 709402 416746 709638
rect 416982 709402 417014 709638
rect 416394 709318 417014 709402
rect 416394 709082 416426 709318
rect 416662 709082 416746 709318
rect 416982 709082 417014 709318
rect 416394 670054 417014 709082
rect 416394 669818 416426 670054
rect 416662 669818 416746 670054
rect 416982 669818 417014 670054
rect 416394 669734 417014 669818
rect 416394 669498 416426 669734
rect 416662 669498 416746 669734
rect 416982 669498 417014 669734
rect 416394 634054 417014 669498
rect 416394 633818 416426 634054
rect 416662 633818 416746 634054
rect 416982 633818 417014 634054
rect 416394 633734 417014 633818
rect 416394 633498 416426 633734
rect 416662 633498 416746 633734
rect 416982 633498 417014 633734
rect 416394 598054 417014 633498
rect 416394 597818 416426 598054
rect 416662 597818 416746 598054
rect 416982 597818 417014 598054
rect 416394 597734 417014 597818
rect 416394 597498 416426 597734
rect 416662 597498 416746 597734
rect 416982 597498 417014 597734
rect 416394 562054 417014 597498
rect 416394 561818 416426 562054
rect 416662 561818 416746 562054
rect 416982 561818 417014 562054
rect 416394 561734 417014 561818
rect 416394 561498 416426 561734
rect 416662 561498 416746 561734
rect 416982 561498 417014 561734
rect 416394 526054 417014 561498
rect 416394 525818 416426 526054
rect 416662 525818 416746 526054
rect 416982 525818 417014 526054
rect 416394 525734 417014 525818
rect 416394 525498 416426 525734
rect 416662 525498 416746 525734
rect 416982 525498 417014 525734
rect 416394 490054 417014 525498
rect 416394 489818 416426 490054
rect 416662 489818 416746 490054
rect 416982 489818 417014 490054
rect 416394 489734 417014 489818
rect 416394 489498 416426 489734
rect 416662 489498 416746 489734
rect 416982 489498 417014 489734
rect 416394 454054 417014 489498
rect 416394 453818 416426 454054
rect 416662 453818 416746 454054
rect 416982 453818 417014 454054
rect 416394 453734 417014 453818
rect 416394 453498 416426 453734
rect 416662 453498 416746 453734
rect 416982 453498 417014 453734
rect 416394 418054 417014 453498
rect 416394 417818 416426 418054
rect 416662 417818 416746 418054
rect 416982 417818 417014 418054
rect 416394 417734 417014 417818
rect 416394 417498 416426 417734
rect 416662 417498 416746 417734
rect 416982 417498 417014 417734
rect 416394 382054 417014 417498
rect 416394 381818 416426 382054
rect 416662 381818 416746 382054
rect 416982 381818 417014 382054
rect 416394 381734 417014 381818
rect 416394 381498 416426 381734
rect 416662 381498 416746 381734
rect 416982 381498 417014 381734
rect 416394 346054 417014 381498
rect 416394 345818 416426 346054
rect 416662 345818 416746 346054
rect 416982 345818 417014 346054
rect 416394 345734 417014 345818
rect 416394 345498 416426 345734
rect 416662 345498 416746 345734
rect 416982 345498 417014 345734
rect 414836 331174 415156 331206
rect 414836 330938 414878 331174
rect 415114 330938 415156 331174
rect 414836 330854 415156 330938
rect 414836 330618 414878 330854
rect 415114 330618 415156 330854
rect 414836 330586 415156 330618
rect 412674 306098 412706 306334
rect 412942 306098 413026 306334
rect 413262 306098 413294 306334
rect 412674 306014 413294 306098
rect 412674 305778 412706 306014
rect 412942 305778 413026 306014
rect 413262 305778 413294 306014
rect 412674 270334 413294 305778
rect 412674 270098 412706 270334
rect 412942 270098 413026 270334
rect 413262 270098 413294 270334
rect 412674 270014 413294 270098
rect 412674 269778 412706 270014
rect 412942 269778 413026 270014
rect 413262 269778 413294 270014
rect 412674 234334 413294 269778
rect 412674 234098 412706 234334
rect 412942 234098 413026 234334
rect 413262 234098 413294 234334
rect 412674 234014 413294 234098
rect 412674 233778 412706 234014
rect 412942 233778 413026 234014
rect 413262 233778 413294 234014
rect 412674 198334 413294 233778
rect 412674 198098 412706 198334
rect 412942 198098 413026 198334
rect 413262 198098 413294 198334
rect 412674 198014 413294 198098
rect 412674 197778 412706 198014
rect 412942 197778 413026 198014
rect 413262 197778 413294 198014
rect 412674 162334 413294 197778
rect 412674 162098 412706 162334
rect 412942 162098 413026 162334
rect 413262 162098 413294 162334
rect 412674 162014 413294 162098
rect 412674 161778 412706 162014
rect 412942 161778 413026 162014
rect 413262 161778 413294 162014
rect 412674 126334 413294 161778
rect 416394 310054 417014 345498
rect 420114 710598 420734 711590
rect 420114 710362 420146 710598
rect 420382 710362 420466 710598
rect 420702 710362 420734 710598
rect 420114 710278 420734 710362
rect 420114 710042 420146 710278
rect 420382 710042 420466 710278
rect 420702 710042 420734 710278
rect 420114 673774 420734 710042
rect 420114 673538 420146 673774
rect 420382 673538 420466 673774
rect 420702 673538 420734 673774
rect 420114 673454 420734 673538
rect 420114 673218 420146 673454
rect 420382 673218 420466 673454
rect 420702 673218 420734 673454
rect 420114 637774 420734 673218
rect 420114 637538 420146 637774
rect 420382 637538 420466 637774
rect 420702 637538 420734 637774
rect 420114 637454 420734 637538
rect 420114 637218 420146 637454
rect 420382 637218 420466 637454
rect 420702 637218 420734 637454
rect 420114 601774 420734 637218
rect 420114 601538 420146 601774
rect 420382 601538 420466 601774
rect 420702 601538 420734 601774
rect 420114 601454 420734 601538
rect 420114 601218 420146 601454
rect 420382 601218 420466 601454
rect 420702 601218 420734 601454
rect 420114 565774 420734 601218
rect 420114 565538 420146 565774
rect 420382 565538 420466 565774
rect 420702 565538 420734 565774
rect 420114 565454 420734 565538
rect 420114 565218 420146 565454
rect 420382 565218 420466 565454
rect 420702 565218 420734 565454
rect 420114 529774 420734 565218
rect 420114 529538 420146 529774
rect 420382 529538 420466 529774
rect 420702 529538 420734 529774
rect 420114 529454 420734 529538
rect 420114 529218 420146 529454
rect 420382 529218 420466 529454
rect 420702 529218 420734 529454
rect 420114 493774 420734 529218
rect 420114 493538 420146 493774
rect 420382 493538 420466 493774
rect 420702 493538 420734 493774
rect 420114 493454 420734 493538
rect 420114 493218 420146 493454
rect 420382 493218 420466 493454
rect 420702 493218 420734 493454
rect 420114 457774 420734 493218
rect 420114 457538 420146 457774
rect 420382 457538 420466 457774
rect 420702 457538 420734 457774
rect 420114 457454 420734 457538
rect 420114 457218 420146 457454
rect 420382 457218 420466 457454
rect 420702 457218 420734 457454
rect 420114 421774 420734 457218
rect 423834 711558 424454 711590
rect 423834 711322 423866 711558
rect 424102 711322 424186 711558
rect 424422 711322 424454 711558
rect 423834 711238 424454 711322
rect 423834 711002 423866 711238
rect 424102 711002 424186 711238
rect 424422 711002 424454 711238
rect 423834 677494 424454 711002
rect 423834 677258 423866 677494
rect 424102 677258 424186 677494
rect 424422 677258 424454 677494
rect 423834 677174 424454 677258
rect 423834 676938 423866 677174
rect 424102 676938 424186 677174
rect 424422 676938 424454 677174
rect 423834 641494 424454 676938
rect 423834 641258 423866 641494
rect 424102 641258 424186 641494
rect 424422 641258 424454 641494
rect 423834 641174 424454 641258
rect 423834 640938 423866 641174
rect 424102 640938 424186 641174
rect 424422 640938 424454 641174
rect 423834 605494 424454 640938
rect 423834 605258 423866 605494
rect 424102 605258 424186 605494
rect 424422 605258 424454 605494
rect 423834 605174 424454 605258
rect 423834 604938 423866 605174
rect 424102 604938 424186 605174
rect 424422 604938 424454 605174
rect 423834 569494 424454 604938
rect 423834 569258 423866 569494
rect 424102 569258 424186 569494
rect 424422 569258 424454 569494
rect 423834 569174 424454 569258
rect 423834 568938 423866 569174
rect 424102 568938 424186 569174
rect 424422 568938 424454 569174
rect 423834 533494 424454 568938
rect 423834 533258 423866 533494
rect 424102 533258 424186 533494
rect 424422 533258 424454 533494
rect 423834 533174 424454 533258
rect 423834 532938 423866 533174
rect 424102 532938 424186 533174
rect 424422 532938 424454 533174
rect 423834 497494 424454 532938
rect 423834 497258 423866 497494
rect 424102 497258 424186 497494
rect 424422 497258 424454 497494
rect 423834 497174 424454 497258
rect 423834 496938 423866 497174
rect 424102 496938 424186 497174
rect 424422 496938 424454 497174
rect 423834 461494 424454 496938
rect 423834 461258 423866 461494
rect 424102 461258 424186 461494
rect 424422 461258 424454 461494
rect 423834 461174 424454 461258
rect 423834 460938 423866 461174
rect 424102 460938 424186 461174
rect 424422 460938 424454 461174
rect 423834 444412 424454 460938
rect 433794 704838 434414 711590
rect 433794 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 434414 704838
rect 433794 704518 434414 704602
rect 433794 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 434414 704518
rect 433794 687454 434414 704282
rect 433794 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 434414 687454
rect 433794 687134 434414 687218
rect 433794 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 434414 687134
rect 433794 651454 434414 686898
rect 433794 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 434414 651454
rect 433794 651134 434414 651218
rect 433794 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 434414 651134
rect 433794 615454 434414 650898
rect 433794 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 434414 615454
rect 433794 615134 434414 615218
rect 433794 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 434414 615134
rect 433794 579454 434414 614898
rect 433794 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 434414 579454
rect 433794 579134 434414 579218
rect 433794 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 434414 579134
rect 433794 543454 434414 578898
rect 433794 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 434414 543454
rect 433794 543134 434414 543218
rect 433794 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 434414 543134
rect 433794 507454 434414 542898
rect 433794 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 434414 507454
rect 433794 507134 434414 507218
rect 433794 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 434414 507134
rect 433794 471454 434414 506898
rect 433794 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 434414 471454
rect 433794 471134 434414 471218
rect 433794 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 434414 471134
rect 433794 442833 434414 470898
rect 437514 705798 438134 711590
rect 437514 705562 437546 705798
rect 437782 705562 437866 705798
rect 438102 705562 438134 705798
rect 437514 705478 438134 705562
rect 437514 705242 437546 705478
rect 437782 705242 437866 705478
rect 438102 705242 438134 705478
rect 437514 691174 438134 705242
rect 437514 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 438134 691174
rect 437514 690854 438134 690938
rect 437514 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 438134 690854
rect 437514 655174 438134 690618
rect 437514 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 438134 655174
rect 437514 654854 438134 654938
rect 437514 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 438134 654854
rect 437514 619174 438134 654618
rect 437514 618938 437546 619174
rect 437782 618938 437866 619174
rect 438102 618938 438134 619174
rect 437514 618854 438134 618938
rect 437514 618618 437546 618854
rect 437782 618618 437866 618854
rect 438102 618618 438134 618854
rect 437514 583174 438134 618618
rect 437514 582938 437546 583174
rect 437782 582938 437866 583174
rect 438102 582938 438134 583174
rect 437514 582854 438134 582938
rect 437514 582618 437546 582854
rect 437782 582618 437866 582854
rect 438102 582618 438134 582854
rect 437514 547174 438134 582618
rect 437514 546938 437546 547174
rect 437782 546938 437866 547174
rect 438102 546938 438134 547174
rect 437514 546854 438134 546938
rect 437514 546618 437546 546854
rect 437782 546618 437866 546854
rect 438102 546618 438134 546854
rect 437514 511174 438134 546618
rect 437514 510938 437546 511174
rect 437782 510938 437866 511174
rect 438102 510938 438134 511174
rect 437514 510854 438134 510938
rect 437514 510618 437546 510854
rect 437782 510618 437866 510854
rect 438102 510618 438134 510854
rect 437514 475174 438134 510618
rect 437514 474938 437546 475174
rect 437782 474938 437866 475174
rect 438102 474938 438134 475174
rect 437514 474854 438134 474938
rect 437514 474618 437546 474854
rect 437782 474618 437866 474854
rect 438102 474618 438134 474854
rect 437514 444412 438134 474618
rect 441234 706758 441854 711590
rect 441234 706522 441266 706758
rect 441502 706522 441586 706758
rect 441822 706522 441854 706758
rect 441234 706438 441854 706522
rect 441234 706202 441266 706438
rect 441502 706202 441586 706438
rect 441822 706202 441854 706438
rect 441234 694894 441854 706202
rect 444954 707718 445574 711590
rect 444954 707482 444986 707718
rect 445222 707482 445306 707718
rect 445542 707482 445574 707718
rect 444954 707398 445574 707482
rect 444954 707162 444986 707398
rect 445222 707162 445306 707398
rect 445542 707162 445574 707398
rect 444235 700364 444301 700365
rect 444235 700300 444236 700364
rect 444300 700300 444301 700364
rect 444235 700299 444301 700300
rect 441234 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 441854 694894
rect 441234 694574 441854 694658
rect 441234 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 441854 694574
rect 441234 658894 441854 694338
rect 441234 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 441854 658894
rect 441234 658574 441854 658658
rect 441234 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 441854 658574
rect 441234 622894 441854 658338
rect 441234 622658 441266 622894
rect 441502 622658 441586 622894
rect 441822 622658 441854 622894
rect 441234 622574 441854 622658
rect 441234 622338 441266 622574
rect 441502 622338 441586 622574
rect 441822 622338 441854 622574
rect 441234 586894 441854 622338
rect 441234 586658 441266 586894
rect 441502 586658 441586 586894
rect 441822 586658 441854 586894
rect 441234 586574 441854 586658
rect 441234 586338 441266 586574
rect 441502 586338 441586 586574
rect 441822 586338 441854 586574
rect 441234 550894 441854 586338
rect 441234 550658 441266 550894
rect 441502 550658 441586 550894
rect 441822 550658 441854 550894
rect 441234 550574 441854 550658
rect 441234 550338 441266 550574
rect 441502 550338 441586 550574
rect 441822 550338 441854 550574
rect 441234 514894 441854 550338
rect 441234 514658 441266 514894
rect 441502 514658 441586 514894
rect 441822 514658 441854 514894
rect 441234 514574 441854 514658
rect 441234 514338 441266 514574
rect 441502 514338 441586 514574
rect 441822 514338 441854 514574
rect 441234 478894 441854 514338
rect 441234 478658 441266 478894
rect 441502 478658 441586 478894
rect 441822 478658 441854 478894
rect 441234 478574 441854 478658
rect 441234 478338 441266 478574
rect 441502 478338 441586 478574
rect 441822 478338 441854 478574
rect 441234 442833 441854 478338
rect 426624 439174 426944 439206
rect 426624 438938 426666 439174
rect 426902 438938 426944 439174
rect 426624 438854 426944 438938
rect 426624 438618 426666 438854
rect 426902 438618 426944 438854
rect 426624 438586 426944 438618
rect 432305 439174 432625 439206
rect 432305 438938 432347 439174
rect 432583 438938 432625 439174
rect 432305 438854 432625 438938
rect 432305 438618 432347 438854
rect 432583 438618 432625 438854
rect 432305 438586 432625 438618
rect 437986 439174 438306 439206
rect 437986 438938 438028 439174
rect 438264 438938 438306 439174
rect 437986 438854 438306 438938
rect 437986 438618 438028 438854
rect 438264 438618 438306 438854
rect 437986 438586 438306 438618
rect 443667 439174 443987 439206
rect 443667 438938 443709 439174
rect 443945 438938 443987 439174
rect 443667 438854 443987 438938
rect 443667 438618 443709 438854
rect 443945 438618 443987 438854
rect 443667 438586 443987 438618
rect 423784 435454 424104 435486
rect 423784 435218 423826 435454
rect 424062 435218 424104 435454
rect 423784 435134 424104 435218
rect 423784 434898 423826 435134
rect 424062 434898 424104 435134
rect 423784 434866 424104 434898
rect 429465 435454 429785 435486
rect 429465 435218 429507 435454
rect 429743 435218 429785 435454
rect 429465 435134 429785 435218
rect 429465 434898 429507 435134
rect 429743 434898 429785 435134
rect 429465 434866 429785 434898
rect 435146 435454 435466 435486
rect 435146 435218 435188 435454
rect 435424 435218 435466 435454
rect 435146 435134 435466 435218
rect 435146 434898 435188 435134
rect 435424 434898 435466 435134
rect 435146 434866 435466 434898
rect 440827 435454 441147 435486
rect 440827 435218 440869 435454
rect 441105 435218 441147 435454
rect 440827 435134 441147 435218
rect 440827 434898 440869 435134
rect 441105 434898 441147 435134
rect 440827 434866 441147 434898
rect 420114 421538 420146 421774
rect 420382 421538 420466 421774
rect 420702 421538 420734 421774
rect 420114 421454 420734 421538
rect 420114 421218 420146 421454
rect 420382 421218 420466 421454
rect 420702 421218 420734 421454
rect 420114 385774 420734 421218
rect 420114 385538 420146 385774
rect 420382 385538 420466 385774
rect 420702 385538 420734 385774
rect 420114 385454 420734 385538
rect 420114 385218 420146 385454
rect 420382 385218 420466 385454
rect 420702 385218 420734 385454
rect 420114 349774 420734 385218
rect 420114 349538 420146 349774
rect 420382 349538 420466 349774
rect 420702 349538 420734 349774
rect 420114 349454 420734 349538
rect 420114 349218 420146 349454
rect 420382 349218 420466 349454
rect 420702 349218 420734 349454
rect 418309 327454 418629 327486
rect 418309 327218 418351 327454
rect 418587 327218 418629 327454
rect 418309 327134 418629 327218
rect 418309 326898 418351 327134
rect 418587 326898 418629 327134
rect 418309 326866 418629 326898
rect 416394 309818 416426 310054
rect 416662 309818 416746 310054
rect 416982 309818 417014 310054
rect 416394 309734 417014 309818
rect 416394 309498 416426 309734
rect 416662 309498 416746 309734
rect 416982 309498 417014 309734
rect 416394 274054 417014 309498
rect 416394 273818 416426 274054
rect 416662 273818 416746 274054
rect 416982 273818 417014 274054
rect 416394 273734 417014 273818
rect 416394 273498 416426 273734
rect 416662 273498 416746 273734
rect 416982 273498 417014 273734
rect 416394 238054 417014 273498
rect 416394 237818 416426 238054
rect 416662 237818 416746 238054
rect 416982 237818 417014 238054
rect 416394 237734 417014 237818
rect 416394 237498 416426 237734
rect 416662 237498 416746 237734
rect 416982 237498 417014 237734
rect 416394 202054 417014 237498
rect 416394 201818 416426 202054
rect 416662 201818 416746 202054
rect 416982 201818 417014 202054
rect 416394 201734 417014 201818
rect 416394 201498 416426 201734
rect 416662 201498 416746 201734
rect 416982 201498 417014 201734
rect 416394 166054 417014 201498
rect 416394 165818 416426 166054
rect 416662 165818 416746 166054
rect 416982 165818 417014 166054
rect 416394 165734 417014 165818
rect 416394 165498 416426 165734
rect 416662 165498 416746 165734
rect 416982 165498 417014 165734
rect 416394 157249 417014 165498
rect 420114 313774 420734 349218
rect 423834 389494 424454 420068
rect 423834 389258 423866 389494
rect 424102 389258 424186 389494
rect 424422 389258 424454 389494
rect 423834 389174 424454 389258
rect 423834 388938 423866 389174
rect 424102 388938 424186 389174
rect 424422 388938 424454 389174
rect 423834 353494 424454 388938
rect 423834 353258 423866 353494
rect 424102 353258 424186 353494
rect 424422 353258 424454 353494
rect 423834 353174 424454 353258
rect 423834 352938 423866 353174
rect 424102 352938 424186 353174
rect 424422 352938 424454 353174
rect 421419 334116 421485 334117
rect 421419 334052 421420 334116
rect 421484 334052 421485 334116
rect 421419 334051 421485 334052
rect 420114 313538 420146 313774
rect 420382 313538 420466 313774
rect 420702 313538 420734 313774
rect 420114 313454 420734 313538
rect 420114 313218 420146 313454
rect 420382 313218 420466 313454
rect 420702 313218 420734 313454
rect 420114 277774 420734 313218
rect 420114 277538 420146 277774
rect 420382 277538 420466 277774
rect 420702 277538 420734 277774
rect 420114 277454 420734 277538
rect 420114 277218 420146 277454
rect 420382 277218 420466 277454
rect 420702 277218 420734 277454
rect 420114 241774 420734 277218
rect 420114 241538 420146 241774
rect 420382 241538 420466 241774
rect 420702 241538 420734 241774
rect 420114 241454 420734 241538
rect 420114 241218 420146 241454
rect 420382 241218 420466 241454
rect 420702 241218 420734 241454
rect 420114 205774 420734 241218
rect 420114 205538 420146 205774
rect 420382 205538 420466 205774
rect 420702 205538 420734 205774
rect 420114 205454 420734 205538
rect 420114 205218 420146 205454
rect 420382 205218 420466 205454
rect 420702 205218 420734 205454
rect 420114 169774 420734 205218
rect 420114 169538 420146 169774
rect 420382 169538 420466 169774
rect 420702 169538 420734 169774
rect 420114 169454 420734 169538
rect 420114 169218 420146 169454
rect 420382 169218 420466 169454
rect 420702 169218 420734 169454
rect 420114 157249 420734 169218
rect 421422 162757 421482 334051
rect 421782 331174 422102 331206
rect 421782 330938 421824 331174
rect 422060 330938 422102 331174
rect 421782 330854 422102 330938
rect 421782 330618 421824 330854
rect 422060 330618 422102 330854
rect 421782 330586 422102 330618
rect 423834 317494 424454 352938
rect 433794 399454 434414 422599
rect 433794 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 434414 399454
rect 433794 399134 434414 399218
rect 433794 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 434414 399134
rect 433794 363454 434414 398898
rect 433794 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 434414 363454
rect 433794 363134 434414 363218
rect 433794 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 434414 363134
rect 428411 334524 428477 334525
rect 428411 334460 428412 334524
rect 428476 334460 428477 334524
rect 428411 334459 428477 334460
rect 425835 334388 425901 334389
rect 425835 334324 425836 334388
rect 425900 334324 425901 334388
rect 425835 334323 425901 334324
rect 425255 327454 425575 327486
rect 425255 327218 425297 327454
rect 425533 327218 425575 327454
rect 425255 327134 425575 327218
rect 425255 326898 425297 327134
rect 425533 326898 425575 327134
rect 425255 326866 425575 326898
rect 423834 317258 423866 317494
rect 424102 317258 424186 317494
rect 424422 317258 424454 317494
rect 423834 317174 424454 317258
rect 423834 316938 423866 317174
rect 424102 316938 424186 317174
rect 424422 316938 424454 317174
rect 423834 281494 424454 316938
rect 423834 281258 423866 281494
rect 424102 281258 424186 281494
rect 424422 281258 424454 281494
rect 423834 281174 424454 281258
rect 423834 280938 423866 281174
rect 424102 280938 424186 281174
rect 424422 280938 424454 281174
rect 423834 245494 424454 280938
rect 423834 245258 423866 245494
rect 424102 245258 424186 245494
rect 424422 245258 424454 245494
rect 423834 245174 424454 245258
rect 423834 244938 423866 245174
rect 424102 244938 424186 245174
rect 424422 244938 424454 245174
rect 423834 209494 424454 244938
rect 423834 209258 423866 209494
rect 424102 209258 424186 209494
rect 424422 209258 424454 209494
rect 423834 209174 424454 209258
rect 423834 208938 423866 209174
rect 424102 208938 424186 209174
rect 424422 208938 424454 209174
rect 423834 173494 424454 208938
rect 423834 173258 423866 173494
rect 424102 173258 424186 173494
rect 424422 173258 424454 173494
rect 423834 173174 424454 173258
rect 423834 172938 423866 173174
rect 424102 172938 424186 173174
rect 424422 172938 424454 173174
rect 421419 162756 421485 162757
rect 421419 162692 421420 162756
rect 421484 162692 421485 162756
rect 421419 162691 421485 162692
rect 423834 157249 424454 172938
rect 425838 162757 425898 334323
rect 428414 162757 428474 334459
rect 428728 331174 429048 331206
rect 428728 330938 428770 331174
rect 429006 330938 429048 331174
rect 428728 330854 429048 330938
rect 428728 330618 428770 330854
rect 429006 330618 429048 330854
rect 428728 330586 429048 330618
rect 433794 327454 434414 362898
rect 433794 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 434414 327454
rect 433794 327134 434414 327218
rect 433794 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 434414 327134
rect 433794 291454 434414 326898
rect 433794 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 434414 291454
rect 433794 291134 434414 291218
rect 433794 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 434414 291134
rect 433794 255454 434414 290898
rect 433794 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 434414 255454
rect 433794 255134 434414 255218
rect 433794 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 434414 255134
rect 433794 219454 434414 254898
rect 433794 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 434414 219454
rect 433794 219134 434414 219218
rect 433794 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 434414 219134
rect 433794 183454 434414 218898
rect 433794 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 434414 183454
rect 433794 183134 434414 183218
rect 433794 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 434414 183134
rect 425835 162756 425901 162757
rect 425835 162692 425836 162756
rect 425900 162692 425901 162756
rect 425835 162691 425901 162692
rect 428411 162756 428477 162757
rect 428411 162692 428412 162756
rect 428476 162692 428477 162756
rect 428411 162691 428477 162692
rect 433794 157249 434414 182898
rect 437514 403174 438134 420068
rect 437514 402938 437546 403174
rect 437782 402938 437866 403174
rect 438102 402938 438134 403174
rect 437514 402854 438134 402938
rect 437514 402618 437546 402854
rect 437782 402618 437866 402854
rect 438102 402618 438134 402854
rect 437514 367174 438134 402618
rect 437514 366938 437546 367174
rect 437782 366938 437866 367174
rect 438102 366938 438134 367174
rect 437514 366854 438134 366938
rect 437514 366618 437546 366854
rect 437782 366618 437866 366854
rect 438102 366618 438134 366854
rect 437514 331174 438134 366618
rect 437514 330938 437546 331174
rect 437782 330938 437866 331174
rect 438102 330938 438134 331174
rect 437514 330854 438134 330938
rect 437514 330618 437546 330854
rect 437782 330618 437866 330854
rect 438102 330618 438134 330854
rect 437514 295174 438134 330618
rect 437514 294938 437546 295174
rect 437782 294938 437866 295174
rect 438102 294938 438134 295174
rect 437514 294854 438134 294938
rect 437514 294618 437546 294854
rect 437782 294618 437866 294854
rect 438102 294618 438134 294854
rect 437514 259174 438134 294618
rect 437514 258938 437546 259174
rect 437782 258938 437866 259174
rect 438102 258938 438134 259174
rect 437514 258854 438134 258938
rect 437514 258618 437546 258854
rect 437782 258618 437866 258854
rect 438102 258618 438134 258854
rect 437514 223174 438134 258618
rect 437514 222938 437546 223174
rect 437782 222938 437866 223174
rect 438102 222938 438134 223174
rect 437514 222854 438134 222938
rect 437514 222618 437546 222854
rect 437782 222618 437866 222854
rect 438102 222618 438134 222854
rect 437514 187174 438134 222618
rect 437514 186938 437546 187174
rect 437782 186938 437866 187174
rect 438102 186938 438134 187174
rect 437514 186854 438134 186938
rect 437514 186618 437546 186854
rect 437782 186618 437866 186854
rect 438102 186618 438134 186854
rect 437514 157249 438134 186618
rect 441234 406894 441854 422599
rect 443499 421972 443565 421973
rect 443499 421908 443500 421972
rect 443564 421908 443565 421972
rect 443499 421907 443565 421908
rect 441234 406658 441266 406894
rect 441502 406658 441586 406894
rect 441822 406658 441854 406894
rect 441234 406574 441854 406658
rect 441234 406338 441266 406574
rect 441502 406338 441586 406574
rect 441822 406338 441854 406574
rect 441234 370894 441854 406338
rect 441234 370658 441266 370894
rect 441502 370658 441586 370894
rect 441822 370658 441854 370894
rect 441234 370574 441854 370658
rect 441234 370338 441266 370574
rect 441502 370338 441586 370574
rect 441822 370338 441854 370574
rect 441234 334894 441854 370338
rect 441234 334658 441266 334894
rect 441502 334658 441586 334894
rect 441822 334658 441854 334894
rect 441234 334574 441854 334658
rect 441234 334338 441266 334574
rect 441502 334338 441586 334574
rect 441822 334338 441854 334574
rect 441234 298894 441854 334338
rect 443502 321061 443562 421907
rect 444051 421836 444117 421837
rect 444051 421772 444052 421836
rect 444116 421772 444117 421836
rect 444051 421771 444117 421772
rect 443499 321060 443565 321061
rect 443499 320996 443500 321060
rect 443564 320996 443565 321060
rect 443499 320995 443565 320996
rect 444054 320109 444114 421771
rect 444238 321333 444298 700299
rect 444954 698614 445574 707162
rect 444954 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 445574 698614
rect 444954 698294 445574 698378
rect 444954 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 445574 698294
rect 444954 662614 445574 698058
rect 448674 708678 449294 711590
rect 448674 708442 448706 708678
rect 448942 708442 449026 708678
rect 449262 708442 449294 708678
rect 448674 708358 449294 708442
rect 448674 708122 448706 708358
rect 448942 708122 449026 708358
rect 449262 708122 449294 708358
rect 446259 686492 446325 686493
rect 446259 686428 446260 686492
rect 446324 686428 446325 686492
rect 446259 686427 446325 686428
rect 444954 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 445574 662614
rect 444954 662294 445574 662378
rect 444954 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 445574 662294
rect 444954 626614 445574 662058
rect 444954 626378 444986 626614
rect 445222 626378 445306 626614
rect 445542 626378 445574 626614
rect 444954 626294 445574 626378
rect 444954 626058 444986 626294
rect 445222 626058 445306 626294
rect 445542 626058 445574 626294
rect 444954 590614 445574 626058
rect 444954 590378 444986 590614
rect 445222 590378 445306 590614
rect 445542 590378 445574 590614
rect 444954 590294 445574 590378
rect 444954 590058 444986 590294
rect 445222 590058 445306 590294
rect 445542 590058 445574 590294
rect 444954 554614 445574 590058
rect 444954 554378 444986 554614
rect 445222 554378 445306 554614
rect 445542 554378 445574 554614
rect 444954 554294 445574 554378
rect 444954 554058 444986 554294
rect 445222 554058 445306 554294
rect 445542 554058 445574 554294
rect 444954 518614 445574 554058
rect 444954 518378 444986 518614
rect 445222 518378 445306 518614
rect 445542 518378 445574 518614
rect 444954 518294 445574 518378
rect 444954 518058 444986 518294
rect 445222 518058 445306 518294
rect 445542 518058 445574 518294
rect 444954 482614 445574 518058
rect 444954 482378 444986 482614
rect 445222 482378 445306 482614
rect 445542 482378 445574 482614
rect 444954 482294 445574 482378
rect 444954 482058 444986 482294
rect 445222 482058 445306 482294
rect 445542 482058 445574 482294
rect 444954 446614 445574 482058
rect 444954 446378 444986 446614
rect 445222 446378 445306 446614
rect 445542 446378 445574 446614
rect 444954 446294 445574 446378
rect 444954 446058 444986 446294
rect 445222 446058 445306 446294
rect 445542 446058 445574 446294
rect 444954 410614 445574 446058
rect 444954 410378 444986 410614
rect 445222 410378 445306 410614
rect 445542 410378 445574 410614
rect 444954 410294 445574 410378
rect 444954 410058 444986 410294
rect 445222 410058 445306 410294
rect 445542 410058 445574 410294
rect 444954 374614 445574 410058
rect 444954 374378 444986 374614
rect 445222 374378 445306 374614
rect 445542 374378 445574 374614
rect 444954 374294 445574 374378
rect 444954 374058 444986 374294
rect 445222 374058 445306 374294
rect 445542 374058 445574 374294
rect 444954 338614 445574 374058
rect 444954 338378 444986 338614
rect 445222 338378 445306 338614
rect 445542 338378 445574 338614
rect 444954 338294 445574 338378
rect 444954 338058 444986 338294
rect 445222 338058 445306 338294
rect 445542 338058 445574 338294
rect 444235 321332 444301 321333
rect 444235 321268 444236 321332
rect 444300 321268 444301 321332
rect 444235 321267 444301 321268
rect 444051 320108 444117 320109
rect 444051 320044 444052 320108
rect 444116 320044 444117 320108
rect 444051 320043 444117 320044
rect 441234 298658 441266 298894
rect 441502 298658 441586 298894
rect 441822 298658 441854 298894
rect 441234 298574 441854 298658
rect 441234 298338 441266 298574
rect 441502 298338 441586 298574
rect 441822 298338 441854 298574
rect 441234 262894 441854 298338
rect 441234 262658 441266 262894
rect 441502 262658 441586 262894
rect 441822 262658 441854 262894
rect 441234 262574 441854 262658
rect 441234 262338 441266 262574
rect 441502 262338 441586 262574
rect 441822 262338 441854 262574
rect 441234 226894 441854 262338
rect 441234 226658 441266 226894
rect 441502 226658 441586 226894
rect 441822 226658 441854 226894
rect 441234 226574 441854 226658
rect 441234 226338 441266 226574
rect 441502 226338 441586 226574
rect 441822 226338 441854 226574
rect 441234 190894 441854 226338
rect 441234 190658 441266 190894
rect 441502 190658 441586 190894
rect 441822 190658 441854 190894
rect 441234 190574 441854 190658
rect 441234 190338 441266 190574
rect 441502 190338 441586 190574
rect 441822 190338 441854 190574
rect 441234 157249 441854 190338
rect 444954 302614 445574 338058
rect 446262 319973 446322 686427
rect 447731 684316 447797 684317
rect 447731 684252 447732 684316
rect 447796 684252 447797 684316
rect 447731 684251 447797 684252
rect 447734 321197 447794 684251
rect 448674 666334 449294 708122
rect 448674 666098 448706 666334
rect 448942 666098 449026 666334
rect 449262 666098 449294 666334
rect 448674 666014 449294 666098
rect 448674 665778 448706 666014
rect 448942 665778 449026 666014
rect 449262 665778 449294 666014
rect 448674 630334 449294 665778
rect 448674 630098 448706 630334
rect 448942 630098 449026 630334
rect 449262 630098 449294 630334
rect 448674 630014 449294 630098
rect 448674 629778 448706 630014
rect 448942 629778 449026 630014
rect 449262 629778 449294 630014
rect 448674 594334 449294 629778
rect 448674 594098 448706 594334
rect 448942 594098 449026 594334
rect 449262 594098 449294 594334
rect 448674 594014 449294 594098
rect 448674 593778 448706 594014
rect 448942 593778 449026 594014
rect 449262 593778 449294 594014
rect 448674 558334 449294 593778
rect 448674 558098 448706 558334
rect 448942 558098 449026 558334
rect 449262 558098 449294 558334
rect 448674 558014 449294 558098
rect 448674 557778 448706 558014
rect 448942 557778 449026 558014
rect 449262 557778 449294 558014
rect 448674 522334 449294 557778
rect 448674 522098 448706 522334
rect 448942 522098 449026 522334
rect 449262 522098 449294 522334
rect 448674 522014 449294 522098
rect 448674 521778 448706 522014
rect 448942 521778 449026 522014
rect 449262 521778 449294 522014
rect 448674 486334 449294 521778
rect 452394 709638 453014 711590
rect 452394 709402 452426 709638
rect 452662 709402 452746 709638
rect 452982 709402 453014 709638
rect 452394 709318 453014 709402
rect 452394 709082 452426 709318
rect 452662 709082 452746 709318
rect 452982 709082 453014 709318
rect 452394 670054 453014 709082
rect 452394 669818 452426 670054
rect 452662 669818 452746 670054
rect 452982 669818 453014 670054
rect 452394 669734 453014 669818
rect 452394 669498 452426 669734
rect 452662 669498 452746 669734
rect 452982 669498 453014 669734
rect 452394 634054 453014 669498
rect 452394 633818 452426 634054
rect 452662 633818 452746 634054
rect 452982 633818 453014 634054
rect 452394 633734 453014 633818
rect 452394 633498 452426 633734
rect 452662 633498 452746 633734
rect 452982 633498 453014 633734
rect 452394 598054 453014 633498
rect 452394 597818 452426 598054
rect 452662 597818 452746 598054
rect 452982 597818 453014 598054
rect 452394 597734 453014 597818
rect 452394 597498 452426 597734
rect 452662 597498 452746 597734
rect 452982 597498 453014 597734
rect 452394 562054 453014 597498
rect 452394 561818 452426 562054
rect 452662 561818 452746 562054
rect 452982 561818 453014 562054
rect 452394 561734 453014 561818
rect 452394 561498 452426 561734
rect 452662 561498 452746 561734
rect 452982 561498 453014 561734
rect 452394 526054 453014 561498
rect 452394 525818 452426 526054
rect 452662 525818 452746 526054
rect 452982 525818 453014 526054
rect 452394 525734 453014 525818
rect 452394 525498 452426 525734
rect 452662 525498 452746 525734
rect 452982 525498 453014 525734
rect 452394 517884 453014 525498
rect 456114 710598 456734 711590
rect 456114 710362 456146 710598
rect 456382 710362 456466 710598
rect 456702 710362 456734 710598
rect 456114 710278 456734 710362
rect 456114 710042 456146 710278
rect 456382 710042 456466 710278
rect 456702 710042 456734 710278
rect 456114 673774 456734 710042
rect 456114 673538 456146 673774
rect 456382 673538 456466 673774
rect 456702 673538 456734 673774
rect 456114 673454 456734 673538
rect 456114 673218 456146 673454
rect 456382 673218 456466 673454
rect 456702 673218 456734 673454
rect 456114 637774 456734 673218
rect 459834 711558 460454 711590
rect 459834 711322 459866 711558
rect 460102 711322 460186 711558
rect 460422 711322 460454 711558
rect 459834 711238 460454 711322
rect 459834 711002 459866 711238
rect 460102 711002 460186 711238
rect 460422 711002 460454 711238
rect 459834 677494 460454 711002
rect 459834 677258 459866 677494
rect 460102 677258 460186 677494
rect 460422 677258 460454 677494
rect 459834 677174 460454 677258
rect 459834 676938 459866 677174
rect 460102 676938 460186 677174
rect 460422 676938 460454 677174
rect 459507 670580 459573 670581
rect 459507 670516 459508 670580
rect 459572 670516 459573 670580
rect 459507 670515 459573 670516
rect 458035 665276 458101 665277
rect 458035 665212 458036 665276
rect 458100 665212 458101 665276
rect 458035 665211 458101 665212
rect 456114 637538 456146 637774
rect 456382 637538 456466 637774
rect 456702 637538 456734 637774
rect 456114 637454 456734 637538
rect 456114 637218 456146 637454
rect 456382 637218 456466 637454
rect 456702 637218 456734 637454
rect 456114 601774 456734 637218
rect 456114 601538 456146 601774
rect 456382 601538 456466 601774
rect 456702 601538 456734 601774
rect 456114 601454 456734 601538
rect 456114 601218 456146 601454
rect 456382 601218 456466 601454
rect 456702 601218 456734 601454
rect 456114 565774 456734 601218
rect 456114 565538 456146 565774
rect 456382 565538 456466 565774
rect 456702 565538 456734 565774
rect 456114 565454 456734 565538
rect 456114 565218 456146 565454
rect 456382 565218 456466 565454
rect 456702 565218 456734 565454
rect 456114 529774 456734 565218
rect 456114 529538 456146 529774
rect 456382 529538 456466 529774
rect 456702 529538 456734 529774
rect 456114 529454 456734 529538
rect 456114 529218 456146 529454
rect 456382 529218 456466 529454
rect 456702 529218 456734 529454
rect 456114 517884 456734 529218
rect 458038 517581 458098 665211
rect 459139 655756 459205 655757
rect 459139 655692 459140 655756
rect 459204 655692 459205 655756
rect 459139 655691 459205 655692
rect 458955 647732 459021 647733
rect 458955 647668 458956 647732
rect 459020 647668 459021 647732
rect 458955 647667 459021 647668
rect 458035 517580 458101 517581
rect 458035 517516 458036 517580
rect 458100 517516 458101 517580
rect 458035 517515 458101 517516
rect 451043 516764 451109 516765
rect 451043 516700 451044 516764
rect 451108 516700 451109 516764
rect 451043 516699 451109 516700
rect 450491 514384 450557 514385
rect 450491 514320 450492 514384
rect 450556 514320 450557 514384
rect 450491 514319 450557 514320
rect 448674 486098 448706 486334
rect 448942 486098 449026 486334
rect 449262 486098 449294 486334
rect 448674 486014 449294 486098
rect 448674 485778 448706 486014
rect 448942 485778 449026 486014
rect 449262 485778 449294 486014
rect 448674 450334 449294 485778
rect 448674 450098 448706 450334
rect 448942 450098 449026 450334
rect 449262 450098 449294 450334
rect 448674 450014 449294 450098
rect 448674 449778 448706 450014
rect 448942 449778 449026 450014
rect 449262 449778 449294 450014
rect 448283 447268 448349 447269
rect 448283 447204 448284 447268
rect 448348 447204 448349 447268
rect 448283 447203 448349 447204
rect 448099 392596 448165 392597
rect 448099 392532 448100 392596
rect 448164 392532 448165 392596
rect 448099 392531 448165 392532
rect 448102 346221 448162 392531
rect 448099 346220 448165 346221
rect 448099 346156 448100 346220
rect 448164 346156 448165 346220
rect 448099 346155 448165 346156
rect 447915 334524 447981 334525
rect 447915 334460 447916 334524
rect 447980 334460 447981 334524
rect 447915 334459 447981 334460
rect 447731 321196 447797 321197
rect 447731 321132 447732 321196
rect 447796 321132 447797 321196
rect 447731 321131 447797 321132
rect 446259 319972 446325 319973
rect 446259 319908 446260 319972
rect 446324 319908 446325 319972
rect 446259 319907 446325 319908
rect 447918 319837 447978 334459
rect 448286 329901 448346 447203
rect 448674 414334 449294 449778
rect 448674 414098 448706 414334
rect 448942 414098 449026 414334
rect 449262 414098 449294 414334
rect 448674 414014 449294 414098
rect 448674 413778 448706 414014
rect 448942 413778 449026 414014
rect 449262 413778 449294 414014
rect 448674 378334 449294 413778
rect 448674 378098 448706 378334
rect 448942 378098 449026 378334
rect 449262 378098 449294 378334
rect 448674 378014 449294 378098
rect 448674 377778 448706 378014
rect 448942 377778 449026 378014
rect 449262 377778 449294 378014
rect 448674 342334 449294 377778
rect 448674 342098 448706 342334
rect 448942 342098 449026 342334
rect 449262 342098 449294 342334
rect 448674 342014 449294 342098
rect 448674 341778 448706 342014
rect 448942 341778 449026 342014
rect 449262 341778 449294 342014
rect 448283 329900 448349 329901
rect 448283 329836 448284 329900
rect 448348 329836 448349 329900
rect 448283 329835 448349 329836
rect 447915 319836 447981 319837
rect 447915 319772 447916 319836
rect 447980 319772 447981 319836
rect 447915 319771 447981 319772
rect 444954 302378 444986 302614
rect 445222 302378 445306 302614
rect 445542 302378 445574 302614
rect 444954 302294 445574 302378
rect 444954 302058 444986 302294
rect 445222 302058 445306 302294
rect 445542 302058 445574 302294
rect 444954 266614 445574 302058
rect 444954 266378 444986 266614
rect 445222 266378 445306 266614
rect 445542 266378 445574 266614
rect 444954 266294 445574 266378
rect 444954 266058 444986 266294
rect 445222 266058 445306 266294
rect 445542 266058 445574 266294
rect 444954 230614 445574 266058
rect 444954 230378 444986 230614
rect 445222 230378 445306 230614
rect 445542 230378 445574 230614
rect 444954 230294 445574 230378
rect 444954 230058 444986 230294
rect 445222 230058 445306 230294
rect 445542 230058 445574 230294
rect 444954 194614 445574 230058
rect 444954 194378 444986 194614
rect 445222 194378 445306 194614
rect 445542 194378 445574 194614
rect 444954 194294 445574 194378
rect 444954 194058 444986 194294
rect 445222 194058 445306 194294
rect 445542 194058 445574 194294
rect 444954 159644 445574 194058
rect 448674 306334 449294 341778
rect 450494 328677 450554 514319
rect 451046 335370 451106 516699
rect 453382 511174 453702 511206
rect 453382 510938 453424 511174
rect 453660 510938 453702 511174
rect 453382 510854 453702 510938
rect 453382 510618 453424 510854
rect 453660 510618 453702 510854
rect 453382 510586 453702 510618
rect 455820 511174 456140 511206
rect 455820 510938 455862 511174
rect 456098 510938 456140 511174
rect 455820 510854 456140 510938
rect 455820 510618 455862 510854
rect 456098 510618 456140 510854
rect 455820 510586 456140 510618
rect 458258 511174 458578 511206
rect 458258 510938 458300 511174
rect 458536 510938 458578 511174
rect 458258 510854 458578 510938
rect 458258 510618 458300 510854
rect 458536 510618 458578 510854
rect 458258 510586 458578 510618
rect 452163 507454 452483 507486
rect 452163 507218 452205 507454
rect 452441 507218 452483 507454
rect 452163 507134 452483 507218
rect 452163 506898 452205 507134
rect 452441 506898 452483 507134
rect 452163 506866 452483 506898
rect 454601 507454 454921 507486
rect 454601 507218 454643 507454
rect 454879 507218 454921 507454
rect 454601 507134 454921 507218
rect 454601 506898 454643 507134
rect 454879 506898 454921 507134
rect 454601 506866 454921 506898
rect 457039 507454 457359 507486
rect 457039 507218 457081 507454
rect 457317 507218 457359 507454
rect 457039 507134 457359 507218
rect 457039 506898 457081 507134
rect 457317 506898 457359 507134
rect 457039 506866 457359 506898
rect 450678 335310 451106 335370
rect 452394 490054 453014 500068
rect 452394 489818 452426 490054
rect 452662 489818 452746 490054
rect 452982 489818 453014 490054
rect 452394 489734 453014 489818
rect 452394 489498 452426 489734
rect 452662 489498 452746 489734
rect 452982 489498 453014 489734
rect 452394 454054 453014 489498
rect 452394 453818 452426 454054
rect 452662 453818 452746 454054
rect 452982 453818 453014 454054
rect 452394 453734 453014 453818
rect 452394 453498 452426 453734
rect 452662 453498 452746 453734
rect 452982 453498 453014 453734
rect 452394 418054 453014 453498
rect 452394 417818 452426 418054
rect 452662 417818 452746 418054
rect 452982 417818 453014 418054
rect 452394 417734 453014 417818
rect 452394 417498 452426 417734
rect 452662 417498 452746 417734
rect 452982 417498 453014 417734
rect 452394 382054 453014 417498
rect 452394 381818 452426 382054
rect 452662 381818 452746 382054
rect 452982 381818 453014 382054
rect 452394 381734 453014 381818
rect 452394 381498 452426 381734
rect 452662 381498 452746 381734
rect 452982 381498 453014 381734
rect 452394 346054 453014 381498
rect 456114 493774 456734 500068
rect 456114 493538 456146 493774
rect 456382 493538 456466 493774
rect 456702 493538 456734 493774
rect 456114 493454 456734 493538
rect 456114 493218 456146 493454
rect 456382 493218 456466 493454
rect 456702 493218 456734 493454
rect 456114 457774 456734 493218
rect 456114 457538 456146 457774
rect 456382 457538 456466 457774
rect 456702 457538 456734 457774
rect 456114 457454 456734 457538
rect 456114 457218 456146 457454
rect 456382 457218 456466 457454
rect 456702 457218 456734 457454
rect 456114 421774 456734 457218
rect 458958 428501 459018 647667
rect 459142 596869 459202 655691
rect 459139 596868 459205 596869
rect 459139 596804 459140 596868
rect 459204 596804 459205 596868
rect 459139 596803 459205 596804
rect 459510 518125 459570 670515
rect 459834 669073 460454 676938
rect 469794 704838 470414 711590
rect 469794 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 470414 704838
rect 469794 704518 470414 704602
rect 469794 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 470414 704518
rect 469794 687454 470414 704282
rect 469794 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 470414 687454
rect 469794 687134 470414 687218
rect 469794 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 470414 687134
rect 469794 669073 470414 686898
rect 473514 705798 474134 711590
rect 473514 705562 473546 705798
rect 473782 705562 473866 705798
rect 474102 705562 474134 705798
rect 473514 705478 474134 705562
rect 473514 705242 473546 705478
rect 473782 705242 473866 705478
rect 474102 705242 474134 705478
rect 473514 691174 474134 705242
rect 473514 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 474134 691174
rect 473514 690854 474134 690938
rect 473514 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 474134 690854
rect 473514 669073 474134 690618
rect 477234 706758 477854 711590
rect 477234 706522 477266 706758
rect 477502 706522 477586 706758
rect 477822 706522 477854 706758
rect 477234 706438 477854 706522
rect 477234 706202 477266 706438
rect 477502 706202 477586 706438
rect 477822 706202 477854 706438
rect 477234 694894 477854 706202
rect 477234 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 477854 694894
rect 477234 694574 477854 694658
rect 477234 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 477854 694574
rect 477234 669073 477854 694338
rect 480954 707718 481574 711590
rect 480954 707482 480986 707718
rect 481222 707482 481306 707718
rect 481542 707482 481574 707718
rect 480954 707398 481574 707482
rect 480954 707162 480986 707398
rect 481222 707162 481306 707398
rect 481542 707162 481574 707398
rect 480954 698614 481574 707162
rect 480954 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 481574 698614
rect 480954 698294 481574 698378
rect 480954 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 481574 698294
rect 480954 669073 481574 698058
rect 488394 709638 489014 711590
rect 488394 709402 488426 709638
rect 488662 709402 488746 709638
rect 488982 709402 489014 709638
rect 488394 709318 489014 709402
rect 488394 709082 488426 709318
rect 488662 709082 488746 709318
rect 488982 709082 489014 709318
rect 488394 670054 489014 709082
rect 488394 669818 488426 670054
rect 488662 669818 488746 670054
rect 488982 669818 489014 670054
rect 488394 669734 489014 669818
rect 488394 669498 488426 669734
rect 488662 669498 488746 669734
rect 488982 669498 489014 669734
rect 488394 669073 489014 669498
rect 492114 710598 492734 711590
rect 492114 710362 492146 710598
rect 492382 710362 492466 710598
rect 492702 710362 492734 710598
rect 492114 710278 492734 710362
rect 492114 710042 492146 710278
rect 492382 710042 492466 710278
rect 492702 710042 492734 710278
rect 492114 673774 492734 710042
rect 492114 673538 492146 673774
rect 492382 673538 492466 673774
rect 492702 673538 492734 673774
rect 492114 673454 492734 673538
rect 492114 673218 492146 673454
rect 492382 673218 492466 673454
rect 492702 673218 492734 673454
rect 492114 669073 492734 673218
rect 495834 711558 496454 711590
rect 495834 711322 495866 711558
rect 496102 711322 496186 711558
rect 496422 711322 496454 711558
rect 495834 711238 496454 711322
rect 495834 711002 495866 711238
rect 496102 711002 496186 711238
rect 496422 711002 496454 711238
rect 495834 677494 496454 711002
rect 495834 677258 495866 677494
rect 496102 677258 496186 677494
rect 496422 677258 496454 677494
rect 495834 677174 496454 677258
rect 495834 676938 495866 677174
rect 496102 676938 496186 677174
rect 496422 676938 496454 677174
rect 495834 669073 496454 676938
rect 505794 704838 506414 711590
rect 505794 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 506414 704838
rect 505794 704518 506414 704602
rect 505794 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 506414 704518
rect 505794 687454 506414 704282
rect 505794 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 506414 687454
rect 505794 687134 506414 687218
rect 505794 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 506414 687134
rect 505794 669073 506414 686898
rect 509514 705798 510134 711590
rect 509514 705562 509546 705798
rect 509782 705562 509866 705798
rect 510102 705562 510134 705798
rect 509514 705478 510134 705562
rect 509514 705242 509546 705478
rect 509782 705242 509866 705478
rect 510102 705242 510134 705478
rect 509514 691174 510134 705242
rect 509514 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 510134 691174
rect 509514 690854 510134 690938
rect 509514 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 510134 690854
rect 509514 669073 510134 690618
rect 513234 706758 513854 711590
rect 513234 706522 513266 706758
rect 513502 706522 513586 706758
rect 513822 706522 513854 706758
rect 513234 706438 513854 706522
rect 513234 706202 513266 706438
rect 513502 706202 513586 706438
rect 513822 706202 513854 706438
rect 513234 694894 513854 706202
rect 513234 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 513854 694894
rect 513234 694574 513854 694658
rect 513234 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 513854 694574
rect 513234 669073 513854 694338
rect 516954 707718 517574 711590
rect 516954 707482 516986 707718
rect 517222 707482 517306 707718
rect 517542 707482 517574 707718
rect 516954 707398 517574 707482
rect 516954 707162 516986 707398
rect 517222 707162 517306 707398
rect 517542 707162 517574 707398
rect 516954 698614 517574 707162
rect 516954 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 517574 698614
rect 516954 698294 517574 698378
rect 516954 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 517574 698294
rect 516954 669073 517574 698058
rect 520674 708678 521294 711590
rect 520674 708442 520706 708678
rect 520942 708442 521026 708678
rect 521262 708442 521294 708678
rect 520674 708358 521294 708442
rect 520674 708122 520706 708358
rect 520942 708122 521026 708358
rect 521262 708122 521294 708358
rect 520674 666334 521294 708122
rect 520674 666098 520706 666334
rect 520942 666098 521026 666334
rect 521262 666098 521294 666334
rect 520674 666014 521294 666098
rect 520674 665778 520706 666014
rect 520942 665778 521026 666014
rect 521262 665778 521294 666014
rect 479568 655174 479888 655206
rect 479568 654938 479610 655174
rect 479846 654938 479888 655174
rect 479568 654854 479888 654938
rect 479568 654618 479610 654854
rect 479846 654618 479888 654854
rect 479568 654586 479888 654618
rect 510288 655174 510608 655206
rect 510288 654938 510330 655174
rect 510566 654938 510608 655174
rect 510288 654854 510608 654938
rect 510288 654618 510330 654854
rect 510566 654618 510608 654854
rect 510288 654586 510608 654618
rect 464208 651454 464528 651486
rect 464208 651218 464250 651454
rect 464486 651218 464528 651454
rect 464208 651134 464528 651218
rect 464208 650898 464250 651134
rect 464486 650898 464528 651134
rect 464208 650866 464528 650898
rect 494928 651454 495248 651486
rect 494928 651218 494970 651454
rect 495206 651218 495248 651454
rect 494928 651134 495248 651218
rect 494928 650898 494970 651134
rect 495206 650898 495248 651134
rect 494928 650866 495248 650898
rect 520674 630334 521294 665778
rect 520674 630098 520706 630334
rect 520942 630098 521026 630334
rect 521262 630098 521294 630334
rect 520674 630014 521294 630098
rect 520674 629778 520706 630014
rect 520942 629778 521026 630014
rect 521262 629778 521294 630014
rect 479568 619174 479888 619206
rect 479568 618938 479610 619174
rect 479846 618938 479888 619174
rect 479568 618854 479888 618938
rect 479568 618618 479610 618854
rect 479846 618618 479888 618854
rect 479568 618586 479888 618618
rect 510288 619174 510608 619206
rect 510288 618938 510330 619174
rect 510566 618938 510608 619174
rect 510288 618854 510608 618938
rect 510288 618618 510330 618854
rect 510566 618618 510608 618854
rect 510288 618586 510608 618618
rect 464208 615454 464528 615486
rect 464208 615218 464250 615454
rect 464486 615218 464528 615454
rect 464208 615134 464528 615218
rect 464208 614898 464250 615134
rect 464486 614898 464528 615134
rect 464208 614866 464528 614898
rect 494928 615454 495248 615486
rect 494928 615218 494970 615454
rect 495206 615218 495248 615454
rect 494928 615134 495248 615218
rect 494928 614898 494970 615134
rect 495206 614898 495248 615134
rect 494928 614866 495248 614898
rect 459834 569494 460454 601103
rect 459834 569258 459866 569494
rect 460102 569258 460186 569494
rect 460422 569258 460454 569494
rect 459834 569174 460454 569258
rect 459834 568938 459866 569174
rect 460102 568938 460186 569174
rect 460422 568938 460454 569174
rect 459834 533494 460454 568938
rect 459834 533258 459866 533494
rect 460102 533258 460186 533494
rect 460422 533258 460454 533494
rect 459834 533174 460454 533258
rect 459834 532938 459866 533174
rect 460102 532938 460186 533174
rect 460422 532938 460454 533174
rect 459507 518124 459573 518125
rect 459507 518060 459508 518124
rect 459572 518060 459573 518124
rect 459507 518059 459573 518060
rect 459834 517884 460454 532938
rect 469794 579454 470414 601103
rect 472019 599588 472085 599589
rect 472019 599524 472020 599588
rect 472084 599524 472085 599588
rect 472019 599523 472085 599524
rect 469794 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 470414 579454
rect 469794 579134 470414 579218
rect 469794 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 470414 579134
rect 469794 543454 470414 578898
rect 469794 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 470414 543454
rect 469794 543134 470414 543218
rect 469794 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 470414 543134
rect 460696 511174 461016 511206
rect 460696 510938 460738 511174
rect 460974 510938 461016 511174
rect 460696 510854 461016 510938
rect 460696 510618 460738 510854
rect 460974 510618 461016 510854
rect 460696 510586 461016 510618
rect 459477 507454 459797 507486
rect 459477 507218 459519 507454
rect 459755 507218 459797 507454
rect 459477 507134 459797 507218
rect 459477 506898 459519 507134
rect 459755 506898 459797 507134
rect 459477 506866 459797 506898
rect 469794 507454 470414 542898
rect 469794 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 470414 507454
rect 469794 507134 470414 507218
rect 469794 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 470414 507134
rect 459834 497494 460454 500068
rect 459834 497258 459866 497494
rect 460102 497258 460186 497494
rect 460422 497258 460454 497494
rect 459834 497174 460454 497258
rect 459834 496938 459866 497174
rect 460102 496938 460186 497174
rect 460422 496938 460454 497174
rect 459834 461494 460454 496938
rect 459834 461258 459866 461494
rect 460102 461258 460186 461494
rect 460422 461258 460454 461494
rect 459834 461174 460454 461258
rect 459834 460938 459866 461174
rect 460102 460938 460186 461174
rect 460422 460938 460454 461174
rect 458955 428500 459021 428501
rect 458955 428436 458956 428500
rect 459020 428436 459021 428500
rect 458955 428435 459021 428436
rect 456114 421538 456146 421774
rect 456382 421538 456466 421774
rect 456702 421538 456734 421774
rect 456114 421454 456734 421538
rect 456114 421218 456146 421454
rect 456382 421218 456466 421454
rect 456702 421218 456734 421454
rect 456114 385774 456734 421218
rect 456114 385538 456146 385774
rect 456382 385538 456466 385774
rect 456702 385538 456734 385774
rect 456114 385454 456734 385538
rect 456114 385218 456146 385454
rect 456382 385218 456466 385454
rect 456702 385218 456734 385454
rect 454208 363454 454528 363486
rect 454208 363218 454250 363454
rect 454486 363218 454528 363454
rect 454208 363134 454528 363218
rect 454208 362898 454250 363134
rect 454486 362898 454528 363134
rect 454208 362866 454528 362898
rect 452394 345818 452426 346054
rect 452662 345818 452746 346054
rect 452982 345818 453014 346054
rect 452394 345734 453014 345818
rect 452394 345498 452426 345734
rect 452662 345498 452746 345734
rect 452982 345498 453014 345734
rect 450678 329221 450738 335310
rect 450675 329220 450741 329221
rect 450675 329156 450676 329220
rect 450740 329156 450741 329220
rect 450675 329155 450741 329156
rect 450491 328676 450557 328677
rect 450491 328612 450492 328676
rect 450556 328612 450557 328676
rect 450491 328611 450557 328612
rect 448674 306098 448706 306334
rect 448942 306098 449026 306334
rect 449262 306098 449294 306334
rect 448674 306014 449294 306098
rect 448674 305778 448706 306014
rect 448942 305778 449026 306014
rect 449262 305778 449294 306014
rect 448674 270334 449294 305778
rect 448674 270098 448706 270334
rect 448942 270098 449026 270334
rect 449262 270098 449294 270334
rect 448674 270014 449294 270098
rect 448674 269778 448706 270014
rect 448942 269778 449026 270014
rect 449262 269778 449294 270014
rect 448674 234334 449294 269778
rect 448674 234098 448706 234334
rect 448942 234098 449026 234334
rect 449262 234098 449294 234334
rect 448674 234014 449294 234098
rect 448674 233778 448706 234014
rect 448942 233778 449026 234014
rect 449262 233778 449294 234014
rect 448674 198334 449294 233778
rect 448674 198098 448706 198334
rect 448942 198098 449026 198334
rect 449262 198098 449294 198334
rect 448674 198014 449294 198098
rect 448674 197778 448706 198014
rect 448942 197778 449026 198014
rect 449262 197778 449294 198014
rect 448674 162334 449294 197778
rect 448674 162098 448706 162334
rect 448942 162098 449026 162334
rect 449262 162098 449294 162334
rect 448674 162014 449294 162098
rect 448674 161778 448706 162014
rect 448942 161778 449026 162014
rect 449262 161778 449294 162014
rect 429568 151174 429888 151206
rect 429568 150938 429610 151174
rect 429846 150938 429888 151174
rect 429568 150854 429888 150938
rect 429568 150618 429610 150854
rect 429846 150618 429888 150854
rect 429568 150586 429888 150618
rect 414208 147454 414528 147486
rect 414208 147218 414250 147454
rect 414486 147218 414528 147454
rect 414208 147134 414528 147218
rect 414208 146898 414250 147134
rect 414486 146898 414528 147134
rect 414208 146866 414528 146898
rect 444928 147454 445248 147486
rect 444928 147218 444970 147454
rect 445206 147218 445248 147454
rect 444928 147134 445248 147218
rect 444928 146898 444970 147134
rect 445206 146898 445248 147134
rect 444928 146866 445248 146898
rect 412674 126098 412706 126334
rect 412942 126098 413026 126334
rect 413262 126098 413294 126334
rect 412674 126014 413294 126098
rect 412674 125778 412706 126014
rect 412942 125778 413026 126014
rect 413262 125778 413294 126014
rect 412674 90334 413294 125778
rect 412674 90098 412706 90334
rect 412942 90098 413026 90334
rect 413262 90098 413294 90334
rect 412674 90014 413294 90098
rect 412674 89778 412706 90014
rect 412942 89778 413026 90014
rect 413262 89778 413294 90014
rect 412674 54334 413294 89778
rect 412674 54098 412706 54334
rect 412942 54098 413026 54334
rect 413262 54098 413294 54334
rect 412674 54014 413294 54098
rect 412674 53778 412706 54014
rect 412942 53778 413026 54014
rect 413262 53778 413294 54014
rect 412674 18334 413294 53778
rect 412674 18098 412706 18334
rect 412942 18098 413026 18334
rect 413262 18098 413294 18334
rect 412674 18014 413294 18098
rect 412674 17778 412706 18014
rect 412942 17778 413026 18014
rect 413262 17778 413294 18014
rect 412674 -4186 413294 17778
rect 412674 -4422 412706 -4186
rect 412942 -4422 413026 -4186
rect 413262 -4422 413294 -4186
rect 412674 -4506 413294 -4422
rect 412674 -4742 412706 -4506
rect 412942 -4742 413026 -4506
rect 413262 -4742 413294 -4506
rect 412674 -7654 413294 -4742
rect 416394 94054 417014 127767
rect 416394 93818 416426 94054
rect 416662 93818 416746 94054
rect 416982 93818 417014 94054
rect 416394 93734 417014 93818
rect 416394 93498 416426 93734
rect 416662 93498 416746 93734
rect 416982 93498 417014 93734
rect 416394 58054 417014 93498
rect 416394 57818 416426 58054
rect 416662 57818 416746 58054
rect 416982 57818 417014 58054
rect 416394 57734 417014 57818
rect 416394 57498 416426 57734
rect 416662 57498 416746 57734
rect 416982 57498 417014 57734
rect 416394 22054 417014 57498
rect 416394 21818 416426 22054
rect 416662 21818 416746 22054
rect 416982 21818 417014 22054
rect 416394 21734 417014 21818
rect 416394 21498 416426 21734
rect 416662 21498 416746 21734
rect 416982 21498 417014 21734
rect 416394 -5146 417014 21498
rect 416394 -5382 416426 -5146
rect 416662 -5382 416746 -5146
rect 416982 -5382 417014 -5146
rect 416394 -5466 417014 -5382
rect 416394 -5702 416426 -5466
rect 416662 -5702 416746 -5466
rect 416982 -5702 417014 -5466
rect 416394 -7654 417014 -5702
rect 420114 97774 420734 127767
rect 420114 97538 420146 97774
rect 420382 97538 420466 97774
rect 420702 97538 420734 97774
rect 420114 97454 420734 97538
rect 420114 97218 420146 97454
rect 420382 97218 420466 97454
rect 420702 97218 420734 97454
rect 420114 61774 420734 97218
rect 420114 61538 420146 61774
rect 420382 61538 420466 61774
rect 420702 61538 420734 61774
rect 420114 61454 420734 61538
rect 420114 61218 420146 61454
rect 420382 61218 420466 61454
rect 420702 61218 420734 61454
rect 420114 25774 420734 61218
rect 420114 25538 420146 25774
rect 420382 25538 420466 25774
rect 420702 25538 420734 25774
rect 420114 25454 420734 25538
rect 420114 25218 420146 25454
rect 420382 25218 420466 25454
rect 420702 25218 420734 25454
rect 420114 -6106 420734 25218
rect 420114 -6342 420146 -6106
rect 420382 -6342 420466 -6106
rect 420702 -6342 420734 -6106
rect 420114 -6426 420734 -6342
rect 420114 -6662 420146 -6426
rect 420382 -6662 420466 -6426
rect 420702 -6662 420734 -6426
rect 420114 -7654 420734 -6662
rect 423834 101494 424454 127767
rect 423834 101258 423866 101494
rect 424102 101258 424186 101494
rect 424422 101258 424454 101494
rect 423834 101174 424454 101258
rect 423834 100938 423866 101174
rect 424102 100938 424186 101174
rect 424422 100938 424454 101174
rect 423834 65494 424454 100938
rect 423834 65258 423866 65494
rect 424102 65258 424186 65494
rect 424422 65258 424454 65494
rect 423834 65174 424454 65258
rect 423834 64938 423866 65174
rect 424102 64938 424186 65174
rect 424422 64938 424454 65174
rect 423834 29494 424454 64938
rect 423834 29258 423866 29494
rect 424102 29258 424186 29494
rect 424422 29258 424454 29494
rect 423834 29174 424454 29258
rect 423834 28938 423866 29174
rect 424102 28938 424186 29174
rect 424422 28938 424454 29174
rect 423834 -7066 424454 28938
rect 423834 -7302 423866 -7066
rect 424102 -7302 424186 -7066
rect 424422 -7302 424454 -7066
rect 423834 -7386 424454 -7302
rect 423834 -7622 423866 -7386
rect 424102 -7622 424186 -7386
rect 424422 -7622 424454 -7386
rect 423834 -7654 424454 -7622
rect 433794 111454 434414 127767
rect 433794 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 434414 111454
rect 433794 111134 434414 111218
rect 433794 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 434414 111134
rect 433794 75454 434414 110898
rect 433794 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 434414 75454
rect 433794 75134 434414 75218
rect 433794 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 434414 75134
rect 433794 39454 434414 74898
rect 433794 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 434414 39454
rect 433794 39134 434414 39218
rect 433794 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 434414 39134
rect 433794 3454 434414 38898
rect 433794 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 434414 3454
rect 433794 3134 434414 3218
rect 433794 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 434414 3134
rect 433794 -346 434414 2898
rect 433794 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 434414 -346
rect 433794 -666 434414 -582
rect 433794 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 434414 -666
rect 433794 -7654 434414 -902
rect 437514 115174 438134 127767
rect 437514 114938 437546 115174
rect 437782 114938 437866 115174
rect 438102 114938 438134 115174
rect 437514 114854 438134 114938
rect 437514 114618 437546 114854
rect 437782 114618 437866 114854
rect 438102 114618 438134 114854
rect 437514 79174 438134 114618
rect 437514 78938 437546 79174
rect 437782 78938 437866 79174
rect 438102 78938 438134 79174
rect 437514 78854 438134 78938
rect 437514 78618 437546 78854
rect 437782 78618 437866 78854
rect 438102 78618 438134 78854
rect 437514 43174 438134 78618
rect 437514 42938 437546 43174
rect 437782 42938 437866 43174
rect 438102 42938 438134 43174
rect 437514 42854 438134 42938
rect 437514 42618 437546 42854
rect 437782 42618 437866 42854
rect 438102 42618 438134 42854
rect 437514 7174 438134 42618
rect 437514 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 438134 7174
rect 437514 6854 438134 6938
rect 437514 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 438134 6854
rect 437514 -1306 438134 6618
rect 437514 -1542 437546 -1306
rect 437782 -1542 437866 -1306
rect 438102 -1542 438134 -1306
rect 437514 -1626 438134 -1542
rect 437514 -1862 437546 -1626
rect 437782 -1862 437866 -1626
rect 438102 -1862 438134 -1626
rect 437514 -7654 438134 -1862
rect 441234 118894 441854 127767
rect 448674 126334 449294 161778
rect 448674 126098 448706 126334
rect 448942 126098 449026 126334
rect 449262 126098 449294 126334
rect 448674 126014 449294 126098
rect 448674 125778 448706 126014
rect 448942 125778 449026 126014
rect 449262 125778 449294 126014
rect 441234 118658 441266 118894
rect 441502 118658 441586 118894
rect 441822 118658 441854 118894
rect 441234 118574 441854 118658
rect 441234 118338 441266 118574
rect 441502 118338 441586 118574
rect 441822 118338 441854 118574
rect 441234 82894 441854 118338
rect 441234 82658 441266 82894
rect 441502 82658 441586 82894
rect 441822 82658 441854 82894
rect 441234 82574 441854 82658
rect 441234 82338 441266 82574
rect 441502 82338 441586 82574
rect 441822 82338 441854 82574
rect 441234 46894 441854 82338
rect 441234 46658 441266 46894
rect 441502 46658 441586 46894
rect 441822 46658 441854 46894
rect 441234 46574 441854 46658
rect 441234 46338 441266 46574
rect 441502 46338 441586 46574
rect 441822 46338 441854 46574
rect 441234 10894 441854 46338
rect 441234 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 441854 10894
rect 441234 10574 441854 10658
rect 441234 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 441854 10574
rect 441234 -2266 441854 10338
rect 441234 -2502 441266 -2266
rect 441502 -2502 441586 -2266
rect 441822 -2502 441854 -2266
rect 441234 -2586 441854 -2502
rect 441234 -2822 441266 -2586
rect 441502 -2822 441586 -2586
rect 441822 -2822 441854 -2586
rect 441234 -7654 441854 -2822
rect 444954 86614 445574 120068
rect 444954 86378 444986 86614
rect 445222 86378 445306 86614
rect 445542 86378 445574 86614
rect 444954 86294 445574 86378
rect 444954 86058 444986 86294
rect 445222 86058 445306 86294
rect 445542 86058 445574 86294
rect 444954 50614 445574 86058
rect 444954 50378 444986 50614
rect 445222 50378 445306 50614
rect 445542 50378 445574 50614
rect 444954 50294 445574 50378
rect 444954 50058 444986 50294
rect 445222 50058 445306 50294
rect 445542 50058 445574 50294
rect 444954 14614 445574 50058
rect 444954 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 445574 14614
rect 444954 14294 445574 14378
rect 444954 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 445574 14294
rect 444954 -3226 445574 14058
rect 444954 -3462 444986 -3226
rect 445222 -3462 445306 -3226
rect 445542 -3462 445574 -3226
rect 444954 -3546 445574 -3462
rect 444954 -3782 444986 -3546
rect 445222 -3782 445306 -3546
rect 445542 -3782 445574 -3546
rect 444954 -7654 445574 -3782
rect 448674 90334 449294 125778
rect 448674 90098 448706 90334
rect 448942 90098 449026 90334
rect 449262 90098 449294 90334
rect 448674 90014 449294 90098
rect 448674 89778 448706 90014
rect 448942 89778 449026 90014
rect 449262 89778 449294 90014
rect 448674 54334 449294 89778
rect 448674 54098 448706 54334
rect 448942 54098 449026 54334
rect 449262 54098 449294 54334
rect 448674 54014 449294 54098
rect 448674 53778 448706 54014
rect 448942 53778 449026 54014
rect 449262 53778 449294 54014
rect 448674 18334 449294 53778
rect 448674 18098 448706 18334
rect 448942 18098 449026 18334
rect 449262 18098 449294 18334
rect 448674 18014 449294 18098
rect 448674 17778 448706 18014
rect 448942 17778 449026 18014
rect 449262 17778 449294 18014
rect 448674 -4186 449294 17778
rect 448674 -4422 448706 -4186
rect 448942 -4422 449026 -4186
rect 449262 -4422 449294 -4186
rect 448674 -4506 449294 -4422
rect 448674 -4742 448706 -4506
rect 448942 -4742 449026 -4506
rect 449262 -4742 449294 -4506
rect 448674 -7654 449294 -4742
rect 452394 310054 453014 345498
rect 456114 349774 456734 385218
rect 456114 349538 456146 349774
rect 456382 349538 456466 349774
rect 456702 349538 456734 349774
rect 456114 349454 456734 349538
rect 456114 349218 456146 349454
rect 456382 349218 456466 349454
rect 456702 349218 456734 349454
rect 454208 327454 454528 327486
rect 454208 327218 454250 327454
rect 454486 327218 454528 327454
rect 454208 327134 454528 327218
rect 454208 326898 454250 327134
rect 454486 326898 454528 327134
rect 454208 326866 454528 326898
rect 452394 309818 452426 310054
rect 452662 309818 452746 310054
rect 452982 309818 453014 310054
rect 452394 309734 453014 309818
rect 452394 309498 452426 309734
rect 452662 309498 452746 309734
rect 452982 309498 453014 309734
rect 452394 274054 453014 309498
rect 452394 273818 452426 274054
rect 452662 273818 452746 274054
rect 452982 273818 453014 274054
rect 452394 273734 453014 273818
rect 452394 273498 452426 273734
rect 452662 273498 452746 273734
rect 452982 273498 453014 273734
rect 452394 238054 453014 273498
rect 452394 237818 452426 238054
rect 452662 237818 452746 238054
rect 452982 237818 453014 238054
rect 452394 237734 453014 237818
rect 452394 237498 452426 237734
rect 452662 237498 452746 237734
rect 452982 237498 453014 237734
rect 452394 202054 453014 237498
rect 452394 201818 452426 202054
rect 452662 201818 452746 202054
rect 452982 201818 453014 202054
rect 452394 201734 453014 201818
rect 452394 201498 452426 201734
rect 452662 201498 452746 201734
rect 452982 201498 453014 201734
rect 452394 166054 453014 201498
rect 452394 165818 452426 166054
rect 452662 165818 452746 166054
rect 452982 165818 453014 166054
rect 452394 165734 453014 165818
rect 452394 165498 452426 165734
rect 452662 165498 452746 165734
rect 452982 165498 453014 165734
rect 452394 130054 453014 165498
rect 452394 129818 452426 130054
rect 452662 129818 452746 130054
rect 452982 129818 453014 130054
rect 452394 129734 453014 129818
rect 452394 129498 452426 129734
rect 452662 129498 452746 129734
rect 452982 129498 453014 129734
rect 452394 94054 453014 129498
rect 452394 93818 452426 94054
rect 452662 93818 452746 94054
rect 452982 93818 453014 94054
rect 452394 93734 453014 93818
rect 452394 93498 452426 93734
rect 452662 93498 452746 93734
rect 452982 93498 453014 93734
rect 452394 58054 453014 93498
rect 452394 57818 452426 58054
rect 452662 57818 452746 58054
rect 452982 57818 453014 58054
rect 452394 57734 453014 57818
rect 452394 57498 452426 57734
rect 452662 57498 452746 57734
rect 452982 57498 453014 57734
rect 452394 22054 453014 57498
rect 452394 21818 452426 22054
rect 452662 21818 452746 22054
rect 452982 21818 453014 22054
rect 452394 21734 453014 21818
rect 452394 21498 452426 21734
rect 452662 21498 452746 21734
rect 452982 21498 453014 21734
rect 452394 -5146 453014 21498
rect 452394 -5382 452426 -5146
rect 452662 -5382 452746 -5146
rect 452982 -5382 453014 -5146
rect 452394 -5466 453014 -5382
rect 452394 -5702 452426 -5466
rect 452662 -5702 452746 -5466
rect 452982 -5702 453014 -5466
rect 452394 -7654 453014 -5702
rect 456114 313774 456734 349218
rect 459834 425494 460454 460938
rect 459834 425258 459866 425494
rect 460102 425258 460186 425494
rect 460422 425258 460454 425494
rect 459834 425174 460454 425258
rect 459834 424938 459866 425174
rect 460102 424938 460186 425174
rect 460422 424938 460454 425174
rect 459834 389494 460454 424938
rect 459834 389258 459866 389494
rect 460102 389258 460186 389494
rect 460422 389258 460454 389494
rect 459834 389174 460454 389258
rect 459834 388938 459866 389174
rect 460102 388938 460186 389174
rect 460422 388938 460454 389174
rect 459834 353494 460454 388938
rect 469794 471454 470414 506898
rect 469794 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 470414 471454
rect 469794 471134 470414 471218
rect 469794 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 470414 471134
rect 469794 435454 470414 470898
rect 469794 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 470414 435454
rect 469794 435134 470414 435218
rect 469794 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 470414 435134
rect 469794 399454 470414 434898
rect 469794 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 470414 399454
rect 469794 399134 470414 399218
rect 469794 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 470414 399134
rect 469794 385580 470414 398898
rect 472022 388925 472082 599523
rect 473514 583174 474134 601103
rect 473514 582938 473546 583174
rect 473782 582938 473866 583174
rect 474102 582938 474134 583174
rect 473514 582854 474134 582938
rect 473514 582618 473546 582854
rect 473782 582618 473866 582854
rect 474102 582618 474134 582854
rect 473514 547174 474134 582618
rect 473514 546938 473546 547174
rect 473782 546938 473866 547174
rect 474102 546938 474134 547174
rect 473514 546854 474134 546938
rect 473514 546618 473546 546854
rect 473782 546618 473866 546854
rect 474102 546618 474134 546854
rect 472203 518260 472269 518261
rect 472203 518196 472204 518260
rect 472268 518196 472269 518260
rect 472203 518195 472269 518196
rect 472206 389061 472266 518195
rect 473514 511174 474134 546618
rect 477234 586894 477854 601103
rect 478827 596868 478893 596869
rect 478827 596804 478828 596868
rect 478892 596804 478893 596868
rect 478827 596803 478893 596804
rect 477234 586658 477266 586894
rect 477502 586658 477586 586894
rect 477822 586658 477854 586894
rect 477234 586574 477854 586658
rect 477234 586338 477266 586574
rect 477502 586338 477586 586574
rect 477822 586338 477854 586574
rect 477234 550894 477854 586338
rect 477234 550658 477266 550894
rect 477502 550658 477586 550894
rect 477822 550658 477854 550894
rect 477234 550574 477854 550658
rect 477234 550338 477266 550574
rect 477502 550338 477586 550574
rect 477822 550338 477854 550574
rect 474411 543012 474477 543013
rect 474411 542948 474412 543012
rect 474476 542948 474477 543012
rect 474411 542947 474477 542948
rect 473514 510938 473546 511174
rect 473782 510938 473866 511174
rect 474102 510938 474134 511174
rect 473514 510854 474134 510938
rect 473514 510618 473546 510854
rect 473782 510618 473866 510854
rect 474102 510618 474134 510854
rect 473514 475174 474134 510618
rect 473514 474938 473546 475174
rect 473782 474938 473866 475174
rect 474102 474938 474134 475174
rect 473514 474854 474134 474938
rect 473514 474618 473546 474854
rect 473782 474618 473866 474854
rect 474102 474618 474134 474854
rect 473514 453692 474134 474618
rect 473416 435454 473736 435486
rect 473416 435218 473458 435454
rect 473694 435218 473736 435454
rect 473416 435134 473736 435218
rect 473416 434898 473458 435134
rect 473694 434898 473736 435134
rect 473416 434866 473736 434898
rect 474414 389061 474474 542947
rect 477234 514894 477854 550338
rect 477234 514658 477266 514894
rect 477502 514658 477586 514894
rect 477822 514658 477854 514894
rect 477234 514574 477854 514658
rect 477234 514338 477266 514574
rect 477502 514338 477586 514574
rect 477822 514338 477854 514574
rect 477234 478894 477854 514338
rect 477234 478658 477266 478894
rect 477502 478658 477586 478894
rect 477822 478658 477854 478894
rect 477234 478574 477854 478658
rect 477234 478338 477266 478574
rect 477502 478338 477586 478574
rect 477822 478338 477854 478574
rect 477234 442894 477854 478338
rect 477234 442658 477266 442894
rect 477502 442658 477586 442894
rect 477822 442658 477854 442894
rect 477234 442574 477854 442658
rect 477234 442338 477266 442574
rect 477502 442338 477586 442574
rect 477822 442338 477854 442574
rect 475888 439174 476208 439206
rect 475888 438938 475930 439174
rect 476166 438938 476208 439174
rect 475888 438854 476208 438938
rect 475888 438618 475930 438854
rect 476166 438618 476208 438854
rect 475888 438586 476208 438618
rect 477234 406894 477854 442338
rect 478361 435454 478681 435486
rect 478361 435218 478403 435454
rect 478639 435218 478681 435454
rect 478361 435134 478681 435218
rect 478361 434898 478403 435134
rect 478639 434898 478681 435134
rect 478361 434866 478681 434898
rect 477234 406658 477266 406894
rect 477502 406658 477586 406894
rect 477822 406658 477854 406894
rect 477234 406574 477854 406658
rect 477234 406338 477266 406574
rect 477502 406338 477586 406574
rect 477822 406338 477854 406574
rect 472203 389060 472269 389061
rect 472203 388996 472204 389060
rect 472268 388996 472269 389060
rect 472203 388995 472269 388996
rect 474411 389060 474477 389061
rect 474411 388996 474412 389060
rect 474476 388996 474477 389060
rect 474411 388995 474477 388996
rect 472019 388924 472085 388925
rect 472019 388860 472020 388924
rect 472084 388860 472085 388924
rect 472019 388859 472085 388860
rect 477234 385225 477854 406338
rect 478830 389061 478890 596803
rect 480954 590614 481574 601103
rect 480954 590378 480986 590614
rect 481222 590378 481306 590614
rect 481542 590378 481574 590614
rect 480954 590294 481574 590378
rect 480954 590058 480986 590294
rect 481222 590058 481306 590294
rect 481542 590058 481574 590294
rect 480954 554614 481574 590058
rect 480954 554378 480986 554614
rect 481222 554378 481306 554614
rect 481542 554378 481574 554614
rect 480954 554294 481574 554378
rect 480954 554058 480986 554294
rect 481222 554058 481306 554294
rect 481542 554058 481574 554294
rect 480954 518614 481574 554058
rect 480954 518378 480986 518614
rect 481222 518378 481306 518614
rect 481542 518378 481574 518614
rect 480954 518294 481574 518378
rect 480954 518058 480986 518294
rect 481222 518058 481306 518294
rect 481542 518058 481574 518294
rect 480954 482614 481574 518058
rect 484674 594334 485294 601103
rect 484674 594098 484706 594334
rect 484942 594098 485026 594334
rect 485262 594098 485294 594334
rect 484674 594014 485294 594098
rect 484674 593778 484706 594014
rect 484942 593778 485026 594014
rect 485262 593778 485294 594014
rect 484674 558334 485294 593778
rect 484674 558098 484706 558334
rect 484942 558098 485026 558334
rect 485262 558098 485294 558334
rect 484674 558014 485294 558098
rect 484674 557778 484706 558014
rect 484942 557778 485026 558014
rect 485262 557778 485294 558014
rect 484674 522334 485294 557778
rect 484674 522098 484706 522334
rect 484942 522098 485026 522334
rect 485262 522098 485294 522334
rect 484674 522014 485294 522098
rect 484674 521778 484706 522014
rect 484942 521778 485026 522014
rect 485262 521778 485294 522014
rect 484674 517884 485294 521778
rect 488394 598054 489014 601103
rect 488394 597818 488426 598054
rect 488662 597818 488746 598054
rect 488982 597818 489014 598054
rect 488394 597734 489014 597818
rect 488394 597498 488426 597734
rect 488662 597498 488746 597734
rect 488982 597498 489014 597734
rect 488394 562054 489014 597498
rect 488394 561818 488426 562054
rect 488662 561818 488746 562054
rect 488982 561818 489014 562054
rect 488394 561734 489014 561818
rect 488394 561498 488426 561734
rect 488662 561498 488746 561734
rect 488982 561498 489014 561734
rect 488394 526054 489014 561498
rect 488394 525818 488426 526054
rect 488662 525818 488746 526054
rect 488982 525818 489014 526054
rect 488394 525734 489014 525818
rect 488394 525498 488426 525734
rect 488662 525498 488746 525734
rect 488982 525498 489014 525734
rect 488394 517884 489014 525498
rect 492114 565774 492734 601103
rect 492114 565538 492146 565774
rect 492382 565538 492466 565774
rect 492702 565538 492734 565774
rect 492114 565454 492734 565538
rect 492114 565218 492146 565454
rect 492382 565218 492466 565454
rect 492702 565218 492734 565454
rect 492114 529774 492734 565218
rect 492114 529538 492146 529774
rect 492382 529538 492466 529774
rect 492702 529538 492734 529774
rect 492114 529454 492734 529538
rect 492114 529218 492146 529454
rect 492382 529218 492466 529454
rect 492702 529218 492734 529454
rect 482691 517580 482757 517581
rect 482691 517516 482692 517580
rect 482756 517516 482757 517580
rect 482691 517515 482757 517516
rect 482163 507454 482483 507486
rect 482163 507218 482205 507454
rect 482441 507218 482483 507454
rect 482163 507134 482483 507218
rect 482163 506898 482205 507134
rect 482441 506898 482483 507134
rect 482163 506866 482483 506898
rect 480954 482378 480986 482614
rect 481222 482378 481306 482614
rect 481542 482378 481574 482614
rect 480954 482294 481574 482378
rect 480954 482058 480986 482294
rect 481222 482058 481306 482294
rect 481542 482058 481574 482294
rect 480954 453692 481574 482058
rect 482694 462909 482754 517515
rect 483382 511174 483702 511206
rect 483382 510938 483424 511174
rect 483660 510938 483702 511174
rect 483382 510854 483702 510938
rect 483382 510618 483424 510854
rect 483660 510618 483702 510854
rect 483382 510586 483702 510618
rect 485820 511174 486140 511206
rect 485820 510938 485862 511174
rect 486098 510938 486140 511174
rect 485820 510854 486140 510938
rect 485820 510618 485862 510854
rect 486098 510618 486140 510854
rect 485820 510586 486140 510618
rect 488258 511174 488578 511206
rect 488258 510938 488300 511174
rect 488536 510938 488578 511174
rect 488258 510854 488578 510938
rect 488258 510618 488300 510854
rect 488536 510618 488578 510854
rect 488258 510586 488578 510618
rect 490696 511174 491016 511206
rect 490696 510938 490738 511174
rect 490974 510938 491016 511174
rect 490696 510854 491016 510938
rect 490696 510618 490738 510854
rect 490974 510618 491016 510854
rect 490696 510586 491016 510618
rect 484601 507454 484921 507486
rect 484601 507218 484643 507454
rect 484879 507218 484921 507454
rect 484601 507134 484921 507218
rect 484601 506898 484643 507134
rect 484879 506898 484921 507134
rect 484601 506866 484921 506898
rect 487039 507454 487359 507486
rect 487039 507218 487081 507454
rect 487317 507218 487359 507454
rect 487039 507134 487359 507218
rect 487039 506898 487081 507134
rect 487317 506898 487359 507134
rect 487039 506866 487359 506898
rect 489477 507454 489797 507486
rect 489477 507218 489519 507454
rect 489755 507218 489797 507454
rect 489477 507134 489797 507218
rect 489477 506898 489519 507134
rect 489755 506898 489797 507134
rect 489477 506866 489797 506898
rect 484674 486334 485294 500068
rect 484674 486098 484706 486334
rect 484942 486098 485026 486334
rect 485262 486098 485294 486334
rect 484674 486014 485294 486098
rect 484674 485778 484706 486014
rect 484942 485778 485026 486014
rect 485262 485778 485294 486014
rect 482691 462908 482757 462909
rect 482691 462844 482692 462908
rect 482756 462844 482757 462908
rect 482691 462843 482757 462844
rect 484674 450334 485294 485778
rect 488394 490054 489014 500068
rect 489315 496908 489381 496909
rect 489315 496844 489316 496908
rect 489380 496844 489381 496908
rect 489315 496843 489381 496844
rect 488394 489818 488426 490054
rect 488662 489818 488746 490054
rect 488982 489818 489014 490054
rect 488394 489734 489014 489818
rect 488394 489498 488426 489734
rect 488662 489498 488746 489734
rect 488982 489498 489014 489734
rect 488394 454007 489014 489498
rect 488394 453771 488426 454007
rect 488662 453771 488746 454007
rect 488982 453771 489014 454007
rect 488394 453692 489014 453771
rect 484674 450098 484706 450334
rect 484942 450098 485026 450334
rect 485262 450098 485294 450334
rect 484674 450014 485294 450098
rect 484674 449778 484706 450014
rect 484942 449778 485026 450014
rect 485262 449778 485294 450014
rect 480833 439174 481153 439206
rect 480833 438938 480875 439174
rect 481111 438938 481153 439174
rect 480833 438854 481153 438938
rect 480833 438618 480875 438854
rect 481111 438618 481153 438854
rect 480833 438586 481153 438618
rect 483306 435454 483626 435486
rect 483306 435218 483348 435454
rect 483584 435218 483626 435454
rect 483306 435134 483626 435218
rect 483306 434898 483348 435134
rect 483584 434898 483626 435134
rect 483306 434866 483626 434898
rect 484674 414334 485294 449778
rect 485778 439174 486098 439206
rect 485778 438938 485820 439174
rect 486056 438938 486098 439174
rect 485778 438854 486098 438938
rect 485778 438618 485820 438854
rect 486056 438618 486098 438854
rect 485778 438586 486098 438618
rect 488251 435454 488571 435486
rect 488251 435218 488293 435454
rect 488529 435218 488571 435454
rect 488251 435134 488571 435218
rect 488251 434898 488293 435134
rect 488529 434898 488571 435134
rect 488251 434866 488571 434898
rect 484674 414098 484706 414334
rect 484942 414098 485026 414334
rect 485262 414098 485294 414334
rect 484674 414014 485294 414098
rect 484674 413778 484706 414014
rect 484942 413778 485026 414014
rect 485262 413778 485294 414014
rect 478827 389060 478893 389061
rect 478827 388996 478828 389060
rect 478892 388996 478893 389060
rect 478827 388995 478893 388996
rect 484674 385580 485294 413778
rect 489318 387021 489378 496843
rect 492114 493774 492734 529218
rect 492114 493538 492146 493774
rect 492382 493538 492466 493774
rect 492702 493538 492734 493774
rect 492114 493454 492734 493538
rect 492114 493218 492146 493454
rect 492382 493218 492466 493454
rect 492702 493218 492734 493454
rect 492114 457774 492734 493218
rect 492114 457538 492146 457774
rect 492382 457538 492466 457774
rect 492702 457538 492734 457774
rect 492114 457454 492734 457538
rect 492114 457218 492146 457454
rect 492382 457218 492466 457454
rect 492702 457218 492734 457454
rect 490723 439174 491043 439206
rect 490723 438938 490765 439174
rect 491001 438938 491043 439174
rect 490723 438854 491043 438938
rect 490723 438618 490765 438854
rect 491001 438618 491043 438854
rect 490723 438586 491043 438618
rect 492114 421774 492734 457218
rect 492114 421538 492146 421774
rect 492382 421538 492466 421774
rect 492702 421538 492734 421774
rect 492114 421454 492734 421538
rect 492114 421218 492146 421454
rect 492382 421218 492466 421454
rect 492702 421218 492734 421454
rect 489315 387020 489381 387021
rect 489315 386956 489316 387020
rect 489380 386956 489381 387020
rect 489315 386955 489381 386956
rect 492114 385225 492734 421218
rect 495834 569494 496454 601103
rect 495834 569258 495866 569494
rect 496102 569258 496186 569494
rect 496422 569258 496454 569494
rect 495834 569174 496454 569258
rect 495834 568938 495866 569174
rect 496102 568938 496186 569174
rect 496422 568938 496454 569174
rect 495834 533494 496454 568938
rect 495834 533258 495866 533494
rect 496102 533258 496186 533494
rect 496422 533258 496454 533494
rect 495834 533174 496454 533258
rect 495834 532938 495866 533174
rect 496102 532938 496186 533174
rect 496422 532938 496454 533174
rect 495834 497494 496454 532938
rect 495834 497258 495866 497494
rect 496102 497258 496186 497494
rect 496422 497258 496454 497494
rect 495834 497174 496454 497258
rect 495834 496938 495866 497174
rect 496102 496938 496186 497174
rect 496422 496938 496454 497174
rect 495834 461494 496454 496938
rect 495834 461258 495866 461494
rect 496102 461258 496186 461494
rect 496422 461258 496454 461494
rect 495834 461174 496454 461258
rect 495834 460938 495866 461174
rect 496102 460938 496186 461174
rect 496422 460938 496454 461174
rect 495834 425494 496454 460938
rect 495834 425258 495866 425494
rect 496102 425258 496186 425494
rect 496422 425258 496454 425494
rect 495834 425174 496454 425258
rect 495834 424938 495866 425174
rect 496102 424938 496186 425174
rect 496422 424938 496454 425174
rect 495834 389494 496454 424938
rect 495834 389258 495866 389494
rect 496102 389258 496186 389494
rect 496422 389258 496454 389494
rect 495834 389174 496454 389258
rect 495834 388938 495866 389174
rect 496102 388938 496186 389174
rect 496422 388938 496454 389174
rect 469568 367174 469888 367206
rect 469568 366938 469610 367174
rect 469846 366938 469888 367174
rect 469568 366854 469888 366938
rect 469568 366618 469610 366854
rect 469846 366618 469888 366854
rect 469568 366586 469888 366618
rect 484928 363454 485248 363486
rect 484928 363218 484970 363454
rect 485206 363218 485248 363454
rect 484928 363134 485248 363218
rect 484928 362898 484970 363134
rect 485206 362898 485248 363134
rect 484928 362866 485248 362898
rect 459834 353258 459866 353494
rect 460102 353258 460186 353494
rect 460422 353258 460454 353494
rect 459834 353174 460454 353258
rect 459834 352938 459866 353174
rect 460102 352938 460186 353174
rect 460422 352938 460454 353174
rect 458771 320788 458837 320789
rect 458771 320724 458772 320788
rect 458836 320724 458837 320788
rect 458771 320723 458837 320724
rect 456114 313538 456146 313774
rect 456382 313538 456466 313774
rect 456702 313538 456734 313774
rect 456114 313454 456734 313538
rect 456114 313218 456146 313454
rect 456382 313218 456466 313454
rect 456702 313218 456734 313454
rect 456114 277774 456734 313218
rect 456114 277538 456146 277774
rect 456382 277538 456466 277774
rect 456702 277538 456734 277774
rect 456114 277454 456734 277538
rect 456114 277218 456146 277454
rect 456382 277218 456466 277454
rect 456702 277218 456734 277454
rect 456114 241774 456734 277218
rect 456114 241538 456146 241774
rect 456382 241538 456466 241774
rect 456702 241538 456734 241774
rect 456114 241454 456734 241538
rect 456114 241218 456146 241454
rect 456382 241218 456466 241454
rect 456702 241218 456734 241454
rect 456114 205774 456734 241218
rect 456114 205538 456146 205774
rect 456382 205538 456466 205774
rect 456702 205538 456734 205774
rect 456114 205454 456734 205538
rect 456114 205218 456146 205454
rect 456382 205218 456466 205454
rect 456702 205218 456734 205454
rect 456114 169774 456734 205218
rect 456114 169538 456146 169774
rect 456382 169538 456466 169774
rect 456702 169538 456734 169774
rect 456114 169454 456734 169538
rect 456114 169218 456146 169454
rect 456382 169218 456466 169454
rect 456702 169218 456734 169454
rect 456114 133774 456734 169218
rect 456114 133538 456146 133774
rect 456382 133538 456466 133774
rect 456702 133538 456734 133774
rect 456114 133454 456734 133538
rect 456114 133218 456146 133454
rect 456382 133218 456466 133454
rect 456702 133218 456734 133454
rect 456114 97774 456734 133218
rect 456114 97538 456146 97774
rect 456382 97538 456466 97774
rect 456702 97538 456734 97774
rect 456114 97454 456734 97538
rect 456114 97218 456146 97454
rect 456382 97218 456466 97454
rect 456702 97218 456734 97454
rect 456114 61774 456734 97218
rect 456114 61538 456146 61774
rect 456382 61538 456466 61774
rect 456702 61538 456734 61774
rect 456114 61454 456734 61538
rect 456114 61218 456146 61454
rect 456382 61218 456466 61454
rect 456702 61218 456734 61454
rect 456114 25774 456734 61218
rect 456114 25538 456146 25774
rect 456382 25538 456466 25774
rect 456702 25538 456734 25774
rect 456114 25454 456734 25538
rect 456114 25218 456146 25454
rect 456382 25218 456466 25454
rect 456702 25218 456734 25454
rect 456114 -6106 456734 25218
rect 458774 3365 458834 320723
rect 459834 317494 460454 352938
rect 495834 353494 496454 388938
rect 505794 579454 506414 601103
rect 505794 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 506414 579454
rect 505794 579134 506414 579218
rect 505794 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 506414 579134
rect 505794 543454 506414 578898
rect 505794 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 506414 543454
rect 505794 543134 506414 543218
rect 505794 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 506414 543134
rect 505794 507454 506414 542898
rect 505794 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 506414 507454
rect 505794 507134 506414 507218
rect 505794 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 506414 507134
rect 505794 471454 506414 506898
rect 505794 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 506414 471454
rect 505794 471134 506414 471218
rect 505794 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 506414 471134
rect 505794 435454 506414 470898
rect 505794 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 506414 435454
rect 505794 435134 506414 435218
rect 505794 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 506414 435134
rect 505794 399454 506414 434898
rect 505794 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 506414 399454
rect 505794 399134 506414 399218
rect 505794 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 506414 399134
rect 500288 367174 500608 367206
rect 500288 366938 500330 367174
rect 500566 366938 500608 367174
rect 500288 366854 500608 366938
rect 500288 366618 500330 366854
rect 500566 366618 500608 366854
rect 500288 366586 500608 366618
rect 495834 353258 495866 353494
rect 496102 353258 496186 353494
rect 496422 353258 496454 353494
rect 495834 353174 496454 353258
rect 495834 352938 495866 353174
rect 496102 352938 496186 353174
rect 496422 352938 496454 353174
rect 469568 331174 469888 331206
rect 469568 330938 469610 331174
rect 469846 330938 469888 331174
rect 469568 330854 469888 330938
rect 469568 330618 469610 330854
rect 469846 330618 469888 330854
rect 469568 330586 469888 330618
rect 484928 327454 485248 327486
rect 484928 327218 484970 327454
rect 485206 327218 485248 327454
rect 484928 327134 485248 327218
rect 484928 326898 484970 327134
rect 485206 326898 485248 327134
rect 484928 326866 485248 326898
rect 459834 317258 459866 317494
rect 460102 317258 460186 317494
rect 460422 317258 460454 317494
rect 459834 317174 460454 317258
rect 459834 316938 459866 317174
rect 460102 316938 460186 317174
rect 460422 316938 460454 317174
rect 459834 281494 460454 316938
rect 459834 281258 459866 281494
rect 460102 281258 460186 281494
rect 460422 281258 460454 281494
rect 459834 281174 460454 281258
rect 459834 280938 459866 281174
rect 460102 280938 460186 281174
rect 460422 280938 460454 281174
rect 459834 245494 460454 280938
rect 477234 298894 477854 322287
rect 477234 298658 477266 298894
rect 477502 298658 477586 298894
rect 477822 298658 477854 298894
rect 477234 298574 477854 298658
rect 477234 298338 477266 298574
rect 477502 298338 477586 298574
rect 477822 298338 477854 298574
rect 477234 262894 477854 298338
rect 477234 262658 477266 262894
rect 477502 262658 477586 262894
rect 477822 262658 477854 262894
rect 477234 262574 477854 262658
rect 477234 262338 477266 262574
rect 477502 262338 477586 262574
rect 477822 262338 477854 262574
rect 477234 259417 477854 262338
rect 480954 302614 481574 322287
rect 480954 302378 480986 302614
rect 481222 302378 481306 302614
rect 481542 302378 481574 302614
rect 480954 302294 481574 302378
rect 480954 302058 480986 302294
rect 481222 302058 481306 302294
rect 481542 302058 481574 302294
rect 480954 266614 481574 302058
rect 480954 266378 480986 266614
rect 481222 266378 481306 266614
rect 481542 266378 481574 266614
rect 480954 266294 481574 266378
rect 480954 266058 480986 266294
rect 481222 266058 481306 266294
rect 481542 266058 481574 266294
rect 480954 259417 481574 266058
rect 484674 306334 485294 322068
rect 484674 306098 484706 306334
rect 484942 306098 485026 306334
rect 485262 306098 485294 306334
rect 484674 306014 485294 306098
rect 484674 305778 484706 306014
rect 484942 305778 485026 306014
rect 485262 305778 485294 306014
rect 484674 270334 485294 305778
rect 484674 270098 484706 270334
rect 484942 270098 485026 270334
rect 485262 270098 485294 270334
rect 484674 270014 485294 270098
rect 484674 269778 484706 270014
rect 484942 269778 485026 270014
rect 485262 269778 485294 270014
rect 484674 259417 485294 269778
rect 488394 310054 489014 322287
rect 488394 309818 488426 310054
rect 488662 309818 488746 310054
rect 488982 309818 489014 310054
rect 488394 309734 489014 309818
rect 488394 309498 488426 309734
rect 488662 309498 488746 309734
rect 488982 309498 489014 309734
rect 488394 274054 489014 309498
rect 488394 273818 488426 274054
rect 488662 273818 488746 274054
rect 488982 273818 489014 274054
rect 488394 273734 489014 273818
rect 488394 273498 488426 273734
rect 488662 273498 488746 273734
rect 488982 273498 489014 273734
rect 488394 259417 489014 273498
rect 492114 313774 492734 322287
rect 492114 313538 492146 313774
rect 492382 313538 492466 313774
rect 492702 313538 492734 313774
rect 492114 313454 492734 313538
rect 492114 313218 492146 313454
rect 492382 313218 492466 313454
rect 492702 313218 492734 313454
rect 492114 277774 492734 313218
rect 492114 277538 492146 277774
rect 492382 277538 492466 277774
rect 492702 277538 492734 277774
rect 492114 277454 492734 277538
rect 492114 277218 492146 277454
rect 492382 277218 492466 277454
rect 492702 277218 492734 277454
rect 492114 259417 492734 277218
rect 495834 317494 496454 352938
rect 505794 363454 506414 398898
rect 505794 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 506414 363454
rect 505794 363134 506414 363218
rect 505794 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 506414 363134
rect 500288 331174 500608 331206
rect 500288 330938 500330 331174
rect 500566 330938 500608 331174
rect 500288 330854 500608 330938
rect 500288 330618 500330 330854
rect 500566 330618 500608 330854
rect 500288 330586 500608 330618
rect 495834 317258 495866 317494
rect 496102 317258 496186 317494
rect 496422 317258 496454 317494
rect 495834 317174 496454 317258
rect 495834 316938 495866 317174
rect 496102 316938 496186 317174
rect 496422 316938 496454 317174
rect 495834 281494 496454 316938
rect 495834 281258 495866 281494
rect 496102 281258 496186 281494
rect 496422 281258 496454 281494
rect 495834 281174 496454 281258
rect 495834 280938 495866 281174
rect 496102 280938 496186 281174
rect 496422 280938 496454 281174
rect 495834 259417 496454 280938
rect 505794 327454 506414 362898
rect 505794 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 506414 327454
rect 505794 327134 506414 327218
rect 505794 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 506414 327134
rect 505794 291454 506414 326898
rect 505794 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 506414 291454
rect 505794 291134 506414 291218
rect 505794 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 506414 291134
rect 505794 259417 506414 290898
rect 509514 583174 510134 601103
rect 509514 582938 509546 583174
rect 509782 582938 509866 583174
rect 510102 582938 510134 583174
rect 509514 582854 510134 582938
rect 509514 582618 509546 582854
rect 509782 582618 509866 582854
rect 510102 582618 510134 582854
rect 509514 547174 510134 582618
rect 509514 546938 509546 547174
rect 509782 546938 509866 547174
rect 510102 546938 510134 547174
rect 509514 546854 510134 546938
rect 509514 546618 509546 546854
rect 509782 546618 509866 546854
rect 510102 546618 510134 546854
rect 509514 511174 510134 546618
rect 509514 510938 509546 511174
rect 509782 510938 509866 511174
rect 510102 510938 510134 511174
rect 509514 510854 510134 510938
rect 509514 510618 509546 510854
rect 509782 510618 509866 510854
rect 510102 510618 510134 510854
rect 509514 475174 510134 510618
rect 509514 474938 509546 475174
rect 509782 474938 509866 475174
rect 510102 474938 510134 475174
rect 509514 474854 510134 474938
rect 509514 474618 509546 474854
rect 509782 474618 509866 474854
rect 510102 474618 510134 474854
rect 509514 439174 510134 474618
rect 509514 438938 509546 439174
rect 509782 438938 509866 439174
rect 510102 438938 510134 439174
rect 509514 438854 510134 438938
rect 509514 438618 509546 438854
rect 509782 438618 509866 438854
rect 510102 438618 510134 438854
rect 509514 403174 510134 438618
rect 509514 402938 509546 403174
rect 509782 402938 509866 403174
rect 510102 402938 510134 403174
rect 509514 402854 510134 402938
rect 509514 402618 509546 402854
rect 509782 402618 509866 402854
rect 510102 402618 510134 402854
rect 509514 367174 510134 402618
rect 509514 366938 509546 367174
rect 509782 366938 509866 367174
rect 510102 366938 510134 367174
rect 509514 366854 510134 366938
rect 509514 366618 509546 366854
rect 509782 366618 509866 366854
rect 510102 366618 510134 366854
rect 509514 331174 510134 366618
rect 513234 586894 513854 601103
rect 513234 586658 513266 586894
rect 513502 586658 513586 586894
rect 513822 586658 513854 586894
rect 513234 586574 513854 586658
rect 513234 586338 513266 586574
rect 513502 586338 513586 586574
rect 513822 586338 513854 586574
rect 513234 550894 513854 586338
rect 513234 550658 513266 550894
rect 513502 550658 513586 550894
rect 513822 550658 513854 550894
rect 513234 550574 513854 550658
rect 513234 550338 513266 550574
rect 513502 550338 513586 550574
rect 513822 550338 513854 550574
rect 513234 514894 513854 550338
rect 513234 514658 513266 514894
rect 513502 514658 513586 514894
rect 513822 514658 513854 514894
rect 513234 514574 513854 514658
rect 513234 514338 513266 514574
rect 513502 514338 513586 514574
rect 513822 514338 513854 514574
rect 513234 478894 513854 514338
rect 513234 478658 513266 478894
rect 513502 478658 513586 478894
rect 513822 478658 513854 478894
rect 513234 478574 513854 478658
rect 513234 478338 513266 478574
rect 513502 478338 513586 478574
rect 513822 478338 513854 478574
rect 513234 442894 513854 478338
rect 513234 442658 513266 442894
rect 513502 442658 513586 442894
rect 513822 442658 513854 442894
rect 513234 442574 513854 442658
rect 513234 442338 513266 442574
rect 513502 442338 513586 442574
rect 513822 442338 513854 442574
rect 513234 406894 513854 442338
rect 513234 406658 513266 406894
rect 513502 406658 513586 406894
rect 513822 406658 513854 406894
rect 513234 406574 513854 406658
rect 513234 406338 513266 406574
rect 513502 406338 513586 406574
rect 513822 406338 513854 406574
rect 513234 370894 513854 406338
rect 513234 370658 513266 370894
rect 513502 370658 513586 370894
rect 513822 370658 513854 370894
rect 513234 370574 513854 370658
rect 513234 370338 513266 370574
rect 513502 370338 513586 370574
rect 513822 370338 513854 370574
rect 510659 342820 510725 342821
rect 510659 342756 510660 342820
rect 510724 342756 510725 342820
rect 510659 342755 510725 342756
rect 509514 330938 509546 331174
rect 509782 330938 509866 331174
rect 510102 330938 510134 331174
rect 509514 330854 510134 330938
rect 509514 330618 509546 330854
rect 509782 330618 509866 330854
rect 510102 330618 510134 330854
rect 509514 295174 510134 330618
rect 510291 325956 510357 325957
rect 510291 325892 510292 325956
rect 510356 325892 510357 325956
rect 510291 325891 510357 325892
rect 510294 322693 510354 325891
rect 510475 323780 510541 323781
rect 510475 323716 510476 323780
rect 510540 323716 510541 323780
rect 510475 323715 510541 323716
rect 510291 322692 510357 322693
rect 510291 322628 510292 322692
rect 510356 322628 510357 322692
rect 510291 322627 510357 322628
rect 510478 305965 510538 323715
rect 510475 305964 510541 305965
rect 510475 305900 510476 305964
rect 510540 305900 510541 305964
rect 510475 305899 510541 305900
rect 510662 305829 510722 342755
rect 513234 334894 513854 370338
rect 513234 334658 513266 334894
rect 513502 334658 513586 334894
rect 513822 334658 513854 334894
rect 513234 334574 513854 334658
rect 513234 334338 513266 334574
rect 513502 334338 513586 334574
rect 513822 334338 513854 334574
rect 510843 331940 510909 331941
rect 510843 331876 510844 331940
rect 510908 331876 510909 331940
rect 510843 331875 510909 331876
rect 510659 305828 510725 305829
rect 510659 305764 510660 305828
rect 510724 305764 510725 305828
rect 510659 305763 510725 305764
rect 509514 294938 509546 295174
rect 509782 294938 509866 295174
rect 510102 294938 510134 295174
rect 509514 294854 510134 294938
rect 509514 294618 509546 294854
rect 509782 294618 509866 294854
rect 510102 294618 510134 294854
rect 509514 259417 510134 294618
rect 510846 294541 510906 331875
rect 511211 327588 511277 327589
rect 511211 327524 511212 327588
rect 511276 327524 511277 327588
rect 511211 327523 511277 327524
rect 511027 324324 511093 324325
rect 511027 324260 511028 324324
rect 511092 324260 511093 324324
rect 511027 324259 511093 324260
rect 511030 305693 511090 324259
rect 511214 321469 511274 327523
rect 511211 321468 511277 321469
rect 511211 321404 511212 321468
rect 511276 321404 511277 321468
rect 511211 321403 511277 321404
rect 511027 305692 511093 305693
rect 511027 305628 511028 305692
rect 511092 305628 511093 305692
rect 511027 305627 511093 305628
rect 513234 298894 513854 334338
rect 516954 590614 517574 601103
rect 516954 590378 516986 590614
rect 517222 590378 517306 590614
rect 517542 590378 517574 590614
rect 516954 590294 517574 590378
rect 516954 590058 516986 590294
rect 517222 590058 517306 590294
rect 517542 590058 517574 590294
rect 516954 554614 517574 590058
rect 516954 554378 516986 554614
rect 517222 554378 517306 554614
rect 517542 554378 517574 554614
rect 516954 554294 517574 554378
rect 516954 554058 516986 554294
rect 517222 554058 517306 554294
rect 517542 554058 517574 554294
rect 516954 518614 517574 554058
rect 516954 518378 516986 518614
rect 517222 518378 517306 518614
rect 517542 518378 517574 518614
rect 516954 518294 517574 518378
rect 516954 518058 516986 518294
rect 517222 518058 517306 518294
rect 517542 518058 517574 518294
rect 516954 482614 517574 518058
rect 516954 482378 516986 482614
rect 517222 482378 517306 482614
rect 517542 482378 517574 482614
rect 516954 482294 517574 482378
rect 516954 482058 516986 482294
rect 517222 482058 517306 482294
rect 517542 482058 517574 482294
rect 516954 446614 517574 482058
rect 516954 446378 516986 446614
rect 517222 446378 517306 446614
rect 517542 446378 517574 446614
rect 516954 446294 517574 446378
rect 516954 446058 516986 446294
rect 517222 446058 517306 446294
rect 517542 446058 517574 446294
rect 516954 410614 517574 446058
rect 516954 410378 516986 410614
rect 517222 410378 517306 410614
rect 517542 410378 517574 410614
rect 516954 410294 517574 410378
rect 516954 410058 516986 410294
rect 517222 410058 517306 410294
rect 517542 410058 517574 410294
rect 516954 374614 517574 410058
rect 516954 374378 516986 374614
rect 517222 374378 517306 374614
rect 517542 374378 517574 374614
rect 516954 374294 517574 374378
rect 516954 374058 516986 374294
rect 517222 374058 517306 374294
rect 517542 374058 517574 374294
rect 516954 338614 517574 374058
rect 520674 594334 521294 629778
rect 520674 594098 520706 594334
rect 520942 594098 521026 594334
rect 521262 594098 521294 594334
rect 520674 594014 521294 594098
rect 520674 593778 520706 594014
rect 520942 593778 521026 594014
rect 521262 593778 521294 594014
rect 520674 558334 521294 593778
rect 520674 558098 520706 558334
rect 520942 558098 521026 558334
rect 521262 558098 521294 558334
rect 520674 558014 521294 558098
rect 520674 557778 520706 558014
rect 520942 557778 521026 558014
rect 521262 557778 521294 558014
rect 520674 522334 521294 557778
rect 520674 522098 520706 522334
rect 520942 522098 521026 522334
rect 521262 522098 521294 522334
rect 520674 522014 521294 522098
rect 520674 521778 520706 522014
rect 520942 521778 521026 522014
rect 521262 521778 521294 522014
rect 520674 486334 521294 521778
rect 520674 486098 520706 486334
rect 520942 486098 521026 486334
rect 521262 486098 521294 486334
rect 520674 486014 521294 486098
rect 520674 485778 520706 486014
rect 520942 485778 521026 486014
rect 521262 485778 521294 486014
rect 520674 450334 521294 485778
rect 520674 450098 520706 450334
rect 520942 450098 521026 450334
rect 521262 450098 521294 450334
rect 520674 450014 521294 450098
rect 520674 449778 520706 450014
rect 520942 449778 521026 450014
rect 521262 449778 521294 450014
rect 520674 414334 521294 449778
rect 520674 414098 520706 414334
rect 520942 414098 521026 414334
rect 521262 414098 521294 414334
rect 520674 414014 521294 414098
rect 520674 413778 520706 414014
rect 520942 413778 521026 414014
rect 521262 413778 521294 414014
rect 520674 378334 521294 413778
rect 520674 378098 520706 378334
rect 520942 378098 521026 378334
rect 521262 378098 521294 378334
rect 520674 378014 521294 378098
rect 520674 377778 520706 378014
rect 520942 377778 521026 378014
rect 521262 377778 521294 378014
rect 520674 342334 521294 377778
rect 520674 342098 520706 342334
rect 520942 342098 521026 342334
rect 521262 342098 521294 342334
rect 520674 342014 521294 342098
rect 520674 341778 520706 342014
rect 520942 341778 521026 342014
rect 521262 341778 521294 342014
rect 517835 339556 517901 339557
rect 517835 339492 517836 339556
rect 517900 339492 517901 339556
rect 517835 339491 517901 339492
rect 516954 338378 516986 338614
rect 517222 338378 517306 338614
rect 517542 338378 517574 338614
rect 516954 338294 517574 338378
rect 516954 338058 516986 338294
rect 517222 338058 517306 338294
rect 517542 338058 517574 338294
rect 515259 331396 515325 331397
rect 515259 331332 515260 331396
rect 515324 331332 515325 331396
rect 515259 331331 515325 331332
rect 515075 329764 515141 329765
rect 515075 329700 515076 329764
rect 515140 329700 515141 329764
rect 515075 329699 515141 329700
rect 514155 327044 514221 327045
rect 514155 326980 514156 327044
rect 514220 326980 514221 327044
rect 514155 326979 514221 326980
rect 514158 300525 514218 326979
rect 514891 324868 514957 324869
rect 514891 324804 514892 324868
rect 514956 324804 514957 324868
rect 514891 324803 514957 324804
rect 514155 300524 514221 300525
rect 514155 300460 514156 300524
rect 514220 300460 514221 300524
rect 514155 300459 514221 300460
rect 514894 300389 514954 324803
rect 515078 316709 515138 329699
rect 515075 316708 515141 316709
rect 515075 316644 515076 316708
rect 515140 316644 515141 316708
rect 515075 316643 515141 316644
rect 515262 300661 515322 331331
rect 516954 302614 517574 338058
rect 516954 302378 516986 302614
rect 517222 302378 517306 302614
rect 517542 302378 517574 302614
rect 516954 302294 517574 302378
rect 516954 302058 516986 302294
rect 517222 302058 517306 302294
rect 517542 302058 517574 302294
rect 515259 300660 515325 300661
rect 515259 300596 515260 300660
rect 515324 300596 515325 300660
rect 515259 300595 515325 300596
rect 514891 300388 514957 300389
rect 514891 300324 514892 300388
rect 514956 300324 514957 300388
rect 514891 300323 514957 300324
rect 513234 298658 513266 298894
rect 513502 298658 513586 298894
rect 513822 298658 513854 298894
rect 513234 298574 513854 298658
rect 513234 298338 513266 298574
rect 513502 298338 513586 298574
rect 513822 298338 513854 298574
rect 510843 294540 510909 294541
rect 510843 294476 510844 294540
rect 510908 294476 510909 294540
rect 510843 294475 510909 294476
rect 513234 262894 513854 298338
rect 513234 262658 513266 262894
rect 513502 262658 513586 262894
rect 513822 262658 513854 262894
rect 513234 262574 513854 262658
rect 513234 262338 513266 262574
rect 513502 262338 513586 262574
rect 513822 262338 513854 262574
rect 513234 259417 513854 262338
rect 516954 266614 517574 302058
rect 517838 300117 517898 339491
rect 518019 334660 518085 334661
rect 518019 334596 518020 334660
rect 518084 334596 518085 334660
rect 518019 334595 518085 334596
rect 518022 300253 518082 334595
rect 518939 329900 519005 329901
rect 518939 329836 518940 329900
rect 519004 329836 519005 329900
rect 518939 329835 519005 329836
rect 518019 300252 518085 300253
rect 518019 300188 518020 300252
rect 518084 300188 518085 300252
rect 518019 300187 518085 300188
rect 517835 300116 517901 300117
rect 517835 300052 517836 300116
rect 517900 300052 517901 300116
rect 517835 300051 517901 300052
rect 518942 291821 519002 329835
rect 520674 306334 521294 341778
rect 520674 306098 520706 306334
rect 520942 306098 521026 306334
rect 521262 306098 521294 306334
rect 520674 306014 521294 306098
rect 520674 305778 520706 306014
rect 520942 305778 521026 306014
rect 521262 305778 521294 306014
rect 518939 291820 519005 291821
rect 518939 291756 518940 291820
rect 519004 291756 519005 291820
rect 518939 291755 519005 291756
rect 516954 266378 516986 266614
rect 517222 266378 517306 266614
rect 517542 266378 517574 266614
rect 516954 266294 517574 266378
rect 516954 266058 516986 266294
rect 517222 266058 517306 266294
rect 517542 266058 517574 266294
rect 516954 259417 517574 266058
rect 520674 270334 521294 305778
rect 520674 270098 520706 270334
rect 520942 270098 521026 270334
rect 521262 270098 521294 270334
rect 520674 270014 521294 270098
rect 520674 269778 520706 270014
rect 520942 269778 521026 270014
rect 521262 269778 521294 270014
rect 520674 259417 521294 269778
rect 524394 709638 525014 711590
rect 524394 709402 524426 709638
rect 524662 709402 524746 709638
rect 524982 709402 525014 709638
rect 524394 709318 525014 709402
rect 524394 709082 524426 709318
rect 524662 709082 524746 709318
rect 524982 709082 525014 709318
rect 524394 670054 525014 709082
rect 528114 710598 528734 711590
rect 528114 710362 528146 710598
rect 528382 710362 528466 710598
rect 528702 710362 528734 710598
rect 528114 710278 528734 710362
rect 528114 710042 528146 710278
rect 528382 710042 528466 710278
rect 528702 710042 528734 710278
rect 527219 699820 527285 699821
rect 527219 699756 527220 699820
rect 527284 699756 527285 699820
rect 527219 699755 527285 699756
rect 524394 669818 524426 670054
rect 524662 669818 524746 670054
rect 524982 669818 525014 670054
rect 524394 669734 525014 669818
rect 524394 669498 524426 669734
rect 524662 669498 524746 669734
rect 524982 669498 525014 669734
rect 524394 634054 525014 669498
rect 525648 651454 525968 651486
rect 525648 651218 525690 651454
rect 525926 651218 525968 651454
rect 525648 651134 525968 651218
rect 525648 650898 525690 651134
rect 525926 650898 525968 651134
rect 525648 650866 525968 650898
rect 524394 633818 524426 634054
rect 524662 633818 524746 634054
rect 524982 633818 525014 634054
rect 524394 633734 525014 633818
rect 524394 633498 524426 633734
rect 524662 633498 524746 633734
rect 524982 633498 525014 633734
rect 524394 598054 525014 633498
rect 525648 615454 525968 615486
rect 525648 615218 525690 615454
rect 525926 615218 525968 615454
rect 525648 615134 525968 615218
rect 525648 614898 525690 615134
rect 525926 614898 525968 615134
rect 525648 614866 525968 614898
rect 524394 597818 524426 598054
rect 524662 597818 524746 598054
rect 524982 597818 525014 598054
rect 524394 597734 525014 597818
rect 524394 597498 524426 597734
rect 524662 597498 524746 597734
rect 524982 597498 525014 597734
rect 524394 562054 525014 597498
rect 524394 561818 524426 562054
rect 524662 561818 524746 562054
rect 524982 561818 525014 562054
rect 524394 561734 525014 561818
rect 524394 561498 524426 561734
rect 524662 561498 524746 561734
rect 524982 561498 525014 561734
rect 524394 526054 525014 561498
rect 524394 525818 524426 526054
rect 524662 525818 524746 526054
rect 524982 525818 525014 526054
rect 524394 525734 525014 525818
rect 524394 525498 524426 525734
rect 524662 525498 524746 525734
rect 524982 525498 525014 525734
rect 524394 490054 525014 525498
rect 527222 502349 527282 699755
rect 528114 673774 528734 710042
rect 531834 711558 532454 711590
rect 531834 711322 531866 711558
rect 532102 711322 532186 711558
rect 532422 711322 532454 711558
rect 531834 711238 532454 711322
rect 531834 711002 531866 711238
rect 532102 711002 532186 711238
rect 532422 711002 532454 711238
rect 530531 700364 530597 700365
rect 530531 700300 530532 700364
rect 530596 700300 530597 700364
rect 530531 700299 530597 700300
rect 528114 673538 528146 673774
rect 528382 673538 528466 673774
rect 528702 673538 528734 673774
rect 528114 673454 528734 673538
rect 528114 673218 528146 673454
rect 528382 673218 528466 673454
rect 528702 673218 528734 673454
rect 528114 637774 528734 673218
rect 528114 637538 528146 637774
rect 528382 637538 528466 637774
rect 528702 637538 528734 637774
rect 528114 637454 528734 637538
rect 528114 637218 528146 637454
rect 528382 637218 528466 637454
rect 528702 637218 528734 637454
rect 528114 601774 528734 637218
rect 528114 601538 528146 601774
rect 528382 601538 528466 601774
rect 528702 601538 528734 601774
rect 528114 601454 528734 601538
rect 528114 601218 528146 601454
rect 528382 601218 528466 601454
rect 528702 601218 528734 601454
rect 528114 565774 528734 601218
rect 528114 565538 528146 565774
rect 528382 565538 528466 565774
rect 528702 565538 528734 565774
rect 528114 565454 528734 565538
rect 528114 565218 528146 565454
rect 528382 565218 528466 565454
rect 528702 565218 528734 565454
rect 528114 529774 528734 565218
rect 528114 529538 528146 529774
rect 528382 529538 528466 529774
rect 528702 529538 528734 529774
rect 528114 529454 528734 529538
rect 528114 529218 528146 529454
rect 528382 529218 528466 529454
rect 528702 529218 528734 529454
rect 527219 502348 527285 502349
rect 527219 502284 527220 502348
rect 527284 502284 527285 502348
rect 527219 502283 527285 502284
rect 524394 489818 524426 490054
rect 524662 489818 524746 490054
rect 524982 489818 525014 490054
rect 524394 489734 525014 489818
rect 524394 489498 524426 489734
rect 524662 489498 524746 489734
rect 524982 489498 525014 489734
rect 524394 454054 525014 489498
rect 524394 453818 524426 454054
rect 524662 453818 524746 454054
rect 524982 453818 525014 454054
rect 524394 453734 525014 453818
rect 524394 453498 524426 453734
rect 524662 453498 524746 453734
rect 524982 453498 525014 453734
rect 524394 418054 525014 453498
rect 528114 493774 528734 529218
rect 528114 493538 528146 493774
rect 528382 493538 528466 493774
rect 528702 493538 528734 493774
rect 528114 493454 528734 493538
rect 528114 493218 528146 493454
rect 528382 493218 528466 493454
rect 528702 493218 528734 493454
rect 528114 457774 528734 493218
rect 528114 457538 528146 457774
rect 528382 457538 528466 457774
rect 528702 457538 528734 457774
rect 528114 457454 528734 457538
rect 528114 457218 528146 457454
rect 528382 457218 528466 457454
rect 528702 457218 528734 457454
rect 525164 435454 525484 435486
rect 525164 435218 525206 435454
rect 525442 435218 525484 435454
rect 525164 435134 525484 435218
rect 525164 434898 525206 435134
rect 525442 434898 525484 435134
rect 525164 434866 525484 434898
rect 524394 417818 524426 418054
rect 524662 417818 524746 418054
rect 524982 417818 525014 418054
rect 524394 417734 525014 417818
rect 524394 417498 524426 417734
rect 524662 417498 524746 417734
rect 524982 417498 525014 417734
rect 524394 382054 525014 417498
rect 524394 381818 524426 382054
rect 524662 381818 524746 382054
rect 524982 381818 525014 382054
rect 524394 381734 525014 381818
rect 524394 381498 524426 381734
rect 524662 381498 524746 381734
rect 524982 381498 525014 381734
rect 524394 346054 525014 381498
rect 524394 345818 524426 346054
rect 524662 345818 524746 346054
rect 524982 345818 525014 346054
rect 524394 345734 525014 345818
rect 524394 345498 524426 345734
rect 524662 345498 524746 345734
rect 524982 345498 525014 345734
rect 524394 310054 525014 345498
rect 524394 309818 524426 310054
rect 524662 309818 524746 310054
rect 524982 309818 525014 310054
rect 524394 309734 525014 309818
rect 524394 309498 524426 309734
rect 524662 309498 524746 309734
rect 524982 309498 525014 309734
rect 524394 274054 525014 309498
rect 524394 273818 524426 274054
rect 524662 273818 524746 274054
rect 524982 273818 525014 274054
rect 524394 273734 525014 273818
rect 524394 273498 524426 273734
rect 524662 273498 524746 273734
rect 524982 273498 525014 273734
rect 524394 259417 525014 273498
rect 528114 421774 528734 457218
rect 529384 439174 529704 439206
rect 529384 438938 529426 439174
rect 529662 438938 529704 439174
rect 529384 438854 529704 438938
rect 529384 438618 529426 438854
rect 529662 438618 529704 438854
rect 529384 438586 529704 438618
rect 528114 421538 528146 421774
rect 528382 421538 528466 421774
rect 528702 421538 528734 421774
rect 528114 421454 528734 421538
rect 528114 421218 528146 421454
rect 528382 421218 528466 421454
rect 528702 421218 528734 421454
rect 528114 385774 528734 421218
rect 528114 385538 528146 385774
rect 528382 385538 528466 385774
rect 528702 385538 528734 385774
rect 528114 385454 528734 385538
rect 528114 385218 528146 385454
rect 528382 385218 528466 385454
rect 528702 385218 528734 385454
rect 528114 349774 528734 385218
rect 528114 349538 528146 349774
rect 528382 349538 528466 349774
rect 528702 349538 528734 349774
rect 528114 349454 528734 349538
rect 528114 349218 528146 349454
rect 528382 349218 528466 349454
rect 528702 349218 528734 349454
rect 528114 313774 528734 349218
rect 530534 321333 530594 700299
rect 531834 677494 532454 711002
rect 531834 677258 531866 677494
rect 532102 677258 532186 677494
rect 532422 677258 532454 677494
rect 531834 677174 532454 677258
rect 531834 676938 531866 677174
rect 532102 676938 532186 677174
rect 532422 676938 532454 677174
rect 531834 641494 532454 676938
rect 531834 641258 531866 641494
rect 532102 641258 532186 641494
rect 532422 641258 532454 641494
rect 531834 641174 532454 641258
rect 531834 640938 531866 641174
rect 532102 640938 532186 641174
rect 532422 640938 532454 641174
rect 531834 605494 532454 640938
rect 531834 605258 531866 605494
rect 532102 605258 532186 605494
rect 532422 605258 532454 605494
rect 531834 605174 532454 605258
rect 531834 604938 531866 605174
rect 532102 604938 532186 605174
rect 532422 604938 532454 605174
rect 531834 569494 532454 604938
rect 531834 569258 531866 569494
rect 532102 569258 532186 569494
rect 532422 569258 532454 569494
rect 531834 569174 532454 569258
rect 531834 568938 531866 569174
rect 532102 568938 532186 569174
rect 532422 568938 532454 569174
rect 531834 533494 532454 568938
rect 531834 533258 531866 533494
rect 532102 533258 532186 533494
rect 532422 533258 532454 533494
rect 531834 533174 532454 533258
rect 531834 532938 531866 533174
rect 532102 532938 532186 533174
rect 532422 532938 532454 533174
rect 531834 497494 532454 532938
rect 531834 497258 531866 497494
rect 532102 497258 532186 497494
rect 532422 497258 532454 497494
rect 531834 497174 532454 497258
rect 531834 496938 531866 497174
rect 532102 496938 532186 497174
rect 532422 496938 532454 497174
rect 531834 461494 532454 496938
rect 531834 461258 531866 461494
rect 532102 461258 532186 461494
rect 532422 461258 532454 461494
rect 531834 461174 532454 461258
rect 531834 460938 531866 461174
rect 532102 460938 532186 461174
rect 532422 460938 532454 461174
rect 531834 425494 532454 460938
rect 541794 704838 542414 711590
rect 541794 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 542414 704838
rect 541794 704518 542414 704602
rect 541794 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 542414 704518
rect 541794 687454 542414 704282
rect 541794 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 542414 687454
rect 541794 687134 542414 687218
rect 541794 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 542414 687134
rect 541794 651454 542414 686898
rect 541794 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 542414 651454
rect 541794 651134 542414 651218
rect 541794 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 542414 651134
rect 541794 615454 542414 650898
rect 541794 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 542414 615454
rect 541794 615134 542414 615218
rect 541794 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 542414 615134
rect 541794 579454 542414 614898
rect 541794 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 542414 579454
rect 541794 579134 542414 579218
rect 541794 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 542414 579134
rect 541794 543454 542414 578898
rect 541794 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 542414 543454
rect 541794 543134 542414 543218
rect 541794 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 542414 543134
rect 541794 507454 542414 542898
rect 541794 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 542414 507454
rect 541794 507134 542414 507218
rect 541794 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 542414 507134
rect 541794 471454 542414 506898
rect 541794 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 542414 471454
rect 541794 471134 542414 471218
rect 541794 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 542414 471134
rect 541794 460836 542414 470898
rect 545514 705798 546134 711590
rect 545514 705562 545546 705798
rect 545782 705562 545866 705798
rect 546102 705562 546134 705798
rect 545514 705478 546134 705562
rect 545514 705242 545546 705478
rect 545782 705242 545866 705478
rect 546102 705242 546134 705478
rect 545514 691174 546134 705242
rect 545514 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 546134 691174
rect 545514 690854 546134 690938
rect 545514 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 546134 690854
rect 545514 655174 546134 690618
rect 545514 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 546134 655174
rect 545514 654854 546134 654938
rect 545514 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 546134 654854
rect 545514 619174 546134 654618
rect 545514 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 546134 619174
rect 545514 618854 546134 618938
rect 545514 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 546134 618854
rect 545514 583174 546134 618618
rect 545514 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 546134 583174
rect 545514 582854 546134 582938
rect 545514 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 546134 582854
rect 545514 547174 546134 582618
rect 545514 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 546134 547174
rect 545514 546854 546134 546938
rect 545514 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 546134 546854
rect 545514 511174 546134 546618
rect 545514 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 546134 511174
rect 545514 510854 546134 510938
rect 545514 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 546134 510854
rect 545514 475174 546134 510618
rect 545514 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 546134 475174
rect 545514 474854 546134 474938
rect 545514 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 546134 474854
rect 537825 439174 538145 439206
rect 537825 438938 537867 439174
rect 538103 438938 538145 439174
rect 537825 438854 538145 438938
rect 537825 438618 537867 438854
rect 538103 438618 538145 438854
rect 537825 438586 538145 438618
rect 545514 439174 546134 474618
rect 549234 706758 549854 711590
rect 549234 706522 549266 706758
rect 549502 706522 549586 706758
rect 549822 706522 549854 706758
rect 549234 706438 549854 706522
rect 549234 706202 549266 706438
rect 549502 706202 549586 706438
rect 549822 706202 549854 706438
rect 549234 694894 549854 706202
rect 549234 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 549854 694894
rect 549234 694574 549854 694658
rect 549234 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 549854 694574
rect 549234 658894 549854 694338
rect 549234 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 549854 658894
rect 549234 658574 549854 658658
rect 549234 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 549854 658574
rect 549234 622894 549854 658338
rect 549234 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 549854 622894
rect 549234 622574 549854 622658
rect 549234 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 549854 622574
rect 549234 586894 549854 622338
rect 549234 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 549854 586894
rect 549234 586574 549854 586658
rect 549234 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 549854 586574
rect 549234 550894 549854 586338
rect 549234 550658 549266 550894
rect 549502 550658 549586 550894
rect 549822 550658 549854 550894
rect 549234 550574 549854 550658
rect 549234 550338 549266 550574
rect 549502 550338 549586 550574
rect 549822 550338 549854 550574
rect 549234 514894 549854 550338
rect 549234 514658 549266 514894
rect 549502 514658 549586 514894
rect 549822 514658 549854 514894
rect 549234 514574 549854 514658
rect 549234 514338 549266 514574
rect 549502 514338 549586 514574
rect 549822 514338 549854 514574
rect 549234 478894 549854 514338
rect 549234 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 549854 478894
rect 549234 478574 549854 478658
rect 549234 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 549854 478574
rect 549234 442894 549854 478338
rect 549234 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 549854 442894
rect 549234 442574 549854 442658
rect 549234 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 549854 442574
rect 545514 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 546134 439174
rect 545514 438854 546134 438938
rect 545514 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 546134 438854
rect 533605 435454 533925 435486
rect 533605 435218 533647 435454
rect 533883 435218 533925 435454
rect 533605 435134 533925 435218
rect 533605 434898 533647 435134
rect 533883 434898 533925 435134
rect 533605 434866 533925 434898
rect 542046 435454 542366 435486
rect 542046 435218 542088 435454
rect 542324 435218 542366 435454
rect 542046 435134 542366 435218
rect 542046 434898 542088 435134
rect 542324 434898 542366 435134
rect 542046 434866 542366 434898
rect 531834 425258 531866 425494
rect 532102 425258 532186 425494
rect 532422 425258 532454 425494
rect 531834 425174 532454 425258
rect 531834 424938 531866 425174
rect 532102 424938 532186 425174
rect 532422 424938 532454 425174
rect 531834 389494 532454 424938
rect 531834 389258 531866 389494
rect 532102 389258 532186 389494
rect 532422 389258 532454 389494
rect 531834 389174 532454 389258
rect 531834 388938 531866 389174
rect 532102 388938 532186 389174
rect 532422 388938 532454 389174
rect 531834 353494 532454 388938
rect 531834 353258 531866 353494
rect 532102 353258 532186 353494
rect 532422 353258 532454 353494
rect 531834 353174 532454 353258
rect 531834 352938 531866 353174
rect 532102 352938 532186 353174
rect 532422 352938 532454 353174
rect 530531 321332 530597 321333
rect 530531 321268 530532 321332
rect 530596 321268 530597 321332
rect 530531 321267 530597 321268
rect 528114 313538 528146 313774
rect 528382 313538 528466 313774
rect 528702 313538 528734 313774
rect 528114 313454 528734 313538
rect 528114 313218 528146 313454
rect 528382 313218 528466 313454
rect 528702 313218 528734 313454
rect 528114 277774 528734 313218
rect 528114 277538 528146 277774
rect 528382 277538 528466 277774
rect 528702 277538 528734 277774
rect 528114 277454 528734 277538
rect 528114 277218 528146 277454
rect 528382 277218 528466 277454
rect 528702 277218 528734 277454
rect 528114 259417 528734 277218
rect 531834 317494 532454 352938
rect 531834 317258 531866 317494
rect 532102 317258 532186 317494
rect 532422 317258 532454 317494
rect 531834 317174 532454 317258
rect 531834 316938 531866 317174
rect 532102 316938 532186 317174
rect 532422 316938 532454 317174
rect 531834 281494 532454 316938
rect 531834 281258 531866 281494
rect 532102 281258 532186 281494
rect 532422 281258 532454 281494
rect 531834 281174 532454 281258
rect 531834 280938 531866 281174
rect 532102 280938 532186 281174
rect 532422 280938 532454 281174
rect 479568 259174 479888 259206
rect 479568 258938 479610 259174
rect 479846 258938 479888 259174
rect 479568 258854 479888 258938
rect 479568 258618 479610 258854
rect 479846 258618 479888 258854
rect 479568 258586 479888 258618
rect 510288 259174 510608 259206
rect 510288 258938 510330 259174
rect 510566 258938 510608 259174
rect 510288 258854 510608 258938
rect 510288 258618 510330 258854
rect 510566 258618 510608 258854
rect 510288 258586 510608 258618
rect 464208 255454 464528 255486
rect 464208 255218 464250 255454
rect 464486 255218 464528 255454
rect 464208 255134 464528 255218
rect 464208 254898 464250 255134
rect 464486 254898 464528 255134
rect 464208 254866 464528 254898
rect 494928 255454 495248 255486
rect 494928 255218 494970 255454
rect 495206 255218 495248 255454
rect 494928 255134 495248 255218
rect 494928 254898 494970 255134
rect 495206 254898 495248 255134
rect 494928 254866 495248 254898
rect 525648 255454 525968 255486
rect 525648 255218 525690 255454
rect 525926 255218 525968 255454
rect 525648 255134 525968 255218
rect 525648 254898 525690 255134
rect 525926 254898 525968 255134
rect 525648 254866 525968 254898
rect 459834 245258 459866 245494
rect 460102 245258 460186 245494
rect 460422 245258 460454 245494
rect 459834 245174 460454 245258
rect 459834 244938 459866 245174
rect 460102 244938 460186 245174
rect 460422 244938 460454 245174
rect 459834 209494 460454 244938
rect 531834 245494 532454 280938
rect 541794 399454 542414 425068
rect 541794 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 542414 399454
rect 541794 399134 542414 399218
rect 541794 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 542414 399134
rect 541794 363454 542414 398898
rect 541794 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 542414 363454
rect 541794 363134 542414 363218
rect 541794 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 542414 363134
rect 541794 327454 542414 362898
rect 541794 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 542414 327454
rect 541794 327134 542414 327218
rect 541794 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 542414 327134
rect 541794 291454 542414 326898
rect 545514 403174 546134 438618
rect 546266 439174 546586 439206
rect 546266 438938 546308 439174
rect 546544 438938 546586 439174
rect 546266 438854 546586 438938
rect 546266 438618 546308 438854
rect 546544 438618 546586 438854
rect 546266 438586 546586 438618
rect 545514 402938 545546 403174
rect 545782 402938 545866 403174
rect 546102 402938 546134 403174
rect 545514 402854 546134 402938
rect 545514 402618 545546 402854
rect 545782 402618 545866 402854
rect 546102 402618 546134 402854
rect 545514 367174 546134 402618
rect 545514 366938 545546 367174
rect 545782 366938 545866 367174
rect 546102 366938 546134 367174
rect 545514 366854 546134 366938
rect 545514 366618 545546 366854
rect 545782 366618 545866 366854
rect 546102 366618 546134 366854
rect 545514 331174 546134 366618
rect 545514 330938 545546 331174
rect 545782 330938 545866 331174
rect 546102 330938 546134 331174
rect 545514 330854 546134 330938
rect 545514 330618 545546 330854
rect 545782 330618 545866 330854
rect 546102 330618 546134 330854
rect 542675 311132 542741 311133
rect 542675 311068 542676 311132
rect 542740 311068 542741 311132
rect 542675 311067 542741 311068
rect 541794 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 542414 291454
rect 541794 291134 542414 291218
rect 541794 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 542414 291134
rect 538259 278084 538325 278085
rect 538259 278020 538260 278084
rect 538324 278020 538325 278084
rect 538259 278019 538325 278020
rect 531834 245258 531866 245494
rect 532102 245258 532186 245494
rect 532422 245258 532454 245494
rect 531834 245174 532454 245258
rect 531834 244938 531866 245174
rect 532102 244938 532186 245174
rect 532422 244938 532454 245174
rect 479568 223174 479888 223206
rect 479568 222938 479610 223174
rect 479846 222938 479888 223174
rect 479568 222854 479888 222938
rect 479568 222618 479610 222854
rect 479846 222618 479888 222854
rect 479568 222586 479888 222618
rect 510288 223174 510608 223206
rect 510288 222938 510330 223174
rect 510566 222938 510608 223174
rect 510288 222854 510608 222938
rect 510288 222618 510330 222854
rect 510566 222618 510608 222854
rect 510288 222586 510608 222618
rect 464208 219454 464528 219486
rect 464208 219218 464250 219454
rect 464486 219218 464528 219454
rect 464208 219134 464528 219218
rect 464208 218898 464250 219134
rect 464486 218898 464528 219134
rect 464208 218866 464528 218898
rect 494928 219454 495248 219486
rect 494928 219218 494970 219454
rect 495206 219218 495248 219454
rect 494928 219134 495248 219218
rect 494928 218898 494970 219134
rect 495206 218898 495248 219134
rect 494928 218866 495248 218898
rect 525648 219454 525968 219486
rect 525648 219218 525690 219454
rect 525926 219218 525968 219454
rect 525648 219134 525968 219218
rect 525648 218898 525690 219134
rect 525926 218898 525968 219134
rect 525648 218866 525968 218898
rect 459834 209258 459866 209494
rect 460102 209258 460186 209494
rect 460422 209258 460454 209494
rect 459834 209174 460454 209258
rect 459834 208938 459866 209174
rect 460102 208938 460186 209174
rect 460422 208938 460454 209174
rect 459834 173494 460454 208938
rect 531834 209494 532454 244938
rect 531834 209258 531866 209494
rect 532102 209258 532186 209494
rect 532422 209258 532454 209494
rect 531834 209174 532454 209258
rect 531834 208938 531866 209174
rect 532102 208938 532186 209174
rect 532422 208938 532454 209174
rect 459834 173258 459866 173494
rect 460102 173258 460186 173494
rect 460422 173258 460454 173494
rect 459834 173174 460454 173258
rect 459834 172938 459866 173174
rect 460102 172938 460186 173174
rect 460422 172938 460454 173174
rect 459834 137494 460454 172938
rect 459834 137258 459866 137494
rect 460102 137258 460186 137494
rect 460422 137258 460454 137494
rect 459834 137174 460454 137258
rect 459834 136938 459866 137174
rect 460102 136938 460186 137174
rect 460422 136938 460454 137174
rect 459834 101494 460454 136938
rect 459834 101258 459866 101494
rect 460102 101258 460186 101494
rect 460422 101258 460454 101494
rect 459834 101174 460454 101258
rect 459834 100938 459866 101174
rect 460102 100938 460186 101174
rect 460422 100938 460454 101174
rect 459834 65494 460454 100938
rect 459834 65258 459866 65494
rect 460102 65258 460186 65494
rect 460422 65258 460454 65494
rect 459834 65174 460454 65258
rect 459834 64938 459866 65174
rect 460102 64938 460186 65174
rect 460422 64938 460454 65174
rect 459834 29494 460454 64938
rect 459834 29258 459866 29494
rect 460102 29258 460186 29494
rect 460422 29258 460454 29494
rect 459834 29174 460454 29258
rect 459834 28938 459866 29174
rect 460102 28938 460186 29174
rect 460422 28938 460454 29174
rect 458771 3364 458837 3365
rect 458771 3300 458772 3364
rect 458836 3300 458837 3364
rect 458771 3299 458837 3300
rect 456114 -6342 456146 -6106
rect 456382 -6342 456466 -6106
rect 456702 -6342 456734 -6106
rect 456114 -6426 456734 -6342
rect 456114 -6662 456146 -6426
rect 456382 -6662 456466 -6426
rect 456702 -6662 456734 -6426
rect 456114 -7654 456734 -6662
rect 459834 -7066 460454 28938
rect 459834 -7302 459866 -7066
rect 460102 -7302 460186 -7066
rect 460422 -7302 460454 -7066
rect 459834 -7386 460454 -7302
rect 459834 -7622 459866 -7386
rect 460102 -7622 460186 -7386
rect 460422 -7622 460454 -7386
rect 459834 -7654 460454 -7622
rect 469794 183454 470414 201919
rect 469794 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 470414 183454
rect 469794 183134 470414 183218
rect 469794 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 470414 183134
rect 469794 147454 470414 182898
rect 469794 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 470414 147454
rect 469794 147134 470414 147218
rect 469794 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 470414 147134
rect 469794 111454 470414 146898
rect 469794 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 470414 111454
rect 469794 111134 470414 111218
rect 469794 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 470414 111134
rect 469794 75454 470414 110898
rect 469794 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 470414 75454
rect 469794 75134 470414 75218
rect 469794 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 470414 75134
rect 469794 39454 470414 74898
rect 469794 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 470414 39454
rect 469794 39134 470414 39218
rect 469794 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 470414 39134
rect 469794 3454 470414 38898
rect 469794 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 470414 3454
rect 469794 3134 470414 3218
rect 469794 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 470414 3134
rect 469794 -346 470414 2898
rect 469794 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 470414 -346
rect 469794 -666 470414 -582
rect 469794 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 470414 -666
rect 469794 -7654 470414 -902
rect 473514 187174 474134 201919
rect 473514 186938 473546 187174
rect 473782 186938 473866 187174
rect 474102 186938 474134 187174
rect 473514 186854 474134 186938
rect 473514 186618 473546 186854
rect 473782 186618 473866 186854
rect 474102 186618 474134 186854
rect 473514 151174 474134 186618
rect 473514 150938 473546 151174
rect 473782 150938 473866 151174
rect 474102 150938 474134 151174
rect 473514 150854 474134 150938
rect 473514 150618 473546 150854
rect 473782 150618 473866 150854
rect 474102 150618 474134 150854
rect 473514 115174 474134 150618
rect 473514 114938 473546 115174
rect 473782 114938 473866 115174
rect 474102 114938 474134 115174
rect 473514 114854 474134 114938
rect 473514 114618 473546 114854
rect 473782 114618 473866 114854
rect 474102 114618 474134 114854
rect 473514 79174 474134 114618
rect 473514 78938 473546 79174
rect 473782 78938 473866 79174
rect 474102 78938 474134 79174
rect 473514 78854 474134 78938
rect 473514 78618 473546 78854
rect 473782 78618 473866 78854
rect 474102 78618 474134 78854
rect 473514 43174 474134 78618
rect 473514 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 474134 43174
rect 473514 42854 474134 42938
rect 473514 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 474134 42854
rect 473514 7174 474134 42618
rect 473514 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 474134 7174
rect 473514 6854 474134 6938
rect 473514 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 474134 6854
rect 473514 -1306 474134 6618
rect 473514 -1542 473546 -1306
rect 473782 -1542 473866 -1306
rect 474102 -1542 474134 -1306
rect 473514 -1626 474134 -1542
rect 473514 -1862 473546 -1626
rect 473782 -1862 473866 -1626
rect 474102 -1862 474134 -1626
rect 473514 -7654 474134 -1862
rect 477234 190894 477854 201919
rect 477234 190658 477266 190894
rect 477502 190658 477586 190894
rect 477822 190658 477854 190894
rect 477234 190574 477854 190658
rect 477234 190338 477266 190574
rect 477502 190338 477586 190574
rect 477822 190338 477854 190574
rect 477234 154894 477854 190338
rect 477234 154658 477266 154894
rect 477502 154658 477586 154894
rect 477822 154658 477854 154894
rect 477234 154574 477854 154658
rect 477234 154338 477266 154574
rect 477502 154338 477586 154574
rect 477822 154338 477854 154574
rect 477234 118894 477854 154338
rect 477234 118658 477266 118894
rect 477502 118658 477586 118894
rect 477822 118658 477854 118894
rect 477234 118574 477854 118658
rect 477234 118338 477266 118574
rect 477502 118338 477586 118574
rect 477822 118338 477854 118574
rect 477234 82894 477854 118338
rect 477234 82658 477266 82894
rect 477502 82658 477586 82894
rect 477822 82658 477854 82894
rect 477234 82574 477854 82658
rect 477234 82338 477266 82574
rect 477502 82338 477586 82574
rect 477822 82338 477854 82574
rect 477234 46894 477854 82338
rect 477234 46658 477266 46894
rect 477502 46658 477586 46894
rect 477822 46658 477854 46894
rect 477234 46574 477854 46658
rect 477234 46338 477266 46574
rect 477502 46338 477586 46574
rect 477822 46338 477854 46574
rect 477234 10894 477854 46338
rect 477234 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 477854 10894
rect 477234 10574 477854 10658
rect 477234 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 477854 10574
rect 477234 -2266 477854 10338
rect 477234 -2502 477266 -2266
rect 477502 -2502 477586 -2266
rect 477822 -2502 477854 -2266
rect 477234 -2586 477854 -2502
rect 477234 -2822 477266 -2586
rect 477502 -2822 477586 -2586
rect 477822 -2822 477854 -2586
rect 477234 -7654 477854 -2822
rect 480954 194614 481574 201919
rect 480954 194378 480986 194614
rect 481222 194378 481306 194614
rect 481542 194378 481574 194614
rect 480954 194294 481574 194378
rect 480954 194058 480986 194294
rect 481222 194058 481306 194294
rect 481542 194058 481574 194294
rect 480954 158614 481574 194058
rect 480954 158378 480986 158614
rect 481222 158378 481306 158614
rect 481542 158378 481574 158614
rect 480954 158294 481574 158378
rect 480954 158058 480986 158294
rect 481222 158058 481306 158294
rect 481542 158058 481574 158294
rect 480954 122614 481574 158058
rect 480954 122378 480986 122614
rect 481222 122378 481306 122614
rect 481542 122378 481574 122614
rect 480954 122294 481574 122378
rect 480954 122058 480986 122294
rect 481222 122058 481306 122294
rect 481542 122058 481574 122294
rect 480954 86614 481574 122058
rect 484674 198334 485294 201919
rect 484674 198098 484706 198334
rect 484942 198098 485026 198334
rect 485262 198098 485294 198334
rect 484674 198014 485294 198098
rect 484674 197778 484706 198014
rect 484942 197778 485026 198014
rect 485262 197778 485294 198014
rect 484674 162334 485294 197778
rect 484674 162098 484706 162334
rect 484942 162098 485026 162334
rect 485262 162098 485294 162334
rect 484674 162014 485294 162098
rect 484674 161778 484706 162014
rect 484942 161778 485026 162014
rect 485262 161778 485294 162014
rect 484674 126334 485294 161778
rect 488394 166054 489014 201919
rect 488394 165818 488426 166054
rect 488662 165818 488746 166054
rect 488982 165818 489014 166054
rect 488394 165734 489014 165818
rect 488394 165498 488426 165734
rect 488662 165498 488746 165734
rect 488982 165498 489014 165734
rect 488394 139281 489014 165498
rect 505794 183454 506414 201919
rect 505794 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 506414 183454
rect 505794 183134 506414 183218
rect 505794 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 506414 183134
rect 505794 147454 506414 182898
rect 505794 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 506414 147454
rect 505794 147134 506414 147218
rect 505794 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 506414 147134
rect 505794 139281 506414 146898
rect 509514 187174 510134 201919
rect 509514 186938 509546 187174
rect 509782 186938 509866 187174
rect 510102 186938 510134 187174
rect 509514 186854 510134 186938
rect 509514 186618 509546 186854
rect 509782 186618 509866 186854
rect 510102 186618 510134 186854
rect 509514 151174 510134 186618
rect 509514 150938 509546 151174
rect 509782 150938 509866 151174
rect 510102 150938 510134 151174
rect 509514 150854 510134 150938
rect 509514 150618 509546 150854
rect 509782 150618 509866 150854
rect 510102 150618 510134 150854
rect 509514 139281 510134 150618
rect 513234 190894 513854 201919
rect 513234 190658 513266 190894
rect 513502 190658 513586 190894
rect 513822 190658 513854 190894
rect 513234 190574 513854 190658
rect 513234 190338 513266 190574
rect 513502 190338 513586 190574
rect 513822 190338 513854 190574
rect 513234 154894 513854 190338
rect 513234 154658 513266 154894
rect 513502 154658 513586 154894
rect 513822 154658 513854 154894
rect 513234 154574 513854 154658
rect 513234 154338 513266 154574
rect 513502 154338 513586 154574
rect 513822 154338 513854 154574
rect 513234 139281 513854 154338
rect 516954 194614 517574 201919
rect 516954 194378 516986 194614
rect 517222 194378 517306 194614
rect 517542 194378 517574 194614
rect 516954 194294 517574 194378
rect 516954 194058 516986 194294
rect 517222 194058 517306 194294
rect 517542 194058 517574 194294
rect 516954 158614 517574 194058
rect 516954 158378 516986 158614
rect 517222 158378 517306 158614
rect 517542 158378 517574 158614
rect 516954 158294 517574 158378
rect 516954 158058 516986 158294
rect 517222 158058 517306 158294
rect 517542 158058 517574 158294
rect 516954 139281 517574 158058
rect 520674 198334 521294 201919
rect 520674 198098 520706 198334
rect 520942 198098 521026 198334
rect 521262 198098 521294 198334
rect 520674 198014 521294 198098
rect 520674 197778 520706 198014
rect 520942 197778 521026 198014
rect 521262 197778 521294 198014
rect 520674 162334 521294 197778
rect 520674 162098 520706 162334
rect 520942 162098 521026 162334
rect 521262 162098 521294 162334
rect 520674 162014 521294 162098
rect 520674 161778 520706 162014
rect 520942 161778 521026 162014
rect 521262 161778 521294 162014
rect 520674 139281 521294 161778
rect 524394 166054 525014 201919
rect 524394 165818 524426 166054
rect 524662 165818 524746 166054
rect 524982 165818 525014 166054
rect 524394 165734 525014 165818
rect 524394 165498 524426 165734
rect 524662 165498 524746 165734
rect 524982 165498 525014 165734
rect 524394 139281 525014 165498
rect 531834 173494 532454 208938
rect 531834 173258 531866 173494
rect 532102 173258 532186 173494
rect 532422 173258 532454 173494
rect 531834 173174 532454 173258
rect 531834 172938 531866 173174
rect 532102 172938 532186 173174
rect 532422 172938 532454 173174
rect 531834 139281 532454 172938
rect 538262 151830 538322 278019
rect 541794 255454 542414 290898
rect 541794 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 542414 255454
rect 541794 255134 542414 255218
rect 541794 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 542414 255134
rect 541794 219454 542414 254898
rect 541794 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 542414 219454
rect 541794 219134 542414 219218
rect 541794 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 542414 219134
rect 541794 183454 542414 218898
rect 541794 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 542414 183454
rect 541794 183134 542414 183218
rect 541794 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 542414 183134
rect 538262 151770 539426 151830
rect 539366 127261 539426 151770
rect 541794 147454 542414 182898
rect 541794 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 542414 147454
rect 541794 147134 542414 147218
rect 541794 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 542414 147134
rect 539363 127260 539429 127261
rect 539363 127196 539364 127260
rect 539428 127196 539429 127260
rect 539363 127195 539429 127196
rect 484674 126098 484706 126334
rect 484942 126098 485026 126334
rect 485262 126098 485294 126334
rect 484674 126014 485294 126098
rect 484674 125778 484706 126014
rect 484942 125778 485026 126014
rect 485262 125778 485294 126014
rect 484208 111454 484528 111486
rect 484208 111218 484250 111454
rect 484486 111218 484528 111454
rect 484208 111134 484528 111218
rect 484208 110898 484250 111134
rect 484486 110898 484528 111134
rect 484208 110866 484528 110898
rect 480954 86378 480986 86614
rect 481222 86378 481306 86614
rect 481542 86378 481574 86614
rect 480954 86294 481574 86378
rect 480954 86058 480986 86294
rect 481222 86058 481306 86294
rect 481542 86058 481574 86294
rect 480954 50614 481574 86058
rect 480954 50378 480986 50614
rect 481222 50378 481306 50614
rect 481542 50378 481574 50614
rect 480954 50294 481574 50378
rect 480954 50058 480986 50294
rect 481222 50058 481306 50294
rect 481542 50058 481574 50294
rect 480954 14614 481574 50058
rect 480954 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 481574 14614
rect 480954 14294 481574 14378
rect 480954 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 481574 14294
rect 480954 -3226 481574 14058
rect 480954 -3462 480986 -3226
rect 481222 -3462 481306 -3226
rect 481542 -3462 481574 -3226
rect 480954 -3546 481574 -3462
rect 480954 -3782 480986 -3546
rect 481222 -3782 481306 -3546
rect 481542 -3782 481574 -3546
rect 480954 -7654 481574 -3782
rect 484674 90334 485294 125778
rect 499568 115174 499888 115206
rect 499568 114938 499610 115174
rect 499846 114938 499888 115174
rect 499568 114854 499888 114938
rect 499568 114618 499610 114854
rect 499846 114618 499888 114854
rect 499568 114586 499888 114618
rect 530288 115174 530608 115206
rect 530288 114938 530330 115174
rect 530566 114938 530608 115174
rect 530288 114854 530608 114938
rect 530288 114618 530330 114854
rect 530566 114618 530608 114854
rect 530288 114586 530608 114618
rect 514928 111454 515248 111486
rect 514928 111218 514970 111454
rect 515206 111218 515248 111454
rect 514928 111134 515248 111218
rect 514928 110898 514970 111134
rect 515206 110898 515248 111134
rect 514928 110866 515248 110898
rect 541794 111454 542414 146898
rect 541794 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 542414 111454
rect 541794 111134 542414 111218
rect 541794 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 542414 111134
rect 484674 90098 484706 90334
rect 484942 90098 485026 90334
rect 485262 90098 485294 90334
rect 484674 90014 485294 90098
rect 484674 89778 484706 90014
rect 484942 89778 485026 90014
rect 485262 89778 485294 90014
rect 484674 54334 485294 89778
rect 484674 54098 484706 54334
rect 484942 54098 485026 54334
rect 485262 54098 485294 54334
rect 484674 54014 485294 54098
rect 484674 53778 484706 54014
rect 484942 53778 485026 54014
rect 485262 53778 485294 54014
rect 484674 18334 485294 53778
rect 484674 18098 484706 18334
rect 484942 18098 485026 18334
rect 485262 18098 485294 18334
rect 484674 18014 485294 18098
rect 484674 17778 484706 18014
rect 484942 17778 485026 18014
rect 485262 17778 485294 18014
rect 484674 -4186 485294 17778
rect 484674 -4422 484706 -4186
rect 484942 -4422 485026 -4186
rect 485262 -4422 485294 -4186
rect 484674 -4506 485294 -4422
rect 484674 -4742 484706 -4506
rect 484942 -4742 485026 -4506
rect 485262 -4742 485294 -4506
rect 484674 -7654 485294 -4742
rect 488394 58054 489014 82599
rect 488394 57818 488426 58054
rect 488662 57818 488746 58054
rect 488982 57818 489014 58054
rect 488394 57734 489014 57818
rect 488394 57498 488426 57734
rect 488662 57498 488746 57734
rect 488982 57498 489014 57734
rect 488394 22054 489014 57498
rect 488394 21818 488426 22054
rect 488662 21818 488746 22054
rect 488982 21818 489014 22054
rect 488394 21734 489014 21818
rect 488394 21498 488426 21734
rect 488662 21498 488746 21734
rect 488982 21498 489014 21734
rect 488394 -5146 489014 21498
rect 488394 -5382 488426 -5146
rect 488662 -5382 488746 -5146
rect 488982 -5382 489014 -5146
rect 488394 -5466 489014 -5382
rect 488394 -5702 488426 -5466
rect 488662 -5702 488746 -5466
rect 488982 -5702 489014 -5466
rect 488394 -7654 489014 -5702
rect 492114 61774 492734 82599
rect 492114 61538 492146 61774
rect 492382 61538 492466 61774
rect 492702 61538 492734 61774
rect 492114 61454 492734 61538
rect 492114 61218 492146 61454
rect 492382 61218 492466 61454
rect 492702 61218 492734 61454
rect 492114 25774 492734 61218
rect 492114 25538 492146 25774
rect 492382 25538 492466 25774
rect 492702 25538 492734 25774
rect 492114 25454 492734 25538
rect 492114 25218 492146 25454
rect 492382 25218 492466 25454
rect 492702 25218 492734 25454
rect 492114 -6106 492734 25218
rect 492114 -6342 492146 -6106
rect 492382 -6342 492466 -6106
rect 492702 -6342 492734 -6106
rect 492114 -6426 492734 -6342
rect 492114 -6662 492146 -6426
rect 492382 -6662 492466 -6426
rect 492702 -6662 492734 -6426
rect 492114 -7654 492734 -6662
rect 495834 65494 496454 82599
rect 495834 65258 495866 65494
rect 496102 65258 496186 65494
rect 496422 65258 496454 65494
rect 495834 65174 496454 65258
rect 495834 64938 495866 65174
rect 496102 64938 496186 65174
rect 496422 64938 496454 65174
rect 495834 29494 496454 64938
rect 495834 29258 495866 29494
rect 496102 29258 496186 29494
rect 496422 29258 496454 29494
rect 495834 29174 496454 29258
rect 495834 28938 495866 29174
rect 496102 28938 496186 29174
rect 496422 28938 496454 29174
rect 495834 -7066 496454 28938
rect 495834 -7302 495866 -7066
rect 496102 -7302 496186 -7066
rect 496422 -7302 496454 -7066
rect 495834 -7386 496454 -7302
rect 495834 -7622 495866 -7386
rect 496102 -7622 496186 -7386
rect 496422 -7622 496454 -7386
rect 495834 -7654 496454 -7622
rect 505794 75454 506414 82599
rect 505794 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 506414 75454
rect 505794 75134 506414 75218
rect 505794 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 506414 75134
rect 505794 39454 506414 74898
rect 505794 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 506414 39454
rect 505794 39134 506414 39218
rect 505794 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 506414 39134
rect 505794 3454 506414 38898
rect 505794 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 506414 3454
rect 505794 3134 506414 3218
rect 505794 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 506414 3134
rect 505794 -346 506414 2898
rect 505794 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 506414 -346
rect 505794 -666 506414 -582
rect 505794 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 506414 -666
rect 505794 -7654 506414 -902
rect 509514 79174 510134 82599
rect 509514 78938 509546 79174
rect 509782 78938 509866 79174
rect 510102 78938 510134 79174
rect 509514 78854 510134 78938
rect 509514 78618 509546 78854
rect 509782 78618 509866 78854
rect 510102 78618 510134 78854
rect 509514 43174 510134 78618
rect 509514 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 510134 43174
rect 509514 42854 510134 42938
rect 509514 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 510134 42854
rect 509514 7174 510134 42618
rect 509514 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 510134 7174
rect 509514 6854 510134 6938
rect 509514 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 510134 6854
rect 509514 -1306 510134 6618
rect 509514 -1542 509546 -1306
rect 509782 -1542 509866 -1306
rect 510102 -1542 510134 -1306
rect 509514 -1626 510134 -1542
rect 509514 -1862 509546 -1626
rect 509782 -1862 509866 -1626
rect 510102 -1862 510134 -1626
rect 509514 -7654 510134 -1862
rect 513234 46894 513854 82599
rect 513234 46658 513266 46894
rect 513502 46658 513586 46894
rect 513822 46658 513854 46894
rect 513234 46574 513854 46658
rect 513234 46338 513266 46574
rect 513502 46338 513586 46574
rect 513822 46338 513854 46574
rect 513234 10894 513854 46338
rect 513234 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 513854 10894
rect 513234 10574 513854 10658
rect 513234 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 513854 10574
rect 513234 -2266 513854 10338
rect 513234 -2502 513266 -2266
rect 513502 -2502 513586 -2266
rect 513822 -2502 513854 -2266
rect 513234 -2586 513854 -2502
rect 513234 -2822 513266 -2586
rect 513502 -2822 513586 -2586
rect 513822 -2822 513854 -2586
rect 513234 -7654 513854 -2822
rect 516954 50614 517574 82599
rect 516954 50378 516986 50614
rect 517222 50378 517306 50614
rect 517542 50378 517574 50614
rect 516954 50294 517574 50378
rect 516954 50058 516986 50294
rect 517222 50058 517306 50294
rect 517542 50058 517574 50294
rect 516954 14614 517574 50058
rect 516954 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 517574 14614
rect 516954 14294 517574 14378
rect 516954 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 517574 14294
rect 516954 -3226 517574 14058
rect 516954 -3462 516986 -3226
rect 517222 -3462 517306 -3226
rect 517542 -3462 517574 -3226
rect 516954 -3546 517574 -3462
rect 516954 -3782 516986 -3546
rect 517222 -3782 517306 -3546
rect 517542 -3782 517574 -3546
rect 516954 -7654 517574 -3782
rect 520674 54334 521294 82599
rect 520674 54098 520706 54334
rect 520942 54098 521026 54334
rect 521262 54098 521294 54334
rect 520674 54014 521294 54098
rect 520674 53778 520706 54014
rect 520942 53778 521026 54014
rect 521262 53778 521294 54014
rect 520674 18334 521294 53778
rect 520674 18098 520706 18334
rect 520942 18098 521026 18334
rect 521262 18098 521294 18334
rect 520674 18014 521294 18098
rect 520674 17778 520706 18014
rect 520942 17778 521026 18014
rect 521262 17778 521294 18014
rect 520674 -4186 521294 17778
rect 520674 -4422 520706 -4186
rect 520942 -4422 521026 -4186
rect 521262 -4422 521294 -4186
rect 520674 -4506 521294 -4422
rect 520674 -4742 520706 -4506
rect 520942 -4742 521026 -4506
rect 521262 -4742 521294 -4506
rect 520674 -7654 521294 -4742
rect 524394 58054 525014 82599
rect 524394 57818 524426 58054
rect 524662 57818 524746 58054
rect 524982 57818 525014 58054
rect 524394 57734 525014 57818
rect 524394 57498 524426 57734
rect 524662 57498 524746 57734
rect 524982 57498 525014 57734
rect 524394 22054 525014 57498
rect 524394 21818 524426 22054
rect 524662 21818 524746 22054
rect 524982 21818 525014 22054
rect 524394 21734 525014 21818
rect 524394 21498 524426 21734
rect 524662 21498 524746 21734
rect 524982 21498 525014 21734
rect 524394 -5146 525014 21498
rect 524394 -5382 524426 -5146
rect 524662 -5382 524746 -5146
rect 524982 -5382 525014 -5146
rect 524394 -5466 525014 -5382
rect 524394 -5702 524426 -5466
rect 524662 -5702 524746 -5466
rect 524982 -5702 525014 -5466
rect 524394 -7654 525014 -5702
rect 528114 61774 528734 82599
rect 528114 61538 528146 61774
rect 528382 61538 528466 61774
rect 528702 61538 528734 61774
rect 528114 61454 528734 61538
rect 528114 61218 528146 61454
rect 528382 61218 528466 61454
rect 528702 61218 528734 61454
rect 528114 25774 528734 61218
rect 528114 25538 528146 25774
rect 528382 25538 528466 25774
rect 528702 25538 528734 25774
rect 528114 25454 528734 25538
rect 528114 25218 528146 25454
rect 528382 25218 528466 25454
rect 528702 25218 528734 25454
rect 528114 -6106 528734 25218
rect 528114 -6342 528146 -6106
rect 528382 -6342 528466 -6106
rect 528702 -6342 528734 -6106
rect 528114 -6426 528734 -6342
rect 528114 -6662 528146 -6426
rect 528382 -6662 528466 -6426
rect 528702 -6662 528734 -6426
rect 528114 -7654 528734 -6662
rect 531834 65494 532454 82599
rect 531834 65258 531866 65494
rect 532102 65258 532186 65494
rect 532422 65258 532454 65494
rect 531834 65174 532454 65258
rect 531834 64938 531866 65174
rect 532102 64938 532186 65174
rect 532422 64938 532454 65174
rect 531834 29494 532454 64938
rect 531834 29258 531866 29494
rect 532102 29258 532186 29494
rect 532422 29258 532454 29494
rect 531834 29174 532454 29258
rect 531834 28938 531866 29174
rect 532102 28938 532186 29174
rect 532422 28938 532454 29174
rect 531834 -7066 532454 28938
rect 531834 -7302 531866 -7066
rect 532102 -7302 532186 -7066
rect 532422 -7302 532454 -7066
rect 531834 -7386 532454 -7302
rect 531834 -7622 531866 -7386
rect 532102 -7622 532186 -7386
rect 532422 -7622 532454 -7386
rect 531834 -7654 532454 -7622
rect 541794 75454 542414 110898
rect 542678 88501 542738 311067
rect 545514 295174 546134 330618
rect 545514 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 546134 295174
rect 545514 294854 546134 294938
rect 545514 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 546134 294854
rect 545514 259174 546134 294618
rect 545514 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 546134 259174
rect 545514 258854 546134 258938
rect 545514 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 546134 258854
rect 545514 223174 546134 258618
rect 545514 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 546134 223174
rect 545514 222854 546134 222938
rect 545514 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 546134 222854
rect 545514 187174 546134 222618
rect 545514 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 546134 187174
rect 545514 186854 546134 186938
rect 545514 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 546134 186854
rect 545514 151174 546134 186618
rect 545514 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 546134 151174
rect 545514 150854 546134 150938
rect 545514 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 546134 150854
rect 545514 115174 546134 150618
rect 545514 114938 545546 115174
rect 545782 114938 545866 115174
rect 546102 114938 546134 115174
rect 545514 114854 546134 114938
rect 545514 114618 545546 114854
rect 545782 114618 545866 114854
rect 546102 114618 546134 114854
rect 542675 88500 542741 88501
rect 542675 88436 542676 88500
rect 542740 88436 542741 88500
rect 542675 88435 542741 88436
rect 541794 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 542414 75454
rect 541794 75134 542414 75218
rect 541794 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 542414 75134
rect 541794 39454 542414 74898
rect 545514 79174 546134 114618
rect 545514 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 546134 79174
rect 545514 78854 546134 78938
rect 545514 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 546134 78854
rect 545514 51692 546134 78618
rect 549234 406894 549854 442338
rect 552954 707718 553574 711590
rect 552954 707482 552986 707718
rect 553222 707482 553306 707718
rect 553542 707482 553574 707718
rect 552954 707398 553574 707482
rect 552954 707162 552986 707398
rect 553222 707162 553306 707398
rect 553542 707162 553574 707398
rect 552954 698614 553574 707162
rect 552954 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 553574 698614
rect 552954 698294 553574 698378
rect 552954 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 553574 698294
rect 552954 662614 553574 698058
rect 552954 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 553574 662614
rect 552954 662294 553574 662378
rect 552954 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 553574 662294
rect 552954 626614 553574 662058
rect 552954 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 553574 626614
rect 552954 626294 553574 626378
rect 552954 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 553574 626294
rect 552954 590614 553574 626058
rect 552954 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 553574 590614
rect 552954 590294 553574 590378
rect 552954 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 553574 590294
rect 552954 554614 553574 590058
rect 552954 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 553574 554614
rect 552954 554294 553574 554378
rect 552954 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 553574 554294
rect 552954 518614 553574 554058
rect 552954 518378 552986 518614
rect 553222 518378 553306 518614
rect 553542 518378 553574 518614
rect 552954 518294 553574 518378
rect 552954 518058 552986 518294
rect 553222 518058 553306 518294
rect 553542 518058 553574 518294
rect 552954 482614 553574 518058
rect 552954 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 553574 482614
rect 552954 482294 553574 482378
rect 552954 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 553574 482294
rect 552954 446614 553574 482058
rect 552954 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 553574 446614
rect 552954 446294 553574 446378
rect 552954 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 553574 446294
rect 550487 435454 550807 435486
rect 550487 435218 550529 435454
rect 550765 435218 550807 435454
rect 550487 435134 550807 435218
rect 550487 434898 550529 435134
rect 550765 434898 550807 435134
rect 550487 434866 550807 434898
rect 549234 406658 549266 406894
rect 549502 406658 549586 406894
rect 549822 406658 549854 406894
rect 549234 406574 549854 406658
rect 549234 406338 549266 406574
rect 549502 406338 549586 406574
rect 549822 406338 549854 406574
rect 549234 370894 549854 406338
rect 552954 410614 553574 446058
rect 556674 708678 557294 711590
rect 556674 708442 556706 708678
rect 556942 708442 557026 708678
rect 557262 708442 557294 708678
rect 556674 708358 557294 708442
rect 556674 708122 556706 708358
rect 556942 708122 557026 708358
rect 557262 708122 557294 708358
rect 556674 666334 557294 708122
rect 560394 709638 561014 711590
rect 560394 709402 560426 709638
rect 560662 709402 560746 709638
rect 560982 709402 561014 709638
rect 560394 709318 561014 709402
rect 560394 709082 560426 709318
rect 560662 709082 560746 709318
rect 560982 709082 561014 709318
rect 558131 699820 558197 699821
rect 558131 699756 558132 699820
rect 558196 699756 558197 699820
rect 558131 699755 558197 699756
rect 556674 666098 556706 666334
rect 556942 666098 557026 666334
rect 557262 666098 557294 666334
rect 556674 666014 557294 666098
rect 556674 665778 556706 666014
rect 556942 665778 557026 666014
rect 557262 665778 557294 666014
rect 556674 630334 557294 665778
rect 556674 630098 556706 630334
rect 556942 630098 557026 630334
rect 557262 630098 557294 630334
rect 556674 630014 557294 630098
rect 556674 629778 556706 630014
rect 556942 629778 557026 630014
rect 557262 629778 557294 630014
rect 556674 594334 557294 629778
rect 556674 594098 556706 594334
rect 556942 594098 557026 594334
rect 557262 594098 557294 594334
rect 556674 594014 557294 594098
rect 556674 593778 556706 594014
rect 556942 593778 557026 594014
rect 557262 593778 557294 594014
rect 556674 558334 557294 593778
rect 556674 558098 556706 558334
rect 556942 558098 557026 558334
rect 557262 558098 557294 558334
rect 556674 558014 557294 558098
rect 556674 557778 556706 558014
rect 556942 557778 557026 558014
rect 557262 557778 557294 558014
rect 556674 522334 557294 557778
rect 556674 522098 556706 522334
rect 556942 522098 557026 522334
rect 557262 522098 557294 522334
rect 556674 522014 557294 522098
rect 556674 521778 556706 522014
rect 556942 521778 557026 522014
rect 557262 521778 557294 522014
rect 556674 486334 557294 521778
rect 556674 486098 556706 486334
rect 556942 486098 557026 486334
rect 557262 486098 557294 486334
rect 556674 486014 557294 486098
rect 556674 485778 556706 486014
rect 556942 485778 557026 486014
rect 557262 485778 557294 486014
rect 556674 450334 557294 485778
rect 556674 450098 556706 450334
rect 556942 450098 557026 450334
rect 557262 450098 557294 450334
rect 556674 450014 557294 450098
rect 556674 449778 556706 450014
rect 556942 449778 557026 450014
rect 557262 449778 557294 450014
rect 554707 439174 555027 439206
rect 554707 438938 554749 439174
rect 554985 438938 555027 439174
rect 554707 438854 555027 438938
rect 554707 438618 554749 438854
rect 554985 438618 555027 438854
rect 554707 438586 555027 438618
rect 552954 410378 552986 410614
rect 553222 410378 553306 410614
rect 553542 410378 553574 410614
rect 552954 410294 553574 410378
rect 552954 410058 552986 410294
rect 553222 410058 553306 410294
rect 553542 410058 553574 410294
rect 552954 377884 553574 410058
rect 556674 414334 557294 449778
rect 556674 414098 556706 414334
rect 556942 414098 557026 414334
rect 557262 414098 557294 414334
rect 556674 414014 557294 414098
rect 556674 413778 556706 414014
rect 556942 413778 557026 414014
rect 557262 413778 557294 414014
rect 556674 378243 557294 413778
rect 556674 378007 556706 378243
rect 556942 378007 557026 378243
rect 557262 378007 557294 378243
rect 556674 377884 557294 378007
rect 549234 370658 549266 370894
rect 549502 370658 549586 370894
rect 549822 370658 549854 370894
rect 549234 370574 549854 370658
rect 549234 370338 549266 370574
rect 549502 370338 549586 370574
rect 549822 370338 549854 370574
rect 549234 334894 549854 370338
rect 554876 367174 555196 367206
rect 554876 366938 554918 367174
rect 555154 366938 555196 367174
rect 554876 366854 555196 366938
rect 554876 366618 554918 366854
rect 555154 366618 555196 366854
rect 554876 366586 555196 366618
rect 552910 363454 553230 363486
rect 552910 363218 552952 363454
rect 553188 363218 553230 363454
rect 552910 363134 553230 363218
rect 552910 362898 552952 363134
rect 553188 362898 553230 363134
rect 552910 362866 553230 362898
rect 556843 363454 557163 363486
rect 556843 363218 556885 363454
rect 557121 363218 557163 363454
rect 556843 363134 557163 363218
rect 556843 362898 556885 363134
rect 557121 362898 557163 363134
rect 556843 362866 557163 362898
rect 549234 334658 549266 334894
rect 549502 334658 549586 334894
rect 549822 334658 549854 334894
rect 549234 334574 549854 334658
rect 549234 334338 549266 334574
rect 549502 334338 549586 334574
rect 549822 334338 549854 334574
rect 549234 298894 549854 334338
rect 549234 298658 549266 298894
rect 549502 298658 549586 298894
rect 549822 298658 549854 298894
rect 549234 298574 549854 298658
rect 549234 298338 549266 298574
rect 549502 298338 549586 298574
rect 549822 298338 549854 298574
rect 549234 262894 549854 298338
rect 549234 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 549854 262894
rect 549234 262574 549854 262658
rect 549234 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 549854 262574
rect 549234 226894 549854 262338
rect 549234 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 549854 226894
rect 549234 226574 549854 226658
rect 549234 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 549854 226574
rect 549234 190894 549854 226338
rect 549234 190658 549266 190894
rect 549502 190658 549586 190894
rect 549822 190658 549854 190894
rect 549234 190574 549854 190658
rect 549234 190338 549266 190574
rect 549502 190338 549586 190574
rect 549822 190338 549854 190574
rect 549234 154894 549854 190338
rect 549234 154658 549266 154894
rect 549502 154658 549586 154894
rect 549822 154658 549854 154894
rect 549234 154574 549854 154658
rect 549234 154338 549266 154574
rect 549502 154338 549586 154574
rect 549822 154338 549854 154574
rect 549234 118894 549854 154338
rect 549234 118658 549266 118894
rect 549502 118658 549586 118894
rect 549822 118658 549854 118894
rect 549234 118574 549854 118658
rect 549234 118338 549266 118574
rect 549502 118338 549586 118574
rect 549822 118338 549854 118574
rect 549234 82894 549854 118338
rect 549234 82658 549266 82894
rect 549502 82658 549586 82894
rect 549822 82658 549854 82894
rect 549234 82574 549854 82658
rect 549234 82338 549266 82574
rect 549502 82338 549586 82574
rect 549822 82338 549854 82574
rect 549234 46894 549854 82338
rect 552954 338614 553574 360068
rect 552954 338378 552986 338614
rect 553222 338378 553306 338614
rect 553542 338378 553574 338614
rect 552954 338294 553574 338378
rect 552954 338058 552986 338294
rect 553222 338058 553306 338294
rect 553542 338058 553574 338294
rect 552954 302614 553574 338058
rect 552954 302378 552986 302614
rect 553222 302378 553306 302614
rect 553542 302378 553574 302614
rect 552954 302294 553574 302378
rect 552954 302058 552986 302294
rect 553222 302058 553306 302294
rect 553542 302058 553574 302294
rect 552954 266614 553574 302058
rect 552954 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 553574 266614
rect 552954 266294 553574 266378
rect 552954 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 553574 266294
rect 552954 230614 553574 266058
rect 552954 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 553574 230614
rect 552954 230294 553574 230378
rect 552954 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 553574 230294
rect 552954 194614 553574 230058
rect 552954 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 553574 194614
rect 552954 194294 553574 194378
rect 552954 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 553574 194294
rect 552954 158614 553574 194058
rect 552954 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 553574 158614
rect 552954 158294 553574 158378
rect 552954 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 553574 158294
rect 552954 122614 553574 158058
rect 552954 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 553574 122614
rect 552954 122294 553574 122378
rect 552954 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 553574 122294
rect 552954 86614 553574 122058
rect 552954 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 553574 86614
rect 552954 86294 553574 86378
rect 552954 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 553574 86294
rect 552954 51692 553574 86058
rect 556674 342334 557294 360068
rect 556674 342098 556706 342334
rect 556942 342098 557026 342334
rect 557262 342098 557294 342334
rect 556674 342014 557294 342098
rect 556674 341778 556706 342014
rect 556942 341778 557026 342014
rect 557262 341778 557294 342014
rect 556674 306334 557294 341778
rect 558134 320653 558194 699755
rect 560394 670054 561014 709082
rect 560394 669818 560426 670054
rect 560662 669818 560746 670054
rect 560982 669818 561014 670054
rect 560394 669734 561014 669818
rect 560394 669498 560426 669734
rect 560662 669498 560746 669734
rect 560982 669498 561014 669734
rect 560394 634054 561014 669498
rect 560394 633818 560426 634054
rect 560662 633818 560746 634054
rect 560982 633818 561014 634054
rect 560394 633734 561014 633818
rect 560394 633498 560426 633734
rect 560662 633498 560746 633734
rect 560982 633498 561014 633734
rect 560394 598054 561014 633498
rect 560394 597818 560426 598054
rect 560662 597818 560746 598054
rect 560982 597818 561014 598054
rect 560394 597734 561014 597818
rect 560394 597498 560426 597734
rect 560662 597498 560746 597734
rect 560982 597498 561014 597734
rect 560394 562054 561014 597498
rect 560394 561818 560426 562054
rect 560662 561818 560746 562054
rect 560982 561818 561014 562054
rect 560394 561734 561014 561818
rect 560394 561498 560426 561734
rect 560662 561498 560746 561734
rect 560982 561498 561014 561734
rect 560394 526054 561014 561498
rect 560394 525818 560426 526054
rect 560662 525818 560746 526054
rect 560982 525818 561014 526054
rect 560394 525734 561014 525818
rect 560394 525498 560426 525734
rect 560662 525498 560746 525734
rect 560982 525498 561014 525734
rect 560394 490054 561014 525498
rect 560394 489818 560426 490054
rect 560662 489818 560746 490054
rect 560982 489818 561014 490054
rect 560394 489734 561014 489818
rect 560394 489498 560426 489734
rect 560662 489498 560746 489734
rect 560982 489498 561014 489734
rect 560394 454054 561014 489498
rect 560394 453818 560426 454054
rect 560662 453818 560746 454054
rect 560982 453818 561014 454054
rect 560394 453734 561014 453818
rect 560394 453498 560426 453734
rect 560662 453498 560746 453734
rect 560982 453498 561014 453734
rect 560394 418054 561014 453498
rect 560394 417818 560426 418054
rect 560662 417818 560746 418054
rect 560982 417818 561014 418054
rect 560394 417734 561014 417818
rect 560394 417498 560426 417734
rect 560662 417498 560746 417734
rect 560982 417498 561014 417734
rect 560394 382054 561014 417498
rect 560394 381818 560426 382054
rect 560662 381818 560746 382054
rect 560982 381818 561014 382054
rect 560394 381734 561014 381818
rect 560394 381498 560426 381734
rect 560662 381498 560746 381734
rect 560982 381498 561014 381734
rect 560394 377884 561014 381498
rect 564114 710598 564734 711590
rect 564114 710362 564146 710598
rect 564382 710362 564466 710598
rect 564702 710362 564734 710598
rect 564114 710278 564734 710362
rect 564114 710042 564146 710278
rect 564382 710042 564466 710278
rect 564702 710042 564734 710278
rect 564114 673774 564734 710042
rect 564114 673538 564146 673774
rect 564382 673538 564466 673774
rect 564702 673538 564734 673774
rect 564114 673454 564734 673538
rect 564114 673218 564146 673454
rect 564382 673218 564466 673454
rect 564702 673218 564734 673454
rect 564114 637774 564734 673218
rect 564114 637538 564146 637774
rect 564382 637538 564466 637774
rect 564702 637538 564734 637774
rect 564114 637454 564734 637538
rect 564114 637218 564146 637454
rect 564382 637218 564466 637454
rect 564702 637218 564734 637454
rect 564114 601774 564734 637218
rect 564114 601538 564146 601774
rect 564382 601538 564466 601774
rect 564702 601538 564734 601774
rect 564114 601454 564734 601538
rect 564114 601218 564146 601454
rect 564382 601218 564466 601454
rect 564702 601218 564734 601454
rect 564114 565774 564734 601218
rect 564114 565538 564146 565774
rect 564382 565538 564466 565774
rect 564702 565538 564734 565774
rect 564114 565454 564734 565538
rect 564114 565218 564146 565454
rect 564382 565218 564466 565454
rect 564702 565218 564734 565454
rect 564114 529774 564734 565218
rect 564114 529538 564146 529774
rect 564382 529538 564466 529774
rect 564702 529538 564734 529774
rect 564114 529454 564734 529538
rect 564114 529218 564146 529454
rect 564382 529218 564466 529454
rect 564702 529218 564734 529454
rect 564114 493774 564734 529218
rect 564114 493538 564146 493774
rect 564382 493538 564466 493774
rect 564702 493538 564734 493774
rect 564114 493454 564734 493538
rect 564114 493218 564146 493454
rect 564382 493218 564466 493454
rect 564702 493218 564734 493454
rect 564114 457774 564734 493218
rect 564114 457538 564146 457774
rect 564382 457538 564466 457774
rect 564702 457538 564734 457774
rect 564114 457454 564734 457538
rect 564114 457218 564146 457454
rect 564382 457218 564466 457454
rect 564702 457218 564734 457454
rect 564114 421774 564734 457218
rect 564114 421538 564146 421774
rect 564382 421538 564466 421774
rect 564702 421538 564734 421774
rect 564114 421454 564734 421538
rect 564114 421218 564146 421454
rect 564382 421218 564466 421454
rect 564702 421218 564734 421454
rect 564114 385774 564734 421218
rect 564114 385538 564146 385774
rect 564382 385538 564466 385774
rect 564702 385538 564734 385774
rect 564114 385454 564734 385538
rect 564114 385218 564146 385454
rect 564382 385218 564466 385454
rect 564702 385218 564734 385454
rect 564114 377884 564734 385218
rect 567834 711558 568454 711590
rect 567834 711322 567866 711558
rect 568102 711322 568186 711558
rect 568422 711322 568454 711558
rect 567834 711238 568454 711322
rect 567834 711002 567866 711238
rect 568102 711002 568186 711238
rect 568422 711002 568454 711238
rect 567834 677494 568454 711002
rect 567834 677258 567866 677494
rect 568102 677258 568186 677494
rect 568422 677258 568454 677494
rect 567834 677174 568454 677258
rect 567834 676938 567866 677174
rect 568102 676938 568186 677174
rect 568422 676938 568454 677174
rect 567834 641494 568454 676938
rect 567834 641258 567866 641494
rect 568102 641258 568186 641494
rect 568422 641258 568454 641494
rect 567834 641174 568454 641258
rect 567834 640938 567866 641174
rect 568102 640938 568186 641174
rect 568422 640938 568454 641174
rect 567834 605494 568454 640938
rect 567834 605258 567866 605494
rect 568102 605258 568186 605494
rect 568422 605258 568454 605494
rect 567834 605174 568454 605258
rect 567834 604938 567866 605174
rect 568102 604938 568186 605174
rect 568422 604938 568454 605174
rect 567834 569494 568454 604938
rect 567834 569258 567866 569494
rect 568102 569258 568186 569494
rect 568422 569258 568454 569494
rect 567834 569174 568454 569258
rect 567834 568938 567866 569174
rect 568102 568938 568186 569174
rect 568422 568938 568454 569174
rect 567834 533494 568454 568938
rect 567834 533258 567866 533494
rect 568102 533258 568186 533494
rect 568422 533258 568454 533494
rect 567834 533174 568454 533258
rect 567834 532938 567866 533174
rect 568102 532938 568186 533174
rect 568422 532938 568454 533174
rect 567834 497494 568454 532938
rect 567834 497258 567866 497494
rect 568102 497258 568186 497494
rect 568422 497258 568454 497494
rect 567834 497174 568454 497258
rect 567834 496938 567866 497174
rect 568102 496938 568186 497174
rect 568422 496938 568454 497174
rect 567834 461494 568454 496938
rect 567834 461258 567866 461494
rect 568102 461258 568186 461494
rect 568422 461258 568454 461494
rect 567834 461174 568454 461258
rect 567834 460938 567866 461174
rect 568102 460938 568186 461174
rect 568422 460938 568454 461174
rect 567834 425494 568454 460938
rect 567834 425258 567866 425494
rect 568102 425258 568186 425494
rect 568422 425258 568454 425494
rect 567834 425174 568454 425258
rect 567834 424938 567866 425174
rect 568102 424938 568186 425174
rect 568422 424938 568454 425174
rect 567834 389494 568454 424938
rect 567834 389258 567866 389494
rect 568102 389258 568186 389494
rect 568422 389258 568454 389494
rect 567834 389174 568454 389258
rect 567834 388938 567866 389174
rect 568102 388938 568186 389174
rect 568422 388938 568454 389174
rect 558809 367174 559129 367206
rect 558809 366938 558851 367174
rect 559087 366938 559129 367174
rect 558809 366854 559129 366938
rect 558809 366618 558851 366854
rect 559087 366618 559129 366854
rect 558809 366586 559129 366618
rect 562742 367174 563062 367206
rect 562742 366938 562784 367174
rect 563020 366938 563062 367174
rect 562742 366854 563062 366938
rect 562742 366618 562784 366854
rect 563020 366618 563062 366854
rect 562742 366586 563062 366618
rect 566675 367174 566995 367206
rect 566675 366938 566717 367174
rect 566953 366938 566995 367174
rect 566675 366854 566995 366938
rect 566675 366618 566717 366854
rect 566953 366618 566995 366854
rect 566675 366586 566995 366618
rect 560776 363454 561096 363486
rect 560776 363218 560818 363454
rect 561054 363218 561096 363454
rect 560776 363134 561096 363218
rect 560776 362898 560818 363134
rect 561054 362898 561096 363134
rect 560776 362866 561096 362898
rect 564709 363454 565029 363486
rect 564709 363218 564751 363454
rect 564987 363218 565029 363454
rect 564709 363134 565029 363218
rect 564709 362898 564751 363134
rect 564987 362898 565029 363134
rect 564709 362866 565029 362898
rect 560394 346054 561014 360068
rect 560394 345818 560426 346054
rect 560662 345818 560746 346054
rect 560982 345818 561014 346054
rect 560394 345734 561014 345818
rect 560394 345498 560426 345734
rect 560662 345498 560746 345734
rect 560982 345498 561014 345734
rect 558131 320652 558197 320653
rect 558131 320588 558132 320652
rect 558196 320588 558197 320652
rect 558131 320587 558197 320588
rect 556674 306098 556706 306334
rect 556942 306098 557026 306334
rect 557262 306098 557294 306334
rect 556674 306014 557294 306098
rect 556674 305778 556706 306014
rect 556942 305778 557026 306014
rect 557262 305778 557294 306014
rect 556674 270334 557294 305778
rect 556674 270098 556706 270334
rect 556942 270098 557026 270334
rect 557262 270098 557294 270334
rect 556674 270014 557294 270098
rect 556674 269778 556706 270014
rect 556942 269778 557026 270014
rect 557262 269778 557294 270014
rect 556674 234334 557294 269778
rect 556674 234098 556706 234334
rect 556942 234098 557026 234334
rect 557262 234098 557294 234334
rect 556674 234014 557294 234098
rect 556674 233778 556706 234014
rect 556942 233778 557026 234014
rect 557262 233778 557294 234014
rect 556674 198334 557294 233778
rect 556674 198098 556706 198334
rect 556942 198098 557026 198334
rect 557262 198098 557294 198334
rect 556674 198014 557294 198098
rect 556674 197778 556706 198014
rect 556942 197778 557026 198014
rect 557262 197778 557294 198014
rect 556674 162334 557294 197778
rect 556674 162098 556706 162334
rect 556942 162098 557026 162334
rect 557262 162098 557294 162334
rect 556674 162014 557294 162098
rect 556674 161778 556706 162014
rect 556942 161778 557026 162014
rect 557262 161778 557294 162014
rect 556674 126334 557294 161778
rect 556674 126098 556706 126334
rect 556942 126098 557026 126334
rect 557262 126098 557294 126334
rect 556674 126014 557294 126098
rect 556674 125778 556706 126014
rect 556942 125778 557026 126014
rect 557262 125778 557294 126014
rect 556674 90334 557294 125778
rect 556674 90098 556706 90334
rect 556942 90098 557026 90334
rect 557262 90098 557294 90334
rect 556674 90014 557294 90098
rect 556674 89778 556706 90014
rect 556942 89778 557026 90014
rect 557262 89778 557294 90014
rect 556674 54334 557294 89778
rect 556674 54098 556706 54334
rect 556942 54098 557026 54334
rect 557262 54098 557294 54334
rect 556674 54014 557294 54098
rect 556674 53778 556706 54014
rect 556942 53778 557026 54014
rect 557262 53778 557294 54014
rect 549234 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 549854 46894
rect 549234 46574 549854 46658
rect 549234 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 549854 46574
rect 545888 43174 546208 43206
rect 545888 42938 545930 43174
rect 546166 42938 546208 43174
rect 545888 42854 546208 42938
rect 545888 42618 545930 42854
rect 546166 42618 546208 42854
rect 545888 42586 546208 42618
rect 541794 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 542414 39454
rect 541794 39134 542414 39218
rect 541794 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 542414 39134
rect 541794 3454 542414 38898
rect 543416 39454 543736 39486
rect 543416 39218 543458 39454
rect 543694 39218 543736 39454
rect 543416 39134 543736 39218
rect 543416 38898 543458 39134
rect 543694 38898 543736 39134
rect 543416 38866 543736 38898
rect 548361 39454 548681 39486
rect 548361 39218 548403 39454
rect 548639 39218 548681 39454
rect 548361 39134 548681 39218
rect 548361 38898 548403 39134
rect 548639 38898 548681 39134
rect 548361 38866 548681 38898
rect 541794 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 542414 3454
rect 541794 3134 542414 3218
rect 541794 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 542414 3134
rect 541794 -346 542414 2898
rect 541794 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 542414 -346
rect 541794 -666 542414 -582
rect 541794 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 542414 -666
rect 541794 -7654 542414 -902
rect 545514 7174 546134 30068
rect 545514 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 546134 7174
rect 545514 6854 546134 6938
rect 545514 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 546134 6854
rect 545514 -1306 546134 6618
rect 545514 -1542 545546 -1306
rect 545782 -1542 545866 -1306
rect 546102 -1542 546134 -1306
rect 545514 -1626 546134 -1542
rect 545514 -1862 545546 -1626
rect 545782 -1862 545866 -1626
rect 546102 -1862 546134 -1626
rect 545514 -7654 546134 -1862
rect 549234 10894 549854 46338
rect 550833 43174 551153 43206
rect 550833 42938 550875 43174
rect 551111 42938 551153 43174
rect 550833 42854 551153 42938
rect 550833 42618 550875 42854
rect 551111 42618 551153 42854
rect 550833 42586 551153 42618
rect 555778 43174 556098 43206
rect 555778 42938 555820 43174
rect 556056 42938 556098 43174
rect 555778 42854 556098 42938
rect 555778 42618 555820 42854
rect 556056 42618 556098 42854
rect 555778 42586 556098 42618
rect 553306 39454 553626 39486
rect 553306 39218 553348 39454
rect 553584 39218 553626 39454
rect 553306 39134 553626 39218
rect 553306 38898 553348 39134
rect 553584 38898 553626 39134
rect 553306 38866 553626 38898
rect 549234 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 549854 10894
rect 549234 10574 549854 10658
rect 549234 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 549854 10574
rect 549234 -2266 549854 10338
rect 549234 -2502 549266 -2266
rect 549502 -2502 549586 -2266
rect 549822 -2502 549854 -2266
rect 549234 -2586 549854 -2502
rect 549234 -2822 549266 -2586
rect 549502 -2822 549586 -2586
rect 549822 -2822 549854 -2586
rect 549234 -7654 549854 -2822
rect 552954 14614 553574 30068
rect 552954 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 553574 14614
rect 552954 14294 553574 14378
rect 552954 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 553574 14294
rect 552954 -3226 553574 14058
rect 552954 -3462 552986 -3226
rect 553222 -3462 553306 -3226
rect 553542 -3462 553574 -3226
rect 552954 -3546 553574 -3462
rect 552954 -3782 552986 -3546
rect 553222 -3782 553306 -3546
rect 553542 -3782 553574 -3546
rect 552954 -7654 553574 -3782
rect 556674 18334 557294 53778
rect 560394 310054 561014 345498
rect 560394 309818 560426 310054
rect 560662 309818 560746 310054
rect 560982 309818 561014 310054
rect 560394 309734 561014 309818
rect 560394 309498 560426 309734
rect 560662 309498 560746 309734
rect 560982 309498 561014 309734
rect 560394 274054 561014 309498
rect 560394 273818 560426 274054
rect 560662 273818 560746 274054
rect 560982 273818 561014 274054
rect 560394 273734 561014 273818
rect 560394 273498 560426 273734
rect 560662 273498 560746 273734
rect 560982 273498 561014 273734
rect 560394 238054 561014 273498
rect 560394 237818 560426 238054
rect 560662 237818 560746 238054
rect 560982 237818 561014 238054
rect 560394 237734 561014 237818
rect 560394 237498 560426 237734
rect 560662 237498 560746 237734
rect 560982 237498 561014 237734
rect 560394 202054 561014 237498
rect 560394 201818 560426 202054
rect 560662 201818 560746 202054
rect 560982 201818 561014 202054
rect 560394 201734 561014 201818
rect 560394 201498 560426 201734
rect 560662 201498 560746 201734
rect 560982 201498 561014 201734
rect 560394 166054 561014 201498
rect 560394 165818 560426 166054
rect 560662 165818 560746 166054
rect 560982 165818 561014 166054
rect 560394 165734 561014 165818
rect 560394 165498 560426 165734
rect 560662 165498 560746 165734
rect 560982 165498 561014 165734
rect 560394 130054 561014 165498
rect 560394 129818 560426 130054
rect 560662 129818 560746 130054
rect 560982 129818 561014 130054
rect 560394 129734 561014 129818
rect 560394 129498 560426 129734
rect 560662 129498 560746 129734
rect 560982 129498 561014 129734
rect 560394 94054 561014 129498
rect 560394 93818 560426 94054
rect 560662 93818 560746 94054
rect 560982 93818 561014 94054
rect 560394 93734 561014 93818
rect 560394 93498 560426 93734
rect 560662 93498 560746 93734
rect 560982 93498 561014 93734
rect 560394 58054 561014 93498
rect 560394 57818 560426 58054
rect 560662 57818 560746 58054
rect 560982 57818 561014 58054
rect 560394 57734 561014 57818
rect 560394 57498 560426 57734
rect 560662 57498 560746 57734
rect 560982 57498 561014 57734
rect 560394 51692 561014 57498
rect 564114 349774 564734 360068
rect 564114 349538 564146 349774
rect 564382 349538 564466 349774
rect 564702 349538 564734 349774
rect 564114 349454 564734 349538
rect 564114 349218 564146 349454
rect 564382 349218 564466 349454
rect 564702 349218 564734 349454
rect 564114 313774 564734 349218
rect 564114 313538 564146 313774
rect 564382 313538 564466 313774
rect 564702 313538 564734 313774
rect 564114 313454 564734 313538
rect 564114 313218 564146 313454
rect 564382 313218 564466 313454
rect 564702 313218 564734 313454
rect 564114 277774 564734 313218
rect 564114 277538 564146 277774
rect 564382 277538 564466 277774
rect 564702 277538 564734 277774
rect 564114 277454 564734 277538
rect 564114 277218 564146 277454
rect 564382 277218 564466 277454
rect 564702 277218 564734 277454
rect 564114 241774 564734 277218
rect 564114 241538 564146 241774
rect 564382 241538 564466 241774
rect 564702 241538 564734 241774
rect 564114 241454 564734 241538
rect 564114 241218 564146 241454
rect 564382 241218 564466 241454
rect 564702 241218 564734 241454
rect 564114 205774 564734 241218
rect 564114 205538 564146 205774
rect 564382 205538 564466 205774
rect 564702 205538 564734 205774
rect 564114 205454 564734 205538
rect 564114 205218 564146 205454
rect 564382 205218 564466 205454
rect 564702 205218 564734 205454
rect 564114 169774 564734 205218
rect 564114 169538 564146 169774
rect 564382 169538 564466 169774
rect 564702 169538 564734 169774
rect 564114 169454 564734 169538
rect 564114 169218 564146 169454
rect 564382 169218 564466 169454
rect 564702 169218 564734 169454
rect 564114 133774 564734 169218
rect 564114 133538 564146 133774
rect 564382 133538 564466 133774
rect 564702 133538 564734 133774
rect 564114 133454 564734 133538
rect 564114 133218 564146 133454
rect 564382 133218 564466 133454
rect 564702 133218 564734 133454
rect 564114 97774 564734 133218
rect 564114 97538 564146 97774
rect 564382 97538 564466 97774
rect 564702 97538 564734 97774
rect 564114 97454 564734 97538
rect 564114 97218 564146 97454
rect 564382 97218 564466 97454
rect 564702 97218 564734 97454
rect 564114 61774 564734 97218
rect 564114 61538 564146 61774
rect 564382 61538 564466 61774
rect 564702 61538 564734 61774
rect 564114 61454 564734 61538
rect 564114 61218 564146 61454
rect 564382 61218 564466 61454
rect 564702 61218 564734 61454
rect 560723 43174 561043 43206
rect 560723 42938 560765 43174
rect 561001 42938 561043 43174
rect 560723 42854 561043 42938
rect 560723 42618 560765 42854
rect 561001 42618 561043 42854
rect 560723 42586 561043 42618
rect 558251 39454 558571 39486
rect 558251 39218 558293 39454
rect 558529 39218 558571 39454
rect 558251 39134 558571 39218
rect 558251 38898 558293 39134
rect 558529 38898 558571 39134
rect 558251 38866 558571 38898
rect 556674 18098 556706 18334
rect 556942 18098 557026 18334
rect 557262 18098 557294 18334
rect 556674 18014 557294 18098
rect 556674 17778 556706 18014
rect 556942 17778 557026 18014
rect 557262 17778 557294 18014
rect 556674 -4186 557294 17778
rect 556674 -4422 556706 -4186
rect 556942 -4422 557026 -4186
rect 557262 -4422 557294 -4186
rect 556674 -4506 557294 -4422
rect 556674 -4742 556706 -4506
rect 556942 -4742 557026 -4506
rect 557262 -4742 557294 -4506
rect 556674 -7654 557294 -4742
rect 560394 22054 561014 30068
rect 560394 21818 560426 22054
rect 560662 21818 560746 22054
rect 560982 21818 561014 22054
rect 560394 21734 561014 21818
rect 560394 21498 560426 21734
rect 560662 21498 560746 21734
rect 560982 21498 561014 21734
rect 560394 -5146 561014 21498
rect 560394 -5382 560426 -5146
rect 560662 -5382 560746 -5146
rect 560982 -5382 561014 -5146
rect 560394 -5466 561014 -5382
rect 560394 -5702 560426 -5466
rect 560662 -5702 560746 -5466
rect 560982 -5702 561014 -5466
rect 560394 -7654 561014 -5702
rect 564114 25774 564734 61218
rect 564114 25538 564146 25774
rect 564382 25538 564466 25774
rect 564702 25538 564734 25774
rect 564114 25454 564734 25538
rect 564114 25218 564146 25454
rect 564382 25218 564466 25454
rect 564702 25218 564734 25454
rect 564114 -6106 564734 25218
rect 564114 -6342 564146 -6106
rect 564382 -6342 564466 -6106
rect 564702 -6342 564734 -6106
rect 564114 -6426 564734 -6342
rect 564114 -6662 564146 -6426
rect 564382 -6662 564466 -6426
rect 564702 -6662 564734 -6426
rect 564114 -7654 564734 -6662
rect 567834 353494 568454 388938
rect 567834 353258 567866 353494
rect 568102 353258 568186 353494
rect 568422 353258 568454 353494
rect 567834 353174 568454 353258
rect 567834 352938 567866 353174
rect 568102 352938 568186 353174
rect 568422 352938 568454 353174
rect 567834 317494 568454 352938
rect 567834 317258 567866 317494
rect 568102 317258 568186 317494
rect 568422 317258 568454 317494
rect 567834 317174 568454 317258
rect 567834 316938 567866 317174
rect 568102 316938 568186 317174
rect 568422 316938 568454 317174
rect 567834 281494 568454 316938
rect 567834 281258 567866 281494
rect 568102 281258 568186 281494
rect 568422 281258 568454 281494
rect 567834 281174 568454 281258
rect 567834 280938 567866 281174
rect 568102 280938 568186 281174
rect 568422 280938 568454 281174
rect 567834 245494 568454 280938
rect 567834 245258 567866 245494
rect 568102 245258 568186 245494
rect 568422 245258 568454 245494
rect 567834 245174 568454 245258
rect 567834 244938 567866 245174
rect 568102 244938 568186 245174
rect 568422 244938 568454 245174
rect 567834 209494 568454 244938
rect 567834 209258 567866 209494
rect 568102 209258 568186 209494
rect 568422 209258 568454 209494
rect 567834 209174 568454 209258
rect 567834 208938 567866 209174
rect 568102 208938 568186 209174
rect 568422 208938 568454 209174
rect 567834 173494 568454 208938
rect 567834 173258 567866 173494
rect 568102 173258 568186 173494
rect 568422 173258 568454 173494
rect 567834 173174 568454 173258
rect 567834 172938 567866 173174
rect 568102 172938 568186 173174
rect 568422 172938 568454 173174
rect 567834 137494 568454 172938
rect 567834 137258 567866 137494
rect 568102 137258 568186 137494
rect 568422 137258 568454 137494
rect 567834 137174 568454 137258
rect 567834 136938 567866 137174
rect 568102 136938 568186 137174
rect 568422 136938 568454 137174
rect 567834 101494 568454 136938
rect 567834 101258 567866 101494
rect 568102 101258 568186 101494
rect 568422 101258 568454 101494
rect 567834 101174 568454 101258
rect 567834 100938 567866 101174
rect 568102 100938 568186 101174
rect 568422 100938 568454 101174
rect 567834 65494 568454 100938
rect 567834 65258 567866 65494
rect 568102 65258 568186 65494
rect 568422 65258 568454 65494
rect 567834 65174 568454 65258
rect 567834 64938 567866 65174
rect 568102 64938 568186 65174
rect 568422 64938 568454 65174
rect 567834 29494 568454 64938
rect 567834 29258 567866 29494
rect 568102 29258 568186 29494
rect 568422 29258 568454 29494
rect 567834 29174 568454 29258
rect 567834 28938 567866 29174
rect 568102 28938 568186 29174
rect 568422 28938 568454 29174
rect 567834 -7066 568454 28938
rect 567834 -7302 567866 -7066
rect 568102 -7302 568186 -7066
rect 568422 -7302 568454 -7066
rect 567834 -7386 568454 -7302
rect 567834 -7622 567866 -7386
rect 568102 -7622 568186 -7386
rect 568422 -7622 568454 -7386
rect 567834 -7654 568454 -7622
rect 577794 704838 578414 711590
rect 577794 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 578414 704838
rect 577794 704518 578414 704602
rect 577794 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 578414 704518
rect 577794 687454 578414 704282
rect 577794 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 578414 687454
rect 577794 687134 578414 687218
rect 577794 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 578414 687134
rect 577794 651454 578414 686898
rect 577794 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 578414 651454
rect 577794 651134 578414 651218
rect 577794 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 578414 651134
rect 577794 615454 578414 650898
rect 577794 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 578414 615454
rect 577794 615134 578414 615218
rect 577794 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 578414 615134
rect 577794 579454 578414 614898
rect 577794 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 578414 579454
rect 577794 579134 578414 579218
rect 577794 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 578414 579134
rect 577794 543454 578414 578898
rect 577794 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 578414 543454
rect 577794 543134 578414 543218
rect 577794 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 578414 543134
rect 577794 507454 578414 542898
rect 577794 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 578414 507454
rect 577794 507134 578414 507218
rect 577794 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 578414 507134
rect 577794 471454 578414 506898
rect 577794 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 578414 471454
rect 577794 471134 578414 471218
rect 577794 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 578414 471134
rect 577794 435454 578414 470898
rect 577794 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 578414 435454
rect 577794 435134 578414 435218
rect 577794 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 578414 435134
rect 577794 399454 578414 434898
rect 577794 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 578414 399454
rect 577794 399134 578414 399218
rect 577794 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 578414 399134
rect 577794 363454 578414 398898
rect 577794 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 578414 363454
rect 577794 363134 578414 363218
rect 577794 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 578414 363134
rect 577794 327454 578414 362898
rect 577794 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 578414 327454
rect 577794 327134 578414 327218
rect 577794 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 578414 327134
rect 577794 291454 578414 326898
rect 577794 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 578414 291454
rect 577794 291134 578414 291218
rect 577794 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 578414 291134
rect 577794 255454 578414 290898
rect 577794 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 578414 255454
rect 577794 255134 578414 255218
rect 577794 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 578414 255134
rect 577794 219454 578414 254898
rect 577794 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 578414 219454
rect 577794 219134 578414 219218
rect 577794 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 578414 219134
rect 577794 183454 578414 218898
rect 577794 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 578414 183454
rect 577794 183134 578414 183218
rect 577794 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 578414 183134
rect 577794 147454 578414 182898
rect 577794 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 578414 147454
rect 577794 147134 578414 147218
rect 577794 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 578414 147134
rect 577794 111454 578414 146898
rect 577794 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 578414 111454
rect 577794 111134 578414 111218
rect 577794 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 578414 111134
rect 577794 75454 578414 110898
rect 577794 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 578414 75454
rect 577794 75134 578414 75218
rect 577794 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 578414 75134
rect 577794 39454 578414 74898
rect 577794 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 578414 39454
rect 577794 39134 578414 39218
rect 577794 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 578414 39134
rect 577794 3454 578414 38898
rect 577794 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 578414 3454
rect 577794 3134 578414 3218
rect 577794 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 578414 3134
rect 577794 -346 578414 2898
rect 577794 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 578414 -346
rect 577794 -666 578414 -582
rect 577794 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 578414 -666
rect 577794 -7654 578414 -902
rect 581514 705798 582134 711590
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 581514 705562 581546 705798
rect 581782 705562 581866 705798
rect 582102 705562 582134 705798
rect 581514 705478 582134 705562
rect 581514 705242 581546 705478
rect 581782 705242 581866 705478
rect 582102 705242 582134 705478
rect 581514 691174 582134 705242
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 581514 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 582134 691174
rect 581514 690854 582134 690938
rect 581514 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 582134 690854
rect 581514 655174 582134 690618
rect 581514 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 582134 655174
rect 581514 654854 582134 654938
rect 581514 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 582134 654854
rect 581514 619174 582134 654618
rect 581514 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 582134 619174
rect 581514 618854 582134 618938
rect 581514 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 582134 618854
rect 581514 583174 582134 618618
rect 581514 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 582134 583174
rect 581514 582854 582134 582938
rect 581514 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 582134 582854
rect 581514 547174 582134 582618
rect 581514 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 582134 547174
rect 581514 546854 582134 546938
rect 581514 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 582134 546854
rect 581514 511174 582134 546618
rect 581514 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 582134 511174
rect 581514 510854 582134 510938
rect 581514 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 582134 510854
rect 581514 475174 582134 510618
rect 581514 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 582134 475174
rect 581514 474854 582134 474938
rect 581514 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 582134 474854
rect 581514 439174 582134 474618
rect 581514 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 582134 439174
rect 581514 438854 582134 438938
rect 581514 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 582134 438854
rect 581514 403174 582134 438618
rect 581514 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 582134 403174
rect 581514 402854 582134 402938
rect 581514 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 582134 402854
rect 581514 367174 582134 402618
rect 581514 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 582134 367174
rect 581514 366854 582134 366938
rect 581514 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 582134 366854
rect 581514 331174 582134 366618
rect 581514 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 582134 331174
rect 581514 330854 582134 330938
rect 581514 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 582134 330854
rect 581514 295174 582134 330618
rect 581514 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 582134 295174
rect 581514 294854 582134 294938
rect 581514 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 582134 294854
rect 581514 259174 582134 294618
rect 581514 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 582134 259174
rect 581514 258854 582134 258938
rect 581514 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 582134 258854
rect 581514 223174 582134 258618
rect 581514 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 582134 223174
rect 581514 222854 582134 222938
rect 581514 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 582134 222854
rect 581514 187174 582134 222618
rect 581514 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 582134 187174
rect 581514 186854 582134 186938
rect 581514 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 582134 186854
rect 581514 151174 582134 186618
rect 581514 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 582134 151174
rect 581514 150854 582134 150938
rect 581514 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 582134 150854
rect 581514 115174 582134 150618
rect 581514 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 582134 115174
rect 581514 114854 582134 114938
rect 581514 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 582134 114854
rect 581514 79174 582134 114618
rect 581514 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 582134 79174
rect 581514 78854 582134 78938
rect 581514 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 582134 78854
rect 581514 43174 582134 78618
rect 581514 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 582134 43174
rect 581514 42854 582134 42938
rect 581514 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 582134 42854
rect 581514 7174 582134 42618
rect 581514 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 582134 7174
rect 581514 6854 582134 6938
rect 581514 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 582134 6854
rect 581514 -1306 582134 6618
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 687454 585930 704282
rect 585310 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 585930 687454
rect 585310 687134 585930 687218
rect 585310 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 585930 687134
rect 585310 651454 585930 686898
rect 585310 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 585930 651454
rect 585310 651134 585930 651218
rect 585310 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 585930 651134
rect 585310 615454 585930 650898
rect 585310 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 585930 615454
rect 585310 615134 585930 615218
rect 585310 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 585930 615134
rect 585310 579454 585930 614898
rect 585310 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 585930 579454
rect 585310 579134 585930 579218
rect 585310 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 585930 579134
rect 585310 543454 585930 578898
rect 585310 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 585930 543454
rect 585310 543134 585930 543218
rect 585310 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 585930 543134
rect 585310 507454 585930 542898
rect 585310 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 585930 507454
rect 585310 507134 585930 507218
rect 585310 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 585930 507134
rect 585310 471454 585930 506898
rect 585310 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 585930 471454
rect 585310 471134 585930 471218
rect 585310 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 585930 471134
rect 585310 435454 585930 470898
rect 585310 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 585930 435454
rect 585310 435134 585930 435218
rect 585310 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 585930 435134
rect 585310 399454 585930 434898
rect 585310 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 585930 399454
rect 585310 399134 585930 399218
rect 585310 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 585930 399134
rect 585310 363454 585930 398898
rect 585310 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 585930 363454
rect 585310 363134 585930 363218
rect 585310 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 585930 363134
rect 585310 327454 585930 362898
rect 585310 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 585930 327454
rect 585310 327134 585930 327218
rect 585310 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 585930 327134
rect 585310 291454 585930 326898
rect 585310 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 585930 291454
rect 585310 291134 585930 291218
rect 585310 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 585930 291134
rect 585310 255454 585930 290898
rect 585310 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 585930 255454
rect 585310 255134 585930 255218
rect 585310 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 585930 255134
rect 585310 219454 585930 254898
rect 585310 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 585930 219454
rect 585310 219134 585930 219218
rect 585310 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 585930 219134
rect 585310 183454 585930 218898
rect 585310 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 585930 183454
rect 585310 183134 585930 183218
rect 585310 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 585930 183134
rect 585310 147454 585930 182898
rect 585310 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 585930 147454
rect 585310 147134 585930 147218
rect 585310 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 585930 147134
rect 585310 111454 585930 146898
rect 585310 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 585930 111454
rect 585310 111134 585930 111218
rect 585310 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 585930 111134
rect 585310 75454 585930 110898
rect 585310 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 585930 75454
rect 585310 75134 585930 75218
rect 585310 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 585930 75134
rect 585310 39454 585930 74898
rect 585310 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 585930 39454
rect 585310 39134 585930 39218
rect 585310 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 585930 39134
rect 585310 3454 585930 38898
rect 585310 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 585930 3454
rect 585310 3134 585930 3218
rect 585310 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 585930 3134
rect 585310 -346 585930 2898
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 691174 586890 705242
rect 586270 690938 586302 691174
rect 586538 690938 586622 691174
rect 586858 690938 586890 691174
rect 586270 690854 586890 690938
rect 586270 690618 586302 690854
rect 586538 690618 586622 690854
rect 586858 690618 586890 690854
rect 586270 655174 586890 690618
rect 586270 654938 586302 655174
rect 586538 654938 586622 655174
rect 586858 654938 586890 655174
rect 586270 654854 586890 654938
rect 586270 654618 586302 654854
rect 586538 654618 586622 654854
rect 586858 654618 586890 654854
rect 586270 619174 586890 654618
rect 586270 618938 586302 619174
rect 586538 618938 586622 619174
rect 586858 618938 586890 619174
rect 586270 618854 586890 618938
rect 586270 618618 586302 618854
rect 586538 618618 586622 618854
rect 586858 618618 586890 618854
rect 586270 583174 586890 618618
rect 586270 582938 586302 583174
rect 586538 582938 586622 583174
rect 586858 582938 586890 583174
rect 586270 582854 586890 582938
rect 586270 582618 586302 582854
rect 586538 582618 586622 582854
rect 586858 582618 586890 582854
rect 586270 547174 586890 582618
rect 586270 546938 586302 547174
rect 586538 546938 586622 547174
rect 586858 546938 586890 547174
rect 586270 546854 586890 546938
rect 586270 546618 586302 546854
rect 586538 546618 586622 546854
rect 586858 546618 586890 546854
rect 586270 511174 586890 546618
rect 586270 510938 586302 511174
rect 586538 510938 586622 511174
rect 586858 510938 586890 511174
rect 586270 510854 586890 510938
rect 586270 510618 586302 510854
rect 586538 510618 586622 510854
rect 586858 510618 586890 510854
rect 586270 475174 586890 510618
rect 586270 474938 586302 475174
rect 586538 474938 586622 475174
rect 586858 474938 586890 475174
rect 586270 474854 586890 474938
rect 586270 474618 586302 474854
rect 586538 474618 586622 474854
rect 586858 474618 586890 474854
rect 586270 439174 586890 474618
rect 586270 438938 586302 439174
rect 586538 438938 586622 439174
rect 586858 438938 586890 439174
rect 586270 438854 586890 438938
rect 586270 438618 586302 438854
rect 586538 438618 586622 438854
rect 586858 438618 586890 438854
rect 586270 403174 586890 438618
rect 586270 402938 586302 403174
rect 586538 402938 586622 403174
rect 586858 402938 586890 403174
rect 586270 402854 586890 402938
rect 586270 402618 586302 402854
rect 586538 402618 586622 402854
rect 586858 402618 586890 402854
rect 586270 367174 586890 402618
rect 586270 366938 586302 367174
rect 586538 366938 586622 367174
rect 586858 366938 586890 367174
rect 586270 366854 586890 366938
rect 586270 366618 586302 366854
rect 586538 366618 586622 366854
rect 586858 366618 586890 366854
rect 586270 331174 586890 366618
rect 586270 330938 586302 331174
rect 586538 330938 586622 331174
rect 586858 330938 586890 331174
rect 586270 330854 586890 330938
rect 586270 330618 586302 330854
rect 586538 330618 586622 330854
rect 586858 330618 586890 330854
rect 586270 295174 586890 330618
rect 586270 294938 586302 295174
rect 586538 294938 586622 295174
rect 586858 294938 586890 295174
rect 586270 294854 586890 294938
rect 586270 294618 586302 294854
rect 586538 294618 586622 294854
rect 586858 294618 586890 294854
rect 586270 259174 586890 294618
rect 586270 258938 586302 259174
rect 586538 258938 586622 259174
rect 586858 258938 586890 259174
rect 586270 258854 586890 258938
rect 586270 258618 586302 258854
rect 586538 258618 586622 258854
rect 586858 258618 586890 258854
rect 586270 223174 586890 258618
rect 586270 222938 586302 223174
rect 586538 222938 586622 223174
rect 586858 222938 586890 223174
rect 586270 222854 586890 222938
rect 586270 222618 586302 222854
rect 586538 222618 586622 222854
rect 586858 222618 586890 222854
rect 586270 187174 586890 222618
rect 586270 186938 586302 187174
rect 586538 186938 586622 187174
rect 586858 186938 586890 187174
rect 586270 186854 586890 186938
rect 586270 186618 586302 186854
rect 586538 186618 586622 186854
rect 586858 186618 586890 186854
rect 586270 151174 586890 186618
rect 586270 150938 586302 151174
rect 586538 150938 586622 151174
rect 586858 150938 586890 151174
rect 586270 150854 586890 150938
rect 586270 150618 586302 150854
rect 586538 150618 586622 150854
rect 586858 150618 586890 150854
rect 586270 115174 586890 150618
rect 586270 114938 586302 115174
rect 586538 114938 586622 115174
rect 586858 114938 586890 115174
rect 586270 114854 586890 114938
rect 586270 114618 586302 114854
rect 586538 114618 586622 114854
rect 586858 114618 586890 114854
rect 586270 79174 586890 114618
rect 586270 78938 586302 79174
rect 586538 78938 586622 79174
rect 586858 78938 586890 79174
rect 586270 78854 586890 78938
rect 586270 78618 586302 78854
rect 586538 78618 586622 78854
rect 586858 78618 586890 78854
rect 586270 43174 586890 78618
rect 586270 42938 586302 43174
rect 586538 42938 586622 43174
rect 586858 42938 586890 43174
rect 586270 42854 586890 42938
rect 586270 42618 586302 42854
rect 586538 42618 586622 42854
rect 586858 42618 586890 42854
rect 586270 7174 586890 42618
rect 586270 6938 586302 7174
rect 586538 6938 586622 7174
rect 586858 6938 586890 7174
rect 586270 6854 586890 6938
rect 586270 6618 586302 6854
rect 586538 6618 586622 6854
rect 586858 6618 586890 6854
rect 581514 -1542 581546 -1306
rect 581782 -1542 581866 -1306
rect 582102 -1542 582134 -1306
rect 581514 -1626 582134 -1542
rect 581514 -1862 581546 -1626
rect 581782 -1862 581866 -1626
rect 582102 -1862 582134 -1626
rect 581514 -7654 582134 -1862
rect 586270 -1306 586890 6618
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 694894 587850 706202
rect 587230 694658 587262 694894
rect 587498 694658 587582 694894
rect 587818 694658 587850 694894
rect 587230 694574 587850 694658
rect 587230 694338 587262 694574
rect 587498 694338 587582 694574
rect 587818 694338 587850 694574
rect 587230 658894 587850 694338
rect 587230 658658 587262 658894
rect 587498 658658 587582 658894
rect 587818 658658 587850 658894
rect 587230 658574 587850 658658
rect 587230 658338 587262 658574
rect 587498 658338 587582 658574
rect 587818 658338 587850 658574
rect 587230 622894 587850 658338
rect 587230 622658 587262 622894
rect 587498 622658 587582 622894
rect 587818 622658 587850 622894
rect 587230 622574 587850 622658
rect 587230 622338 587262 622574
rect 587498 622338 587582 622574
rect 587818 622338 587850 622574
rect 587230 586894 587850 622338
rect 587230 586658 587262 586894
rect 587498 586658 587582 586894
rect 587818 586658 587850 586894
rect 587230 586574 587850 586658
rect 587230 586338 587262 586574
rect 587498 586338 587582 586574
rect 587818 586338 587850 586574
rect 587230 550894 587850 586338
rect 587230 550658 587262 550894
rect 587498 550658 587582 550894
rect 587818 550658 587850 550894
rect 587230 550574 587850 550658
rect 587230 550338 587262 550574
rect 587498 550338 587582 550574
rect 587818 550338 587850 550574
rect 587230 514894 587850 550338
rect 587230 514658 587262 514894
rect 587498 514658 587582 514894
rect 587818 514658 587850 514894
rect 587230 514574 587850 514658
rect 587230 514338 587262 514574
rect 587498 514338 587582 514574
rect 587818 514338 587850 514574
rect 587230 478894 587850 514338
rect 587230 478658 587262 478894
rect 587498 478658 587582 478894
rect 587818 478658 587850 478894
rect 587230 478574 587850 478658
rect 587230 478338 587262 478574
rect 587498 478338 587582 478574
rect 587818 478338 587850 478574
rect 587230 442894 587850 478338
rect 587230 442658 587262 442894
rect 587498 442658 587582 442894
rect 587818 442658 587850 442894
rect 587230 442574 587850 442658
rect 587230 442338 587262 442574
rect 587498 442338 587582 442574
rect 587818 442338 587850 442574
rect 587230 406894 587850 442338
rect 587230 406658 587262 406894
rect 587498 406658 587582 406894
rect 587818 406658 587850 406894
rect 587230 406574 587850 406658
rect 587230 406338 587262 406574
rect 587498 406338 587582 406574
rect 587818 406338 587850 406574
rect 587230 370894 587850 406338
rect 587230 370658 587262 370894
rect 587498 370658 587582 370894
rect 587818 370658 587850 370894
rect 587230 370574 587850 370658
rect 587230 370338 587262 370574
rect 587498 370338 587582 370574
rect 587818 370338 587850 370574
rect 587230 334894 587850 370338
rect 587230 334658 587262 334894
rect 587498 334658 587582 334894
rect 587818 334658 587850 334894
rect 587230 334574 587850 334658
rect 587230 334338 587262 334574
rect 587498 334338 587582 334574
rect 587818 334338 587850 334574
rect 587230 298894 587850 334338
rect 587230 298658 587262 298894
rect 587498 298658 587582 298894
rect 587818 298658 587850 298894
rect 587230 298574 587850 298658
rect 587230 298338 587262 298574
rect 587498 298338 587582 298574
rect 587818 298338 587850 298574
rect 587230 262894 587850 298338
rect 587230 262658 587262 262894
rect 587498 262658 587582 262894
rect 587818 262658 587850 262894
rect 587230 262574 587850 262658
rect 587230 262338 587262 262574
rect 587498 262338 587582 262574
rect 587818 262338 587850 262574
rect 587230 226894 587850 262338
rect 587230 226658 587262 226894
rect 587498 226658 587582 226894
rect 587818 226658 587850 226894
rect 587230 226574 587850 226658
rect 587230 226338 587262 226574
rect 587498 226338 587582 226574
rect 587818 226338 587850 226574
rect 587230 190894 587850 226338
rect 587230 190658 587262 190894
rect 587498 190658 587582 190894
rect 587818 190658 587850 190894
rect 587230 190574 587850 190658
rect 587230 190338 587262 190574
rect 587498 190338 587582 190574
rect 587818 190338 587850 190574
rect 587230 154894 587850 190338
rect 587230 154658 587262 154894
rect 587498 154658 587582 154894
rect 587818 154658 587850 154894
rect 587230 154574 587850 154658
rect 587230 154338 587262 154574
rect 587498 154338 587582 154574
rect 587818 154338 587850 154574
rect 587230 118894 587850 154338
rect 587230 118658 587262 118894
rect 587498 118658 587582 118894
rect 587818 118658 587850 118894
rect 587230 118574 587850 118658
rect 587230 118338 587262 118574
rect 587498 118338 587582 118574
rect 587818 118338 587850 118574
rect 587230 82894 587850 118338
rect 587230 82658 587262 82894
rect 587498 82658 587582 82894
rect 587818 82658 587850 82894
rect 587230 82574 587850 82658
rect 587230 82338 587262 82574
rect 587498 82338 587582 82574
rect 587818 82338 587850 82574
rect 587230 46894 587850 82338
rect 587230 46658 587262 46894
rect 587498 46658 587582 46894
rect 587818 46658 587850 46894
rect 587230 46574 587850 46658
rect 587230 46338 587262 46574
rect 587498 46338 587582 46574
rect 587818 46338 587850 46574
rect 587230 10894 587850 46338
rect 587230 10658 587262 10894
rect 587498 10658 587582 10894
rect 587818 10658 587850 10894
rect 587230 10574 587850 10658
rect 587230 10338 587262 10574
rect 587498 10338 587582 10574
rect 587818 10338 587850 10574
rect 587230 -2266 587850 10338
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 698614 588810 707162
rect 588190 698378 588222 698614
rect 588458 698378 588542 698614
rect 588778 698378 588810 698614
rect 588190 698294 588810 698378
rect 588190 698058 588222 698294
rect 588458 698058 588542 698294
rect 588778 698058 588810 698294
rect 588190 662614 588810 698058
rect 588190 662378 588222 662614
rect 588458 662378 588542 662614
rect 588778 662378 588810 662614
rect 588190 662294 588810 662378
rect 588190 662058 588222 662294
rect 588458 662058 588542 662294
rect 588778 662058 588810 662294
rect 588190 626614 588810 662058
rect 588190 626378 588222 626614
rect 588458 626378 588542 626614
rect 588778 626378 588810 626614
rect 588190 626294 588810 626378
rect 588190 626058 588222 626294
rect 588458 626058 588542 626294
rect 588778 626058 588810 626294
rect 588190 590614 588810 626058
rect 588190 590378 588222 590614
rect 588458 590378 588542 590614
rect 588778 590378 588810 590614
rect 588190 590294 588810 590378
rect 588190 590058 588222 590294
rect 588458 590058 588542 590294
rect 588778 590058 588810 590294
rect 588190 554614 588810 590058
rect 588190 554378 588222 554614
rect 588458 554378 588542 554614
rect 588778 554378 588810 554614
rect 588190 554294 588810 554378
rect 588190 554058 588222 554294
rect 588458 554058 588542 554294
rect 588778 554058 588810 554294
rect 588190 518614 588810 554058
rect 588190 518378 588222 518614
rect 588458 518378 588542 518614
rect 588778 518378 588810 518614
rect 588190 518294 588810 518378
rect 588190 518058 588222 518294
rect 588458 518058 588542 518294
rect 588778 518058 588810 518294
rect 588190 482614 588810 518058
rect 588190 482378 588222 482614
rect 588458 482378 588542 482614
rect 588778 482378 588810 482614
rect 588190 482294 588810 482378
rect 588190 482058 588222 482294
rect 588458 482058 588542 482294
rect 588778 482058 588810 482294
rect 588190 446614 588810 482058
rect 588190 446378 588222 446614
rect 588458 446378 588542 446614
rect 588778 446378 588810 446614
rect 588190 446294 588810 446378
rect 588190 446058 588222 446294
rect 588458 446058 588542 446294
rect 588778 446058 588810 446294
rect 588190 410614 588810 446058
rect 588190 410378 588222 410614
rect 588458 410378 588542 410614
rect 588778 410378 588810 410614
rect 588190 410294 588810 410378
rect 588190 410058 588222 410294
rect 588458 410058 588542 410294
rect 588778 410058 588810 410294
rect 588190 374614 588810 410058
rect 588190 374378 588222 374614
rect 588458 374378 588542 374614
rect 588778 374378 588810 374614
rect 588190 374294 588810 374378
rect 588190 374058 588222 374294
rect 588458 374058 588542 374294
rect 588778 374058 588810 374294
rect 588190 338614 588810 374058
rect 588190 338378 588222 338614
rect 588458 338378 588542 338614
rect 588778 338378 588810 338614
rect 588190 338294 588810 338378
rect 588190 338058 588222 338294
rect 588458 338058 588542 338294
rect 588778 338058 588810 338294
rect 588190 302614 588810 338058
rect 588190 302378 588222 302614
rect 588458 302378 588542 302614
rect 588778 302378 588810 302614
rect 588190 302294 588810 302378
rect 588190 302058 588222 302294
rect 588458 302058 588542 302294
rect 588778 302058 588810 302294
rect 588190 266614 588810 302058
rect 588190 266378 588222 266614
rect 588458 266378 588542 266614
rect 588778 266378 588810 266614
rect 588190 266294 588810 266378
rect 588190 266058 588222 266294
rect 588458 266058 588542 266294
rect 588778 266058 588810 266294
rect 588190 230614 588810 266058
rect 588190 230378 588222 230614
rect 588458 230378 588542 230614
rect 588778 230378 588810 230614
rect 588190 230294 588810 230378
rect 588190 230058 588222 230294
rect 588458 230058 588542 230294
rect 588778 230058 588810 230294
rect 588190 194614 588810 230058
rect 588190 194378 588222 194614
rect 588458 194378 588542 194614
rect 588778 194378 588810 194614
rect 588190 194294 588810 194378
rect 588190 194058 588222 194294
rect 588458 194058 588542 194294
rect 588778 194058 588810 194294
rect 588190 158614 588810 194058
rect 588190 158378 588222 158614
rect 588458 158378 588542 158614
rect 588778 158378 588810 158614
rect 588190 158294 588810 158378
rect 588190 158058 588222 158294
rect 588458 158058 588542 158294
rect 588778 158058 588810 158294
rect 588190 122614 588810 158058
rect 588190 122378 588222 122614
rect 588458 122378 588542 122614
rect 588778 122378 588810 122614
rect 588190 122294 588810 122378
rect 588190 122058 588222 122294
rect 588458 122058 588542 122294
rect 588778 122058 588810 122294
rect 588190 86614 588810 122058
rect 588190 86378 588222 86614
rect 588458 86378 588542 86614
rect 588778 86378 588810 86614
rect 588190 86294 588810 86378
rect 588190 86058 588222 86294
rect 588458 86058 588542 86294
rect 588778 86058 588810 86294
rect 588190 50614 588810 86058
rect 588190 50378 588222 50614
rect 588458 50378 588542 50614
rect 588778 50378 588810 50614
rect 588190 50294 588810 50378
rect 588190 50058 588222 50294
rect 588458 50058 588542 50294
rect 588778 50058 588810 50294
rect 588190 14614 588810 50058
rect 588190 14378 588222 14614
rect 588458 14378 588542 14614
rect 588778 14378 588810 14614
rect 588190 14294 588810 14378
rect 588190 14058 588222 14294
rect 588458 14058 588542 14294
rect 588778 14058 588810 14294
rect 588190 -3226 588810 14058
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 666334 589770 708122
rect 589150 666098 589182 666334
rect 589418 666098 589502 666334
rect 589738 666098 589770 666334
rect 589150 666014 589770 666098
rect 589150 665778 589182 666014
rect 589418 665778 589502 666014
rect 589738 665778 589770 666014
rect 589150 630334 589770 665778
rect 589150 630098 589182 630334
rect 589418 630098 589502 630334
rect 589738 630098 589770 630334
rect 589150 630014 589770 630098
rect 589150 629778 589182 630014
rect 589418 629778 589502 630014
rect 589738 629778 589770 630014
rect 589150 594334 589770 629778
rect 589150 594098 589182 594334
rect 589418 594098 589502 594334
rect 589738 594098 589770 594334
rect 589150 594014 589770 594098
rect 589150 593778 589182 594014
rect 589418 593778 589502 594014
rect 589738 593778 589770 594014
rect 589150 558334 589770 593778
rect 589150 558098 589182 558334
rect 589418 558098 589502 558334
rect 589738 558098 589770 558334
rect 589150 558014 589770 558098
rect 589150 557778 589182 558014
rect 589418 557778 589502 558014
rect 589738 557778 589770 558014
rect 589150 522334 589770 557778
rect 589150 522098 589182 522334
rect 589418 522098 589502 522334
rect 589738 522098 589770 522334
rect 589150 522014 589770 522098
rect 589150 521778 589182 522014
rect 589418 521778 589502 522014
rect 589738 521778 589770 522014
rect 589150 486334 589770 521778
rect 589150 486098 589182 486334
rect 589418 486098 589502 486334
rect 589738 486098 589770 486334
rect 589150 486014 589770 486098
rect 589150 485778 589182 486014
rect 589418 485778 589502 486014
rect 589738 485778 589770 486014
rect 589150 450334 589770 485778
rect 589150 450098 589182 450334
rect 589418 450098 589502 450334
rect 589738 450098 589770 450334
rect 589150 450014 589770 450098
rect 589150 449778 589182 450014
rect 589418 449778 589502 450014
rect 589738 449778 589770 450014
rect 589150 414334 589770 449778
rect 589150 414098 589182 414334
rect 589418 414098 589502 414334
rect 589738 414098 589770 414334
rect 589150 414014 589770 414098
rect 589150 413778 589182 414014
rect 589418 413778 589502 414014
rect 589738 413778 589770 414014
rect 589150 378334 589770 413778
rect 589150 378098 589182 378334
rect 589418 378098 589502 378334
rect 589738 378098 589770 378334
rect 589150 378014 589770 378098
rect 589150 377778 589182 378014
rect 589418 377778 589502 378014
rect 589738 377778 589770 378014
rect 589150 342334 589770 377778
rect 589150 342098 589182 342334
rect 589418 342098 589502 342334
rect 589738 342098 589770 342334
rect 589150 342014 589770 342098
rect 589150 341778 589182 342014
rect 589418 341778 589502 342014
rect 589738 341778 589770 342014
rect 589150 306334 589770 341778
rect 589150 306098 589182 306334
rect 589418 306098 589502 306334
rect 589738 306098 589770 306334
rect 589150 306014 589770 306098
rect 589150 305778 589182 306014
rect 589418 305778 589502 306014
rect 589738 305778 589770 306014
rect 589150 270334 589770 305778
rect 589150 270098 589182 270334
rect 589418 270098 589502 270334
rect 589738 270098 589770 270334
rect 589150 270014 589770 270098
rect 589150 269778 589182 270014
rect 589418 269778 589502 270014
rect 589738 269778 589770 270014
rect 589150 234334 589770 269778
rect 589150 234098 589182 234334
rect 589418 234098 589502 234334
rect 589738 234098 589770 234334
rect 589150 234014 589770 234098
rect 589150 233778 589182 234014
rect 589418 233778 589502 234014
rect 589738 233778 589770 234014
rect 589150 198334 589770 233778
rect 589150 198098 589182 198334
rect 589418 198098 589502 198334
rect 589738 198098 589770 198334
rect 589150 198014 589770 198098
rect 589150 197778 589182 198014
rect 589418 197778 589502 198014
rect 589738 197778 589770 198014
rect 589150 162334 589770 197778
rect 589150 162098 589182 162334
rect 589418 162098 589502 162334
rect 589738 162098 589770 162334
rect 589150 162014 589770 162098
rect 589150 161778 589182 162014
rect 589418 161778 589502 162014
rect 589738 161778 589770 162014
rect 589150 126334 589770 161778
rect 589150 126098 589182 126334
rect 589418 126098 589502 126334
rect 589738 126098 589770 126334
rect 589150 126014 589770 126098
rect 589150 125778 589182 126014
rect 589418 125778 589502 126014
rect 589738 125778 589770 126014
rect 589150 90334 589770 125778
rect 589150 90098 589182 90334
rect 589418 90098 589502 90334
rect 589738 90098 589770 90334
rect 589150 90014 589770 90098
rect 589150 89778 589182 90014
rect 589418 89778 589502 90014
rect 589738 89778 589770 90014
rect 589150 54334 589770 89778
rect 589150 54098 589182 54334
rect 589418 54098 589502 54334
rect 589738 54098 589770 54334
rect 589150 54014 589770 54098
rect 589150 53778 589182 54014
rect 589418 53778 589502 54014
rect 589738 53778 589770 54014
rect 589150 18334 589770 53778
rect 589150 18098 589182 18334
rect 589418 18098 589502 18334
rect 589738 18098 589770 18334
rect 589150 18014 589770 18098
rect 589150 17778 589182 18014
rect 589418 17778 589502 18014
rect 589738 17778 589770 18014
rect 589150 -4186 589770 17778
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 670054 590730 709082
rect 590110 669818 590142 670054
rect 590378 669818 590462 670054
rect 590698 669818 590730 670054
rect 590110 669734 590730 669818
rect 590110 669498 590142 669734
rect 590378 669498 590462 669734
rect 590698 669498 590730 669734
rect 590110 634054 590730 669498
rect 590110 633818 590142 634054
rect 590378 633818 590462 634054
rect 590698 633818 590730 634054
rect 590110 633734 590730 633818
rect 590110 633498 590142 633734
rect 590378 633498 590462 633734
rect 590698 633498 590730 633734
rect 590110 598054 590730 633498
rect 590110 597818 590142 598054
rect 590378 597818 590462 598054
rect 590698 597818 590730 598054
rect 590110 597734 590730 597818
rect 590110 597498 590142 597734
rect 590378 597498 590462 597734
rect 590698 597498 590730 597734
rect 590110 562054 590730 597498
rect 590110 561818 590142 562054
rect 590378 561818 590462 562054
rect 590698 561818 590730 562054
rect 590110 561734 590730 561818
rect 590110 561498 590142 561734
rect 590378 561498 590462 561734
rect 590698 561498 590730 561734
rect 590110 526054 590730 561498
rect 590110 525818 590142 526054
rect 590378 525818 590462 526054
rect 590698 525818 590730 526054
rect 590110 525734 590730 525818
rect 590110 525498 590142 525734
rect 590378 525498 590462 525734
rect 590698 525498 590730 525734
rect 590110 490054 590730 525498
rect 590110 489818 590142 490054
rect 590378 489818 590462 490054
rect 590698 489818 590730 490054
rect 590110 489734 590730 489818
rect 590110 489498 590142 489734
rect 590378 489498 590462 489734
rect 590698 489498 590730 489734
rect 590110 454054 590730 489498
rect 590110 453818 590142 454054
rect 590378 453818 590462 454054
rect 590698 453818 590730 454054
rect 590110 453734 590730 453818
rect 590110 453498 590142 453734
rect 590378 453498 590462 453734
rect 590698 453498 590730 453734
rect 590110 418054 590730 453498
rect 590110 417818 590142 418054
rect 590378 417818 590462 418054
rect 590698 417818 590730 418054
rect 590110 417734 590730 417818
rect 590110 417498 590142 417734
rect 590378 417498 590462 417734
rect 590698 417498 590730 417734
rect 590110 382054 590730 417498
rect 590110 381818 590142 382054
rect 590378 381818 590462 382054
rect 590698 381818 590730 382054
rect 590110 381734 590730 381818
rect 590110 381498 590142 381734
rect 590378 381498 590462 381734
rect 590698 381498 590730 381734
rect 590110 346054 590730 381498
rect 590110 345818 590142 346054
rect 590378 345818 590462 346054
rect 590698 345818 590730 346054
rect 590110 345734 590730 345818
rect 590110 345498 590142 345734
rect 590378 345498 590462 345734
rect 590698 345498 590730 345734
rect 590110 310054 590730 345498
rect 590110 309818 590142 310054
rect 590378 309818 590462 310054
rect 590698 309818 590730 310054
rect 590110 309734 590730 309818
rect 590110 309498 590142 309734
rect 590378 309498 590462 309734
rect 590698 309498 590730 309734
rect 590110 274054 590730 309498
rect 590110 273818 590142 274054
rect 590378 273818 590462 274054
rect 590698 273818 590730 274054
rect 590110 273734 590730 273818
rect 590110 273498 590142 273734
rect 590378 273498 590462 273734
rect 590698 273498 590730 273734
rect 590110 238054 590730 273498
rect 590110 237818 590142 238054
rect 590378 237818 590462 238054
rect 590698 237818 590730 238054
rect 590110 237734 590730 237818
rect 590110 237498 590142 237734
rect 590378 237498 590462 237734
rect 590698 237498 590730 237734
rect 590110 202054 590730 237498
rect 590110 201818 590142 202054
rect 590378 201818 590462 202054
rect 590698 201818 590730 202054
rect 590110 201734 590730 201818
rect 590110 201498 590142 201734
rect 590378 201498 590462 201734
rect 590698 201498 590730 201734
rect 590110 166054 590730 201498
rect 590110 165818 590142 166054
rect 590378 165818 590462 166054
rect 590698 165818 590730 166054
rect 590110 165734 590730 165818
rect 590110 165498 590142 165734
rect 590378 165498 590462 165734
rect 590698 165498 590730 165734
rect 590110 130054 590730 165498
rect 590110 129818 590142 130054
rect 590378 129818 590462 130054
rect 590698 129818 590730 130054
rect 590110 129734 590730 129818
rect 590110 129498 590142 129734
rect 590378 129498 590462 129734
rect 590698 129498 590730 129734
rect 590110 94054 590730 129498
rect 590110 93818 590142 94054
rect 590378 93818 590462 94054
rect 590698 93818 590730 94054
rect 590110 93734 590730 93818
rect 590110 93498 590142 93734
rect 590378 93498 590462 93734
rect 590698 93498 590730 93734
rect 590110 58054 590730 93498
rect 590110 57818 590142 58054
rect 590378 57818 590462 58054
rect 590698 57818 590730 58054
rect 590110 57734 590730 57818
rect 590110 57498 590142 57734
rect 590378 57498 590462 57734
rect 590698 57498 590730 57734
rect 590110 22054 590730 57498
rect 590110 21818 590142 22054
rect 590378 21818 590462 22054
rect 590698 21818 590730 22054
rect 590110 21734 590730 21818
rect 590110 21498 590142 21734
rect 590378 21498 590462 21734
rect 590698 21498 590730 21734
rect 590110 -5146 590730 21498
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 673774 591690 710042
rect 591070 673538 591102 673774
rect 591338 673538 591422 673774
rect 591658 673538 591690 673774
rect 591070 673454 591690 673538
rect 591070 673218 591102 673454
rect 591338 673218 591422 673454
rect 591658 673218 591690 673454
rect 591070 637774 591690 673218
rect 591070 637538 591102 637774
rect 591338 637538 591422 637774
rect 591658 637538 591690 637774
rect 591070 637454 591690 637538
rect 591070 637218 591102 637454
rect 591338 637218 591422 637454
rect 591658 637218 591690 637454
rect 591070 601774 591690 637218
rect 591070 601538 591102 601774
rect 591338 601538 591422 601774
rect 591658 601538 591690 601774
rect 591070 601454 591690 601538
rect 591070 601218 591102 601454
rect 591338 601218 591422 601454
rect 591658 601218 591690 601454
rect 591070 565774 591690 601218
rect 591070 565538 591102 565774
rect 591338 565538 591422 565774
rect 591658 565538 591690 565774
rect 591070 565454 591690 565538
rect 591070 565218 591102 565454
rect 591338 565218 591422 565454
rect 591658 565218 591690 565454
rect 591070 529774 591690 565218
rect 591070 529538 591102 529774
rect 591338 529538 591422 529774
rect 591658 529538 591690 529774
rect 591070 529454 591690 529538
rect 591070 529218 591102 529454
rect 591338 529218 591422 529454
rect 591658 529218 591690 529454
rect 591070 493774 591690 529218
rect 591070 493538 591102 493774
rect 591338 493538 591422 493774
rect 591658 493538 591690 493774
rect 591070 493454 591690 493538
rect 591070 493218 591102 493454
rect 591338 493218 591422 493454
rect 591658 493218 591690 493454
rect 591070 457774 591690 493218
rect 591070 457538 591102 457774
rect 591338 457538 591422 457774
rect 591658 457538 591690 457774
rect 591070 457454 591690 457538
rect 591070 457218 591102 457454
rect 591338 457218 591422 457454
rect 591658 457218 591690 457454
rect 591070 421774 591690 457218
rect 591070 421538 591102 421774
rect 591338 421538 591422 421774
rect 591658 421538 591690 421774
rect 591070 421454 591690 421538
rect 591070 421218 591102 421454
rect 591338 421218 591422 421454
rect 591658 421218 591690 421454
rect 591070 385774 591690 421218
rect 591070 385538 591102 385774
rect 591338 385538 591422 385774
rect 591658 385538 591690 385774
rect 591070 385454 591690 385538
rect 591070 385218 591102 385454
rect 591338 385218 591422 385454
rect 591658 385218 591690 385454
rect 591070 349774 591690 385218
rect 591070 349538 591102 349774
rect 591338 349538 591422 349774
rect 591658 349538 591690 349774
rect 591070 349454 591690 349538
rect 591070 349218 591102 349454
rect 591338 349218 591422 349454
rect 591658 349218 591690 349454
rect 591070 313774 591690 349218
rect 591070 313538 591102 313774
rect 591338 313538 591422 313774
rect 591658 313538 591690 313774
rect 591070 313454 591690 313538
rect 591070 313218 591102 313454
rect 591338 313218 591422 313454
rect 591658 313218 591690 313454
rect 591070 277774 591690 313218
rect 591070 277538 591102 277774
rect 591338 277538 591422 277774
rect 591658 277538 591690 277774
rect 591070 277454 591690 277538
rect 591070 277218 591102 277454
rect 591338 277218 591422 277454
rect 591658 277218 591690 277454
rect 591070 241774 591690 277218
rect 591070 241538 591102 241774
rect 591338 241538 591422 241774
rect 591658 241538 591690 241774
rect 591070 241454 591690 241538
rect 591070 241218 591102 241454
rect 591338 241218 591422 241454
rect 591658 241218 591690 241454
rect 591070 205774 591690 241218
rect 591070 205538 591102 205774
rect 591338 205538 591422 205774
rect 591658 205538 591690 205774
rect 591070 205454 591690 205538
rect 591070 205218 591102 205454
rect 591338 205218 591422 205454
rect 591658 205218 591690 205454
rect 591070 169774 591690 205218
rect 591070 169538 591102 169774
rect 591338 169538 591422 169774
rect 591658 169538 591690 169774
rect 591070 169454 591690 169538
rect 591070 169218 591102 169454
rect 591338 169218 591422 169454
rect 591658 169218 591690 169454
rect 591070 133774 591690 169218
rect 591070 133538 591102 133774
rect 591338 133538 591422 133774
rect 591658 133538 591690 133774
rect 591070 133454 591690 133538
rect 591070 133218 591102 133454
rect 591338 133218 591422 133454
rect 591658 133218 591690 133454
rect 591070 97774 591690 133218
rect 591070 97538 591102 97774
rect 591338 97538 591422 97774
rect 591658 97538 591690 97774
rect 591070 97454 591690 97538
rect 591070 97218 591102 97454
rect 591338 97218 591422 97454
rect 591658 97218 591690 97454
rect 591070 61774 591690 97218
rect 591070 61538 591102 61774
rect 591338 61538 591422 61774
rect 591658 61538 591690 61774
rect 591070 61454 591690 61538
rect 591070 61218 591102 61454
rect 591338 61218 591422 61454
rect 591658 61218 591690 61454
rect 591070 25774 591690 61218
rect 591070 25538 591102 25774
rect 591338 25538 591422 25774
rect 591658 25538 591690 25774
rect 591070 25454 591690 25538
rect 591070 25218 591102 25454
rect 591338 25218 591422 25454
rect 591658 25218 591690 25454
rect 591070 -6106 591690 25218
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 677494 592650 711002
rect 592030 677258 592062 677494
rect 592298 677258 592382 677494
rect 592618 677258 592650 677494
rect 592030 677174 592650 677258
rect 592030 676938 592062 677174
rect 592298 676938 592382 677174
rect 592618 676938 592650 677174
rect 592030 641494 592650 676938
rect 592030 641258 592062 641494
rect 592298 641258 592382 641494
rect 592618 641258 592650 641494
rect 592030 641174 592650 641258
rect 592030 640938 592062 641174
rect 592298 640938 592382 641174
rect 592618 640938 592650 641174
rect 592030 605494 592650 640938
rect 592030 605258 592062 605494
rect 592298 605258 592382 605494
rect 592618 605258 592650 605494
rect 592030 605174 592650 605258
rect 592030 604938 592062 605174
rect 592298 604938 592382 605174
rect 592618 604938 592650 605174
rect 592030 569494 592650 604938
rect 592030 569258 592062 569494
rect 592298 569258 592382 569494
rect 592618 569258 592650 569494
rect 592030 569174 592650 569258
rect 592030 568938 592062 569174
rect 592298 568938 592382 569174
rect 592618 568938 592650 569174
rect 592030 533494 592650 568938
rect 592030 533258 592062 533494
rect 592298 533258 592382 533494
rect 592618 533258 592650 533494
rect 592030 533174 592650 533258
rect 592030 532938 592062 533174
rect 592298 532938 592382 533174
rect 592618 532938 592650 533174
rect 592030 497494 592650 532938
rect 592030 497258 592062 497494
rect 592298 497258 592382 497494
rect 592618 497258 592650 497494
rect 592030 497174 592650 497258
rect 592030 496938 592062 497174
rect 592298 496938 592382 497174
rect 592618 496938 592650 497174
rect 592030 461494 592650 496938
rect 592030 461258 592062 461494
rect 592298 461258 592382 461494
rect 592618 461258 592650 461494
rect 592030 461174 592650 461258
rect 592030 460938 592062 461174
rect 592298 460938 592382 461174
rect 592618 460938 592650 461174
rect 592030 425494 592650 460938
rect 592030 425258 592062 425494
rect 592298 425258 592382 425494
rect 592618 425258 592650 425494
rect 592030 425174 592650 425258
rect 592030 424938 592062 425174
rect 592298 424938 592382 425174
rect 592618 424938 592650 425174
rect 592030 389494 592650 424938
rect 592030 389258 592062 389494
rect 592298 389258 592382 389494
rect 592618 389258 592650 389494
rect 592030 389174 592650 389258
rect 592030 388938 592062 389174
rect 592298 388938 592382 389174
rect 592618 388938 592650 389174
rect 592030 353494 592650 388938
rect 592030 353258 592062 353494
rect 592298 353258 592382 353494
rect 592618 353258 592650 353494
rect 592030 353174 592650 353258
rect 592030 352938 592062 353174
rect 592298 352938 592382 353174
rect 592618 352938 592650 353174
rect 592030 317494 592650 352938
rect 592030 317258 592062 317494
rect 592298 317258 592382 317494
rect 592618 317258 592650 317494
rect 592030 317174 592650 317258
rect 592030 316938 592062 317174
rect 592298 316938 592382 317174
rect 592618 316938 592650 317174
rect 592030 281494 592650 316938
rect 592030 281258 592062 281494
rect 592298 281258 592382 281494
rect 592618 281258 592650 281494
rect 592030 281174 592650 281258
rect 592030 280938 592062 281174
rect 592298 280938 592382 281174
rect 592618 280938 592650 281174
rect 592030 245494 592650 280938
rect 592030 245258 592062 245494
rect 592298 245258 592382 245494
rect 592618 245258 592650 245494
rect 592030 245174 592650 245258
rect 592030 244938 592062 245174
rect 592298 244938 592382 245174
rect 592618 244938 592650 245174
rect 592030 209494 592650 244938
rect 592030 209258 592062 209494
rect 592298 209258 592382 209494
rect 592618 209258 592650 209494
rect 592030 209174 592650 209258
rect 592030 208938 592062 209174
rect 592298 208938 592382 209174
rect 592618 208938 592650 209174
rect 592030 173494 592650 208938
rect 592030 173258 592062 173494
rect 592298 173258 592382 173494
rect 592618 173258 592650 173494
rect 592030 173174 592650 173258
rect 592030 172938 592062 173174
rect 592298 172938 592382 173174
rect 592618 172938 592650 173174
rect 592030 137494 592650 172938
rect 592030 137258 592062 137494
rect 592298 137258 592382 137494
rect 592618 137258 592650 137494
rect 592030 137174 592650 137258
rect 592030 136938 592062 137174
rect 592298 136938 592382 137174
rect 592618 136938 592650 137174
rect 592030 101494 592650 136938
rect 592030 101258 592062 101494
rect 592298 101258 592382 101494
rect 592618 101258 592650 101494
rect 592030 101174 592650 101258
rect 592030 100938 592062 101174
rect 592298 100938 592382 101174
rect 592618 100938 592650 101174
rect 592030 65494 592650 100938
rect 592030 65258 592062 65494
rect 592298 65258 592382 65494
rect 592618 65258 592650 65494
rect 592030 65174 592650 65258
rect 592030 64938 592062 65174
rect 592298 64938 592382 65174
rect 592618 64938 592650 65174
rect 592030 29494 592650 64938
rect 592030 29258 592062 29494
rect 592298 29258 592382 29494
rect 592618 29258 592650 29494
rect 592030 29174 592650 29258
rect 592030 28938 592062 29174
rect 592298 28938 592382 29174
rect 592618 28938 592650 29174
rect 592030 -7066 592650 28938
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -8694 677258 -8458 677494
rect -8374 677258 -8138 677494
rect -8694 676938 -8458 677174
rect -8374 676938 -8138 677174
rect -8694 641258 -8458 641494
rect -8374 641258 -8138 641494
rect -8694 640938 -8458 641174
rect -8374 640938 -8138 641174
rect -8694 605258 -8458 605494
rect -8374 605258 -8138 605494
rect -8694 604938 -8458 605174
rect -8374 604938 -8138 605174
rect -8694 569258 -8458 569494
rect -8374 569258 -8138 569494
rect -8694 568938 -8458 569174
rect -8374 568938 -8138 569174
rect -8694 533258 -8458 533494
rect -8374 533258 -8138 533494
rect -8694 532938 -8458 533174
rect -8374 532938 -8138 533174
rect -8694 497258 -8458 497494
rect -8374 497258 -8138 497494
rect -8694 496938 -8458 497174
rect -8374 496938 -8138 497174
rect -8694 461258 -8458 461494
rect -8374 461258 -8138 461494
rect -8694 460938 -8458 461174
rect -8374 460938 -8138 461174
rect -8694 425258 -8458 425494
rect -8374 425258 -8138 425494
rect -8694 424938 -8458 425174
rect -8374 424938 -8138 425174
rect -8694 389258 -8458 389494
rect -8374 389258 -8138 389494
rect -8694 388938 -8458 389174
rect -8374 388938 -8138 389174
rect -8694 353258 -8458 353494
rect -8374 353258 -8138 353494
rect -8694 352938 -8458 353174
rect -8374 352938 -8138 353174
rect -8694 317258 -8458 317494
rect -8374 317258 -8138 317494
rect -8694 316938 -8458 317174
rect -8374 316938 -8138 317174
rect -8694 281258 -8458 281494
rect -8374 281258 -8138 281494
rect -8694 280938 -8458 281174
rect -8374 280938 -8138 281174
rect -8694 245258 -8458 245494
rect -8374 245258 -8138 245494
rect -8694 244938 -8458 245174
rect -8374 244938 -8138 245174
rect -8694 209258 -8458 209494
rect -8374 209258 -8138 209494
rect -8694 208938 -8458 209174
rect -8374 208938 -8138 209174
rect -8694 173258 -8458 173494
rect -8374 173258 -8138 173494
rect -8694 172938 -8458 173174
rect -8374 172938 -8138 173174
rect -8694 137258 -8458 137494
rect -8374 137258 -8138 137494
rect -8694 136938 -8458 137174
rect -8374 136938 -8138 137174
rect -8694 101258 -8458 101494
rect -8374 101258 -8138 101494
rect -8694 100938 -8458 101174
rect -8374 100938 -8138 101174
rect -8694 65258 -8458 65494
rect -8374 65258 -8138 65494
rect -8694 64938 -8458 65174
rect -8374 64938 -8138 65174
rect -8694 29258 -8458 29494
rect -8374 29258 -8138 29494
rect -8694 28938 -8458 29174
rect -8374 28938 -8138 29174
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect -7734 673538 -7498 673774
rect -7414 673538 -7178 673774
rect -7734 673218 -7498 673454
rect -7414 673218 -7178 673454
rect -7734 637538 -7498 637774
rect -7414 637538 -7178 637774
rect -7734 637218 -7498 637454
rect -7414 637218 -7178 637454
rect -7734 601538 -7498 601774
rect -7414 601538 -7178 601774
rect -7734 601218 -7498 601454
rect -7414 601218 -7178 601454
rect -7734 565538 -7498 565774
rect -7414 565538 -7178 565774
rect -7734 565218 -7498 565454
rect -7414 565218 -7178 565454
rect -7734 529538 -7498 529774
rect -7414 529538 -7178 529774
rect -7734 529218 -7498 529454
rect -7414 529218 -7178 529454
rect -7734 493538 -7498 493774
rect -7414 493538 -7178 493774
rect -7734 493218 -7498 493454
rect -7414 493218 -7178 493454
rect -7734 457538 -7498 457774
rect -7414 457538 -7178 457774
rect -7734 457218 -7498 457454
rect -7414 457218 -7178 457454
rect -7734 421538 -7498 421774
rect -7414 421538 -7178 421774
rect -7734 421218 -7498 421454
rect -7414 421218 -7178 421454
rect -7734 385538 -7498 385774
rect -7414 385538 -7178 385774
rect -7734 385218 -7498 385454
rect -7414 385218 -7178 385454
rect -7734 349538 -7498 349774
rect -7414 349538 -7178 349774
rect -7734 349218 -7498 349454
rect -7414 349218 -7178 349454
rect -7734 313538 -7498 313774
rect -7414 313538 -7178 313774
rect -7734 313218 -7498 313454
rect -7414 313218 -7178 313454
rect -7734 277538 -7498 277774
rect -7414 277538 -7178 277774
rect -7734 277218 -7498 277454
rect -7414 277218 -7178 277454
rect -7734 241538 -7498 241774
rect -7414 241538 -7178 241774
rect -7734 241218 -7498 241454
rect -7414 241218 -7178 241454
rect -7734 205538 -7498 205774
rect -7414 205538 -7178 205774
rect -7734 205218 -7498 205454
rect -7414 205218 -7178 205454
rect -7734 169538 -7498 169774
rect -7414 169538 -7178 169774
rect -7734 169218 -7498 169454
rect -7414 169218 -7178 169454
rect -7734 133538 -7498 133774
rect -7414 133538 -7178 133774
rect -7734 133218 -7498 133454
rect -7414 133218 -7178 133454
rect -7734 97538 -7498 97774
rect -7414 97538 -7178 97774
rect -7734 97218 -7498 97454
rect -7414 97218 -7178 97454
rect -7734 61538 -7498 61774
rect -7414 61538 -7178 61774
rect -7734 61218 -7498 61454
rect -7414 61218 -7178 61454
rect -7734 25538 -7498 25774
rect -7414 25538 -7178 25774
rect -7734 25218 -7498 25454
rect -7414 25218 -7178 25454
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -6774 669818 -6538 670054
rect -6454 669818 -6218 670054
rect -6774 669498 -6538 669734
rect -6454 669498 -6218 669734
rect -6774 633818 -6538 634054
rect -6454 633818 -6218 634054
rect -6774 633498 -6538 633734
rect -6454 633498 -6218 633734
rect -6774 597818 -6538 598054
rect -6454 597818 -6218 598054
rect -6774 597498 -6538 597734
rect -6454 597498 -6218 597734
rect -6774 561818 -6538 562054
rect -6454 561818 -6218 562054
rect -6774 561498 -6538 561734
rect -6454 561498 -6218 561734
rect -6774 525818 -6538 526054
rect -6454 525818 -6218 526054
rect -6774 525498 -6538 525734
rect -6454 525498 -6218 525734
rect -6774 489818 -6538 490054
rect -6454 489818 -6218 490054
rect -6774 489498 -6538 489734
rect -6454 489498 -6218 489734
rect -6774 453818 -6538 454054
rect -6454 453818 -6218 454054
rect -6774 453498 -6538 453734
rect -6454 453498 -6218 453734
rect -6774 417818 -6538 418054
rect -6454 417818 -6218 418054
rect -6774 417498 -6538 417734
rect -6454 417498 -6218 417734
rect -6774 381818 -6538 382054
rect -6454 381818 -6218 382054
rect -6774 381498 -6538 381734
rect -6454 381498 -6218 381734
rect -6774 345818 -6538 346054
rect -6454 345818 -6218 346054
rect -6774 345498 -6538 345734
rect -6454 345498 -6218 345734
rect -6774 309818 -6538 310054
rect -6454 309818 -6218 310054
rect -6774 309498 -6538 309734
rect -6454 309498 -6218 309734
rect -6774 273818 -6538 274054
rect -6454 273818 -6218 274054
rect -6774 273498 -6538 273734
rect -6454 273498 -6218 273734
rect -6774 237818 -6538 238054
rect -6454 237818 -6218 238054
rect -6774 237498 -6538 237734
rect -6454 237498 -6218 237734
rect -6774 201818 -6538 202054
rect -6454 201818 -6218 202054
rect -6774 201498 -6538 201734
rect -6454 201498 -6218 201734
rect -6774 165818 -6538 166054
rect -6454 165818 -6218 166054
rect -6774 165498 -6538 165734
rect -6454 165498 -6218 165734
rect -6774 129818 -6538 130054
rect -6454 129818 -6218 130054
rect -6774 129498 -6538 129734
rect -6454 129498 -6218 129734
rect -6774 93818 -6538 94054
rect -6454 93818 -6218 94054
rect -6774 93498 -6538 93734
rect -6454 93498 -6218 93734
rect -6774 57818 -6538 58054
rect -6454 57818 -6218 58054
rect -6774 57498 -6538 57734
rect -6454 57498 -6218 57734
rect -6774 21818 -6538 22054
rect -6454 21818 -6218 22054
rect -6774 21498 -6538 21734
rect -6454 21498 -6218 21734
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect -5814 666098 -5578 666334
rect -5494 666098 -5258 666334
rect -5814 665778 -5578 666014
rect -5494 665778 -5258 666014
rect -5814 630098 -5578 630334
rect -5494 630098 -5258 630334
rect -5814 629778 -5578 630014
rect -5494 629778 -5258 630014
rect -5814 594098 -5578 594334
rect -5494 594098 -5258 594334
rect -5814 593778 -5578 594014
rect -5494 593778 -5258 594014
rect -5814 558098 -5578 558334
rect -5494 558098 -5258 558334
rect -5814 557778 -5578 558014
rect -5494 557778 -5258 558014
rect -5814 522098 -5578 522334
rect -5494 522098 -5258 522334
rect -5814 521778 -5578 522014
rect -5494 521778 -5258 522014
rect -5814 486098 -5578 486334
rect -5494 486098 -5258 486334
rect -5814 485778 -5578 486014
rect -5494 485778 -5258 486014
rect -5814 450098 -5578 450334
rect -5494 450098 -5258 450334
rect -5814 449778 -5578 450014
rect -5494 449778 -5258 450014
rect -5814 414098 -5578 414334
rect -5494 414098 -5258 414334
rect -5814 413778 -5578 414014
rect -5494 413778 -5258 414014
rect -5814 378098 -5578 378334
rect -5494 378098 -5258 378334
rect -5814 377778 -5578 378014
rect -5494 377778 -5258 378014
rect -5814 342098 -5578 342334
rect -5494 342098 -5258 342334
rect -5814 341778 -5578 342014
rect -5494 341778 -5258 342014
rect -5814 306098 -5578 306334
rect -5494 306098 -5258 306334
rect -5814 305778 -5578 306014
rect -5494 305778 -5258 306014
rect -5814 270098 -5578 270334
rect -5494 270098 -5258 270334
rect -5814 269778 -5578 270014
rect -5494 269778 -5258 270014
rect -5814 234098 -5578 234334
rect -5494 234098 -5258 234334
rect -5814 233778 -5578 234014
rect -5494 233778 -5258 234014
rect -5814 198098 -5578 198334
rect -5494 198098 -5258 198334
rect -5814 197778 -5578 198014
rect -5494 197778 -5258 198014
rect -5814 162098 -5578 162334
rect -5494 162098 -5258 162334
rect -5814 161778 -5578 162014
rect -5494 161778 -5258 162014
rect -5814 126098 -5578 126334
rect -5494 126098 -5258 126334
rect -5814 125778 -5578 126014
rect -5494 125778 -5258 126014
rect -5814 90098 -5578 90334
rect -5494 90098 -5258 90334
rect -5814 89778 -5578 90014
rect -5494 89778 -5258 90014
rect -5814 54098 -5578 54334
rect -5494 54098 -5258 54334
rect -5814 53778 -5578 54014
rect -5494 53778 -5258 54014
rect -5814 18098 -5578 18334
rect -5494 18098 -5258 18334
rect -5814 17778 -5578 18014
rect -5494 17778 -5258 18014
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -4854 698378 -4618 698614
rect -4534 698378 -4298 698614
rect -4854 698058 -4618 698294
rect -4534 698058 -4298 698294
rect -4854 662378 -4618 662614
rect -4534 662378 -4298 662614
rect -4854 662058 -4618 662294
rect -4534 662058 -4298 662294
rect -4854 626378 -4618 626614
rect -4534 626378 -4298 626614
rect -4854 626058 -4618 626294
rect -4534 626058 -4298 626294
rect -4854 590378 -4618 590614
rect -4534 590378 -4298 590614
rect -4854 590058 -4618 590294
rect -4534 590058 -4298 590294
rect -4854 554378 -4618 554614
rect -4534 554378 -4298 554614
rect -4854 554058 -4618 554294
rect -4534 554058 -4298 554294
rect -4854 518378 -4618 518614
rect -4534 518378 -4298 518614
rect -4854 518058 -4618 518294
rect -4534 518058 -4298 518294
rect -4854 482378 -4618 482614
rect -4534 482378 -4298 482614
rect -4854 482058 -4618 482294
rect -4534 482058 -4298 482294
rect -4854 446378 -4618 446614
rect -4534 446378 -4298 446614
rect -4854 446058 -4618 446294
rect -4534 446058 -4298 446294
rect -4854 410378 -4618 410614
rect -4534 410378 -4298 410614
rect -4854 410058 -4618 410294
rect -4534 410058 -4298 410294
rect -4854 374378 -4618 374614
rect -4534 374378 -4298 374614
rect -4854 374058 -4618 374294
rect -4534 374058 -4298 374294
rect -4854 338378 -4618 338614
rect -4534 338378 -4298 338614
rect -4854 338058 -4618 338294
rect -4534 338058 -4298 338294
rect -4854 302378 -4618 302614
rect -4534 302378 -4298 302614
rect -4854 302058 -4618 302294
rect -4534 302058 -4298 302294
rect -4854 266378 -4618 266614
rect -4534 266378 -4298 266614
rect -4854 266058 -4618 266294
rect -4534 266058 -4298 266294
rect -4854 230378 -4618 230614
rect -4534 230378 -4298 230614
rect -4854 230058 -4618 230294
rect -4534 230058 -4298 230294
rect -4854 194378 -4618 194614
rect -4534 194378 -4298 194614
rect -4854 194058 -4618 194294
rect -4534 194058 -4298 194294
rect -4854 158378 -4618 158614
rect -4534 158378 -4298 158614
rect -4854 158058 -4618 158294
rect -4534 158058 -4298 158294
rect -4854 122378 -4618 122614
rect -4534 122378 -4298 122614
rect -4854 122058 -4618 122294
rect -4534 122058 -4298 122294
rect -4854 86378 -4618 86614
rect -4534 86378 -4298 86614
rect -4854 86058 -4618 86294
rect -4534 86058 -4298 86294
rect -4854 50378 -4618 50614
rect -4534 50378 -4298 50614
rect -4854 50058 -4618 50294
rect -4534 50058 -4298 50294
rect -4854 14378 -4618 14614
rect -4534 14378 -4298 14614
rect -4854 14058 -4618 14294
rect -4534 14058 -4298 14294
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect -3894 694658 -3658 694894
rect -3574 694658 -3338 694894
rect -3894 694338 -3658 694574
rect -3574 694338 -3338 694574
rect -3894 658658 -3658 658894
rect -3574 658658 -3338 658894
rect -3894 658338 -3658 658574
rect -3574 658338 -3338 658574
rect -3894 622658 -3658 622894
rect -3574 622658 -3338 622894
rect -3894 622338 -3658 622574
rect -3574 622338 -3338 622574
rect -3894 586658 -3658 586894
rect -3574 586658 -3338 586894
rect -3894 586338 -3658 586574
rect -3574 586338 -3338 586574
rect -3894 550658 -3658 550894
rect -3574 550658 -3338 550894
rect -3894 550338 -3658 550574
rect -3574 550338 -3338 550574
rect -3894 514658 -3658 514894
rect -3574 514658 -3338 514894
rect -3894 514338 -3658 514574
rect -3574 514338 -3338 514574
rect -3894 478658 -3658 478894
rect -3574 478658 -3338 478894
rect -3894 478338 -3658 478574
rect -3574 478338 -3338 478574
rect -3894 442658 -3658 442894
rect -3574 442658 -3338 442894
rect -3894 442338 -3658 442574
rect -3574 442338 -3338 442574
rect -3894 406658 -3658 406894
rect -3574 406658 -3338 406894
rect -3894 406338 -3658 406574
rect -3574 406338 -3338 406574
rect -3894 370658 -3658 370894
rect -3574 370658 -3338 370894
rect -3894 370338 -3658 370574
rect -3574 370338 -3338 370574
rect -3894 334658 -3658 334894
rect -3574 334658 -3338 334894
rect -3894 334338 -3658 334574
rect -3574 334338 -3338 334574
rect -3894 298658 -3658 298894
rect -3574 298658 -3338 298894
rect -3894 298338 -3658 298574
rect -3574 298338 -3338 298574
rect -3894 262658 -3658 262894
rect -3574 262658 -3338 262894
rect -3894 262338 -3658 262574
rect -3574 262338 -3338 262574
rect -3894 226658 -3658 226894
rect -3574 226658 -3338 226894
rect -3894 226338 -3658 226574
rect -3574 226338 -3338 226574
rect -3894 190658 -3658 190894
rect -3574 190658 -3338 190894
rect -3894 190338 -3658 190574
rect -3574 190338 -3338 190574
rect -3894 154658 -3658 154894
rect -3574 154658 -3338 154894
rect -3894 154338 -3658 154574
rect -3574 154338 -3338 154574
rect -3894 118658 -3658 118894
rect -3574 118658 -3338 118894
rect -3894 118338 -3658 118574
rect -3574 118338 -3338 118574
rect -3894 82658 -3658 82894
rect -3574 82658 -3338 82894
rect -3894 82338 -3658 82574
rect -3574 82338 -3338 82574
rect -3894 46658 -3658 46894
rect -3574 46658 -3338 46894
rect -3894 46338 -3658 46574
rect -3574 46338 -3338 46574
rect -3894 10658 -3658 10894
rect -3574 10658 -3338 10894
rect -3894 10338 -3658 10574
rect -3574 10338 -3338 10574
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 690938 -2698 691174
rect -2614 690938 -2378 691174
rect -2934 690618 -2698 690854
rect -2614 690618 -2378 690854
rect -2934 654938 -2698 655174
rect -2614 654938 -2378 655174
rect -2934 654618 -2698 654854
rect -2614 654618 -2378 654854
rect -2934 618938 -2698 619174
rect -2614 618938 -2378 619174
rect -2934 618618 -2698 618854
rect -2614 618618 -2378 618854
rect -2934 582938 -2698 583174
rect -2614 582938 -2378 583174
rect -2934 582618 -2698 582854
rect -2614 582618 -2378 582854
rect -2934 546938 -2698 547174
rect -2614 546938 -2378 547174
rect -2934 546618 -2698 546854
rect -2614 546618 -2378 546854
rect -2934 510938 -2698 511174
rect -2614 510938 -2378 511174
rect -2934 510618 -2698 510854
rect -2614 510618 -2378 510854
rect -2934 474938 -2698 475174
rect -2614 474938 -2378 475174
rect -2934 474618 -2698 474854
rect -2614 474618 -2378 474854
rect -2934 438938 -2698 439174
rect -2614 438938 -2378 439174
rect -2934 438618 -2698 438854
rect -2614 438618 -2378 438854
rect -2934 402938 -2698 403174
rect -2614 402938 -2378 403174
rect -2934 402618 -2698 402854
rect -2614 402618 -2378 402854
rect -2934 366938 -2698 367174
rect -2614 366938 -2378 367174
rect -2934 366618 -2698 366854
rect -2614 366618 -2378 366854
rect -2934 330938 -2698 331174
rect -2614 330938 -2378 331174
rect -2934 330618 -2698 330854
rect -2614 330618 -2378 330854
rect -2934 294938 -2698 295174
rect -2614 294938 -2378 295174
rect -2934 294618 -2698 294854
rect -2614 294618 -2378 294854
rect -2934 258938 -2698 259174
rect -2614 258938 -2378 259174
rect -2934 258618 -2698 258854
rect -2614 258618 -2378 258854
rect -2934 222938 -2698 223174
rect -2614 222938 -2378 223174
rect -2934 222618 -2698 222854
rect -2614 222618 -2378 222854
rect -2934 186938 -2698 187174
rect -2614 186938 -2378 187174
rect -2934 186618 -2698 186854
rect -2614 186618 -2378 186854
rect -2934 150938 -2698 151174
rect -2614 150938 -2378 151174
rect -2934 150618 -2698 150854
rect -2614 150618 -2378 150854
rect -2934 114938 -2698 115174
rect -2614 114938 -2378 115174
rect -2934 114618 -2698 114854
rect -2614 114618 -2378 114854
rect -2934 78938 -2698 79174
rect -2614 78938 -2378 79174
rect -2934 78618 -2698 78854
rect -2614 78618 -2378 78854
rect -2934 42938 -2698 43174
rect -2614 42938 -2378 43174
rect -2934 42618 -2698 42854
rect -2614 42618 -2378 42854
rect -2934 6938 -2698 7174
rect -2614 6938 -2378 7174
rect -2934 6618 -2698 6854
rect -2614 6618 -2378 6854
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect -1974 687218 -1738 687454
rect -1654 687218 -1418 687454
rect -1974 686898 -1738 687134
rect -1654 686898 -1418 687134
rect -1974 651218 -1738 651454
rect -1654 651218 -1418 651454
rect -1974 650898 -1738 651134
rect -1654 650898 -1418 651134
rect -1974 615218 -1738 615454
rect -1654 615218 -1418 615454
rect -1974 614898 -1738 615134
rect -1654 614898 -1418 615134
rect -1974 579218 -1738 579454
rect -1654 579218 -1418 579454
rect -1974 578898 -1738 579134
rect -1654 578898 -1418 579134
rect -1974 543218 -1738 543454
rect -1654 543218 -1418 543454
rect -1974 542898 -1738 543134
rect -1654 542898 -1418 543134
rect -1974 507218 -1738 507454
rect -1654 507218 -1418 507454
rect -1974 506898 -1738 507134
rect -1654 506898 -1418 507134
rect -1974 471218 -1738 471454
rect -1654 471218 -1418 471454
rect -1974 470898 -1738 471134
rect -1654 470898 -1418 471134
rect -1974 435218 -1738 435454
rect -1654 435218 -1418 435454
rect -1974 434898 -1738 435134
rect -1654 434898 -1418 435134
rect -1974 399218 -1738 399454
rect -1654 399218 -1418 399454
rect -1974 398898 -1738 399134
rect -1654 398898 -1418 399134
rect -1974 363218 -1738 363454
rect -1654 363218 -1418 363454
rect -1974 362898 -1738 363134
rect -1654 362898 -1418 363134
rect -1974 327218 -1738 327454
rect -1654 327218 -1418 327454
rect -1974 326898 -1738 327134
rect -1654 326898 -1418 327134
rect -1974 291218 -1738 291454
rect -1654 291218 -1418 291454
rect -1974 290898 -1738 291134
rect -1654 290898 -1418 291134
rect -1974 255218 -1738 255454
rect -1654 255218 -1418 255454
rect -1974 254898 -1738 255134
rect -1654 254898 -1418 255134
rect -1974 219218 -1738 219454
rect -1654 219218 -1418 219454
rect -1974 218898 -1738 219134
rect -1654 218898 -1418 219134
rect -1974 183218 -1738 183454
rect -1654 183218 -1418 183454
rect -1974 182898 -1738 183134
rect -1654 182898 -1418 183134
rect -1974 147218 -1738 147454
rect -1654 147218 -1418 147454
rect -1974 146898 -1738 147134
rect -1654 146898 -1418 147134
rect -1974 111218 -1738 111454
rect -1654 111218 -1418 111454
rect -1974 110898 -1738 111134
rect -1654 110898 -1418 111134
rect -1974 75218 -1738 75454
rect -1654 75218 -1418 75454
rect -1974 74898 -1738 75134
rect -1654 74898 -1418 75134
rect -1974 39218 -1738 39454
rect -1654 39218 -1418 39454
rect -1974 38898 -1738 39134
rect -1654 38898 -1418 39134
rect -1974 3218 -1738 3454
rect -1654 3218 -1418 3454
rect -1974 2898 -1738 3134
rect -1654 2898 -1418 3134
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect 1826 704602 2062 704838
rect 2146 704602 2382 704838
rect 1826 704282 2062 704518
rect 2146 704282 2382 704518
rect 1826 687218 2062 687454
rect 2146 687218 2382 687454
rect 1826 686898 2062 687134
rect 2146 686898 2382 687134
rect 5546 705562 5782 705798
rect 5866 705562 6102 705798
rect 5546 705242 5782 705478
rect 5866 705242 6102 705478
rect 5546 690938 5782 691174
rect 5866 690938 6102 691174
rect 5546 690618 5782 690854
rect 5866 690618 6102 690854
rect 1826 651218 2062 651454
rect 2146 651218 2382 651454
rect 1826 650898 2062 651134
rect 2146 650898 2382 651134
rect 1826 615218 2062 615454
rect 2146 615218 2382 615454
rect 1826 614898 2062 615134
rect 2146 614898 2382 615134
rect 5546 654938 5782 655174
rect 5866 654938 6102 655174
rect 5546 654618 5782 654854
rect 5866 654618 6102 654854
rect 5546 618938 5782 619174
rect 5866 618938 6102 619174
rect 5546 618618 5782 618854
rect 5866 618618 6102 618854
rect 1826 579218 2062 579454
rect 2146 579218 2382 579454
rect 1826 578898 2062 579134
rect 2146 578898 2382 579134
rect 1826 543218 2062 543454
rect 2146 543218 2382 543454
rect 1826 542898 2062 543134
rect 2146 542898 2382 543134
rect 1826 507218 2062 507454
rect 2146 507218 2382 507454
rect 1826 506898 2062 507134
rect 2146 506898 2382 507134
rect 1826 471218 2062 471454
rect 2146 471218 2382 471454
rect 1826 470898 2062 471134
rect 2146 470898 2382 471134
rect 1826 435218 2062 435454
rect 2146 435218 2382 435454
rect 1826 434898 2062 435134
rect 2146 434898 2382 435134
rect 1826 399218 2062 399454
rect 2146 399218 2382 399454
rect 1826 398898 2062 399134
rect 2146 398898 2382 399134
rect 1826 363218 2062 363454
rect 2146 363218 2382 363454
rect 1826 362898 2062 363134
rect 2146 362898 2382 363134
rect 1826 327218 2062 327454
rect 2146 327218 2382 327454
rect 1826 326898 2062 327134
rect 2146 326898 2382 327134
rect 1826 291218 2062 291454
rect 2146 291218 2382 291454
rect 1826 290898 2062 291134
rect 2146 290898 2382 291134
rect 1826 255218 2062 255454
rect 2146 255218 2382 255454
rect 1826 254898 2062 255134
rect 2146 254898 2382 255134
rect 1826 219218 2062 219454
rect 2146 219218 2382 219454
rect 1826 218898 2062 219134
rect 2146 218898 2382 219134
rect 1826 183218 2062 183454
rect 2146 183218 2382 183454
rect 1826 182898 2062 183134
rect 2146 182898 2382 183134
rect 1826 147218 2062 147454
rect 2146 147218 2382 147454
rect 1826 146898 2062 147134
rect 2146 146898 2382 147134
rect 5546 582938 5782 583174
rect 5866 582938 6102 583174
rect 5546 582618 5782 582854
rect 5866 582618 6102 582854
rect 5546 546938 5782 547174
rect 5866 546938 6102 547174
rect 5546 546618 5782 546854
rect 5866 546618 6102 546854
rect 5546 510938 5782 511174
rect 5866 510938 6102 511174
rect 5546 510618 5782 510854
rect 5866 510618 6102 510854
rect 5546 474938 5782 475174
rect 5866 474938 6102 475174
rect 5546 474618 5782 474854
rect 5866 474618 6102 474854
rect 5546 438938 5782 439174
rect 5866 438938 6102 439174
rect 5546 438618 5782 438854
rect 5866 438618 6102 438854
rect 5546 402938 5782 403174
rect 5866 402938 6102 403174
rect 5546 402618 5782 402854
rect 5866 402618 6102 402854
rect 5546 366938 5782 367174
rect 5866 366938 6102 367174
rect 5546 366618 5782 366854
rect 5866 366618 6102 366854
rect 5546 330938 5782 331174
rect 5866 330938 6102 331174
rect 5546 330618 5782 330854
rect 5866 330618 6102 330854
rect 5546 294938 5782 295174
rect 5866 294938 6102 295174
rect 5546 294618 5782 294854
rect 5866 294618 6102 294854
rect 5546 258938 5782 259174
rect 5866 258938 6102 259174
rect 5546 258618 5782 258854
rect 5866 258618 6102 258854
rect 5546 222938 5782 223174
rect 5866 222938 6102 223174
rect 5546 222618 5782 222854
rect 5866 222618 6102 222854
rect 5546 186938 5782 187174
rect 5866 186938 6102 187174
rect 5546 186618 5782 186854
rect 5866 186618 6102 186854
rect 5546 150938 5782 151174
rect 5866 150938 6102 151174
rect 5546 150618 5782 150854
rect 5866 150618 6102 150854
rect 1826 111218 2062 111454
rect 2146 111218 2382 111454
rect 1826 110898 2062 111134
rect 2146 110898 2382 111134
rect 5546 114938 5782 115174
rect 5866 114938 6102 115174
rect 5546 114618 5782 114854
rect 5866 114618 6102 114854
rect 1826 75218 2062 75454
rect 2146 75218 2382 75454
rect 1826 74898 2062 75134
rect 2146 74898 2382 75134
rect 5546 78938 5782 79174
rect 5866 78938 6102 79174
rect 5546 78618 5782 78854
rect 5866 78618 6102 78854
rect 1826 39218 2062 39454
rect 2146 39218 2382 39454
rect 1826 38898 2062 39134
rect 2146 38898 2382 39134
rect 1826 3218 2062 3454
rect 2146 3218 2382 3454
rect 1826 2898 2062 3134
rect 2146 2898 2382 3134
rect 1826 -582 2062 -346
rect 2146 -582 2382 -346
rect 1826 -902 2062 -666
rect 2146 -902 2382 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 5546 42938 5782 43174
rect 5866 42938 6102 43174
rect 5546 42618 5782 42854
rect 5866 42618 6102 42854
rect 5546 6938 5782 7174
rect 5866 6938 6102 7174
rect 5546 6618 5782 6854
rect 5866 6618 6102 6854
rect 5546 -1542 5782 -1306
rect 5866 -1542 6102 -1306
rect 5546 -1862 5782 -1626
rect 5866 -1862 6102 -1626
rect 9266 706522 9502 706758
rect 9586 706522 9822 706758
rect 9266 706202 9502 706438
rect 9586 706202 9822 706438
rect 9266 694658 9502 694894
rect 9586 694658 9822 694894
rect 9266 694338 9502 694574
rect 9586 694338 9822 694574
rect 9266 658658 9502 658894
rect 9586 658658 9822 658894
rect 9266 658338 9502 658574
rect 9586 658338 9822 658574
rect 9266 622658 9502 622894
rect 9586 622658 9822 622894
rect 9266 622338 9502 622574
rect 9586 622338 9822 622574
rect 9266 586658 9502 586894
rect 9586 586658 9822 586894
rect 9266 586338 9502 586574
rect 9586 586338 9822 586574
rect 9266 550658 9502 550894
rect 9586 550658 9822 550894
rect 9266 550338 9502 550574
rect 9586 550338 9822 550574
rect 9266 514658 9502 514894
rect 9586 514658 9822 514894
rect 9266 514338 9502 514574
rect 9586 514338 9822 514574
rect 9266 478658 9502 478894
rect 9586 478658 9822 478894
rect 9266 478338 9502 478574
rect 9586 478338 9822 478574
rect 9266 442658 9502 442894
rect 9586 442658 9822 442894
rect 9266 442338 9502 442574
rect 9586 442338 9822 442574
rect 9266 406658 9502 406894
rect 9586 406658 9822 406894
rect 9266 406338 9502 406574
rect 9586 406338 9822 406574
rect 9266 370658 9502 370894
rect 9586 370658 9822 370894
rect 9266 370338 9502 370574
rect 9586 370338 9822 370574
rect 9266 334658 9502 334894
rect 9586 334658 9822 334894
rect 9266 334338 9502 334574
rect 9586 334338 9822 334574
rect 9266 298658 9502 298894
rect 9586 298658 9822 298894
rect 9266 298338 9502 298574
rect 9586 298338 9822 298574
rect 9266 262658 9502 262894
rect 9586 262658 9822 262894
rect 9266 262338 9502 262574
rect 9586 262338 9822 262574
rect 9266 226658 9502 226894
rect 9586 226658 9822 226894
rect 9266 226338 9502 226574
rect 9586 226338 9822 226574
rect 9266 190658 9502 190894
rect 9586 190658 9822 190894
rect 9266 190338 9502 190574
rect 9586 190338 9822 190574
rect 9266 154658 9502 154894
rect 9586 154658 9822 154894
rect 9266 154338 9502 154574
rect 9586 154338 9822 154574
rect 9266 118658 9502 118894
rect 9586 118658 9822 118894
rect 9266 118338 9502 118574
rect 9586 118338 9822 118574
rect 9266 82658 9502 82894
rect 9586 82658 9822 82894
rect 9266 82338 9502 82574
rect 9586 82338 9822 82574
rect 9266 46658 9502 46894
rect 9586 46658 9822 46894
rect 9266 46338 9502 46574
rect 9586 46338 9822 46574
rect 9266 10658 9502 10894
rect 9586 10658 9822 10894
rect 9266 10338 9502 10574
rect 9586 10338 9822 10574
rect 9266 -2502 9502 -2266
rect 9586 -2502 9822 -2266
rect 9266 -2822 9502 -2586
rect 9586 -2822 9822 -2586
rect 12986 707482 13222 707718
rect 13306 707482 13542 707718
rect 12986 707162 13222 707398
rect 13306 707162 13542 707398
rect 12986 698378 13222 698614
rect 13306 698378 13542 698614
rect 12986 698058 13222 698294
rect 13306 698058 13542 698294
rect 12986 662378 13222 662614
rect 13306 662378 13542 662614
rect 12986 662058 13222 662294
rect 13306 662058 13542 662294
rect 12986 626378 13222 626614
rect 13306 626378 13542 626614
rect 12986 626058 13222 626294
rect 13306 626058 13542 626294
rect 12986 590378 13222 590614
rect 13306 590378 13542 590614
rect 12986 590058 13222 590294
rect 13306 590058 13542 590294
rect 12986 554378 13222 554614
rect 13306 554378 13542 554614
rect 12986 554058 13222 554294
rect 13306 554058 13542 554294
rect 12986 518378 13222 518614
rect 13306 518378 13542 518614
rect 12986 518058 13222 518294
rect 13306 518058 13542 518294
rect 12986 482378 13222 482614
rect 13306 482378 13542 482614
rect 12986 482058 13222 482294
rect 13306 482058 13542 482294
rect 12986 446378 13222 446614
rect 13306 446378 13542 446614
rect 12986 446058 13222 446294
rect 13306 446058 13542 446294
rect 12986 410378 13222 410614
rect 13306 410378 13542 410614
rect 12986 410058 13222 410294
rect 13306 410058 13542 410294
rect 12986 374378 13222 374614
rect 13306 374378 13542 374614
rect 12986 374058 13222 374294
rect 13306 374058 13542 374294
rect 12986 338378 13222 338614
rect 13306 338378 13542 338614
rect 12986 338058 13222 338294
rect 13306 338058 13542 338294
rect 12986 302378 13222 302614
rect 13306 302378 13542 302614
rect 12986 302058 13222 302294
rect 13306 302058 13542 302294
rect 12986 266378 13222 266614
rect 13306 266378 13542 266614
rect 12986 266058 13222 266294
rect 13306 266058 13542 266294
rect 12986 230378 13222 230614
rect 13306 230378 13542 230614
rect 12986 230058 13222 230294
rect 13306 230058 13542 230294
rect 12986 194378 13222 194614
rect 13306 194378 13542 194614
rect 12986 194058 13222 194294
rect 13306 194058 13542 194294
rect 12986 158378 13222 158614
rect 13306 158378 13542 158614
rect 12986 158058 13222 158294
rect 13306 158058 13542 158294
rect 12986 122378 13222 122614
rect 13306 122378 13542 122614
rect 12986 122058 13222 122294
rect 13306 122058 13542 122294
rect 12986 86378 13222 86614
rect 13306 86378 13542 86614
rect 12986 86058 13222 86294
rect 13306 86058 13542 86294
rect 12986 50378 13222 50614
rect 13306 50378 13542 50614
rect 12986 50058 13222 50294
rect 13306 50058 13542 50294
rect 12986 14378 13222 14614
rect 13306 14378 13542 14614
rect 12986 14058 13222 14294
rect 13306 14058 13542 14294
rect 12986 -3462 13222 -3226
rect 13306 -3462 13542 -3226
rect 12986 -3782 13222 -3546
rect 13306 -3782 13542 -3546
rect 16706 708442 16942 708678
rect 17026 708442 17262 708678
rect 16706 708122 16942 708358
rect 17026 708122 17262 708358
rect 16706 666098 16942 666334
rect 17026 666098 17262 666334
rect 16706 665778 16942 666014
rect 17026 665778 17262 666014
rect 16706 630098 16942 630334
rect 17026 630098 17262 630334
rect 16706 629778 16942 630014
rect 17026 629778 17262 630014
rect 16706 594098 16942 594334
rect 17026 594098 17262 594334
rect 16706 593778 16942 594014
rect 17026 593778 17262 594014
rect 16706 558098 16942 558334
rect 17026 558098 17262 558334
rect 16706 557778 16942 558014
rect 17026 557778 17262 558014
rect 16706 522098 16942 522334
rect 17026 522098 17262 522334
rect 16706 521778 16942 522014
rect 17026 521778 17262 522014
rect 16706 486098 16942 486334
rect 17026 486098 17262 486334
rect 16706 485778 16942 486014
rect 17026 485778 17262 486014
rect 16706 450098 16942 450334
rect 17026 450098 17262 450334
rect 16706 449778 16942 450014
rect 17026 449778 17262 450014
rect 16706 414098 16942 414334
rect 17026 414098 17262 414334
rect 16706 413778 16942 414014
rect 17026 413778 17262 414014
rect 16706 378098 16942 378334
rect 17026 378098 17262 378334
rect 16706 377778 16942 378014
rect 17026 377778 17262 378014
rect 16706 342098 16942 342334
rect 17026 342098 17262 342334
rect 16706 341778 16942 342014
rect 17026 341778 17262 342014
rect 16706 306098 16942 306334
rect 17026 306098 17262 306334
rect 16706 305778 16942 306014
rect 17026 305778 17262 306014
rect 16706 270098 16942 270334
rect 17026 270098 17262 270334
rect 16706 269778 16942 270014
rect 17026 269778 17262 270014
rect 16706 234098 16942 234334
rect 17026 234098 17262 234334
rect 16706 233778 16942 234014
rect 17026 233778 17262 234014
rect 16706 198098 16942 198334
rect 17026 198098 17262 198334
rect 16706 197778 16942 198014
rect 17026 197778 17262 198014
rect 16706 162098 16942 162334
rect 17026 162098 17262 162334
rect 16706 161778 16942 162014
rect 17026 161778 17262 162014
rect 16706 126098 16942 126334
rect 17026 126098 17262 126334
rect 16706 125778 16942 126014
rect 17026 125778 17262 126014
rect 16706 90098 16942 90334
rect 17026 90098 17262 90334
rect 16706 89778 16942 90014
rect 17026 89778 17262 90014
rect 16706 54098 16942 54334
rect 17026 54098 17262 54334
rect 16706 53778 16942 54014
rect 17026 53778 17262 54014
rect 16706 18098 16942 18334
rect 17026 18098 17262 18334
rect 16706 17778 16942 18014
rect 17026 17778 17262 18014
rect 16706 -4422 16942 -4186
rect 17026 -4422 17262 -4186
rect 16706 -4742 16942 -4506
rect 17026 -4742 17262 -4506
rect 20426 709402 20662 709638
rect 20746 709402 20982 709638
rect 20426 709082 20662 709318
rect 20746 709082 20982 709318
rect 20426 669818 20662 670054
rect 20746 669818 20982 670054
rect 20426 669498 20662 669734
rect 20746 669498 20982 669734
rect 27866 711322 28102 711558
rect 28186 711322 28422 711558
rect 27866 711002 28102 711238
rect 28186 711002 28422 711238
rect 27866 677258 28102 677494
rect 28186 677258 28422 677494
rect 27866 676938 28102 677174
rect 28186 676938 28422 677174
rect 24250 651218 24486 651454
rect 24250 650898 24486 651134
rect 20426 633818 20662 634054
rect 20746 633818 20982 634054
rect 20426 633498 20662 633734
rect 20746 633498 20982 633734
rect 37826 704602 38062 704838
rect 38146 704602 38382 704838
rect 37826 704282 38062 704518
rect 38146 704282 38382 704518
rect 37826 687218 38062 687454
rect 38146 687218 38382 687454
rect 37826 686898 38062 687134
rect 38146 686898 38382 687134
rect 41546 705562 41782 705798
rect 41866 705562 42102 705798
rect 41546 705242 41782 705478
rect 41866 705242 42102 705478
rect 41546 690938 41782 691174
rect 41866 690938 42102 691174
rect 41546 690618 41782 690854
rect 41866 690618 42102 690854
rect 45266 706522 45502 706758
rect 45586 706522 45822 706758
rect 45266 706202 45502 706438
rect 45586 706202 45822 706438
rect 45266 694658 45502 694894
rect 45586 694658 45822 694894
rect 45266 694338 45502 694574
rect 45586 694338 45822 694574
rect 48986 707482 49222 707718
rect 49306 707482 49542 707718
rect 48986 707162 49222 707398
rect 49306 707162 49542 707398
rect 48986 698378 49222 698614
rect 49306 698378 49542 698614
rect 48986 698058 49222 698294
rect 49306 698058 49542 698294
rect 63866 711322 64102 711558
rect 64186 711322 64422 711558
rect 63866 711002 64102 711238
rect 64186 711002 64422 711238
rect 63866 677258 64102 677494
rect 64186 677258 64422 677494
rect 63866 676938 64102 677174
rect 64186 676938 64422 677174
rect 73826 704602 74062 704838
rect 74146 704602 74382 704838
rect 73826 704282 74062 704518
rect 74146 704282 74382 704518
rect 73826 687218 74062 687454
rect 74146 687218 74382 687454
rect 73826 686898 74062 687134
rect 74146 686898 74382 687134
rect 77546 705562 77782 705798
rect 77866 705562 78102 705798
rect 77546 705242 77782 705478
rect 77866 705242 78102 705478
rect 77546 690938 77782 691174
rect 77866 690938 78102 691174
rect 77546 690618 77782 690854
rect 77866 690618 78102 690854
rect 81266 706522 81502 706758
rect 81586 706522 81822 706758
rect 81266 706202 81502 706438
rect 81586 706202 81822 706438
rect 81266 694658 81502 694894
rect 81586 694658 81822 694894
rect 81266 694338 81502 694574
rect 81586 694338 81822 694574
rect 84986 707482 85222 707718
rect 85306 707482 85542 707718
rect 84986 707162 85222 707398
rect 85306 707162 85542 707398
rect 84986 698378 85222 698614
rect 85306 698378 85542 698614
rect 84986 698058 85222 698294
rect 85306 698058 85542 698294
rect 99866 711322 100102 711558
rect 100186 711322 100422 711558
rect 99866 711002 100102 711238
rect 100186 711002 100422 711238
rect 99866 677258 100102 677494
rect 100186 677258 100422 677494
rect 99866 676938 100102 677174
rect 100186 676938 100422 677174
rect 109826 704602 110062 704838
rect 110146 704602 110382 704838
rect 109826 704282 110062 704518
rect 110146 704282 110382 704518
rect 109826 687218 110062 687454
rect 110146 687218 110382 687454
rect 109826 686898 110062 687134
rect 110146 686898 110382 687134
rect 113546 705562 113782 705798
rect 113866 705562 114102 705798
rect 113546 705242 113782 705478
rect 113866 705242 114102 705478
rect 113546 690938 113782 691174
rect 113866 690938 114102 691174
rect 113546 690618 113782 690854
rect 113866 690618 114102 690854
rect 117266 706522 117502 706758
rect 117586 706522 117822 706758
rect 117266 706202 117502 706438
rect 117586 706202 117822 706438
rect 117266 694658 117502 694894
rect 117586 694658 117822 694894
rect 117266 694338 117502 694574
rect 117586 694338 117822 694574
rect 120986 707482 121222 707718
rect 121306 707482 121542 707718
rect 120986 707162 121222 707398
rect 121306 707162 121542 707398
rect 120986 698378 121222 698614
rect 121306 698378 121542 698614
rect 120986 698058 121222 698294
rect 121306 698058 121542 698294
rect 135866 711322 136102 711558
rect 136186 711322 136422 711558
rect 135866 711002 136102 711238
rect 136186 711002 136422 711238
rect 135866 677258 136102 677494
rect 136186 677258 136422 677494
rect 135866 676938 136102 677174
rect 136186 676938 136422 677174
rect 145826 704602 146062 704838
rect 146146 704602 146382 704838
rect 145826 704282 146062 704518
rect 146146 704282 146382 704518
rect 145826 687218 146062 687454
rect 146146 687218 146382 687454
rect 145826 686898 146062 687134
rect 146146 686898 146382 687134
rect 149546 705562 149782 705798
rect 149866 705562 150102 705798
rect 149546 705242 149782 705478
rect 149866 705242 150102 705478
rect 149546 690938 149782 691174
rect 149866 690938 150102 691174
rect 149546 690618 149782 690854
rect 149866 690618 150102 690854
rect 153266 706522 153502 706758
rect 153586 706522 153822 706758
rect 153266 706202 153502 706438
rect 153586 706202 153822 706438
rect 153266 694658 153502 694894
rect 153586 694658 153822 694894
rect 153266 694338 153502 694574
rect 153586 694338 153822 694574
rect 156986 707482 157222 707718
rect 157306 707482 157542 707718
rect 156986 707162 157222 707398
rect 157306 707162 157542 707398
rect 156986 698378 157222 698614
rect 157306 698378 157542 698614
rect 156986 698058 157222 698294
rect 157306 698058 157542 698294
rect 171866 711322 172102 711558
rect 172186 711322 172422 711558
rect 171866 711002 172102 711238
rect 172186 711002 172422 711238
rect 171866 677258 172102 677494
rect 172186 677258 172422 677494
rect 171866 676938 172102 677174
rect 172186 676938 172422 677174
rect 181826 704602 182062 704838
rect 182146 704602 182382 704838
rect 181826 704282 182062 704518
rect 182146 704282 182382 704518
rect 181826 687218 182062 687454
rect 182146 687218 182382 687454
rect 181826 686898 182062 687134
rect 182146 686898 182382 687134
rect 185546 705562 185782 705798
rect 185866 705562 186102 705798
rect 185546 705242 185782 705478
rect 185866 705242 186102 705478
rect 185546 690938 185782 691174
rect 185866 690938 186102 691174
rect 185546 690618 185782 690854
rect 185866 690618 186102 690854
rect 189266 706522 189502 706758
rect 189586 706522 189822 706758
rect 189266 706202 189502 706438
rect 189586 706202 189822 706438
rect 189266 694658 189502 694894
rect 189586 694658 189822 694894
rect 189266 694338 189502 694574
rect 189586 694338 189822 694574
rect 192986 707482 193222 707718
rect 193306 707482 193542 707718
rect 192986 707162 193222 707398
rect 193306 707162 193542 707398
rect 192986 698378 193222 698614
rect 193306 698378 193542 698614
rect 192986 698058 193222 698294
rect 193306 698058 193542 698294
rect 207866 711322 208102 711558
rect 208186 711322 208422 711558
rect 207866 711002 208102 711238
rect 208186 711002 208422 711238
rect 207866 677258 208102 677494
rect 208186 677258 208422 677494
rect 207866 676938 208102 677174
rect 208186 676938 208422 677174
rect 217826 704602 218062 704838
rect 218146 704602 218382 704838
rect 217826 704282 218062 704518
rect 218146 704282 218382 704518
rect 217826 687218 218062 687454
rect 218146 687218 218382 687454
rect 217826 686898 218062 687134
rect 218146 686898 218382 687134
rect 221546 705562 221782 705798
rect 221866 705562 222102 705798
rect 221546 705242 221782 705478
rect 221866 705242 222102 705478
rect 221546 690938 221782 691174
rect 221866 690938 222102 691174
rect 221546 690618 221782 690854
rect 221866 690618 222102 690854
rect 225266 706522 225502 706758
rect 225586 706522 225822 706758
rect 225266 706202 225502 706438
rect 225586 706202 225822 706438
rect 225266 694658 225502 694894
rect 225586 694658 225822 694894
rect 225266 694338 225502 694574
rect 225586 694338 225822 694574
rect 228986 707482 229222 707718
rect 229306 707482 229542 707718
rect 228986 707162 229222 707398
rect 229306 707162 229542 707398
rect 228986 698378 229222 698614
rect 229306 698378 229542 698614
rect 228986 698058 229222 698294
rect 229306 698058 229542 698294
rect 243866 711322 244102 711558
rect 244186 711322 244422 711558
rect 243866 711002 244102 711238
rect 244186 711002 244422 711238
rect 243866 677258 244102 677494
rect 244186 677258 244422 677494
rect 243866 676938 244102 677174
rect 244186 676938 244422 677174
rect 253826 704602 254062 704838
rect 254146 704602 254382 704838
rect 253826 704282 254062 704518
rect 254146 704282 254382 704518
rect 253826 687218 254062 687454
rect 254146 687218 254382 687454
rect 253826 686898 254062 687134
rect 254146 686898 254382 687134
rect 257546 705562 257782 705798
rect 257866 705562 258102 705798
rect 257546 705242 257782 705478
rect 257866 705242 258102 705478
rect 257546 690938 257782 691174
rect 257866 690938 258102 691174
rect 257546 690618 257782 690854
rect 257866 690618 258102 690854
rect 261266 706522 261502 706758
rect 261586 706522 261822 706758
rect 261266 706202 261502 706438
rect 261586 706202 261822 706438
rect 261266 694658 261502 694894
rect 261586 694658 261822 694894
rect 261266 694338 261502 694574
rect 261586 694338 261822 694574
rect 264986 707482 265222 707718
rect 265306 707482 265542 707718
rect 264986 707162 265222 707398
rect 265306 707162 265542 707398
rect 264986 698378 265222 698614
rect 265306 698378 265542 698614
rect 264986 698058 265222 698294
rect 265306 698058 265542 698294
rect 279866 711322 280102 711558
rect 280186 711322 280422 711558
rect 279866 711002 280102 711238
rect 280186 711002 280422 711238
rect 279866 677258 280102 677494
rect 280186 677258 280422 677494
rect 279866 676938 280102 677174
rect 280186 676938 280422 677174
rect 289826 704602 290062 704838
rect 290146 704602 290382 704838
rect 289826 704282 290062 704518
rect 290146 704282 290382 704518
rect 289826 687218 290062 687454
rect 290146 687218 290382 687454
rect 289826 686898 290062 687134
rect 290146 686898 290382 687134
rect 293546 705562 293782 705798
rect 293866 705562 294102 705798
rect 293546 705242 293782 705478
rect 293866 705242 294102 705478
rect 293546 690938 293782 691174
rect 293866 690938 294102 691174
rect 293546 690618 293782 690854
rect 293866 690618 294102 690854
rect 297266 706522 297502 706758
rect 297586 706522 297822 706758
rect 297266 706202 297502 706438
rect 297586 706202 297822 706438
rect 297266 694658 297502 694894
rect 297586 694658 297822 694894
rect 297266 694338 297502 694574
rect 297586 694338 297822 694574
rect 300986 707482 301222 707718
rect 301306 707482 301542 707718
rect 300986 707162 301222 707398
rect 301306 707162 301542 707398
rect 300986 698378 301222 698614
rect 301306 698378 301542 698614
rect 300986 698058 301222 698294
rect 301306 698058 301542 698294
rect 325826 704602 326062 704838
rect 326146 704602 326382 704838
rect 325826 704282 326062 704518
rect 326146 704282 326382 704518
rect 325826 687218 326062 687454
rect 326146 687218 326382 687454
rect 325826 686898 326062 687134
rect 326146 686898 326382 687134
rect 329546 705562 329782 705798
rect 329866 705562 330102 705798
rect 329546 705242 329782 705478
rect 329866 705242 330102 705478
rect 329546 690938 329782 691174
rect 329866 690938 330102 691174
rect 329546 690618 329782 690854
rect 329866 690618 330102 690854
rect 333266 706522 333502 706758
rect 333586 706522 333822 706758
rect 333266 706202 333502 706438
rect 333586 706202 333822 706438
rect 333266 694658 333502 694894
rect 333586 694658 333822 694894
rect 333266 694338 333502 694574
rect 333586 694338 333822 694574
rect 336986 707482 337222 707718
rect 337306 707482 337542 707718
rect 336986 707162 337222 707398
rect 337306 707162 337542 707398
rect 336986 698378 337222 698614
rect 337306 698378 337542 698614
rect 336986 698058 337222 698294
rect 337306 698058 337542 698294
rect 351866 711322 352102 711558
rect 352186 711322 352422 711558
rect 351866 711002 352102 711238
rect 352186 711002 352422 711238
rect 351866 677258 352102 677494
rect 352186 677258 352422 677494
rect 351866 676938 352102 677174
rect 352186 676938 352422 677174
rect 361826 704602 362062 704838
rect 362146 704602 362382 704838
rect 361826 704282 362062 704518
rect 362146 704282 362382 704518
rect 361826 687218 362062 687454
rect 362146 687218 362382 687454
rect 361826 686898 362062 687134
rect 362146 686898 362382 687134
rect 39610 654938 39846 655174
rect 39610 654618 39846 654854
rect 70330 654938 70566 655174
rect 70330 654618 70566 654854
rect 101050 654938 101286 655174
rect 101050 654618 101286 654854
rect 131770 654938 132006 655174
rect 131770 654618 132006 654854
rect 162490 654938 162726 655174
rect 162490 654618 162726 654854
rect 193210 654938 193446 655174
rect 193210 654618 193446 654854
rect 223930 654938 224166 655174
rect 223930 654618 224166 654854
rect 254650 654938 254886 655174
rect 254650 654618 254886 654854
rect 285370 654938 285606 655174
rect 285370 654618 285606 654854
rect 316090 654938 316326 655174
rect 316090 654618 316326 654854
rect 346810 654938 347046 655174
rect 346810 654618 347046 654854
rect 54970 651218 55206 651454
rect 54970 650898 55206 651134
rect 85690 651218 85926 651454
rect 85690 650898 85926 651134
rect 116410 651218 116646 651454
rect 116410 650898 116646 651134
rect 147130 651218 147366 651454
rect 147130 650898 147366 651134
rect 177850 651218 178086 651454
rect 177850 650898 178086 651134
rect 208570 651218 208806 651454
rect 208570 650898 208806 651134
rect 239290 651218 239526 651454
rect 239290 650898 239526 651134
rect 270010 651218 270246 651454
rect 270010 650898 270246 651134
rect 300730 651218 300966 651454
rect 300730 650898 300966 651134
rect 331450 651218 331686 651454
rect 331450 650898 331686 651134
rect 361826 651218 362062 651454
rect 362146 651218 362382 651454
rect 361826 650898 362062 651134
rect 362146 650898 362382 651134
rect 27866 641258 28102 641494
rect 28186 641258 28422 641494
rect 27866 640938 28102 641174
rect 28186 640938 28422 641174
rect 24250 615218 24486 615454
rect 24250 614898 24486 615134
rect 20426 597818 20662 598054
rect 20746 597818 20982 598054
rect 20426 597498 20662 597734
rect 20746 597498 20982 597734
rect 39610 618938 39846 619174
rect 39610 618618 39846 618854
rect 70330 618938 70566 619174
rect 70330 618618 70566 618854
rect 101050 618938 101286 619174
rect 101050 618618 101286 618854
rect 131770 618938 132006 619174
rect 131770 618618 132006 618854
rect 162490 618938 162726 619174
rect 162490 618618 162726 618854
rect 193210 618938 193446 619174
rect 193210 618618 193446 618854
rect 223930 618938 224166 619174
rect 223930 618618 224166 618854
rect 254650 618938 254886 619174
rect 254650 618618 254886 618854
rect 285370 618938 285606 619174
rect 285370 618618 285606 618854
rect 316090 618938 316326 619174
rect 316090 618618 316326 618854
rect 346810 618938 347046 619174
rect 346810 618618 347046 618854
rect 54970 615218 55206 615454
rect 54970 614898 55206 615134
rect 85690 615218 85926 615454
rect 85690 614898 85926 615134
rect 116410 615218 116646 615454
rect 116410 614898 116646 615134
rect 147130 615218 147366 615454
rect 147130 614898 147366 615134
rect 177850 615218 178086 615454
rect 177850 614898 178086 615134
rect 208570 615218 208806 615454
rect 208570 614898 208806 615134
rect 239290 615218 239526 615454
rect 239290 614898 239526 615134
rect 270010 615218 270246 615454
rect 270010 614898 270246 615134
rect 300730 615218 300966 615454
rect 300730 614898 300966 615134
rect 331450 615218 331686 615454
rect 331450 614898 331686 615134
rect 361826 615218 362062 615454
rect 362146 615218 362382 615454
rect 361826 614898 362062 615134
rect 362146 614898 362382 615134
rect 27866 605258 28102 605494
rect 28186 605258 28422 605494
rect 27866 604938 28102 605174
rect 28186 604938 28422 605174
rect 24250 579218 24486 579454
rect 24250 578898 24486 579134
rect 20426 561818 20662 562054
rect 20746 561818 20982 562054
rect 20426 561498 20662 561734
rect 20746 561498 20982 561734
rect 39610 582938 39846 583174
rect 39610 582618 39846 582854
rect 70330 582938 70566 583174
rect 70330 582618 70566 582854
rect 101050 582938 101286 583174
rect 101050 582618 101286 582854
rect 131770 582938 132006 583174
rect 131770 582618 132006 582854
rect 162490 582938 162726 583174
rect 162490 582618 162726 582854
rect 193210 582938 193446 583174
rect 193210 582618 193446 582854
rect 223930 582938 224166 583174
rect 223930 582618 224166 582854
rect 254650 582938 254886 583174
rect 254650 582618 254886 582854
rect 285370 582938 285606 583174
rect 285370 582618 285606 582854
rect 316090 582938 316326 583174
rect 316090 582618 316326 582854
rect 346810 582938 347046 583174
rect 346810 582618 347046 582854
rect 54970 579218 55206 579454
rect 54970 578898 55206 579134
rect 85690 579218 85926 579454
rect 85690 578898 85926 579134
rect 116410 579218 116646 579454
rect 116410 578898 116646 579134
rect 147130 579218 147366 579454
rect 147130 578898 147366 579134
rect 177850 579218 178086 579454
rect 177850 578898 178086 579134
rect 208570 579218 208806 579454
rect 208570 578898 208806 579134
rect 239290 579218 239526 579454
rect 239290 578898 239526 579134
rect 270010 579218 270246 579454
rect 270010 578898 270246 579134
rect 300730 579218 300966 579454
rect 300730 578898 300966 579134
rect 331450 579218 331686 579454
rect 331450 578898 331686 579134
rect 361826 579218 362062 579454
rect 362146 579218 362382 579454
rect 361826 578898 362062 579134
rect 362146 578898 362382 579134
rect 27866 569258 28102 569494
rect 28186 569258 28422 569494
rect 27866 568938 28102 569174
rect 28186 568938 28422 569174
rect 24250 543218 24486 543454
rect 24250 542898 24486 543134
rect 20426 525818 20662 526054
rect 20746 525818 20982 526054
rect 20426 525498 20662 525734
rect 20746 525498 20982 525734
rect 39610 546938 39846 547174
rect 39610 546618 39846 546854
rect 70330 546938 70566 547174
rect 70330 546618 70566 546854
rect 101050 546938 101286 547174
rect 101050 546618 101286 546854
rect 131770 546938 132006 547174
rect 131770 546618 132006 546854
rect 162490 546938 162726 547174
rect 162490 546618 162726 546854
rect 193210 546938 193446 547174
rect 193210 546618 193446 546854
rect 223930 546938 224166 547174
rect 223930 546618 224166 546854
rect 254650 546938 254886 547174
rect 254650 546618 254886 546854
rect 285370 546938 285606 547174
rect 285370 546618 285606 546854
rect 316090 546938 316326 547174
rect 316090 546618 316326 546854
rect 346810 546938 347046 547174
rect 346810 546618 347046 546854
rect 54970 543218 55206 543454
rect 54970 542898 55206 543134
rect 85690 543218 85926 543454
rect 85690 542898 85926 543134
rect 116410 543218 116646 543454
rect 116410 542898 116646 543134
rect 147130 543218 147366 543454
rect 147130 542898 147366 543134
rect 177850 543218 178086 543454
rect 177850 542898 178086 543134
rect 208570 543218 208806 543454
rect 208570 542898 208806 543134
rect 239290 543218 239526 543454
rect 239290 542898 239526 543134
rect 270010 543218 270246 543454
rect 270010 542898 270246 543134
rect 300730 543218 300966 543454
rect 300730 542898 300966 543134
rect 331450 543218 331686 543454
rect 331450 542898 331686 543134
rect 361826 543218 362062 543454
rect 362146 543218 362382 543454
rect 361826 542898 362062 543134
rect 362146 542898 362382 543134
rect 27866 533258 28102 533494
rect 28186 533258 28422 533494
rect 27866 532938 28102 533174
rect 28186 532938 28422 533174
rect 24250 507218 24486 507454
rect 24250 506898 24486 507134
rect 20426 489818 20662 490054
rect 20746 489818 20982 490054
rect 20426 489498 20662 489734
rect 20746 489498 20982 489734
rect 39610 510938 39846 511174
rect 39610 510618 39846 510854
rect 70330 510938 70566 511174
rect 70330 510618 70566 510854
rect 101050 510938 101286 511174
rect 101050 510618 101286 510854
rect 131770 510938 132006 511174
rect 131770 510618 132006 510854
rect 162490 510938 162726 511174
rect 162490 510618 162726 510854
rect 193210 510938 193446 511174
rect 193210 510618 193446 510854
rect 223930 510938 224166 511174
rect 223930 510618 224166 510854
rect 254650 510938 254886 511174
rect 254650 510618 254886 510854
rect 285370 510938 285606 511174
rect 285370 510618 285606 510854
rect 316090 510938 316326 511174
rect 316090 510618 316326 510854
rect 346810 510938 347046 511174
rect 346810 510618 347046 510854
rect 54970 507218 55206 507454
rect 54970 506898 55206 507134
rect 85690 507218 85926 507454
rect 85690 506898 85926 507134
rect 116410 507218 116646 507454
rect 116410 506898 116646 507134
rect 147130 507218 147366 507454
rect 147130 506898 147366 507134
rect 177850 507218 178086 507454
rect 177850 506898 178086 507134
rect 208570 507218 208806 507454
rect 208570 506898 208806 507134
rect 239290 507218 239526 507454
rect 239290 506898 239526 507134
rect 270010 507218 270246 507454
rect 270010 506898 270246 507134
rect 300730 507218 300966 507454
rect 300730 506898 300966 507134
rect 331450 507218 331686 507454
rect 331450 506898 331686 507134
rect 361826 507218 362062 507454
rect 362146 507218 362382 507454
rect 361826 506898 362062 507134
rect 362146 506898 362382 507134
rect 27866 497258 28102 497494
rect 28186 497258 28422 497494
rect 27866 496938 28102 497174
rect 28186 496938 28422 497174
rect 24250 471218 24486 471454
rect 24250 470898 24486 471134
rect 20426 453818 20662 454054
rect 20746 453818 20982 454054
rect 20426 453498 20662 453734
rect 20746 453498 20982 453734
rect 39610 474938 39846 475174
rect 39610 474618 39846 474854
rect 70330 474938 70566 475174
rect 70330 474618 70566 474854
rect 101050 474938 101286 475174
rect 101050 474618 101286 474854
rect 131770 474938 132006 475174
rect 131770 474618 132006 474854
rect 162490 474938 162726 475174
rect 162490 474618 162726 474854
rect 193210 474938 193446 475174
rect 193210 474618 193446 474854
rect 223930 474938 224166 475174
rect 223930 474618 224166 474854
rect 254650 474938 254886 475174
rect 254650 474618 254886 474854
rect 285370 474938 285606 475174
rect 285370 474618 285606 474854
rect 316090 474938 316326 475174
rect 316090 474618 316326 474854
rect 346810 474938 347046 475174
rect 346810 474618 347046 474854
rect 54970 471218 55206 471454
rect 54970 470898 55206 471134
rect 85690 471218 85926 471454
rect 85690 470898 85926 471134
rect 116410 471218 116646 471454
rect 116410 470898 116646 471134
rect 147130 471218 147366 471454
rect 147130 470898 147366 471134
rect 177850 471218 178086 471454
rect 177850 470898 178086 471134
rect 208570 471218 208806 471454
rect 208570 470898 208806 471134
rect 239290 471218 239526 471454
rect 239290 470898 239526 471134
rect 270010 471218 270246 471454
rect 270010 470898 270246 471134
rect 300730 471218 300966 471454
rect 300730 470898 300966 471134
rect 331450 471218 331686 471454
rect 331450 470898 331686 471134
rect 361826 471218 362062 471454
rect 362146 471218 362382 471454
rect 361826 470898 362062 471134
rect 362146 470898 362382 471134
rect 27866 461258 28102 461494
rect 28186 461258 28422 461494
rect 27866 460938 28102 461174
rect 28186 460938 28422 461174
rect 24250 435218 24486 435454
rect 24250 434898 24486 435134
rect 20426 417818 20662 418054
rect 20746 417818 20982 418054
rect 20426 417498 20662 417734
rect 20746 417498 20982 417734
rect 39610 438938 39846 439174
rect 39610 438618 39846 438854
rect 70330 438938 70566 439174
rect 70330 438618 70566 438854
rect 101050 438938 101286 439174
rect 101050 438618 101286 438854
rect 131770 438938 132006 439174
rect 131770 438618 132006 438854
rect 162490 438938 162726 439174
rect 162490 438618 162726 438854
rect 193210 438938 193446 439174
rect 193210 438618 193446 438854
rect 223930 438938 224166 439174
rect 223930 438618 224166 438854
rect 254650 438938 254886 439174
rect 254650 438618 254886 438854
rect 285370 438938 285606 439174
rect 285370 438618 285606 438854
rect 316090 438938 316326 439174
rect 316090 438618 316326 438854
rect 346810 438938 347046 439174
rect 346810 438618 347046 438854
rect 54970 435218 55206 435454
rect 54970 434898 55206 435134
rect 85690 435218 85926 435454
rect 85690 434898 85926 435134
rect 116410 435218 116646 435454
rect 116410 434898 116646 435134
rect 147130 435218 147366 435454
rect 147130 434898 147366 435134
rect 177850 435218 178086 435454
rect 177850 434898 178086 435134
rect 208570 435218 208806 435454
rect 208570 434898 208806 435134
rect 239290 435218 239526 435454
rect 239290 434898 239526 435134
rect 270010 435218 270246 435454
rect 270010 434898 270246 435134
rect 300730 435218 300966 435454
rect 300730 434898 300966 435134
rect 331450 435218 331686 435454
rect 331450 434898 331686 435134
rect 361826 435218 362062 435454
rect 362146 435218 362382 435454
rect 361826 434898 362062 435134
rect 362146 434898 362382 435134
rect 27866 425258 28102 425494
rect 28186 425258 28422 425494
rect 27866 424938 28102 425174
rect 28186 424938 28422 425174
rect 24250 399218 24486 399454
rect 24250 398898 24486 399134
rect 20426 381818 20662 382054
rect 20746 381818 20982 382054
rect 20426 381498 20662 381734
rect 20746 381498 20982 381734
rect 39610 402938 39846 403174
rect 39610 402618 39846 402854
rect 70330 402938 70566 403174
rect 70330 402618 70566 402854
rect 101050 402938 101286 403174
rect 101050 402618 101286 402854
rect 131770 402938 132006 403174
rect 131770 402618 132006 402854
rect 162490 402938 162726 403174
rect 162490 402618 162726 402854
rect 193210 402938 193446 403174
rect 193210 402618 193446 402854
rect 223930 402938 224166 403174
rect 223930 402618 224166 402854
rect 254650 402938 254886 403174
rect 254650 402618 254886 402854
rect 285370 402938 285606 403174
rect 285370 402618 285606 402854
rect 316090 402938 316326 403174
rect 316090 402618 316326 402854
rect 346810 402938 347046 403174
rect 346810 402618 347046 402854
rect 54970 399218 55206 399454
rect 54970 398898 55206 399134
rect 85690 399218 85926 399454
rect 85690 398898 85926 399134
rect 116410 399218 116646 399454
rect 116410 398898 116646 399134
rect 147130 399218 147366 399454
rect 147130 398898 147366 399134
rect 177850 399218 178086 399454
rect 177850 398898 178086 399134
rect 208570 399218 208806 399454
rect 208570 398898 208806 399134
rect 239290 399218 239526 399454
rect 239290 398898 239526 399134
rect 270010 399218 270246 399454
rect 270010 398898 270246 399134
rect 300730 399218 300966 399454
rect 300730 398898 300966 399134
rect 331450 399218 331686 399454
rect 331450 398898 331686 399134
rect 361826 399218 362062 399454
rect 362146 399218 362382 399454
rect 361826 398898 362062 399134
rect 362146 398898 362382 399134
rect 27866 389258 28102 389494
rect 28186 389258 28422 389494
rect 27866 388938 28102 389174
rect 28186 388938 28422 389174
rect 24250 363218 24486 363454
rect 24250 362898 24486 363134
rect 20426 345818 20662 346054
rect 20746 345818 20982 346054
rect 20426 345498 20662 345734
rect 20746 345498 20982 345734
rect 39610 366938 39846 367174
rect 39610 366618 39846 366854
rect 70330 366938 70566 367174
rect 70330 366618 70566 366854
rect 101050 366938 101286 367174
rect 101050 366618 101286 366854
rect 131770 366938 132006 367174
rect 131770 366618 132006 366854
rect 162490 366938 162726 367174
rect 162490 366618 162726 366854
rect 193210 366938 193446 367174
rect 193210 366618 193446 366854
rect 223930 366938 224166 367174
rect 223930 366618 224166 366854
rect 254650 366938 254886 367174
rect 254650 366618 254886 366854
rect 285370 366938 285606 367174
rect 285370 366618 285606 366854
rect 316090 366938 316326 367174
rect 316090 366618 316326 366854
rect 346810 366938 347046 367174
rect 346810 366618 347046 366854
rect 54970 363218 55206 363454
rect 54970 362898 55206 363134
rect 85690 363218 85926 363454
rect 85690 362898 85926 363134
rect 116410 363218 116646 363454
rect 116410 362898 116646 363134
rect 147130 363218 147366 363454
rect 147130 362898 147366 363134
rect 177850 363218 178086 363454
rect 177850 362898 178086 363134
rect 208570 363218 208806 363454
rect 208570 362898 208806 363134
rect 239290 363218 239526 363454
rect 239290 362898 239526 363134
rect 270010 363218 270246 363454
rect 270010 362898 270246 363134
rect 300730 363218 300966 363454
rect 300730 362898 300966 363134
rect 331450 363218 331686 363454
rect 331450 362898 331686 363134
rect 361826 363218 362062 363454
rect 362146 363218 362382 363454
rect 361826 362898 362062 363134
rect 362146 362898 362382 363134
rect 27866 353258 28102 353494
rect 28186 353258 28422 353494
rect 27866 352938 28102 353174
rect 28186 352938 28422 353174
rect 24250 327218 24486 327454
rect 24250 326898 24486 327134
rect 20426 309818 20662 310054
rect 20746 309818 20982 310054
rect 20426 309498 20662 309734
rect 20746 309498 20982 309734
rect 39610 330938 39846 331174
rect 39610 330618 39846 330854
rect 70330 330938 70566 331174
rect 70330 330618 70566 330854
rect 101050 330938 101286 331174
rect 101050 330618 101286 330854
rect 131770 330938 132006 331174
rect 131770 330618 132006 330854
rect 162490 330938 162726 331174
rect 162490 330618 162726 330854
rect 193210 330938 193446 331174
rect 193210 330618 193446 330854
rect 223930 330938 224166 331174
rect 223930 330618 224166 330854
rect 254650 330938 254886 331174
rect 254650 330618 254886 330854
rect 285370 330938 285606 331174
rect 285370 330618 285606 330854
rect 316090 330938 316326 331174
rect 316090 330618 316326 330854
rect 346810 330938 347046 331174
rect 346810 330618 347046 330854
rect 54970 327218 55206 327454
rect 54970 326898 55206 327134
rect 85690 327218 85926 327454
rect 85690 326898 85926 327134
rect 116410 327218 116646 327454
rect 116410 326898 116646 327134
rect 147130 327218 147366 327454
rect 147130 326898 147366 327134
rect 177850 327218 178086 327454
rect 177850 326898 178086 327134
rect 208570 327218 208806 327454
rect 208570 326898 208806 327134
rect 239290 327218 239526 327454
rect 239290 326898 239526 327134
rect 270010 327218 270246 327454
rect 270010 326898 270246 327134
rect 300730 327218 300966 327454
rect 300730 326898 300966 327134
rect 331450 327218 331686 327454
rect 331450 326898 331686 327134
rect 361826 327218 362062 327454
rect 362146 327218 362382 327454
rect 361826 326898 362062 327134
rect 362146 326898 362382 327134
rect 27866 317258 28102 317494
rect 28186 317258 28422 317494
rect 27866 316938 28102 317174
rect 28186 316938 28422 317174
rect 24250 291218 24486 291454
rect 24250 290898 24486 291134
rect 20426 273818 20662 274054
rect 20746 273818 20982 274054
rect 20426 273498 20662 273734
rect 20746 273498 20982 273734
rect 39610 294938 39846 295174
rect 39610 294618 39846 294854
rect 70330 294938 70566 295174
rect 70330 294618 70566 294854
rect 101050 294938 101286 295174
rect 101050 294618 101286 294854
rect 131770 294938 132006 295174
rect 131770 294618 132006 294854
rect 162490 294938 162726 295174
rect 162490 294618 162726 294854
rect 193210 294938 193446 295174
rect 193210 294618 193446 294854
rect 223930 294938 224166 295174
rect 223930 294618 224166 294854
rect 254650 294938 254886 295174
rect 254650 294618 254886 294854
rect 285370 294938 285606 295174
rect 285370 294618 285606 294854
rect 316090 294938 316326 295174
rect 316090 294618 316326 294854
rect 346810 294938 347046 295174
rect 346810 294618 347046 294854
rect 54970 291218 55206 291454
rect 54970 290898 55206 291134
rect 85690 291218 85926 291454
rect 85690 290898 85926 291134
rect 116410 291218 116646 291454
rect 116410 290898 116646 291134
rect 147130 291218 147366 291454
rect 147130 290898 147366 291134
rect 177850 291218 178086 291454
rect 177850 290898 178086 291134
rect 208570 291218 208806 291454
rect 208570 290898 208806 291134
rect 239290 291218 239526 291454
rect 239290 290898 239526 291134
rect 270010 291218 270246 291454
rect 270010 290898 270246 291134
rect 300730 291218 300966 291454
rect 300730 290898 300966 291134
rect 331450 291218 331686 291454
rect 331450 290898 331686 291134
rect 361826 291218 362062 291454
rect 362146 291218 362382 291454
rect 361826 290898 362062 291134
rect 362146 290898 362382 291134
rect 27866 281258 28102 281494
rect 28186 281258 28422 281494
rect 27866 280938 28102 281174
rect 28186 280938 28422 281174
rect 24250 255218 24486 255454
rect 24250 254898 24486 255134
rect 20426 237818 20662 238054
rect 20746 237818 20982 238054
rect 20426 237498 20662 237734
rect 20746 237498 20982 237734
rect 39610 258938 39846 259174
rect 39610 258618 39846 258854
rect 70330 258938 70566 259174
rect 70330 258618 70566 258854
rect 101050 258938 101286 259174
rect 101050 258618 101286 258854
rect 131770 258938 132006 259174
rect 131770 258618 132006 258854
rect 162490 258938 162726 259174
rect 162490 258618 162726 258854
rect 193210 258938 193446 259174
rect 193210 258618 193446 258854
rect 223930 258938 224166 259174
rect 223930 258618 224166 258854
rect 254650 258938 254886 259174
rect 254650 258618 254886 258854
rect 285370 258938 285606 259174
rect 285370 258618 285606 258854
rect 316090 258938 316326 259174
rect 316090 258618 316326 258854
rect 346810 258938 347046 259174
rect 346810 258618 347046 258854
rect 54970 255218 55206 255454
rect 54970 254898 55206 255134
rect 85690 255218 85926 255454
rect 85690 254898 85926 255134
rect 116410 255218 116646 255454
rect 116410 254898 116646 255134
rect 147130 255218 147366 255454
rect 147130 254898 147366 255134
rect 177850 255218 178086 255454
rect 177850 254898 178086 255134
rect 208570 255218 208806 255454
rect 208570 254898 208806 255134
rect 239290 255218 239526 255454
rect 239290 254898 239526 255134
rect 270010 255218 270246 255454
rect 270010 254898 270246 255134
rect 300730 255218 300966 255454
rect 300730 254898 300966 255134
rect 331450 255218 331686 255454
rect 331450 254898 331686 255134
rect 361826 255218 362062 255454
rect 362146 255218 362382 255454
rect 361826 254898 362062 255134
rect 362146 254898 362382 255134
rect 27866 245258 28102 245494
rect 28186 245258 28422 245494
rect 27866 244938 28102 245174
rect 28186 244938 28422 245174
rect 24250 219218 24486 219454
rect 24250 218898 24486 219134
rect 20426 201818 20662 202054
rect 20746 201818 20982 202054
rect 20426 201498 20662 201734
rect 20746 201498 20982 201734
rect 39610 222938 39846 223174
rect 39610 222618 39846 222854
rect 70330 222938 70566 223174
rect 70330 222618 70566 222854
rect 101050 222938 101286 223174
rect 101050 222618 101286 222854
rect 131770 222938 132006 223174
rect 131770 222618 132006 222854
rect 162490 222938 162726 223174
rect 162490 222618 162726 222854
rect 193210 222938 193446 223174
rect 193210 222618 193446 222854
rect 223930 222938 224166 223174
rect 223930 222618 224166 222854
rect 254650 222938 254886 223174
rect 254650 222618 254886 222854
rect 285370 222938 285606 223174
rect 285370 222618 285606 222854
rect 316090 222938 316326 223174
rect 316090 222618 316326 222854
rect 346810 222938 347046 223174
rect 346810 222618 347046 222854
rect 54970 219218 55206 219454
rect 54970 218898 55206 219134
rect 85690 219218 85926 219454
rect 85690 218898 85926 219134
rect 116410 219218 116646 219454
rect 116410 218898 116646 219134
rect 147130 219218 147366 219454
rect 147130 218898 147366 219134
rect 177850 219218 178086 219454
rect 177850 218898 178086 219134
rect 208570 219218 208806 219454
rect 208570 218898 208806 219134
rect 239290 219218 239526 219454
rect 239290 218898 239526 219134
rect 270010 219218 270246 219454
rect 270010 218898 270246 219134
rect 300730 219218 300966 219454
rect 300730 218898 300966 219134
rect 331450 219218 331686 219454
rect 331450 218898 331686 219134
rect 361826 219218 362062 219454
rect 362146 219218 362382 219454
rect 361826 218898 362062 219134
rect 362146 218898 362382 219134
rect 27866 209258 28102 209494
rect 28186 209258 28422 209494
rect 27866 208938 28102 209174
rect 28186 208938 28422 209174
rect 24250 183218 24486 183454
rect 24250 182898 24486 183134
rect 20426 165818 20662 166054
rect 20746 165818 20982 166054
rect 20426 165498 20662 165734
rect 20746 165498 20982 165734
rect 39610 186938 39846 187174
rect 39610 186618 39846 186854
rect 70330 186938 70566 187174
rect 70330 186618 70566 186854
rect 101050 186938 101286 187174
rect 101050 186618 101286 186854
rect 131770 186938 132006 187174
rect 131770 186618 132006 186854
rect 162490 186938 162726 187174
rect 162490 186618 162726 186854
rect 193210 186938 193446 187174
rect 193210 186618 193446 186854
rect 223930 186938 224166 187174
rect 223930 186618 224166 186854
rect 254650 186938 254886 187174
rect 254650 186618 254886 186854
rect 285370 186938 285606 187174
rect 285370 186618 285606 186854
rect 316090 186938 316326 187174
rect 316090 186618 316326 186854
rect 346810 186938 347046 187174
rect 346810 186618 347046 186854
rect 54970 183218 55206 183454
rect 54970 182898 55206 183134
rect 85690 183218 85926 183454
rect 85690 182898 85926 183134
rect 116410 183218 116646 183454
rect 116410 182898 116646 183134
rect 147130 183218 147366 183454
rect 147130 182898 147366 183134
rect 177850 183218 178086 183454
rect 177850 182898 178086 183134
rect 208570 183218 208806 183454
rect 208570 182898 208806 183134
rect 239290 183218 239526 183454
rect 239290 182898 239526 183134
rect 270010 183218 270246 183454
rect 270010 182898 270246 183134
rect 300730 183218 300966 183454
rect 300730 182898 300966 183134
rect 331450 183218 331686 183454
rect 331450 182898 331686 183134
rect 361826 183218 362062 183454
rect 362146 183218 362382 183454
rect 361826 182898 362062 183134
rect 362146 182898 362382 183134
rect 27866 173258 28102 173494
rect 28186 173258 28422 173494
rect 27866 172938 28102 173174
rect 28186 172938 28422 173174
rect 24250 147218 24486 147454
rect 24250 146898 24486 147134
rect 20426 129818 20662 130054
rect 20746 129818 20982 130054
rect 20426 129498 20662 129734
rect 20746 129498 20982 129734
rect 39610 150938 39846 151174
rect 39610 150618 39846 150854
rect 70330 150938 70566 151174
rect 70330 150618 70566 150854
rect 101050 150938 101286 151174
rect 101050 150618 101286 150854
rect 131770 150938 132006 151174
rect 131770 150618 132006 150854
rect 162490 150938 162726 151174
rect 162490 150618 162726 150854
rect 193210 150938 193446 151174
rect 193210 150618 193446 150854
rect 223930 150938 224166 151174
rect 223930 150618 224166 150854
rect 254650 150938 254886 151174
rect 254650 150618 254886 150854
rect 285370 150938 285606 151174
rect 285370 150618 285606 150854
rect 316090 150938 316326 151174
rect 316090 150618 316326 150854
rect 346810 150938 347046 151174
rect 346810 150618 347046 150854
rect 54970 147218 55206 147454
rect 54970 146898 55206 147134
rect 85690 147218 85926 147454
rect 85690 146898 85926 147134
rect 116410 147218 116646 147454
rect 116410 146898 116646 147134
rect 147130 147218 147366 147454
rect 147130 146898 147366 147134
rect 177850 147218 178086 147454
rect 177850 146898 178086 147134
rect 208570 147218 208806 147454
rect 208570 146898 208806 147134
rect 239290 147218 239526 147454
rect 239290 146898 239526 147134
rect 270010 147218 270246 147454
rect 270010 146898 270246 147134
rect 300730 147218 300966 147454
rect 300730 146898 300966 147134
rect 331450 147218 331686 147454
rect 331450 146898 331686 147134
rect 361826 147218 362062 147454
rect 362146 147218 362382 147454
rect 361826 146898 362062 147134
rect 362146 146898 362382 147134
rect 27866 137258 28102 137494
rect 28186 137258 28422 137494
rect 27866 136938 28102 137174
rect 28186 136938 28422 137174
rect 24250 111218 24486 111454
rect 24250 110898 24486 111134
rect 20426 93818 20662 94054
rect 20746 93818 20982 94054
rect 20426 93498 20662 93734
rect 20746 93498 20982 93734
rect 39610 114938 39846 115174
rect 39610 114618 39846 114854
rect 70330 114938 70566 115174
rect 70330 114618 70566 114854
rect 101050 114938 101286 115174
rect 101050 114618 101286 114854
rect 131770 114938 132006 115174
rect 131770 114618 132006 114854
rect 162490 114938 162726 115174
rect 162490 114618 162726 114854
rect 193210 114938 193446 115174
rect 193210 114618 193446 114854
rect 223930 114938 224166 115174
rect 223930 114618 224166 114854
rect 254650 114938 254886 115174
rect 254650 114618 254886 114854
rect 285370 114938 285606 115174
rect 285370 114618 285606 114854
rect 316090 114938 316326 115174
rect 316090 114618 316326 114854
rect 346810 114938 347046 115174
rect 346810 114618 347046 114854
rect 54970 111218 55206 111454
rect 54970 110898 55206 111134
rect 85690 111218 85926 111454
rect 85690 110898 85926 111134
rect 116410 111218 116646 111454
rect 116410 110898 116646 111134
rect 147130 111218 147366 111454
rect 147130 110898 147366 111134
rect 177850 111218 178086 111454
rect 177850 110898 178086 111134
rect 208570 111218 208806 111454
rect 208570 110898 208806 111134
rect 239290 111218 239526 111454
rect 239290 110898 239526 111134
rect 270010 111218 270246 111454
rect 270010 110898 270246 111134
rect 300730 111218 300966 111454
rect 300730 110898 300966 111134
rect 331450 111218 331686 111454
rect 331450 110898 331686 111134
rect 361826 111218 362062 111454
rect 362146 111218 362382 111454
rect 361826 110898 362062 111134
rect 362146 110898 362382 111134
rect 27866 101258 28102 101494
rect 28186 101258 28422 101494
rect 27866 100938 28102 101174
rect 28186 100938 28422 101174
rect 24250 75218 24486 75454
rect 24250 74898 24486 75134
rect 20426 57818 20662 58054
rect 20746 57818 20982 58054
rect 20426 57498 20662 57734
rect 20746 57498 20982 57734
rect 39610 78938 39846 79174
rect 39610 78618 39846 78854
rect 70330 78938 70566 79174
rect 70330 78618 70566 78854
rect 101050 78938 101286 79174
rect 101050 78618 101286 78854
rect 131770 78938 132006 79174
rect 131770 78618 132006 78854
rect 162490 78938 162726 79174
rect 162490 78618 162726 78854
rect 193210 78938 193446 79174
rect 193210 78618 193446 78854
rect 223930 78938 224166 79174
rect 223930 78618 224166 78854
rect 254650 78938 254886 79174
rect 254650 78618 254886 78854
rect 285370 78938 285606 79174
rect 285370 78618 285606 78854
rect 316090 78938 316326 79174
rect 316090 78618 316326 78854
rect 346810 78938 347046 79174
rect 346810 78618 347046 78854
rect 54970 75218 55206 75454
rect 54970 74898 55206 75134
rect 85690 75218 85926 75454
rect 85690 74898 85926 75134
rect 116410 75218 116646 75454
rect 116410 74898 116646 75134
rect 147130 75218 147366 75454
rect 147130 74898 147366 75134
rect 177850 75218 178086 75454
rect 177850 74898 178086 75134
rect 208570 75218 208806 75454
rect 208570 74898 208806 75134
rect 239290 75218 239526 75454
rect 239290 74898 239526 75134
rect 270010 75218 270246 75454
rect 270010 74898 270246 75134
rect 300730 75218 300966 75454
rect 300730 74898 300966 75134
rect 331450 75218 331686 75454
rect 331450 74898 331686 75134
rect 361826 75218 362062 75454
rect 362146 75218 362382 75454
rect 361826 74898 362062 75134
rect 362146 74898 362382 75134
rect 27866 65258 28102 65494
rect 28186 65258 28422 65494
rect 27866 64938 28102 65174
rect 28186 64938 28422 65174
rect 20426 21818 20662 22054
rect 20746 21818 20982 22054
rect 20426 21498 20662 21734
rect 20746 21498 20982 21734
rect 20426 -5382 20662 -5146
rect 20746 -5382 20982 -5146
rect 20426 -5702 20662 -5466
rect 20746 -5702 20982 -5466
rect 24146 25538 24382 25774
rect 24466 25538 24702 25774
rect 24146 25218 24382 25454
rect 24466 25218 24702 25454
rect 24146 -6342 24382 -6106
rect 24466 -6342 24702 -6106
rect 24146 -6662 24382 -6426
rect 24466 -6662 24702 -6426
rect 27866 29258 28102 29494
rect 28186 29258 28422 29494
rect 27866 28938 28102 29174
rect 28186 28938 28422 29174
rect 27866 -7302 28102 -7066
rect 28186 -7302 28422 -7066
rect 27866 -7622 28102 -7386
rect 28186 -7622 28422 -7386
rect 37826 39218 38062 39454
rect 38146 39218 38382 39454
rect 37826 38898 38062 39134
rect 38146 38898 38382 39134
rect 37826 3218 38062 3454
rect 38146 3218 38382 3454
rect 37826 2898 38062 3134
rect 38146 2898 38382 3134
rect 37826 -582 38062 -346
rect 38146 -582 38382 -346
rect 37826 -902 38062 -666
rect 38146 -902 38382 -666
rect 41546 42938 41782 43174
rect 41866 42938 42102 43174
rect 41546 42618 41782 42854
rect 41866 42618 42102 42854
rect 41546 6938 41782 7174
rect 41866 6938 42102 7174
rect 41546 6618 41782 6854
rect 41866 6618 42102 6854
rect 41546 -1542 41782 -1306
rect 41866 -1542 42102 -1306
rect 41546 -1862 41782 -1626
rect 41866 -1862 42102 -1626
rect 45266 46658 45502 46894
rect 45586 46658 45822 46894
rect 45266 46338 45502 46574
rect 45586 46338 45822 46574
rect 45266 10658 45502 10894
rect 45586 10658 45822 10894
rect 45266 10338 45502 10574
rect 45586 10338 45822 10574
rect 45266 -2502 45502 -2266
rect 45586 -2502 45822 -2266
rect 45266 -2822 45502 -2586
rect 45586 -2822 45822 -2586
rect 48986 14378 49222 14614
rect 49306 14378 49542 14614
rect 48986 14058 49222 14294
rect 49306 14058 49542 14294
rect 48986 -3462 49222 -3226
rect 49306 -3462 49542 -3226
rect 48986 -3782 49222 -3546
rect 49306 -3782 49542 -3546
rect 52706 18098 52942 18334
rect 53026 18098 53262 18334
rect 52706 17778 52942 18014
rect 53026 17778 53262 18014
rect 52706 -4422 52942 -4186
rect 53026 -4422 53262 -4186
rect 52706 -4742 52942 -4506
rect 53026 -4742 53262 -4506
rect 56426 21818 56662 22054
rect 56746 21818 56982 22054
rect 56426 21498 56662 21734
rect 56746 21498 56982 21734
rect 56426 -5382 56662 -5146
rect 56746 -5382 56982 -5146
rect 56426 -5702 56662 -5466
rect 56746 -5702 56982 -5466
rect 60146 25538 60382 25774
rect 60466 25538 60702 25774
rect 60146 25218 60382 25454
rect 60466 25218 60702 25454
rect 60146 -6342 60382 -6106
rect 60466 -6342 60702 -6106
rect 60146 -6662 60382 -6426
rect 60466 -6662 60702 -6426
rect 63866 29258 64102 29494
rect 64186 29258 64422 29494
rect 63866 28938 64102 29174
rect 64186 28938 64422 29174
rect 63866 -7302 64102 -7066
rect 64186 -7302 64422 -7066
rect 63866 -7622 64102 -7386
rect 64186 -7622 64422 -7386
rect 73826 39218 74062 39454
rect 74146 39218 74382 39454
rect 73826 38898 74062 39134
rect 74146 38898 74382 39134
rect 73826 3218 74062 3454
rect 74146 3218 74382 3454
rect 73826 2898 74062 3134
rect 74146 2898 74382 3134
rect 73826 -582 74062 -346
rect 74146 -582 74382 -346
rect 73826 -902 74062 -666
rect 74146 -902 74382 -666
rect 77546 42938 77782 43174
rect 77866 42938 78102 43174
rect 77546 42618 77782 42854
rect 77866 42618 78102 42854
rect 77546 6938 77782 7174
rect 77866 6938 78102 7174
rect 77546 6618 77782 6854
rect 77866 6618 78102 6854
rect 77546 -1542 77782 -1306
rect 77866 -1542 78102 -1306
rect 77546 -1862 77782 -1626
rect 77866 -1862 78102 -1626
rect 81266 46658 81502 46894
rect 81586 46658 81822 46894
rect 81266 46338 81502 46574
rect 81586 46338 81822 46574
rect 81266 10658 81502 10894
rect 81586 10658 81822 10894
rect 81266 10338 81502 10574
rect 81586 10338 81822 10574
rect 81266 -2502 81502 -2266
rect 81586 -2502 81822 -2266
rect 81266 -2822 81502 -2586
rect 81586 -2822 81822 -2586
rect 84986 14378 85222 14614
rect 85306 14378 85542 14614
rect 84986 14058 85222 14294
rect 85306 14058 85542 14294
rect 84986 -3462 85222 -3226
rect 85306 -3462 85542 -3226
rect 84986 -3782 85222 -3546
rect 85306 -3782 85542 -3546
rect 88706 18098 88942 18334
rect 89026 18098 89262 18334
rect 88706 17778 88942 18014
rect 89026 17778 89262 18014
rect 88706 -4422 88942 -4186
rect 89026 -4422 89262 -4186
rect 88706 -4742 88942 -4506
rect 89026 -4742 89262 -4506
rect 92426 21818 92662 22054
rect 92746 21818 92982 22054
rect 92426 21498 92662 21734
rect 92746 21498 92982 21734
rect 92426 -5382 92662 -5146
rect 92746 -5382 92982 -5146
rect 92426 -5702 92662 -5466
rect 92746 -5702 92982 -5466
rect 96146 25538 96382 25774
rect 96466 25538 96702 25774
rect 96146 25218 96382 25454
rect 96466 25218 96702 25454
rect 96146 -6342 96382 -6106
rect 96466 -6342 96702 -6106
rect 96146 -6662 96382 -6426
rect 96466 -6662 96702 -6426
rect 99866 29258 100102 29494
rect 100186 29258 100422 29494
rect 99866 28938 100102 29174
rect 100186 28938 100422 29174
rect 99866 -7302 100102 -7066
rect 100186 -7302 100422 -7066
rect 99866 -7622 100102 -7386
rect 100186 -7622 100422 -7386
rect 109826 39218 110062 39454
rect 110146 39218 110382 39454
rect 109826 38898 110062 39134
rect 110146 38898 110382 39134
rect 109826 3218 110062 3454
rect 110146 3218 110382 3454
rect 109826 2898 110062 3134
rect 110146 2898 110382 3134
rect 109826 -582 110062 -346
rect 110146 -582 110382 -346
rect 109826 -902 110062 -666
rect 110146 -902 110382 -666
rect 113546 42938 113782 43174
rect 113866 42938 114102 43174
rect 113546 42618 113782 42854
rect 113866 42618 114102 42854
rect 113546 6938 113782 7174
rect 113866 6938 114102 7174
rect 113546 6618 113782 6854
rect 113866 6618 114102 6854
rect 113546 -1542 113782 -1306
rect 113866 -1542 114102 -1306
rect 113546 -1862 113782 -1626
rect 113866 -1862 114102 -1626
rect 117266 46658 117502 46894
rect 117586 46658 117822 46894
rect 117266 46338 117502 46574
rect 117586 46338 117822 46574
rect 117266 10658 117502 10894
rect 117586 10658 117822 10894
rect 117266 10338 117502 10574
rect 117586 10338 117822 10574
rect 117266 -2502 117502 -2266
rect 117586 -2502 117822 -2266
rect 117266 -2822 117502 -2586
rect 117586 -2822 117822 -2586
rect 120986 14378 121222 14614
rect 121306 14378 121542 14614
rect 120986 14058 121222 14294
rect 121306 14058 121542 14294
rect 120986 -3462 121222 -3226
rect 121306 -3462 121542 -3226
rect 120986 -3782 121222 -3546
rect 121306 -3782 121542 -3546
rect 124706 18098 124942 18334
rect 125026 18098 125262 18334
rect 124706 17778 124942 18014
rect 125026 17778 125262 18014
rect 124706 -4422 124942 -4186
rect 125026 -4422 125262 -4186
rect 124706 -4742 124942 -4506
rect 125026 -4742 125262 -4506
rect 128426 21818 128662 22054
rect 128746 21818 128982 22054
rect 128426 21498 128662 21734
rect 128746 21498 128982 21734
rect 128426 -5382 128662 -5146
rect 128746 -5382 128982 -5146
rect 128426 -5702 128662 -5466
rect 128746 -5702 128982 -5466
rect 132146 25538 132382 25774
rect 132466 25538 132702 25774
rect 132146 25218 132382 25454
rect 132466 25218 132702 25454
rect 132146 -6342 132382 -6106
rect 132466 -6342 132702 -6106
rect 132146 -6662 132382 -6426
rect 132466 -6662 132702 -6426
rect 135866 29258 136102 29494
rect 136186 29258 136422 29494
rect 135866 28938 136102 29174
rect 136186 28938 136422 29174
rect 135866 -7302 136102 -7066
rect 136186 -7302 136422 -7066
rect 135866 -7622 136102 -7386
rect 136186 -7622 136422 -7386
rect 145826 39218 146062 39454
rect 146146 39218 146382 39454
rect 145826 38898 146062 39134
rect 146146 38898 146382 39134
rect 145826 3218 146062 3454
rect 146146 3218 146382 3454
rect 145826 2898 146062 3134
rect 146146 2898 146382 3134
rect 145826 -582 146062 -346
rect 146146 -582 146382 -346
rect 145826 -902 146062 -666
rect 146146 -902 146382 -666
rect 149546 42938 149782 43174
rect 149866 42938 150102 43174
rect 149546 42618 149782 42854
rect 149866 42618 150102 42854
rect 149546 6938 149782 7174
rect 149866 6938 150102 7174
rect 149546 6618 149782 6854
rect 149866 6618 150102 6854
rect 149546 -1542 149782 -1306
rect 149866 -1542 150102 -1306
rect 149546 -1862 149782 -1626
rect 149866 -1862 150102 -1626
rect 153266 46658 153502 46894
rect 153586 46658 153822 46894
rect 153266 46338 153502 46574
rect 153586 46338 153822 46574
rect 153266 10658 153502 10894
rect 153586 10658 153822 10894
rect 153266 10338 153502 10574
rect 153586 10338 153822 10574
rect 153266 -2502 153502 -2266
rect 153586 -2502 153822 -2266
rect 153266 -2822 153502 -2586
rect 153586 -2822 153822 -2586
rect 156986 14378 157222 14614
rect 157306 14378 157542 14614
rect 156986 14058 157222 14294
rect 157306 14058 157542 14294
rect 156986 -3462 157222 -3226
rect 157306 -3462 157542 -3226
rect 156986 -3782 157222 -3546
rect 157306 -3782 157542 -3546
rect 160706 18098 160942 18334
rect 161026 18098 161262 18334
rect 160706 17778 160942 18014
rect 161026 17778 161262 18014
rect 160706 -4422 160942 -4186
rect 161026 -4422 161262 -4186
rect 160706 -4742 160942 -4506
rect 161026 -4742 161262 -4506
rect 164426 21818 164662 22054
rect 164746 21818 164982 22054
rect 164426 21498 164662 21734
rect 164746 21498 164982 21734
rect 164426 -5382 164662 -5146
rect 164746 -5382 164982 -5146
rect 164426 -5702 164662 -5466
rect 164746 -5702 164982 -5466
rect 168146 25538 168382 25774
rect 168466 25538 168702 25774
rect 168146 25218 168382 25454
rect 168466 25218 168702 25454
rect 168146 -6342 168382 -6106
rect 168466 -6342 168702 -6106
rect 168146 -6662 168382 -6426
rect 168466 -6662 168702 -6426
rect 171866 29258 172102 29494
rect 172186 29258 172422 29494
rect 171866 28938 172102 29174
rect 172186 28938 172422 29174
rect 171866 -7302 172102 -7066
rect 172186 -7302 172422 -7066
rect 171866 -7622 172102 -7386
rect 172186 -7622 172422 -7386
rect 181826 39218 182062 39454
rect 182146 39218 182382 39454
rect 181826 38898 182062 39134
rect 182146 38898 182382 39134
rect 181826 3218 182062 3454
rect 182146 3218 182382 3454
rect 181826 2898 182062 3134
rect 182146 2898 182382 3134
rect 181826 -582 182062 -346
rect 182146 -582 182382 -346
rect 181826 -902 182062 -666
rect 182146 -902 182382 -666
rect 185546 42938 185782 43174
rect 185866 42938 186102 43174
rect 185546 42618 185782 42854
rect 185866 42618 186102 42854
rect 185546 6938 185782 7174
rect 185866 6938 186102 7174
rect 185546 6618 185782 6854
rect 185866 6618 186102 6854
rect 185546 -1542 185782 -1306
rect 185866 -1542 186102 -1306
rect 185546 -1862 185782 -1626
rect 185866 -1862 186102 -1626
rect 189266 46658 189502 46894
rect 189586 46658 189822 46894
rect 189266 46338 189502 46574
rect 189586 46338 189822 46574
rect 189266 10658 189502 10894
rect 189586 10658 189822 10894
rect 189266 10338 189502 10574
rect 189586 10338 189822 10574
rect 189266 -2502 189502 -2266
rect 189586 -2502 189822 -2266
rect 189266 -2822 189502 -2586
rect 189586 -2822 189822 -2586
rect 192986 14378 193222 14614
rect 193306 14378 193542 14614
rect 192986 14058 193222 14294
rect 193306 14058 193542 14294
rect 192986 -3462 193222 -3226
rect 193306 -3462 193542 -3226
rect 192986 -3782 193222 -3546
rect 193306 -3782 193542 -3546
rect 196706 18098 196942 18334
rect 197026 18098 197262 18334
rect 196706 17778 196942 18014
rect 197026 17778 197262 18014
rect 196706 -4422 196942 -4186
rect 197026 -4422 197262 -4186
rect 196706 -4742 196942 -4506
rect 197026 -4742 197262 -4506
rect 200426 21818 200662 22054
rect 200746 21818 200982 22054
rect 200426 21498 200662 21734
rect 200746 21498 200982 21734
rect 200426 -5382 200662 -5146
rect 200746 -5382 200982 -5146
rect 200426 -5702 200662 -5466
rect 200746 -5702 200982 -5466
rect 204146 25538 204382 25774
rect 204466 25538 204702 25774
rect 204146 25218 204382 25454
rect 204466 25218 204702 25454
rect 204146 -6342 204382 -6106
rect 204466 -6342 204702 -6106
rect 204146 -6662 204382 -6426
rect 204466 -6662 204702 -6426
rect 207866 29258 208102 29494
rect 208186 29258 208422 29494
rect 207866 28938 208102 29174
rect 208186 28938 208422 29174
rect 207866 -7302 208102 -7066
rect 208186 -7302 208422 -7066
rect 207866 -7622 208102 -7386
rect 208186 -7622 208422 -7386
rect 217826 39218 218062 39454
rect 218146 39218 218382 39454
rect 217826 38898 218062 39134
rect 218146 38898 218382 39134
rect 217826 3218 218062 3454
rect 218146 3218 218382 3454
rect 217826 2898 218062 3134
rect 218146 2898 218382 3134
rect 217826 -582 218062 -346
rect 218146 -582 218382 -346
rect 217826 -902 218062 -666
rect 218146 -902 218382 -666
rect 221546 42938 221782 43174
rect 221866 42938 222102 43174
rect 221546 42618 221782 42854
rect 221866 42618 222102 42854
rect 221546 6938 221782 7174
rect 221866 6938 222102 7174
rect 221546 6618 221782 6854
rect 221866 6618 222102 6854
rect 221546 -1542 221782 -1306
rect 221866 -1542 222102 -1306
rect 221546 -1862 221782 -1626
rect 221866 -1862 222102 -1626
rect 225266 46658 225502 46894
rect 225586 46658 225822 46894
rect 225266 46338 225502 46574
rect 225586 46338 225822 46574
rect 225266 10658 225502 10894
rect 225586 10658 225822 10894
rect 225266 10338 225502 10574
rect 225586 10338 225822 10574
rect 225266 -2502 225502 -2266
rect 225586 -2502 225822 -2266
rect 225266 -2822 225502 -2586
rect 225586 -2822 225822 -2586
rect 228986 14378 229222 14614
rect 229306 14378 229542 14614
rect 228986 14058 229222 14294
rect 229306 14058 229542 14294
rect 228986 -3462 229222 -3226
rect 229306 -3462 229542 -3226
rect 228986 -3782 229222 -3546
rect 229306 -3782 229542 -3546
rect 232706 18098 232942 18334
rect 233026 18098 233262 18334
rect 232706 17778 232942 18014
rect 233026 17778 233262 18014
rect 232706 -4422 232942 -4186
rect 233026 -4422 233262 -4186
rect 232706 -4742 232942 -4506
rect 233026 -4742 233262 -4506
rect 236426 21818 236662 22054
rect 236746 21818 236982 22054
rect 236426 21498 236662 21734
rect 236746 21498 236982 21734
rect 236426 -5382 236662 -5146
rect 236746 -5382 236982 -5146
rect 236426 -5702 236662 -5466
rect 236746 -5702 236982 -5466
rect 240146 25538 240382 25774
rect 240466 25538 240702 25774
rect 240146 25218 240382 25454
rect 240466 25218 240702 25454
rect 240146 -6342 240382 -6106
rect 240466 -6342 240702 -6106
rect 240146 -6662 240382 -6426
rect 240466 -6662 240702 -6426
rect 243866 29258 244102 29494
rect 244186 29258 244422 29494
rect 243866 28938 244102 29174
rect 244186 28938 244422 29174
rect 243866 -7302 244102 -7066
rect 244186 -7302 244422 -7066
rect 243866 -7622 244102 -7386
rect 244186 -7622 244422 -7386
rect 253826 39218 254062 39454
rect 254146 39218 254382 39454
rect 253826 38898 254062 39134
rect 254146 38898 254382 39134
rect 253826 3218 254062 3454
rect 254146 3218 254382 3454
rect 253826 2898 254062 3134
rect 254146 2898 254382 3134
rect 253826 -582 254062 -346
rect 254146 -582 254382 -346
rect 253826 -902 254062 -666
rect 254146 -902 254382 -666
rect 257546 42938 257782 43174
rect 257866 42938 258102 43174
rect 257546 42618 257782 42854
rect 257866 42618 258102 42854
rect 257546 6938 257782 7174
rect 257866 6938 258102 7174
rect 257546 6618 257782 6854
rect 257866 6618 258102 6854
rect 257546 -1542 257782 -1306
rect 257866 -1542 258102 -1306
rect 257546 -1862 257782 -1626
rect 257866 -1862 258102 -1626
rect 261266 46658 261502 46894
rect 261586 46658 261822 46894
rect 261266 46338 261502 46574
rect 261586 46338 261822 46574
rect 261266 10658 261502 10894
rect 261586 10658 261822 10894
rect 261266 10338 261502 10574
rect 261586 10338 261822 10574
rect 261266 -2502 261502 -2266
rect 261586 -2502 261822 -2266
rect 261266 -2822 261502 -2586
rect 261586 -2822 261822 -2586
rect 264986 14378 265222 14614
rect 265306 14378 265542 14614
rect 264986 14058 265222 14294
rect 265306 14058 265542 14294
rect 264986 -3462 265222 -3226
rect 265306 -3462 265542 -3226
rect 264986 -3782 265222 -3546
rect 265306 -3782 265542 -3546
rect 268706 18098 268942 18334
rect 269026 18098 269262 18334
rect 268706 17778 268942 18014
rect 269026 17778 269262 18014
rect 268706 -4422 268942 -4186
rect 269026 -4422 269262 -4186
rect 268706 -4742 268942 -4506
rect 269026 -4742 269262 -4506
rect 272426 21818 272662 22054
rect 272746 21818 272982 22054
rect 272426 21498 272662 21734
rect 272746 21498 272982 21734
rect 272426 -5382 272662 -5146
rect 272746 -5382 272982 -5146
rect 272426 -5702 272662 -5466
rect 272746 -5702 272982 -5466
rect 276146 25538 276382 25774
rect 276466 25538 276702 25774
rect 276146 25218 276382 25454
rect 276466 25218 276702 25454
rect 276146 -6342 276382 -6106
rect 276466 -6342 276702 -6106
rect 276146 -6662 276382 -6426
rect 276466 -6662 276702 -6426
rect 279866 29258 280102 29494
rect 280186 29258 280422 29494
rect 279866 28938 280102 29174
rect 280186 28938 280422 29174
rect 279866 -7302 280102 -7066
rect 280186 -7302 280422 -7066
rect 279866 -7622 280102 -7386
rect 280186 -7622 280422 -7386
rect 289826 39218 290062 39454
rect 290146 39218 290382 39454
rect 289826 38898 290062 39134
rect 290146 38898 290382 39134
rect 289826 3218 290062 3454
rect 290146 3218 290382 3454
rect 289826 2898 290062 3134
rect 290146 2898 290382 3134
rect 289826 -582 290062 -346
rect 290146 -582 290382 -346
rect 289826 -902 290062 -666
rect 290146 -902 290382 -666
rect 293546 42938 293782 43174
rect 293866 42938 294102 43174
rect 293546 42618 293782 42854
rect 293866 42618 294102 42854
rect 293546 6938 293782 7174
rect 293866 6938 294102 7174
rect 293546 6618 293782 6854
rect 293866 6618 294102 6854
rect 293546 -1542 293782 -1306
rect 293866 -1542 294102 -1306
rect 293546 -1862 293782 -1626
rect 293866 -1862 294102 -1626
rect 297266 46658 297502 46894
rect 297586 46658 297822 46894
rect 297266 46338 297502 46574
rect 297586 46338 297822 46574
rect 297266 10658 297502 10894
rect 297586 10658 297822 10894
rect 297266 10338 297502 10574
rect 297586 10338 297822 10574
rect 297266 -2502 297502 -2266
rect 297586 -2502 297822 -2266
rect 297266 -2822 297502 -2586
rect 297586 -2822 297822 -2586
rect 300986 14378 301222 14614
rect 301306 14378 301542 14614
rect 300986 14058 301222 14294
rect 301306 14058 301542 14294
rect 300986 -3462 301222 -3226
rect 301306 -3462 301542 -3226
rect 300986 -3782 301222 -3546
rect 301306 -3782 301542 -3546
rect 304706 18098 304942 18334
rect 305026 18098 305262 18334
rect 304706 17778 304942 18014
rect 305026 17778 305262 18014
rect 304706 -4422 304942 -4186
rect 305026 -4422 305262 -4186
rect 304706 -4742 304942 -4506
rect 305026 -4742 305262 -4506
rect 308426 21818 308662 22054
rect 308746 21818 308982 22054
rect 308426 21498 308662 21734
rect 308746 21498 308982 21734
rect 308426 -5382 308662 -5146
rect 308746 -5382 308982 -5146
rect 308426 -5702 308662 -5466
rect 308746 -5702 308982 -5466
rect 312146 25538 312382 25774
rect 312466 25538 312702 25774
rect 312146 25218 312382 25454
rect 312466 25218 312702 25454
rect 312146 -6342 312382 -6106
rect 312466 -6342 312702 -6106
rect 312146 -6662 312382 -6426
rect 312466 -6662 312702 -6426
rect 315866 29258 316102 29494
rect 316186 29258 316422 29494
rect 315866 28938 316102 29174
rect 316186 28938 316422 29174
rect 315866 -7302 316102 -7066
rect 316186 -7302 316422 -7066
rect 315866 -7622 316102 -7386
rect 316186 -7622 316422 -7386
rect 325826 39218 326062 39454
rect 326146 39218 326382 39454
rect 325826 38898 326062 39134
rect 326146 38898 326382 39134
rect 325826 3218 326062 3454
rect 326146 3218 326382 3454
rect 325826 2898 326062 3134
rect 326146 2898 326382 3134
rect 325826 -582 326062 -346
rect 326146 -582 326382 -346
rect 325826 -902 326062 -666
rect 326146 -902 326382 -666
rect 329546 42938 329782 43174
rect 329866 42938 330102 43174
rect 329546 42618 329782 42854
rect 329866 42618 330102 42854
rect 329546 6938 329782 7174
rect 329866 6938 330102 7174
rect 329546 6618 329782 6854
rect 329866 6618 330102 6854
rect 329546 -1542 329782 -1306
rect 329866 -1542 330102 -1306
rect 329546 -1862 329782 -1626
rect 329866 -1862 330102 -1626
rect 333266 46658 333502 46894
rect 333586 46658 333822 46894
rect 333266 46338 333502 46574
rect 333586 46338 333822 46574
rect 333266 10658 333502 10894
rect 333586 10658 333822 10894
rect 333266 10338 333502 10574
rect 333586 10338 333822 10574
rect 333266 -2502 333502 -2266
rect 333586 -2502 333822 -2266
rect 333266 -2822 333502 -2586
rect 333586 -2822 333822 -2586
rect 336986 14378 337222 14614
rect 337306 14378 337542 14614
rect 336986 14058 337222 14294
rect 337306 14058 337542 14294
rect 336986 -3462 337222 -3226
rect 337306 -3462 337542 -3226
rect 336986 -3782 337222 -3546
rect 337306 -3782 337542 -3546
rect 340706 18098 340942 18334
rect 341026 18098 341262 18334
rect 340706 17778 340942 18014
rect 341026 17778 341262 18014
rect 340706 -4422 340942 -4186
rect 341026 -4422 341262 -4186
rect 340706 -4742 340942 -4506
rect 341026 -4742 341262 -4506
rect 344426 21818 344662 22054
rect 344746 21818 344982 22054
rect 344426 21498 344662 21734
rect 344746 21498 344982 21734
rect 344426 -5382 344662 -5146
rect 344746 -5382 344982 -5146
rect 344426 -5702 344662 -5466
rect 344746 -5702 344982 -5466
rect 348146 25538 348382 25774
rect 348466 25538 348702 25774
rect 348146 25218 348382 25454
rect 348466 25218 348702 25454
rect 348146 -6342 348382 -6106
rect 348466 -6342 348702 -6106
rect 348146 -6662 348382 -6426
rect 348466 -6662 348702 -6426
rect 351866 29258 352102 29494
rect 352186 29258 352422 29494
rect 351866 28938 352102 29174
rect 352186 28938 352422 29174
rect 351866 -7302 352102 -7066
rect 352186 -7302 352422 -7066
rect 351866 -7622 352102 -7386
rect 352186 -7622 352422 -7386
rect 361826 39218 362062 39454
rect 362146 39218 362382 39454
rect 361826 38898 362062 39134
rect 362146 38898 362382 39134
rect 361826 3218 362062 3454
rect 362146 3218 362382 3454
rect 361826 2898 362062 3134
rect 362146 2898 362382 3134
rect 361826 -582 362062 -346
rect 362146 -582 362382 -346
rect 361826 -902 362062 -666
rect 362146 -902 362382 -666
rect 365546 705562 365782 705798
rect 365866 705562 366102 705798
rect 365546 705242 365782 705478
rect 365866 705242 366102 705478
rect 365546 690938 365782 691174
rect 365866 690938 366102 691174
rect 365546 690618 365782 690854
rect 365866 690618 366102 690854
rect 365546 654938 365782 655174
rect 365866 654938 366102 655174
rect 365546 654618 365782 654854
rect 365866 654618 366102 654854
rect 365546 618938 365782 619174
rect 365866 618938 366102 619174
rect 365546 618618 365782 618854
rect 365866 618618 366102 618854
rect 365546 582938 365782 583174
rect 365866 582938 366102 583174
rect 365546 582618 365782 582854
rect 365866 582618 366102 582854
rect 365546 546938 365782 547174
rect 365866 546938 366102 547174
rect 365546 546618 365782 546854
rect 365866 546618 366102 546854
rect 365546 510938 365782 511174
rect 365866 510938 366102 511174
rect 365546 510618 365782 510854
rect 365866 510618 366102 510854
rect 365546 474938 365782 475174
rect 365866 474938 366102 475174
rect 365546 474618 365782 474854
rect 365866 474618 366102 474854
rect 365546 438938 365782 439174
rect 365866 438938 366102 439174
rect 365546 438618 365782 438854
rect 365866 438618 366102 438854
rect 365546 402938 365782 403174
rect 365866 402938 366102 403174
rect 365546 402618 365782 402854
rect 365866 402618 366102 402854
rect 365546 366938 365782 367174
rect 365866 366938 366102 367174
rect 365546 366618 365782 366854
rect 365866 366618 366102 366854
rect 365546 330938 365782 331174
rect 365866 330938 366102 331174
rect 365546 330618 365782 330854
rect 365866 330618 366102 330854
rect 365546 294938 365782 295174
rect 365866 294938 366102 295174
rect 365546 294618 365782 294854
rect 365866 294618 366102 294854
rect 365546 258938 365782 259174
rect 365866 258938 366102 259174
rect 365546 258618 365782 258854
rect 365866 258618 366102 258854
rect 365546 222938 365782 223174
rect 365866 222938 366102 223174
rect 365546 222618 365782 222854
rect 365866 222618 366102 222854
rect 365546 186938 365782 187174
rect 365866 186938 366102 187174
rect 365546 186618 365782 186854
rect 365866 186618 366102 186854
rect 365546 150938 365782 151174
rect 365866 150938 366102 151174
rect 365546 150618 365782 150854
rect 365866 150618 366102 150854
rect 365546 114938 365782 115174
rect 365866 114938 366102 115174
rect 365546 114618 365782 114854
rect 365866 114618 366102 114854
rect 365546 78938 365782 79174
rect 365866 78938 366102 79174
rect 365546 78618 365782 78854
rect 365866 78618 366102 78854
rect 365546 42938 365782 43174
rect 365866 42938 366102 43174
rect 365546 42618 365782 42854
rect 365866 42618 366102 42854
rect 365546 6938 365782 7174
rect 365866 6938 366102 7174
rect 365546 6618 365782 6854
rect 365866 6618 366102 6854
rect 365546 -1542 365782 -1306
rect 365866 -1542 366102 -1306
rect 365546 -1862 365782 -1626
rect 365866 -1862 366102 -1626
rect 369266 706522 369502 706758
rect 369586 706522 369822 706758
rect 369266 706202 369502 706438
rect 369586 706202 369822 706438
rect 369266 694658 369502 694894
rect 369586 694658 369822 694894
rect 369266 694338 369502 694574
rect 369586 694338 369822 694574
rect 369266 658658 369502 658894
rect 369586 658658 369822 658894
rect 369266 658338 369502 658574
rect 369586 658338 369822 658574
rect 369266 622658 369502 622894
rect 369586 622658 369822 622894
rect 369266 622338 369502 622574
rect 369586 622338 369822 622574
rect 369266 586658 369502 586894
rect 369586 586658 369822 586894
rect 369266 586338 369502 586574
rect 369586 586338 369822 586574
rect 369266 550658 369502 550894
rect 369586 550658 369822 550894
rect 369266 550338 369502 550574
rect 369586 550338 369822 550574
rect 369266 514658 369502 514894
rect 369586 514658 369822 514894
rect 369266 514338 369502 514574
rect 369586 514338 369822 514574
rect 369266 478658 369502 478894
rect 369586 478658 369822 478894
rect 369266 478338 369502 478574
rect 369586 478338 369822 478574
rect 369266 442658 369502 442894
rect 369586 442658 369822 442894
rect 369266 442338 369502 442574
rect 369586 442338 369822 442574
rect 369266 406658 369502 406894
rect 369586 406658 369822 406894
rect 369266 406338 369502 406574
rect 369586 406338 369822 406574
rect 369266 370658 369502 370894
rect 369586 370658 369822 370894
rect 369266 370338 369502 370574
rect 369586 370338 369822 370574
rect 369266 334658 369502 334894
rect 369586 334658 369822 334894
rect 369266 334338 369502 334574
rect 369586 334338 369822 334574
rect 369266 298658 369502 298894
rect 369586 298658 369822 298894
rect 369266 298338 369502 298574
rect 369586 298338 369822 298574
rect 369266 262658 369502 262894
rect 369586 262658 369822 262894
rect 369266 262338 369502 262574
rect 369586 262338 369822 262574
rect 369266 226658 369502 226894
rect 369586 226658 369822 226894
rect 369266 226338 369502 226574
rect 369586 226338 369822 226574
rect 369266 190658 369502 190894
rect 369586 190658 369822 190894
rect 369266 190338 369502 190574
rect 369586 190338 369822 190574
rect 369266 154658 369502 154894
rect 369586 154658 369822 154894
rect 369266 154338 369502 154574
rect 369586 154338 369822 154574
rect 369266 118658 369502 118894
rect 369586 118658 369822 118894
rect 369266 118338 369502 118574
rect 369586 118338 369822 118574
rect 369266 82658 369502 82894
rect 369586 82658 369822 82894
rect 369266 82338 369502 82574
rect 369586 82338 369822 82574
rect 369266 46658 369502 46894
rect 369586 46658 369822 46894
rect 369266 46338 369502 46574
rect 369586 46338 369822 46574
rect 369266 10658 369502 10894
rect 369586 10658 369822 10894
rect 369266 10338 369502 10574
rect 369586 10338 369822 10574
rect 369266 -2502 369502 -2266
rect 369586 -2502 369822 -2266
rect 369266 -2822 369502 -2586
rect 369586 -2822 369822 -2586
rect 372986 707482 373222 707718
rect 373306 707482 373542 707718
rect 372986 707162 373222 707398
rect 373306 707162 373542 707398
rect 372986 698378 373222 698614
rect 373306 698378 373542 698614
rect 372986 698058 373222 698294
rect 373306 698058 373542 698294
rect 372986 662378 373222 662614
rect 373306 662378 373542 662614
rect 372986 662058 373222 662294
rect 373306 662058 373542 662294
rect 372986 626378 373222 626614
rect 373306 626378 373542 626614
rect 372986 626058 373222 626294
rect 373306 626058 373542 626294
rect 372986 590378 373222 590614
rect 373306 590378 373542 590614
rect 372986 590058 373222 590294
rect 373306 590058 373542 590294
rect 372986 554378 373222 554614
rect 373306 554378 373542 554614
rect 372986 554058 373222 554294
rect 373306 554058 373542 554294
rect 372986 518378 373222 518614
rect 373306 518378 373542 518614
rect 372986 518058 373222 518294
rect 373306 518058 373542 518294
rect 372986 482378 373222 482614
rect 373306 482378 373542 482614
rect 372986 482058 373222 482294
rect 373306 482058 373542 482294
rect 372986 446378 373222 446614
rect 373306 446378 373542 446614
rect 372986 446058 373222 446294
rect 373306 446058 373542 446294
rect 372986 410378 373222 410614
rect 373306 410378 373542 410614
rect 372986 410058 373222 410294
rect 373306 410058 373542 410294
rect 372986 374378 373222 374614
rect 373306 374378 373542 374614
rect 372986 374058 373222 374294
rect 373306 374058 373542 374294
rect 372986 338378 373222 338614
rect 373306 338378 373542 338614
rect 372986 338058 373222 338294
rect 373306 338058 373542 338294
rect 372986 302378 373222 302614
rect 373306 302378 373542 302614
rect 372986 302058 373222 302294
rect 373306 302058 373542 302294
rect 372986 266378 373222 266614
rect 373306 266378 373542 266614
rect 372986 266058 373222 266294
rect 373306 266058 373542 266294
rect 372986 230378 373222 230614
rect 373306 230378 373542 230614
rect 372986 230058 373222 230294
rect 373306 230058 373542 230294
rect 372986 194378 373222 194614
rect 373306 194378 373542 194614
rect 372986 194058 373222 194294
rect 373306 194058 373542 194294
rect 372986 158378 373222 158614
rect 373306 158378 373542 158614
rect 372986 158058 373222 158294
rect 373306 158058 373542 158294
rect 372986 122378 373222 122614
rect 373306 122378 373542 122614
rect 372986 122058 373222 122294
rect 373306 122058 373542 122294
rect 372986 86378 373222 86614
rect 373306 86378 373542 86614
rect 372986 86058 373222 86294
rect 373306 86058 373542 86294
rect 372986 50378 373222 50614
rect 373306 50378 373542 50614
rect 372986 50058 373222 50294
rect 373306 50058 373542 50294
rect 372986 14378 373222 14614
rect 373306 14378 373542 14614
rect 372986 14058 373222 14294
rect 373306 14058 373542 14294
rect 372986 -3462 373222 -3226
rect 373306 -3462 373542 -3226
rect 372986 -3782 373222 -3546
rect 373306 -3782 373542 -3546
rect 376706 708442 376942 708678
rect 377026 708442 377262 708678
rect 376706 708122 376942 708358
rect 377026 708122 377262 708358
rect 376706 666098 376942 666334
rect 377026 666098 377262 666334
rect 376706 665778 376942 666014
rect 377026 665778 377262 666014
rect 376706 630098 376942 630334
rect 377026 630098 377262 630334
rect 376706 629778 376942 630014
rect 377026 629778 377262 630014
rect 376706 594098 376942 594334
rect 377026 594098 377262 594334
rect 376706 593778 376942 594014
rect 377026 593778 377262 594014
rect 376706 558098 376942 558334
rect 377026 558098 377262 558334
rect 376706 557778 376942 558014
rect 377026 557778 377262 558014
rect 376706 522098 376942 522334
rect 377026 522098 377262 522334
rect 376706 521778 376942 522014
rect 377026 521778 377262 522014
rect 376706 486098 376942 486334
rect 377026 486098 377262 486334
rect 376706 485778 376942 486014
rect 377026 485778 377262 486014
rect 376706 450098 376942 450334
rect 377026 450098 377262 450334
rect 376706 449778 376942 450014
rect 377026 449778 377262 450014
rect 376706 414098 376942 414334
rect 377026 414098 377262 414334
rect 376706 413778 376942 414014
rect 377026 413778 377262 414014
rect 376706 378098 376942 378334
rect 377026 378098 377262 378334
rect 376706 377778 376942 378014
rect 377026 377778 377262 378014
rect 376706 342098 376942 342334
rect 377026 342098 377262 342334
rect 376706 341778 376942 342014
rect 377026 341778 377262 342014
rect 376706 306098 376942 306334
rect 377026 306098 377262 306334
rect 376706 305778 376942 306014
rect 377026 305778 377262 306014
rect 376706 270098 376942 270334
rect 377026 270098 377262 270334
rect 376706 269778 376942 270014
rect 377026 269778 377262 270014
rect 376706 234098 376942 234334
rect 377026 234098 377262 234334
rect 376706 233778 376942 234014
rect 377026 233778 377262 234014
rect 376706 198098 376942 198334
rect 377026 198098 377262 198334
rect 376706 197778 376942 198014
rect 377026 197778 377262 198014
rect 376706 162098 376942 162334
rect 377026 162098 377262 162334
rect 376706 161778 376942 162014
rect 377026 161778 377262 162014
rect 376706 126098 376942 126334
rect 377026 126098 377262 126334
rect 376706 125778 376942 126014
rect 377026 125778 377262 126014
rect 376706 90098 376942 90334
rect 377026 90098 377262 90334
rect 376706 89778 376942 90014
rect 377026 89778 377262 90014
rect 376706 54098 376942 54334
rect 377026 54098 377262 54334
rect 376706 53778 376942 54014
rect 377026 53778 377262 54014
rect 376706 18098 376942 18334
rect 377026 18098 377262 18334
rect 376706 17778 376942 18014
rect 377026 17778 377262 18014
rect 376706 -4422 376942 -4186
rect 377026 -4422 377262 -4186
rect 376706 -4742 376942 -4506
rect 377026 -4742 377262 -4506
rect 380426 709402 380662 709638
rect 380746 709402 380982 709638
rect 380426 709082 380662 709318
rect 380746 709082 380982 709318
rect 380426 669818 380662 670054
rect 380746 669818 380982 670054
rect 380426 669498 380662 669734
rect 380746 669498 380982 669734
rect 380426 633818 380662 634054
rect 380746 633818 380982 634054
rect 380426 633498 380662 633734
rect 380746 633498 380982 633734
rect 380426 597818 380662 598054
rect 380746 597818 380982 598054
rect 380426 597498 380662 597734
rect 380746 597498 380982 597734
rect 380426 561818 380662 562054
rect 380746 561818 380982 562054
rect 380426 561498 380662 561734
rect 380746 561498 380982 561734
rect 380426 525818 380662 526054
rect 380746 525818 380982 526054
rect 380426 525498 380662 525734
rect 380746 525498 380982 525734
rect 380426 489818 380662 490054
rect 380746 489818 380982 490054
rect 380426 489498 380662 489734
rect 380746 489498 380982 489734
rect 380426 453818 380662 454054
rect 380746 453818 380982 454054
rect 380426 453498 380662 453734
rect 380746 453498 380982 453734
rect 380426 417818 380662 418054
rect 380746 417818 380982 418054
rect 380426 417498 380662 417734
rect 380746 417498 380982 417734
rect 380426 381818 380662 382054
rect 380746 381818 380982 382054
rect 380426 381498 380662 381734
rect 380746 381498 380982 381734
rect 380426 345818 380662 346054
rect 380746 345818 380982 346054
rect 380426 345498 380662 345734
rect 380746 345498 380982 345734
rect 380426 309818 380662 310054
rect 380746 309818 380982 310054
rect 380426 309498 380662 309734
rect 380746 309498 380982 309734
rect 380426 273818 380662 274054
rect 380746 273818 380982 274054
rect 380426 273498 380662 273734
rect 380746 273498 380982 273734
rect 380426 237818 380662 238054
rect 380746 237818 380982 238054
rect 380426 237498 380662 237734
rect 380746 237498 380982 237734
rect 380426 201818 380662 202054
rect 380746 201818 380982 202054
rect 380426 201498 380662 201734
rect 380746 201498 380982 201734
rect 380426 165818 380662 166054
rect 380746 165818 380982 166054
rect 380426 165498 380662 165734
rect 380746 165498 380982 165734
rect 380426 129818 380662 130054
rect 380746 129818 380982 130054
rect 380426 129498 380662 129734
rect 380746 129498 380982 129734
rect 380426 93818 380662 94054
rect 380746 93818 380982 94054
rect 380426 93498 380662 93734
rect 380746 93498 380982 93734
rect 380426 57818 380662 58054
rect 380746 57818 380982 58054
rect 380426 57498 380662 57734
rect 380746 57498 380982 57734
rect 380426 21818 380662 22054
rect 380746 21818 380982 22054
rect 380426 21498 380662 21734
rect 380746 21498 380982 21734
rect 380426 -5382 380662 -5146
rect 380746 -5382 380982 -5146
rect 380426 -5702 380662 -5466
rect 380746 -5702 380982 -5466
rect 384146 710362 384382 710598
rect 384466 710362 384702 710598
rect 384146 710042 384382 710278
rect 384466 710042 384702 710278
rect 384146 673538 384382 673774
rect 384466 673538 384702 673774
rect 384146 673218 384382 673454
rect 384466 673218 384702 673454
rect 384146 637538 384382 637774
rect 384466 637538 384702 637774
rect 384146 637218 384382 637454
rect 384466 637218 384702 637454
rect 384146 601538 384382 601774
rect 384466 601538 384702 601774
rect 384146 601218 384382 601454
rect 384466 601218 384702 601454
rect 384146 565538 384382 565774
rect 384466 565538 384702 565774
rect 384146 565218 384382 565454
rect 384466 565218 384702 565454
rect 384146 529538 384382 529774
rect 384466 529538 384702 529774
rect 384146 529218 384382 529454
rect 384466 529218 384702 529454
rect 384146 493538 384382 493774
rect 384466 493538 384702 493774
rect 384146 493218 384382 493454
rect 384466 493218 384702 493454
rect 384146 457538 384382 457774
rect 384466 457538 384702 457774
rect 384146 457218 384382 457454
rect 384466 457218 384702 457454
rect 384146 421538 384382 421774
rect 384466 421538 384702 421774
rect 384146 421218 384382 421454
rect 384466 421218 384702 421454
rect 384146 385538 384382 385774
rect 384466 385538 384702 385774
rect 384146 385218 384382 385454
rect 384466 385218 384702 385454
rect 384146 349538 384382 349774
rect 384466 349538 384702 349774
rect 384146 349218 384382 349454
rect 384466 349218 384702 349454
rect 384146 313538 384382 313774
rect 384466 313538 384702 313774
rect 384146 313218 384382 313454
rect 384466 313218 384702 313454
rect 384146 277538 384382 277774
rect 384466 277538 384702 277774
rect 384146 277218 384382 277454
rect 384466 277218 384702 277454
rect 384146 241538 384382 241774
rect 384466 241538 384702 241774
rect 384146 241218 384382 241454
rect 384466 241218 384702 241454
rect 384146 205538 384382 205774
rect 384466 205538 384702 205774
rect 384146 205218 384382 205454
rect 384466 205218 384702 205454
rect 384146 169538 384382 169774
rect 384466 169538 384702 169774
rect 384146 169218 384382 169454
rect 384466 169218 384702 169454
rect 384146 133538 384382 133774
rect 384466 133538 384702 133774
rect 384146 133218 384382 133454
rect 384466 133218 384702 133454
rect 384146 97538 384382 97774
rect 384466 97538 384702 97774
rect 384146 97218 384382 97454
rect 384466 97218 384702 97454
rect 384146 61538 384382 61774
rect 384466 61538 384702 61774
rect 384146 61218 384382 61454
rect 384466 61218 384702 61454
rect 384146 25538 384382 25774
rect 384466 25538 384702 25774
rect 384146 25218 384382 25454
rect 384466 25218 384702 25454
rect 384146 -6342 384382 -6106
rect 384466 -6342 384702 -6106
rect 384146 -6662 384382 -6426
rect 384466 -6662 384702 -6426
rect 387866 711322 388102 711558
rect 388186 711322 388422 711558
rect 387866 711002 388102 711238
rect 388186 711002 388422 711238
rect 387866 677258 388102 677494
rect 388186 677258 388422 677494
rect 387866 676938 388102 677174
rect 388186 676938 388422 677174
rect 387866 641258 388102 641494
rect 388186 641258 388422 641494
rect 387866 640938 388102 641174
rect 388186 640938 388422 641174
rect 387866 605258 388102 605494
rect 388186 605258 388422 605494
rect 387866 604938 388102 605174
rect 388186 604938 388422 605174
rect 387866 569258 388102 569494
rect 388186 569258 388422 569494
rect 387866 568938 388102 569174
rect 388186 568938 388422 569174
rect 387866 533258 388102 533494
rect 388186 533258 388422 533494
rect 387866 532938 388102 533174
rect 388186 532938 388422 533174
rect 387866 497258 388102 497494
rect 388186 497258 388422 497494
rect 387866 496938 388102 497174
rect 388186 496938 388422 497174
rect 387866 461258 388102 461494
rect 388186 461258 388422 461494
rect 387866 460938 388102 461174
rect 388186 460938 388422 461174
rect 387866 425258 388102 425494
rect 388186 425258 388422 425494
rect 387866 424938 388102 425174
rect 388186 424938 388422 425174
rect 387866 389258 388102 389494
rect 388186 389258 388422 389494
rect 387866 388938 388102 389174
rect 388186 388938 388422 389174
rect 387866 353258 388102 353494
rect 388186 353258 388422 353494
rect 387866 352938 388102 353174
rect 388186 352938 388422 353174
rect 387866 317258 388102 317494
rect 388186 317258 388422 317494
rect 387866 316938 388102 317174
rect 388186 316938 388422 317174
rect 387866 281258 388102 281494
rect 388186 281258 388422 281494
rect 387866 280938 388102 281174
rect 388186 280938 388422 281174
rect 387866 245258 388102 245494
rect 388186 245258 388422 245494
rect 387866 244938 388102 245174
rect 388186 244938 388422 245174
rect 387866 209258 388102 209494
rect 388186 209258 388422 209494
rect 387866 208938 388102 209174
rect 388186 208938 388422 209174
rect 387866 173258 388102 173494
rect 388186 173258 388422 173494
rect 387866 172938 388102 173174
rect 388186 172938 388422 173174
rect 387866 137258 388102 137494
rect 388186 137258 388422 137494
rect 387866 136938 388102 137174
rect 388186 136938 388422 137174
rect 387866 101258 388102 101494
rect 388186 101258 388422 101494
rect 387866 100938 388102 101174
rect 388186 100938 388422 101174
rect 387866 65258 388102 65494
rect 388186 65258 388422 65494
rect 387866 64938 388102 65174
rect 388186 64938 388422 65174
rect 387866 29258 388102 29494
rect 388186 29258 388422 29494
rect 387866 28938 388102 29174
rect 388186 28938 388422 29174
rect 387866 -7302 388102 -7066
rect 388186 -7302 388422 -7066
rect 387866 -7622 388102 -7386
rect 388186 -7622 388422 -7386
rect 397826 704602 398062 704838
rect 398146 704602 398382 704838
rect 397826 704282 398062 704518
rect 398146 704282 398382 704518
rect 397826 687218 398062 687454
rect 398146 687218 398382 687454
rect 397826 686898 398062 687134
rect 398146 686898 398382 687134
rect 397826 651218 398062 651454
rect 398146 651218 398382 651454
rect 397826 650898 398062 651134
rect 398146 650898 398382 651134
rect 397826 615218 398062 615454
rect 398146 615218 398382 615454
rect 397826 614898 398062 615134
rect 398146 614898 398382 615134
rect 397826 579218 398062 579454
rect 398146 579218 398382 579454
rect 397826 578898 398062 579134
rect 398146 578898 398382 579134
rect 397826 543218 398062 543454
rect 398146 543218 398382 543454
rect 397826 542898 398062 543134
rect 398146 542898 398382 543134
rect 397826 507218 398062 507454
rect 398146 507218 398382 507454
rect 397826 506898 398062 507134
rect 398146 506898 398382 507134
rect 397826 471218 398062 471454
rect 398146 471218 398382 471454
rect 397826 470898 398062 471134
rect 398146 470898 398382 471134
rect 397826 435218 398062 435454
rect 398146 435218 398382 435454
rect 397826 434898 398062 435134
rect 398146 434898 398382 435134
rect 397826 399218 398062 399454
rect 398146 399218 398382 399454
rect 397826 398898 398062 399134
rect 398146 398898 398382 399134
rect 397826 363218 398062 363454
rect 398146 363218 398382 363454
rect 397826 362898 398062 363134
rect 398146 362898 398382 363134
rect 397826 327218 398062 327454
rect 398146 327218 398382 327454
rect 397826 326898 398062 327134
rect 398146 326898 398382 327134
rect 397826 291218 398062 291454
rect 398146 291218 398382 291454
rect 397826 290898 398062 291134
rect 398146 290898 398382 291134
rect 397826 255218 398062 255454
rect 398146 255218 398382 255454
rect 397826 254898 398062 255134
rect 398146 254898 398382 255134
rect 397826 219218 398062 219454
rect 398146 219218 398382 219454
rect 397826 218898 398062 219134
rect 398146 218898 398382 219134
rect 397826 183218 398062 183454
rect 398146 183218 398382 183454
rect 397826 182898 398062 183134
rect 398146 182898 398382 183134
rect 397826 147218 398062 147454
rect 398146 147218 398382 147454
rect 397826 146898 398062 147134
rect 398146 146898 398382 147134
rect 397826 111218 398062 111454
rect 398146 111218 398382 111454
rect 397826 110898 398062 111134
rect 398146 110898 398382 111134
rect 397826 75218 398062 75454
rect 398146 75218 398382 75454
rect 397826 74898 398062 75134
rect 398146 74898 398382 75134
rect 397826 39218 398062 39454
rect 398146 39218 398382 39454
rect 397826 38898 398062 39134
rect 398146 38898 398382 39134
rect 397826 3218 398062 3454
rect 398146 3218 398382 3454
rect 397826 2898 398062 3134
rect 398146 2898 398382 3134
rect 397826 -582 398062 -346
rect 398146 -582 398382 -346
rect 397826 -902 398062 -666
rect 398146 -902 398382 -666
rect 401546 705562 401782 705798
rect 401866 705562 402102 705798
rect 401546 705242 401782 705478
rect 401866 705242 402102 705478
rect 401546 690938 401782 691174
rect 401866 690938 402102 691174
rect 401546 690618 401782 690854
rect 401866 690618 402102 690854
rect 401546 654938 401782 655174
rect 401866 654938 402102 655174
rect 401546 654618 401782 654854
rect 401866 654618 402102 654854
rect 401546 618938 401782 619174
rect 401866 618938 402102 619174
rect 401546 618618 401782 618854
rect 401866 618618 402102 618854
rect 401546 582938 401782 583174
rect 401866 582938 402102 583174
rect 401546 582618 401782 582854
rect 401866 582618 402102 582854
rect 401546 546938 401782 547174
rect 401866 546938 402102 547174
rect 401546 546618 401782 546854
rect 401866 546618 402102 546854
rect 401546 510938 401782 511174
rect 401866 510938 402102 511174
rect 401546 510618 401782 510854
rect 401866 510618 402102 510854
rect 401546 474938 401782 475174
rect 401866 474938 402102 475174
rect 401546 474618 401782 474854
rect 401866 474618 402102 474854
rect 401546 438938 401782 439174
rect 401866 438938 402102 439174
rect 401546 438618 401782 438854
rect 401866 438618 402102 438854
rect 401546 402938 401782 403174
rect 401866 402938 402102 403174
rect 401546 402618 401782 402854
rect 401866 402618 402102 402854
rect 401546 366938 401782 367174
rect 401866 366938 402102 367174
rect 401546 366618 401782 366854
rect 401866 366618 402102 366854
rect 401546 330938 401782 331174
rect 401866 330938 402102 331174
rect 401546 330618 401782 330854
rect 401866 330618 402102 330854
rect 405266 706522 405502 706758
rect 405586 706522 405822 706758
rect 405266 706202 405502 706438
rect 405586 706202 405822 706438
rect 405266 694658 405502 694894
rect 405586 694658 405822 694894
rect 405266 694338 405502 694574
rect 405586 694338 405822 694574
rect 405266 658658 405502 658894
rect 405586 658658 405822 658894
rect 405266 658338 405502 658574
rect 405586 658338 405822 658574
rect 405266 622658 405502 622894
rect 405586 622658 405822 622894
rect 405266 622338 405502 622574
rect 405586 622338 405822 622574
rect 405266 586658 405502 586894
rect 405586 586658 405822 586894
rect 405266 586338 405502 586574
rect 405586 586338 405822 586574
rect 405266 550658 405502 550894
rect 405586 550658 405822 550894
rect 405266 550338 405502 550574
rect 405586 550338 405822 550574
rect 405266 514658 405502 514894
rect 405586 514658 405822 514894
rect 405266 514338 405502 514574
rect 405586 514338 405822 514574
rect 405266 478658 405502 478894
rect 405586 478658 405822 478894
rect 405266 478338 405502 478574
rect 405586 478338 405822 478574
rect 405266 442658 405502 442894
rect 405586 442658 405822 442894
rect 405266 442338 405502 442574
rect 405586 442338 405822 442574
rect 405266 406658 405502 406894
rect 405586 406658 405822 406894
rect 405266 406338 405502 406574
rect 405586 406338 405822 406574
rect 405266 370658 405502 370894
rect 405586 370658 405822 370894
rect 405266 370338 405502 370574
rect 405586 370338 405822 370574
rect 405266 334658 405502 334894
rect 405586 334658 405822 334894
rect 405266 334338 405502 334574
rect 405586 334338 405822 334574
rect 404459 327218 404695 327454
rect 404459 326898 404695 327134
rect 401546 294938 401782 295174
rect 401866 294938 402102 295174
rect 401546 294618 401782 294854
rect 401866 294618 402102 294854
rect 401546 258938 401782 259174
rect 401866 258938 402102 259174
rect 401546 258618 401782 258854
rect 401866 258618 402102 258854
rect 401546 222938 401782 223174
rect 401866 222938 402102 223174
rect 401546 222618 401782 222854
rect 401866 222618 402102 222854
rect 401546 186938 401782 187174
rect 401866 186938 402102 187174
rect 401546 186618 401782 186854
rect 401866 186618 402102 186854
rect 401546 150938 401782 151174
rect 401866 150938 402102 151174
rect 401546 150618 401782 150854
rect 401866 150618 402102 150854
rect 401546 114938 401782 115174
rect 401866 114938 402102 115174
rect 401546 114618 401782 114854
rect 401866 114618 402102 114854
rect 401546 78938 401782 79174
rect 401866 78938 402102 79174
rect 401546 78618 401782 78854
rect 401866 78618 402102 78854
rect 401546 42938 401782 43174
rect 401866 42938 402102 43174
rect 401546 42618 401782 42854
rect 401866 42618 402102 42854
rect 401546 6938 401782 7174
rect 401866 6938 402102 7174
rect 401546 6618 401782 6854
rect 401866 6618 402102 6854
rect 401546 -1542 401782 -1306
rect 401866 -1542 402102 -1306
rect 401546 -1862 401782 -1626
rect 401866 -1862 402102 -1626
rect 408986 707482 409222 707718
rect 409306 707482 409542 707718
rect 408986 707162 409222 707398
rect 409306 707162 409542 707398
rect 408986 698378 409222 698614
rect 409306 698378 409542 698614
rect 408986 698058 409222 698294
rect 409306 698058 409542 698294
rect 408986 662378 409222 662614
rect 409306 662378 409542 662614
rect 408986 662058 409222 662294
rect 409306 662058 409542 662294
rect 408986 626378 409222 626614
rect 409306 626378 409542 626614
rect 408986 626058 409222 626294
rect 409306 626058 409542 626294
rect 408986 590378 409222 590614
rect 409306 590378 409542 590614
rect 408986 590058 409222 590294
rect 409306 590058 409542 590294
rect 408986 554378 409222 554614
rect 409306 554378 409542 554614
rect 408986 554058 409222 554294
rect 409306 554058 409542 554294
rect 408986 518378 409222 518614
rect 409306 518378 409542 518614
rect 408986 518058 409222 518294
rect 409306 518058 409542 518294
rect 408986 482378 409222 482614
rect 409306 482378 409542 482614
rect 408986 482058 409222 482294
rect 409306 482058 409542 482294
rect 408986 446378 409222 446614
rect 409306 446378 409542 446614
rect 408986 446058 409222 446294
rect 409306 446058 409542 446294
rect 408986 410378 409222 410614
rect 409306 410378 409542 410614
rect 408986 410058 409222 410294
rect 409306 410058 409542 410294
rect 408986 374378 409222 374614
rect 409306 374378 409542 374614
rect 408986 374058 409222 374294
rect 409306 374058 409542 374294
rect 408986 338378 409222 338614
rect 409306 338378 409542 338614
rect 408986 338058 409222 338294
rect 409306 338058 409542 338294
rect 407932 330938 408168 331174
rect 407932 330618 408168 330854
rect 405266 298658 405502 298894
rect 405586 298658 405822 298894
rect 405266 298338 405502 298574
rect 405586 298338 405822 298574
rect 405266 262658 405502 262894
rect 405586 262658 405822 262894
rect 405266 262338 405502 262574
rect 405586 262338 405822 262574
rect 405266 226658 405502 226894
rect 405586 226658 405822 226894
rect 405266 226338 405502 226574
rect 405586 226338 405822 226574
rect 405266 190658 405502 190894
rect 405586 190658 405822 190894
rect 405266 190338 405502 190574
rect 405586 190338 405822 190574
rect 405266 154658 405502 154894
rect 405586 154658 405822 154894
rect 405266 154338 405502 154574
rect 405586 154338 405822 154574
rect 405266 118658 405502 118894
rect 405586 118658 405822 118894
rect 405266 118338 405502 118574
rect 405586 118338 405822 118574
rect 405266 82658 405502 82894
rect 405586 82658 405822 82894
rect 405266 82338 405502 82574
rect 405586 82338 405822 82574
rect 405266 46658 405502 46894
rect 405586 46658 405822 46894
rect 405266 46338 405502 46574
rect 405586 46338 405822 46574
rect 405266 10658 405502 10894
rect 405586 10658 405822 10894
rect 405266 10338 405502 10574
rect 405586 10338 405822 10574
rect 405266 -2502 405502 -2266
rect 405586 -2502 405822 -2266
rect 405266 -2822 405502 -2586
rect 405586 -2822 405822 -2586
rect 412706 708442 412942 708678
rect 413026 708442 413262 708678
rect 412706 708122 412942 708358
rect 413026 708122 413262 708358
rect 412706 666098 412942 666334
rect 413026 666098 413262 666334
rect 412706 665778 412942 666014
rect 413026 665778 413262 666014
rect 412706 630098 412942 630334
rect 413026 630098 413262 630334
rect 412706 629778 412942 630014
rect 413026 629778 413262 630014
rect 412706 594098 412942 594334
rect 413026 594098 413262 594334
rect 412706 593778 412942 594014
rect 413026 593778 413262 594014
rect 412706 558098 412942 558334
rect 413026 558098 413262 558334
rect 412706 557778 412942 558014
rect 413026 557778 413262 558014
rect 412706 522098 412942 522334
rect 413026 522098 413262 522334
rect 412706 521778 412942 522014
rect 413026 521778 413262 522014
rect 412706 486098 412942 486334
rect 413026 486098 413262 486334
rect 412706 485778 412942 486014
rect 413026 485778 413262 486014
rect 412706 450098 412942 450334
rect 413026 450098 413262 450334
rect 412706 449778 412942 450014
rect 413026 449778 413262 450014
rect 412706 414098 412942 414334
rect 413026 414098 413262 414334
rect 412706 413778 412942 414014
rect 413026 413778 413262 414014
rect 412706 378098 412942 378334
rect 413026 378098 413262 378334
rect 412706 377778 412942 378014
rect 413026 377778 413262 378014
rect 412706 342098 412942 342334
rect 413026 342098 413262 342334
rect 412706 341778 412942 342014
rect 413026 341778 413262 342014
rect 411405 327218 411641 327454
rect 411405 326898 411641 327134
rect 408986 302378 409222 302614
rect 409306 302378 409542 302614
rect 408986 302058 409222 302294
rect 409306 302058 409542 302294
rect 408986 266378 409222 266614
rect 409306 266378 409542 266614
rect 408986 266058 409222 266294
rect 409306 266058 409542 266294
rect 408986 230378 409222 230614
rect 409306 230378 409542 230614
rect 408986 230058 409222 230294
rect 409306 230058 409542 230294
rect 408986 194378 409222 194614
rect 409306 194378 409542 194614
rect 408986 194058 409222 194294
rect 409306 194058 409542 194294
rect 408986 158378 409222 158614
rect 409306 158378 409542 158614
rect 408986 158058 409222 158294
rect 409306 158058 409542 158294
rect 408986 122378 409222 122614
rect 409306 122378 409542 122614
rect 408986 122058 409222 122294
rect 409306 122058 409542 122294
rect 408986 86378 409222 86614
rect 409306 86378 409542 86614
rect 408986 86058 409222 86294
rect 409306 86058 409542 86294
rect 408986 50378 409222 50614
rect 409306 50378 409542 50614
rect 408986 50058 409222 50294
rect 409306 50058 409542 50294
rect 408986 14378 409222 14614
rect 409306 14378 409542 14614
rect 408986 14058 409222 14294
rect 409306 14058 409542 14294
rect 408986 -3462 409222 -3226
rect 409306 -3462 409542 -3226
rect 408986 -3782 409222 -3546
rect 409306 -3782 409542 -3546
rect 416426 709402 416662 709638
rect 416746 709402 416982 709638
rect 416426 709082 416662 709318
rect 416746 709082 416982 709318
rect 416426 669818 416662 670054
rect 416746 669818 416982 670054
rect 416426 669498 416662 669734
rect 416746 669498 416982 669734
rect 416426 633818 416662 634054
rect 416746 633818 416982 634054
rect 416426 633498 416662 633734
rect 416746 633498 416982 633734
rect 416426 597818 416662 598054
rect 416746 597818 416982 598054
rect 416426 597498 416662 597734
rect 416746 597498 416982 597734
rect 416426 561818 416662 562054
rect 416746 561818 416982 562054
rect 416426 561498 416662 561734
rect 416746 561498 416982 561734
rect 416426 525818 416662 526054
rect 416746 525818 416982 526054
rect 416426 525498 416662 525734
rect 416746 525498 416982 525734
rect 416426 489818 416662 490054
rect 416746 489818 416982 490054
rect 416426 489498 416662 489734
rect 416746 489498 416982 489734
rect 416426 453818 416662 454054
rect 416746 453818 416982 454054
rect 416426 453498 416662 453734
rect 416746 453498 416982 453734
rect 416426 417818 416662 418054
rect 416746 417818 416982 418054
rect 416426 417498 416662 417734
rect 416746 417498 416982 417734
rect 416426 381818 416662 382054
rect 416746 381818 416982 382054
rect 416426 381498 416662 381734
rect 416746 381498 416982 381734
rect 416426 345818 416662 346054
rect 416746 345818 416982 346054
rect 416426 345498 416662 345734
rect 416746 345498 416982 345734
rect 414878 330938 415114 331174
rect 414878 330618 415114 330854
rect 412706 306098 412942 306334
rect 413026 306098 413262 306334
rect 412706 305778 412942 306014
rect 413026 305778 413262 306014
rect 412706 270098 412942 270334
rect 413026 270098 413262 270334
rect 412706 269778 412942 270014
rect 413026 269778 413262 270014
rect 412706 234098 412942 234334
rect 413026 234098 413262 234334
rect 412706 233778 412942 234014
rect 413026 233778 413262 234014
rect 412706 198098 412942 198334
rect 413026 198098 413262 198334
rect 412706 197778 412942 198014
rect 413026 197778 413262 198014
rect 412706 162098 412942 162334
rect 413026 162098 413262 162334
rect 412706 161778 412942 162014
rect 413026 161778 413262 162014
rect 420146 710362 420382 710598
rect 420466 710362 420702 710598
rect 420146 710042 420382 710278
rect 420466 710042 420702 710278
rect 420146 673538 420382 673774
rect 420466 673538 420702 673774
rect 420146 673218 420382 673454
rect 420466 673218 420702 673454
rect 420146 637538 420382 637774
rect 420466 637538 420702 637774
rect 420146 637218 420382 637454
rect 420466 637218 420702 637454
rect 420146 601538 420382 601774
rect 420466 601538 420702 601774
rect 420146 601218 420382 601454
rect 420466 601218 420702 601454
rect 420146 565538 420382 565774
rect 420466 565538 420702 565774
rect 420146 565218 420382 565454
rect 420466 565218 420702 565454
rect 420146 529538 420382 529774
rect 420466 529538 420702 529774
rect 420146 529218 420382 529454
rect 420466 529218 420702 529454
rect 420146 493538 420382 493774
rect 420466 493538 420702 493774
rect 420146 493218 420382 493454
rect 420466 493218 420702 493454
rect 420146 457538 420382 457774
rect 420466 457538 420702 457774
rect 420146 457218 420382 457454
rect 420466 457218 420702 457454
rect 423866 711322 424102 711558
rect 424186 711322 424422 711558
rect 423866 711002 424102 711238
rect 424186 711002 424422 711238
rect 423866 677258 424102 677494
rect 424186 677258 424422 677494
rect 423866 676938 424102 677174
rect 424186 676938 424422 677174
rect 423866 641258 424102 641494
rect 424186 641258 424422 641494
rect 423866 640938 424102 641174
rect 424186 640938 424422 641174
rect 423866 605258 424102 605494
rect 424186 605258 424422 605494
rect 423866 604938 424102 605174
rect 424186 604938 424422 605174
rect 423866 569258 424102 569494
rect 424186 569258 424422 569494
rect 423866 568938 424102 569174
rect 424186 568938 424422 569174
rect 423866 533258 424102 533494
rect 424186 533258 424422 533494
rect 423866 532938 424102 533174
rect 424186 532938 424422 533174
rect 423866 497258 424102 497494
rect 424186 497258 424422 497494
rect 423866 496938 424102 497174
rect 424186 496938 424422 497174
rect 423866 461258 424102 461494
rect 424186 461258 424422 461494
rect 423866 460938 424102 461174
rect 424186 460938 424422 461174
rect 433826 704602 434062 704838
rect 434146 704602 434382 704838
rect 433826 704282 434062 704518
rect 434146 704282 434382 704518
rect 433826 687218 434062 687454
rect 434146 687218 434382 687454
rect 433826 686898 434062 687134
rect 434146 686898 434382 687134
rect 433826 651218 434062 651454
rect 434146 651218 434382 651454
rect 433826 650898 434062 651134
rect 434146 650898 434382 651134
rect 433826 615218 434062 615454
rect 434146 615218 434382 615454
rect 433826 614898 434062 615134
rect 434146 614898 434382 615134
rect 433826 579218 434062 579454
rect 434146 579218 434382 579454
rect 433826 578898 434062 579134
rect 434146 578898 434382 579134
rect 433826 543218 434062 543454
rect 434146 543218 434382 543454
rect 433826 542898 434062 543134
rect 434146 542898 434382 543134
rect 433826 507218 434062 507454
rect 434146 507218 434382 507454
rect 433826 506898 434062 507134
rect 434146 506898 434382 507134
rect 433826 471218 434062 471454
rect 434146 471218 434382 471454
rect 433826 470898 434062 471134
rect 434146 470898 434382 471134
rect 437546 705562 437782 705798
rect 437866 705562 438102 705798
rect 437546 705242 437782 705478
rect 437866 705242 438102 705478
rect 437546 690938 437782 691174
rect 437866 690938 438102 691174
rect 437546 690618 437782 690854
rect 437866 690618 438102 690854
rect 437546 654938 437782 655174
rect 437866 654938 438102 655174
rect 437546 654618 437782 654854
rect 437866 654618 438102 654854
rect 437546 618938 437782 619174
rect 437866 618938 438102 619174
rect 437546 618618 437782 618854
rect 437866 618618 438102 618854
rect 437546 582938 437782 583174
rect 437866 582938 438102 583174
rect 437546 582618 437782 582854
rect 437866 582618 438102 582854
rect 437546 546938 437782 547174
rect 437866 546938 438102 547174
rect 437546 546618 437782 546854
rect 437866 546618 438102 546854
rect 437546 510938 437782 511174
rect 437866 510938 438102 511174
rect 437546 510618 437782 510854
rect 437866 510618 438102 510854
rect 437546 474938 437782 475174
rect 437866 474938 438102 475174
rect 437546 474618 437782 474854
rect 437866 474618 438102 474854
rect 441266 706522 441502 706758
rect 441586 706522 441822 706758
rect 441266 706202 441502 706438
rect 441586 706202 441822 706438
rect 444986 707482 445222 707718
rect 445306 707482 445542 707718
rect 444986 707162 445222 707398
rect 445306 707162 445542 707398
rect 441266 694658 441502 694894
rect 441586 694658 441822 694894
rect 441266 694338 441502 694574
rect 441586 694338 441822 694574
rect 441266 658658 441502 658894
rect 441586 658658 441822 658894
rect 441266 658338 441502 658574
rect 441586 658338 441822 658574
rect 441266 622658 441502 622894
rect 441586 622658 441822 622894
rect 441266 622338 441502 622574
rect 441586 622338 441822 622574
rect 441266 586658 441502 586894
rect 441586 586658 441822 586894
rect 441266 586338 441502 586574
rect 441586 586338 441822 586574
rect 441266 550658 441502 550894
rect 441586 550658 441822 550894
rect 441266 550338 441502 550574
rect 441586 550338 441822 550574
rect 441266 514658 441502 514894
rect 441586 514658 441822 514894
rect 441266 514338 441502 514574
rect 441586 514338 441822 514574
rect 441266 478658 441502 478894
rect 441586 478658 441822 478894
rect 441266 478338 441502 478574
rect 441586 478338 441822 478574
rect 426666 438938 426902 439174
rect 426666 438618 426902 438854
rect 432347 438938 432583 439174
rect 432347 438618 432583 438854
rect 438028 438938 438264 439174
rect 438028 438618 438264 438854
rect 443709 438938 443945 439174
rect 443709 438618 443945 438854
rect 423826 435218 424062 435454
rect 423826 434898 424062 435134
rect 429507 435218 429743 435454
rect 429507 434898 429743 435134
rect 435188 435218 435424 435454
rect 435188 434898 435424 435134
rect 440869 435218 441105 435454
rect 440869 434898 441105 435134
rect 420146 421538 420382 421774
rect 420466 421538 420702 421774
rect 420146 421218 420382 421454
rect 420466 421218 420702 421454
rect 420146 385538 420382 385774
rect 420466 385538 420702 385774
rect 420146 385218 420382 385454
rect 420466 385218 420702 385454
rect 420146 349538 420382 349774
rect 420466 349538 420702 349774
rect 420146 349218 420382 349454
rect 420466 349218 420702 349454
rect 418351 327218 418587 327454
rect 418351 326898 418587 327134
rect 416426 309818 416662 310054
rect 416746 309818 416982 310054
rect 416426 309498 416662 309734
rect 416746 309498 416982 309734
rect 416426 273818 416662 274054
rect 416746 273818 416982 274054
rect 416426 273498 416662 273734
rect 416746 273498 416982 273734
rect 416426 237818 416662 238054
rect 416746 237818 416982 238054
rect 416426 237498 416662 237734
rect 416746 237498 416982 237734
rect 416426 201818 416662 202054
rect 416746 201818 416982 202054
rect 416426 201498 416662 201734
rect 416746 201498 416982 201734
rect 416426 165818 416662 166054
rect 416746 165818 416982 166054
rect 416426 165498 416662 165734
rect 416746 165498 416982 165734
rect 423866 389258 424102 389494
rect 424186 389258 424422 389494
rect 423866 388938 424102 389174
rect 424186 388938 424422 389174
rect 423866 353258 424102 353494
rect 424186 353258 424422 353494
rect 423866 352938 424102 353174
rect 424186 352938 424422 353174
rect 420146 313538 420382 313774
rect 420466 313538 420702 313774
rect 420146 313218 420382 313454
rect 420466 313218 420702 313454
rect 420146 277538 420382 277774
rect 420466 277538 420702 277774
rect 420146 277218 420382 277454
rect 420466 277218 420702 277454
rect 420146 241538 420382 241774
rect 420466 241538 420702 241774
rect 420146 241218 420382 241454
rect 420466 241218 420702 241454
rect 420146 205538 420382 205774
rect 420466 205538 420702 205774
rect 420146 205218 420382 205454
rect 420466 205218 420702 205454
rect 420146 169538 420382 169774
rect 420466 169538 420702 169774
rect 420146 169218 420382 169454
rect 420466 169218 420702 169454
rect 421824 330938 422060 331174
rect 421824 330618 422060 330854
rect 433826 399218 434062 399454
rect 434146 399218 434382 399454
rect 433826 398898 434062 399134
rect 434146 398898 434382 399134
rect 433826 363218 434062 363454
rect 434146 363218 434382 363454
rect 433826 362898 434062 363134
rect 434146 362898 434382 363134
rect 425297 327218 425533 327454
rect 425297 326898 425533 327134
rect 423866 317258 424102 317494
rect 424186 317258 424422 317494
rect 423866 316938 424102 317174
rect 424186 316938 424422 317174
rect 423866 281258 424102 281494
rect 424186 281258 424422 281494
rect 423866 280938 424102 281174
rect 424186 280938 424422 281174
rect 423866 245258 424102 245494
rect 424186 245258 424422 245494
rect 423866 244938 424102 245174
rect 424186 244938 424422 245174
rect 423866 209258 424102 209494
rect 424186 209258 424422 209494
rect 423866 208938 424102 209174
rect 424186 208938 424422 209174
rect 423866 173258 424102 173494
rect 424186 173258 424422 173494
rect 423866 172938 424102 173174
rect 424186 172938 424422 173174
rect 428770 330938 429006 331174
rect 428770 330618 429006 330854
rect 433826 327218 434062 327454
rect 434146 327218 434382 327454
rect 433826 326898 434062 327134
rect 434146 326898 434382 327134
rect 433826 291218 434062 291454
rect 434146 291218 434382 291454
rect 433826 290898 434062 291134
rect 434146 290898 434382 291134
rect 433826 255218 434062 255454
rect 434146 255218 434382 255454
rect 433826 254898 434062 255134
rect 434146 254898 434382 255134
rect 433826 219218 434062 219454
rect 434146 219218 434382 219454
rect 433826 218898 434062 219134
rect 434146 218898 434382 219134
rect 433826 183218 434062 183454
rect 434146 183218 434382 183454
rect 433826 182898 434062 183134
rect 434146 182898 434382 183134
rect 437546 402938 437782 403174
rect 437866 402938 438102 403174
rect 437546 402618 437782 402854
rect 437866 402618 438102 402854
rect 437546 366938 437782 367174
rect 437866 366938 438102 367174
rect 437546 366618 437782 366854
rect 437866 366618 438102 366854
rect 437546 330938 437782 331174
rect 437866 330938 438102 331174
rect 437546 330618 437782 330854
rect 437866 330618 438102 330854
rect 437546 294938 437782 295174
rect 437866 294938 438102 295174
rect 437546 294618 437782 294854
rect 437866 294618 438102 294854
rect 437546 258938 437782 259174
rect 437866 258938 438102 259174
rect 437546 258618 437782 258854
rect 437866 258618 438102 258854
rect 437546 222938 437782 223174
rect 437866 222938 438102 223174
rect 437546 222618 437782 222854
rect 437866 222618 438102 222854
rect 437546 186938 437782 187174
rect 437866 186938 438102 187174
rect 437546 186618 437782 186854
rect 437866 186618 438102 186854
rect 441266 406658 441502 406894
rect 441586 406658 441822 406894
rect 441266 406338 441502 406574
rect 441586 406338 441822 406574
rect 441266 370658 441502 370894
rect 441586 370658 441822 370894
rect 441266 370338 441502 370574
rect 441586 370338 441822 370574
rect 441266 334658 441502 334894
rect 441586 334658 441822 334894
rect 441266 334338 441502 334574
rect 441586 334338 441822 334574
rect 444986 698378 445222 698614
rect 445306 698378 445542 698614
rect 444986 698058 445222 698294
rect 445306 698058 445542 698294
rect 448706 708442 448942 708678
rect 449026 708442 449262 708678
rect 448706 708122 448942 708358
rect 449026 708122 449262 708358
rect 444986 662378 445222 662614
rect 445306 662378 445542 662614
rect 444986 662058 445222 662294
rect 445306 662058 445542 662294
rect 444986 626378 445222 626614
rect 445306 626378 445542 626614
rect 444986 626058 445222 626294
rect 445306 626058 445542 626294
rect 444986 590378 445222 590614
rect 445306 590378 445542 590614
rect 444986 590058 445222 590294
rect 445306 590058 445542 590294
rect 444986 554378 445222 554614
rect 445306 554378 445542 554614
rect 444986 554058 445222 554294
rect 445306 554058 445542 554294
rect 444986 518378 445222 518614
rect 445306 518378 445542 518614
rect 444986 518058 445222 518294
rect 445306 518058 445542 518294
rect 444986 482378 445222 482614
rect 445306 482378 445542 482614
rect 444986 482058 445222 482294
rect 445306 482058 445542 482294
rect 444986 446378 445222 446614
rect 445306 446378 445542 446614
rect 444986 446058 445222 446294
rect 445306 446058 445542 446294
rect 444986 410378 445222 410614
rect 445306 410378 445542 410614
rect 444986 410058 445222 410294
rect 445306 410058 445542 410294
rect 444986 374378 445222 374614
rect 445306 374378 445542 374614
rect 444986 374058 445222 374294
rect 445306 374058 445542 374294
rect 444986 338378 445222 338614
rect 445306 338378 445542 338614
rect 444986 338058 445222 338294
rect 445306 338058 445542 338294
rect 441266 298658 441502 298894
rect 441586 298658 441822 298894
rect 441266 298338 441502 298574
rect 441586 298338 441822 298574
rect 441266 262658 441502 262894
rect 441586 262658 441822 262894
rect 441266 262338 441502 262574
rect 441586 262338 441822 262574
rect 441266 226658 441502 226894
rect 441586 226658 441822 226894
rect 441266 226338 441502 226574
rect 441586 226338 441822 226574
rect 441266 190658 441502 190894
rect 441586 190658 441822 190894
rect 441266 190338 441502 190574
rect 441586 190338 441822 190574
rect 448706 666098 448942 666334
rect 449026 666098 449262 666334
rect 448706 665778 448942 666014
rect 449026 665778 449262 666014
rect 448706 630098 448942 630334
rect 449026 630098 449262 630334
rect 448706 629778 448942 630014
rect 449026 629778 449262 630014
rect 448706 594098 448942 594334
rect 449026 594098 449262 594334
rect 448706 593778 448942 594014
rect 449026 593778 449262 594014
rect 448706 558098 448942 558334
rect 449026 558098 449262 558334
rect 448706 557778 448942 558014
rect 449026 557778 449262 558014
rect 448706 522098 448942 522334
rect 449026 522098 449262 522334
rect 448706 521778 448942 522014
rect 449026 521778 449262 522014
rect 452426 709402 452662 709638
rect 452746 709402 452982 709638
rect 452426 709082 452662 709318
rect 452746 709082 452982 709318
rect 452426 669818 452662 670054
rect 452746 669818 452982 670054
rect 452426 669498 452662 669734
rect 452746 669498 452982 669734
rect 452426 633818 452662 634054
rect 452746 633818 452982 634054
rect 452426 633498 452662 633734
rect 452746 633498 452982 633734
rect 452426 597818 452662 598054
rect 452746 597818 452982 598054
rect 452426 597498 452662 597734
rect 452746 597498 452982 597734
rect 452426 561818 452662 562054
rect 452746 561818 452982 562054
rect 452426 561498 452662 561734
rect 452746 561498 452982 561734
rect 452426 525818 452662 526054
rect 452746 525818 452982 526054
rect 452426 525498 452662 525734
rect 452746 525498 452982 525734
rect 456146 710362 456382 710598
rect 456466 710362 456702 710598
rect 456146 710042 456382 710278
rect 456466 710042 456702 710278
rect 456146 673538 456382 673774
rect 456466 673538 456702 673774
rect 456146 673218 456382 673454
rect 456466 673218 456702 673454
rect 459866 711322 460102 711558
rect 460186 711322 460422 711558
rect 459866 711002 460102 711238
rect 460186 711002 460422 711238
rect 459866 677258 460102 677494
rect 460186 677258 460422 677494
rect 459866 676938 460102 677174
rect 460186 676938 460422 677174
rect 456146 637538 456382 637774
rect 456466 637538 456702 637774
rect 456146 637218 456382 637454
rect 456466 637218 456702 637454
rect 456146 601538 456382 601774
rect 456466 601538 456702 601774
rect 456146 601218 456382 601454
rect 456466 601218 456702 601454
rect 456146 565538 456382 565774
rect 456466 565538 456702 565774
rect 456146 565218 456382 565454
rect 456466 565218 456702 565454
rect 456146 529538 456382 529774
rect 456466 529538 456702 529774
rect 456146 529218 456382 529454
rect 456466 529218 456702 529454
rect 448706 486098 448942 486334
rect 449026 486098 449262 486334
rect 448706 485778 448942 486014
rect 449026 485778 449262 486014
rect 448706 450098 448942 450334
rect 449026 450098 449262 450334
rect 448706 449778 448942 450014
rect 449026 449778 449262 450014
rect 448706 414098 448942 414334
rect 449026 414098 449262 414334
rect 448706 413778 448942 414014
rect 449026 413778 449262 414014
rect 448706 378098 448942 378334
rect 449026 378098 449262 378334
rect 448706 377778 448942 378014
rect 449026 377778 449262 378014
rect 448706 342098 448942 342334
rect 449026 342098 449262 342334
rect 448706 341778 448942 342014
rect 449026 341778 449262 342014
rect 444986 302378 445222 302614
rect 445306 302378 445542 302614
rect 444986 302058 445222 302294
rect 445306 302058 445542 302294
rect 444986 266378 445222 266614
rect 445306 266378 445542 266614
rect 444986 266058 445222 266294
rect 445306 266058 445542 266294
rect 444986 230378 445222 230614
rect 445306 230378 445542 230614
rect 444986 230058 445222 230294
rect 445306 230058 445542 230294
rect 444986 194378 445222 194614
rect 445306 194378 445542 194614
rect 444986 194058 445222 194294
rect 445306 194058 445542 194294
rect 453424 510938 453660 511174
rect 453424 510618 453660 510854
rect 455862 510938 456098 511174
rect 455862 510618 456098 510854
rect 458300 510938 458536 511174
rect 458300 510618 458536 510854
rect 452205 507218 452441 507454
rect 452205 506898 452441 507134
rect 454643 507218 454879 507454
rect 454643 506898 454879 507134
rect 457081 507218 457317 507454
rect 457081 506898 457317 507134
rect 452426 489818 452662 490054
rect 452746 489818 452982 490054
rect 452426 489498 452662 489734
rect 452746 489498 452982 489734
rect 452426 453818 452662 454054
rect 452746 453818 452982 454054
rect 452426 453498 452662 453734
rect 452746 453498 452982 453734
rect 452426 417818 452662 418054
rect 452746 417818 452982 418054
rect 452426 417498 452662 417734
rect 452746 417498 452982 417734
rect 452426 381818 452662 382054
rect 452746 381818 452982 382054
rect 452426 381498 452662 381734
rect 452746 381498 452982 381734
rect 456146 493538 456382 493774
rect 456466 493538 456702 493774
rect 456146 493218 456382 493454
rect 456466 493218 456702 493454
rect 456146 457538 456382 457774
rect 456466 457538 456702 457774
rect 456146 457218 456382 457454
rect 456466 457218 456702 457454
rect 469826 704602 470062 704838
rect 470146 704602 470382 704838
rect 469826 704282 470062 704518
rect 470146 704282 470382 704518
rect 469826 687218 470062 687454
rect 470146 687218 470382 687454
rect 469826 686898 470062 687134
rect 470146 686898 470382 687134
rect 473546 705562 473782 705798
rect 473866 705562 474102 705798
rect 473546 705242 473782 705478
rect 473866 705242 474102 705478
rect 473546 690938 473782 691174
rect 473866 690938 474102 691174
rect 473546 690618 473782 690854
rect 473866 690618 474102 690854
rect 477266 706522 477502 706758
rect 477586 706522 477822 706758
rect 477266 706202 477502 706438
rect 477586 706202 477822 706438
rect 477266 694658 477502 694894
rect 477586 694658 477822 694894
rect 477266 694338 477502 694574
rect 477586 694338 477822 694574
rect 480986 707482 481222 707718
rect 481306 707482 481542 707718
rect 480986 707162 481222 707398
rect 481306 707162 481542 707398
rect 480986 698378 481222 698614
rect 481306 698378 481542 698614
rect 480986 698058 481222 698294
rect 481306 698058 481542 698294
rect 488426 709402 488662 709638
rect 488746 709402 488982 709638
rect 488426 709082 488662 709318
rect 488746 709082 488982 709318
rect 488426 669818 488662 670054
rect 488746 669818 488982 670054
rect 488426 669498 488662 669734
rect 488746 669498 488982 669734
rect 492146 710362 492382 710598
rect 492466 710362 492702 710598
rect 492146 710042 492382 710278
rect 492466 710042 492702 710278
rect 492146 673538 492382 673774
rect 492466 673538 492702 673774
rect 492146 673218 492382 673454
rect 492466 673218 492702 673454
rect 495866 711322 496102 711558
rect 496186 711322 496422 711558
rect 495866 711002 496102 711238
rect 496186 711002 496422 711238
rect 495866 677258 496102 677494
rect 496186 677258 496422 677494
rect 495866 676938 496102 677174
rect 496186 676938 496422 677174
rect 505826 704602 506062 704838
rect 506146 704602 506382 704838
rect 505826 704282 506062 704518
rect 506146 704282 506382 704518
rect 505826 687218 506062 687454
rect 506146 687218 506382 687454
rect 505826 686898 506062 687134
rect 506146 686898 506382 687134
rect 509546 705562 509782 705798
rect 509866 705562 510102 705798
rect 509546 705242 509782 705478
rect 509866 705242 510102 705478
rect 509546 690938 509782 691174
rect 509866 690938 510102 691174
rect 509546 690618 509782 690854
rect 509866 690618 510102 690854
rect 513266 706522 513502 706758
rect 513586 706522 513822 706758
rect 513266 706202 513502 706438
rect 513586 706202 513822 706438
rect 513266 694658 513502 694894
rect 513586 694658 513822 694894
rect 513266 694338 513502 694574
rect 513586 694338 513822 694574
rect 516986 707482 517222 707718
rect 517306 707482 517542 707718
rect 516986 707162 517222 707398
rect 517306 707162 517542 707398
rect 516986 698378 517222 698614
rect 517306 698378 517542 698614
rect 516986 698058 517222 698294
rect 517306 698058 517542 698294
rect 520706 708442 520942 708678
rect 521026 708442 521262 708678
rect 520706 708122 520942 708358
rect 521026 708122 521262 708358
rect 520706 666098 520942 666334
rect 521026 666098 521262 666334
rect 520706 665778 520942 666014
rect 521026 665778 521262 666014
rect 479610 654938 479846 655174
rect 479610 654618 479846 654854
rect 510330 654938 510566 655174
rect 510330 654618 510566 654854
rect 464250 651218 464486 651454
rect 464250 650898 464486 651134
rect 494970 651218 495206 651454
rect 494970 650898 495206 651134
rect 520706 630098 520942 630334
rect 521026 630098 521262 630334
rect 520706 629778 520942 630014
rect 521026 629778 521262 630014
rect 479610 618938 479846 619174
rect 479610 618618 479846 618854
rect 510330 618938 510566 619174
rect 510330 618618 510566 618854
rect 464250 615218 464486 615454
rect 464250 614898 464486 615134
rect 494970 615218 495206 615454
rect 494970 614898 495206 615134
rect 459866 569258 460102 569494
rect 460186 569258 460422 569494
rect 459866 568938 460102 569174
rect 460186 568938 460422 569174
rect 459866 533258 460102 533494
rect 460186 533258 460422 533494
rect 459866 532938 460102 533174
rect 460186 532938 460422 533174
rect 469826 579218 470062 579454
rect 470146 579218 470382 579454
rect 469826 578898 470062 579134
rect 470146 578898 470382 579134
rect 469826 543218 470062 543454
rect 470146 543218 470382 543454
rect 469826 542898 470062 543134
rect 470146 542898 470382 543134
rect 460738 510938 460974 511174
rect 460738 510618 460974 510854
rect 459519 507218 459755 507454
rect 459519 506898 459755 507134
rect 469826 507218 470062 507454
rect 470146 507218 470382 507454
rect 469826 506898 470062 507134
rect 470146 506898 470382 507134
rect 459866 497258 460102 497494
rect 460186 497258 460422 497494
rect 459866 496938 460102 497174
rect 460186 496938 460422 497174
rect 459866 461258 460102 461494
rect 460186 461258 460422 461494
rect 459866 460938 460102 461174
rect 460186 460938 460422 461174
rect 456146 421538 456382 421774
rect 456466 421538 456702 421774
rect 456146 421218 456382 421454
rect 456466 421218 456702 421454
rect 456146 385538 456382 385774
rect 456466 385538 456702 385774
rect 456146 385218 456382 385454
rect 456466 385218 456702 385454
rect 454250 363218 454486 363454
rect 454250 362898 454486 363134
rect 452426 345818 452662 346054
rect 452746 345818 452982 346054
rect 452426 345498 452662 345734
rect 452746 345498 452982 345734
rect 448706 306098 448942 306334
rect 449026 306098 449262 306334
rect 448706 305778 448942 306014
rect 449026 305778 449262 306014
rect 448706 270098 448942 270334
rect 449026 270098 449262 270334
rect 448706 269778 448942 270014
rect 449026 269778 449262 270014
rect 448706 234098 448942 234334
rect 449026 234098 449262 234334
rect 448706 233778 448942 234014
rect 449026 233778 449262 234014
rect 448706 198098 448942 198334
rect 449026 198098 449262 198334
rect 448706 197778 448942 198014
rect 449026 197778 449262 198014
rect 448706 162098 448942 162334
rect 449026 162098 449262 162334
rect 448706 161778 448942 162014
rect 449026 161778 449262 162014
rect 429610 150938 429846 151174
rect 429610 150618 429846 150854
rect 414250 147218 414486 147454
rect 414250 146898 414486 147134
rect 444970 147218 445206 147454
rect 444970 146898 445206 147134
rect 412706 126098 412942 126334
rect 413026 126098 413262 126334
rect 412706 125778 412942 126014
rect 413026 125778 413262 126014
rect 412706 90098 412942 90334
rect 413026 90098 413262 90334
rect 412706 89778 412942 90014
rect 413026 89778 413262 90014
rect 412706 54098 412942 54334
rect 413026 54098 413262 54334
rect 412706 53778 412942 54014
rect 413026 53778 413262 54014
rect 412706 18098 412942 18334
rect 413026 18098 413262 18334
rect 412706 17778 412942 18014
rect 413026 17778 413262 18014
rect 412706 -4422 412942 -4186
rect 413026 -4422 413262 -4186
rect 412706 -4742 412942 -4506
rect 413026 -4742 413262 -4506
rect 416426 93818 416662 94054
rect 416746 93818 416982 94054
rect 416426 93498 416662 93734
rect 416746 93498 416982 93734
rect 416426 57818 416662 58054
rect 416746 57818 416982 58054
rect 416426 57498 416662 57734
rect 416746 57498 416982 57734
rect 416426 21818 416662 22054
rect 416746 21818 416982 22054
rect 416426 21498 416662 21734
rect 416746 21498 416982 21734
rect 416426 -5382 416662 -5146
rect 416746 -5382 416982 -5146
rect 416426 -5702 416662 -5466
rect 416746 -5702 416982 -5466
rect 420146 97538 420382 97774
rect 420466 97538 420702 97774
rect 420146 97218 420382 97454
rect 420466 97218 420702 97454
rect 420146 61538 420382 61774
rect 420466 61538 420702 61774
rect 420146 61218 420382 61454
rect 420466 61218 420702 61454
rect 420146 25538 420382 25774
rect 420466 25538 420702 25774
rect 420146 25218 420382 25454
rect 420466 25218 420702 25454
rect 420146 -6342 420382 -6106
rect 420466 -6342 420702 -6106
rect 420146 -6662 420382 -6426
rect 420466 -6662 420702 -6426
rect 423866 101258 424102 101494
rect 424186 101258 424422 101494
rect 423866 100938 424102 101174
rect 424186 100938 424422 101174
rect 423866 65258 424102 65494
rect 424186 65258 424422 65494
rect 423866 64938 424102 65174
rect 424186 64938 424422 65174
rect 423866 29258 424102 29494
rect 424186 29258 424422 29494
rect 423866 28938 424102 29174
rect 424186 28938 424422 29174
rect 423866 -7302 424102 -7066
rect 424186 -7302 424422 -7066
rect 423866 -7622 424102 -7386
rect 424186 -7622 424422 -7386
rect 433826 111218 434062 111454
rect 434146 111218 434382 111454
rect 433826 110898 434062 111134
rect 434146 110898 434382 111134
rect 433826 75218 434062 75454
rect 434146 75218 434382 75454
rect 433826 74898 434062 75134
rect 434146 74898 434382 75134
rect 433826 39218 434062 39454
rect 434146 39218 434382 39454
rect 433826 38898 434062 39134
rect 434146 38898 434382 39134
rect 433826 3218 434062 3454
rect 434146 3218 434382 3454
rect 433826 2898 434062 3134
rect 434146 2898 434382 3134
rect 433826 -582 434062 -346
rect 434146 -582 434382 -346
rect 433826 -902 434062 -666
rect 434146 -902 434382 -666
rect 437546 114938 437782 115174
rect 437866 114938 438102 115174
rect 437546 114618 437782 114854
rect 437866 114618 438102 114854
rect 437546 78938 437782 79174
rect 437866 78938 438102 79174
rect 437546 78618 437782 78854
rect 437866 78618 438102 78854
rect 437546 42938 437782 43174
rect 437866 42938 438102 43174
rect 437546 42618 437782 42854
rect 437866 42618 438102 42854
rect 437546 6938 437782 7174
rect 437866 6938 438102 7174
rect 437546 6618 437782 6854
rect 437866 6618 438102 6854
rect 437546 -1542 437782 -1306
rect 437866 -1542 438102 -1306
rect 437546 -1862 437782 -1626
rect 437866 -1862 438102 -1626
rect 448706 126098 448942 126334
rect 449026 126098 449262 126334
rect 448706 125778 448942 126014
rect 449026 125778 449262 126014
rect 441266 118658 441502 118894
rect 441586 118658 441822 118894
rect 441266 118338 441502 118574
rect 441586 118338 441822 118574
rect 441266 82658 441502 82894
rect 441586 82658 441822 82894
rect 441266 82338 441502 82574
rect 441586 82338 441822 82574
rect 441266 46658 441502 46894
rect 441586 46658 441822 46894
rect 441266 46338 441502 46574
rect 441586 46338 441822 46574
rect 441266 10658 441502 10894
rect 441586 10658 441822 10894
rect 441266 10338 441502 10574
rect 441586 10338 441822 10574
rect 441266 -2502 441502 -2266
rect 441586 -2502 441822 -2266
rect 441266 -2822 441502 -2586
rect 441586 -2822 441822 -2586
rect 444986 86378 445222 86614
rect 445306 86378 445542 86614
rect 444986 86058 445222 86294
rect 445306 86058 445542 86294
rect 444986 50378 445222 50614
rect 445306 50378 445542 50614
rect 444986 50058 445222 50294
rect 445306 50058 445542 50294
rect 444986 14378 445222 14614
rect 445306 14378 445542 14614
rect 444986 14058 445222 14294
rect 445306 14058 445542 14294
rect 444986 -3462 445222 -3226
rect 445306 -3462 445542 -3226
rect 444986 -3782 445222 -3546
rect 445306 -3782 445542 -3546
rect 448706 90098 448942 90334
rect 449026 90098 449262 90334
rect 448706 89778 448942 90014
rect 449026 89778 449262 90014
rect 448706 54098 448942 54334
rect 449026 54098 449262 54334
rect 448706 53778 448942 54014
rect 449026 53778 449262 54014
rect 448706 18098 448942 18334
rect 449026 18098 449262 18334
rect 448706 17778 448942 18014
rect 449026 17778 449262 18014
rect 448706 -4422 448942 -4186
rect 449026 -4422 449262 -4186
rect 448706 -4742 448942 -4506
rect 449026 -4742 449262 -4506
rect 456146 349538 456382 349774
rect 456466 349538 456702 349774
rect 456146 349218 456382 349454
rect 456466 349218 456702 349454
rect 454250 327218 454486 327454
rect 454250 326898 454486 327134
rect 452426 309818 452662 310054
rect 452746 309818 452982 310054
rect 452426 309498 452662 309734
rect 452746 309498 452982 309734
rect 452426 273818 452662 274054
rect 452746 273818 452982 274054
rect 452426 273498 452662 273734
rect 452746 273498 452982 273734
rect 452426 237818 452662 238054
rect 452746 237818 452982 238054
rect 452426 237498 452662 237734
rect 452746 237498 452982 237734
rect 452426 201818 452662 202054
rect 452746 201818 452982 202054
rect 452426 201498 452662 201734
rect 452746 201498 452982 201734
rect 452426 165818 452662 166054
rect 452746 165818 452982 166054
rect 452426 165498 452662 165734
rect 452746 165498 452982 165734
rect 452426 129818 452662 130054
rect 452746 129818 452982 130054
rect 452426 129498 452662 129734
rect 452746 129498 452982 129734
rect 452426 93818 452662 94054
rect 452746 93818 452982 94054
rect 452426 93498 452662 93734
rect 452746 93498 452982 93734
rect 452426 57818 452662 58054
rect 452746 57818 452982 58054
rect 452426 57498 452662 57734
rect 452746 57498 452982 57734
rect 452426 21818 452662 22054
rect 452746 21818 452982 22054
rect 452426 21498 452662 21734
rect 452746 21498 452982 21734
rect 452426 -5382 452662 -5146
rect 452746 -5382 452982 -5146
rect 452426 -5702 452662 -5466
rect 452746 -5702 452982 -5466
rect 459866 425258 460102 425494
rect 460186 425258 460422 425494
rect 459866 424938 460102 425174
rect 460186 424938 460422 425174
rect 459866 389258 460102 389494
rect 460186 389258 460422 389494
rect 459866 388938 460102 389174
rect 460186 388938 460422 389174
rect 469826 471218 470062 471454
rect 470146 471218 470382 471454
rect 469826 470898 470062 471134
rect 470146 470898 470382 471134
rect 469826 435218 470062 435454
rect 470146 435218 470382 435454
rect 469826 434898 470062 435134
rect 470146 434898 470382 435134
rect 469826 399218 470062 399454
rect 470146 399218 470382 399454
rect 469826 398898 470062 399134
rect 470146 398898 470382 399134
rect 473546 582938 473782 583174
rect 473866 582938 474102 583174
rect 473546 582618 473782 582854
rect 473866 582618 474102 582854
rect 473546 546938 473782 547174
rect 473866 546938 474102 547174
rect 473546 546618 473782 546854
rect 473866 546618 474102 546854
rect 477266 586658 477502 586894
rect 477586 586658 477822 586894
rect 477266 586338 477502 586574
rect 477586 586338 477822 586574
rect 477266 550658 477502 550894
rect 477586 550658 477822 550894
rect 477266 550338 477502 550574
rect 477586 550338 477822 550574
rect 473546 510938 473782 511174
rect 473866 510938 474102 511174
rect 473546 510618 473782 510854
rect 473866 510618 474102 510854
rect 473546 474938 473782 475174
rect 473866 474938 474102 475174
rect 473546 474618 473782 474854
rect 473866 474618 474102 474854
rect 473458 435218 473694 435454
rect 473458 434898 473694 435134
rect 477266 514658 477502 514894
rect 477586 514658 477822 514894
rect 477266 514338 477502 514574
rect 477586 514338 477822 514574
rect 477266 478658 477502 478894
rect 477586 478658 477822 478894
rect 477266 478338 477502 478574
rect 477586 478338 477822 478574
rect 477266 442658 477502 442894
rect 477586 442658 477822 442894
rect 477266 442338 477502 442574
rect 477586 442338 477822 442574
rect 475930 438938 476166 439174
rect 475930 438618 476166 438854
rect 478403 435218 478639 435454
rect 478403 434898 478639 435134
rect 477266 406658 477502 406894
rect 477586 406658 477822 406894
rect 477266 406338 477502 406574
rect 477586 406338 477822 406574
rect 480986 590378 481222 590614
rect 481306 590378 481542 590614
rect 480986 590058 481222 590294
rect 481306 590058 481542 590294
rect 480986 554378 481222 554614
rect 481306 554378 481542 554614
rect 480986 554058 481222 554294
rect 481306 554058 481542 554294
rect 480986 518378 481222 518614
rect 481306 518378 481542 518614
rect 480986 518058 481222 518294
rect 481306 518058 481542 518294
rect 484706 594098 484942 594334
rect 485026 594098 485262 594334
rect 484706 593778 484942 594014
rect 485026 593778 485262 594014
rect 484706 558098 484942 558334
rect 485026 558098 485262 558334
rect 484706 557778 484942 558014
rect 485026 557778 485262 558014
rect 484706 522098 484942 522334
rect 485026 522098 485262 522334
rect 484706 521778 484942 522014
rect 485026 521778 485262 522014
rect 488426 597818 488662 598054
rect 488746 597818 488982 598054
rect 488426 597498 488662 597734
rect 488746 597498 488982 597734
rect 488426 561818 488662 562054
rect 488746 561818 488982 562054
rect 488426 561498 488662 561734
rect 488746 561498 488982 561734
rect 488426 525818 488662 526054
rect 488746 525818 488982 526054
rect 488426 525498 488662 525734
rect 488746 525498 488982 525734
rect 492146 565538 492382 565774
rect 492466 565538 492702 565774
rect 492146 565218 492382 565454
rect 492466 565218 492702 565454
rect 492146 529538 492382 529774
rect 492466 529538 492702 529774
rect 492146 529218 492382 529454
rect 492466 529218 492702 529454
rect 482205 507218 482441 507454
rect 482205 506898 482441 507134
rect 480986 482378 481222 482614
rect 481306 482378 481542 482614
rect 480986 482058 481222 482294
rect 481306 482058 481542 482294
rect 483424 510938 483660 511174
rect 483424 510618 483660 510854
rect 485862 510938 486098 511174
rect 485862 510618 486098 510854
rect 488300 510938 488536 511174
rect 488300 510618 488536 510854
rect 490738 510938 490974 511174
rect 490738 510618 490974 510854
rect 484643 507218 484879 507454
rect 484643 506898 484879 507134
rect 487081 507218 487317 507454
rect 487081 506898 487317 507134
rect 489519 507218 489755 507454
rect 489519 506898 489755 507134
rect 484706 486098 484942 486334
rect 485026 486098 485262 486334
rect 484706 485778 484942 486014
rect 485026 485778 485262 486014
rect 488426 489818 488662 490054
rect 488746 489818 488982 490054
rect 488426 489498 488662 489734
rect 488746 489498 488982 489734
rect 488426 453771 488662 454007
rect 488746 453771 488982 454007
rect 484706 450098 484942 450334
rect 485026 450098 485262 450334
rect 484706 449778 484942 450014
rect 485026 449778 485262 450014
rect 480875 438938 481111 439174
rect 480875 438618 481111 438854
rect 483348 435218 483584 435454
rect 483348 434898 483584 435134
rect 485820 438938 486056 439174
rect 485820 438618 486056 438854
rect 488293 435218 488529 435454
rect 488293 434898 488529 435134
rect 484706 414098 484942 414334
rect 485026 414098 485262 414334
rect 484706 413778 484942 414014
rect 485026 413778 485262 414014
rect 492146 493538 492382 493774
rect 492466 493538 492702 493774
rect 492146 493218 492382 493454
rect 492466 493218 492702 493454
rect 492146 457538 492382 457774
rect 492466 457538 492702 457774
rect 492146 457218 492382 457454
rect 492466 457218 492702 457454
rect 490765 438938 491001 439174
rect 490765 438618 491001 438854
rect 492146 421538 492382 421774
rect 492466 421538 492702 421774
rect 492146 421218 492382 421454
rect 492466 421218 492702 421454
rect 495866 569258 496102 569494
rect 496186 569258 496422 569494
rect 495866 568938 496102 569174
rect 496186 568938 496422 569174
rect 495866 533258 496102 533494
rect 496186 533258 496422 533494
rect 495866 532938 496102 533174
rect 496186 532938 496422 533174
rect 495866 497258 496102 497494
rect 496186 497258 496422 497494
rect 495866 496938 496102 497174
rect 496186 496938 496422 497174
rect 495866 461258 496102 461494
rect 496186 461258 496422 461494
rect 495866 460938 496102 461174
rect 496186 460938 496422 461174
rect 495866 425258 496102 425494
rect 496186 425258 496422 425494
rect 495866 424938 496102 425174
rect 496186 424938 496422 425174
rect 495866 389258 496102 389494
rect 496186 389258 496422 389494
rect 495866 388938 496102 389174
rect 496186 388938 496422 389174
rect 469610 366938 469846 367174
rect 469610 366618 469846 366854
rect 484970 363218 485206 363454
rect 484970 362898 485206 363134
rect 459866 353258 460102 353494
rect 460186 353258 460422 353494
rect 459866 352938 460102 353174
rect 460186 352938 460422 353174
rect 456146 313538 456382 313774
rect 456466 313538 456702 313774
rect 456146 313218 456382 313454
rect 456466 313218 456702 313454
rect 456146 277538 456382 277774
rect 456466 277538 456702 277774
rect 456146 277218 456382 277454
rect 456466 277218 456702 277454
rect 456146 241538 456382 241774
rect 456466 241538 456702 241774
rect 456146 241218 456382 241454
rect 456466 241218 456702 241454
rect 456146 205538 456382 205774
rect 456466 205538 456702 205774
rect 456146 205218 456382 205454
rect 456466 205218 456702 205454
rect 456146 169538 456382 169774
rect 456466 169538 456702 169774
rect 456146 169218 456382 169454
rect 456466 169218 456702 169454
rect 456146 133538 456382 133774
rect 456466 133538 456702 133774
rect 456146 133218 456382 133454
rect 456466 133218 456702 133454
rect 456146 97538 456382 97774
rect 456466 97538 456702 97774
rect 456146 97218 456382 97454
rect 456466 97218 456702 97454
rect 456146 61538 456382 61774
rect 456466 61538 456702 61774
rect 456146 61218 456382 61454
rect 456466 61218 456702 61454
rect 456146 25538 456382 25774
rect 456466 25538 456702 25774
rect 456146 25218 456382 25454
rect 456466 25218 456702 25454
rect 505826 579218 506062 579454
rect 506146 579218 506382 579454
rect 505826 578898 506062 579134
rect 506146 578898 506382 579134
rect 505826 543218 506062 543454
rect 506146 543218 506382 543454
rect 505826 542898 506062 543134
rect 506146 542898 506382 543134
rect 505826 507218 506062 507454
rect 506146 507218 506382 507454
rect 505826 506898 506062 507134
rect 506146 506898 506382 507134
rect 505826 471218 506062 471454
rect 506146 471218 506382 471454
rect 505826 470898 506062 471134
rect 506146 470898 506382 471134
rect 505826 435218 506062 435454
rect 506146 435218 506382 435454
rect 505826 434898 506062 435134
rect 506146 434898 506382 435134
rect 505826 399218 506062 399454
rect 506146 399218 506382 399454
rect 505826 398898 506062 399134
rect 506146 398898 506382 399134
rect 500330 366938 500566 367174
rect 500330 366618 500566 366854
rect 495866 353258 496102 353494
rect 496186 353258 496422 353494
rect 495866 352938 496102 353174
rect 496186 352938 496422 353174
rect 469610 330938 469846 331174
rect 469610 330618 469846 330854
rect 484970 327218 485206 327454
rect 484970 326898 485206 327134
rect 459866 317258 460102 317494
rect 460186 317258 460422 317494
rect 459866 316938 460102 317174
rect 460186 316938 460422 317174
rect 459866 281258 460102 281494
rect 460186 281258 460422 281494
rect 459866 280938 460102 281174
rect 460186 280938 460422 281174
rect 477266 298658 477502 298894
rect 477586 298658 477822 298894
rect 477266 298338 477502 298574
rect 477586 298338 477822 298574
rect 477266 262658 477502 262894
rect 477586 262658 477822 262894
rect 477266 262338 477502 262574
rect 477586 262338 477822 262574
rect 480986 302378 481222 302614
rect 481306 302378 481542 302614
rect 480986 302058 481222 302294
rect 481306 302058 481542 302294
rect 480986 266378 481222 266614
rect 481306 266378 481542 266614
rect 480986 266058 481222 266294
rect 481306 266058 481542 266294
rect 484706 306098 484942 306334
rect 485026 306098 485262 306334
rect 484706 305778 484942 306014
rect 485026 305778 485262 306014
rect 484706 270098 484942 270334
rect 485026 270098 485262 270334
rect 484706 269778 484942 270014
rect 485026 269778 485262 270014
rect 488426 309818 488662 310054
rect 488746 309818 488982 310054
rect 488426 309498 488662 309734
rect 488746 309498 488982 309734
rect 488426 273818 488662 274054
rect 488746 273818 488982 274054
rect 488426 273498 488662 273734
rect 488746 273498 488982 273734
rect 492146 313538 492382 313774
rect 492466 313538 492702 313774
rect 492146 313218 492382 313454
rect 492466 313218 492702 313454
rect 492146 277538 492382 277774
rect 492466 277538 492702 277774
rect 492146 277218 492382 277454
rect 492466 277218 492702 277454
rect 505826 363218 506062 363454
rect 506146 363218 506382 363454
rect 505826 362898 506062 363134
rect 506146 362898 506382 363134
rect 500330 330938 500566 331174
rect 500330 330618 500566 330854
rect 495866 317258 496102 317494
rect 496186 317258 496422 317494
rect 495866 316938 496102 317174
rect 496186 316938 496422 317174
rect 495866 281258 496102 281494
rect 496186 281258 496422 281494
rect 495866 280938 496102 281174
rect 496186 280938 496422 281174
rect 505826 327218 506062 327454
rect 506146 327218 506382 327454
rect 505826 326898 506062 327134
rect 506146 326898 506382 327134
rect 505826 291218 506062 291454
rect 506146 291218 506382 291454
rect 505826 290898 506062 291134
rect 506146 290898 506382 291134
rect 509546 582938 509782 583174
rect 509866 582938 510102 583174
rect 509546 582618 509782 582854
rect 509866 582618 510102 582854
rect 509546 546938 509782 547174
rect 509866 546938 510102 547174
rect 509546 546618 509782 546854
rect 509866 546618 510102 546854
rect 509546 510938 509782 511174
rect 509866 510938 510102 511174
rect 509546 510618 509782 510854
rect 509866 510618 510102 510854
rect 509546 474938 509782 475174
rect 509866 474938 510102 475174
rect 509546 474618 509782 474854
rect 509866 474618 510102 474854
rect 509546 438938 509782 439174
rect 509866 438938 510102 439174
rect 509546 438618 509782 438854
rect 509866 438618 510102 438854
rect 509546 402938 509782 403174
rect 509866 402938 510102 403174
rect 509546 402618 509782 402854
rect 509866 402618 510102 402854
rect 509546 366938 509782 367174
rect 509866 366938 510102 367174
rect 509546 366618 509782 366854
rect 509866 366618 510102 366854
rect 513266 586658 513502 586894
rect 513586 586658 513822 586894
rect 513266 586338 513502 586574
rect 513586 586338 513822 586574
rect 513266 550658 513502 550894
rect 513586 550658 513822 550894
rect 513266 550338 513502 550574
rect 513586 550338 513822 550574
rect 513266 514658 513502 514894
rect 513586 514658 513822 514894
rect 513266 514338 513502 514574
rect 513586 514338 513822 514574
rect 513266 478658 513502 478894
rect 513586 478658 513822 478894
rect 513266 478338 513502 478574
rect 513586 478338 513822 478574
rect 513266 442658 513502 442894
rect 513586 442658 513822 442894
rect 513266 442338 513502 442574
rect 513586 442338 513822 442574
rect 513266 406658 513502 406894
rect 513586 406658 513822 406894
rect 513266 406338 513502 406574
rect 513586 406338 513822 406574
rect 513266 370658 513502 370894
rect 513586 370658 513822 370894
rect 513266 370338 513502 370574
rect 513586 370338 513822 370574
rect 509546 330938 509782 331174
rect 509866 330938 510102 331174
rect 509546 330618 509782 330854
rect 509866 330618 510102 330854
rect 513266 334658 513502 334894
rect 513586 334658 513822 334894
rect 513266 334338 513502 334574
rect 513586 334338 513822 334574
rect 509546 294938 509782 295174
rect 509866 294938 510102 295174
rect 509546 294618 509782 294854
rect 509866 294618 510102 294854
rect 516986 590378 517222 590614
rect 517306 590378 517542 590614
rect 516986 590058 517222 590294
rect 517306 590058 517542 590294
rect 516986 554378 517222 554614
rect 517306 554378 517542 554614
rect 516986 554058 517222 554294
rect 517306 554058 517542 554294
rect 516986 518378 517222 518614
rect 517306 518378 517542 518614
rect 516986 518058 517222 518294
rect 517306 518058 517542 518294
rect 516986 482378 517222 482614
rect 517306 482378 517542 482614
rect 516986 482058 517222 482294
rect 517306 482058 517542 482294
rect 516986 446378 517222 446614
rect 517306 446378 517542 446614
rect 516986 446058 517222 446294
rect 517306 446058 517542 446294
rect 516986 410378 517222 410614
rect 517306 410378 517542 410614
rect 516986 410058 517222 410294
rect 517306 410058 517542 410294
rect 516986 374378 517222 374614
rect 517306 374378 517542 374614
rect 516986 374058 517222 374294
rect 517306 374058 517542 374294
rect 520706 594098 520942 594334
rect 521026 594098 521262 594334
rect 520706 593778 520942 594014
rect 521026 593778 521262 594014
rect 520706 558098 520942 558334
rect 521026 558098 521262 558334
rect 520706 557778 520942 558014
rect 521026 557778 521262 558014
rect 520706 522098 520942 522334
rect 521026 522098 521262 522334
rect 520706 521778 520942 522014
rect 521026 521778 521262 522014
rect 520706 486098 520942 486334
rect 521026 486098 521262 486334
rect 520706 485778 520942 486014
rect 521026 485778 521262 486014
rect 520706 450098 520942 450334
rect 521026 450098 521262 450334
rect 520706 449778 520942 450014
rect 521026 449778 521262 450014
rect 520706 414098 520942 414334
rect 521026 414098 521262 414334
rect 520706 413778 520942 414014
rect 521026 413778 521262 414014
rect 520706 378098 520942 378334
rect 521026 378098 521262 378334
rect 520706 377778 520942 378014
rect 521026 377778 521262 378014
rect 520706 342098 520942 342334
rect 521026 342098 521262 342334
rect 520706 341778 520942 342014
rect 521026 341778 521262 342014
rect 516986 338378 517222 338614
rect 517306 338378 517542 338614
rect 516986 338058 517222 338294
rect 517306 338058 517542 338294
rect 516986 302378 517222 302614
rect 517306 302378 517542 302614
rect 516986 302058 517222 302294
rect 517306 302058 517542 302294
rect 513266 298658 513502 298894
rect 513586 298658 513822 298894
rect 513266 298338 513502 298574
rect 513586 298338 513822 298574
rect 513266 262658 513502 262894
rect 513586 262658 513822 262894
rect 513266 262338 513502 262574
rect 513586 262338 513822 262574
rect 520706 306098 520942 306334
rect 521026 306098 521262 306334
rect 520706 305778 520942 306014
rect 521026 305778 521262 306014
rect 516986 266378 517222 266614
rect 517306 266378 517542 266614
rect 516986 266058 517222 266294
rect 517306 266058 517542 266294
rect 520706 270098 520942 270334
rect 521026 270098 521262 270334
rect 520706 269778 520942 270014
rect 521026 269778 521262 270014
rect 524426 709402 524662 709638
rect 524746 709402 524982 709638
rect 524426 709082 524662 709318
rect 524746 709082 524982 709318
rect 528146 710362 528382 710598
rect 528466 710362 528702 710598
rect 528146 710042 528382 710278
rect 528466 710042 528702 710278
rect 524426 669818 524662 670054
rect 524746 669818 524982 670054
rect 524426 669498 524662 669734
rect 524746 669498 524982 669734
rect 525690 651218 525926 651454
rect 525690 650898 525926 651134
rect 524426 633818 524662 634054
rect 524746 633818 524982 634054
rect 524426 633498 524662 633734
rect 524746 633498 524982 633734
rect 525690 615218 525926 615454
rect 525690 614898 525926 615134
rect 524426 597818 524662 598054
rect 524746 597818 524982 598054
rect 524426 597498 524662 597734
rect 524746 597498 524982 597734
rect 524426 561818 524662 562054
rect 524746 561818 524982 562054
rect 524426 561498 524662 561734
rect 524746 561498 524982 561734
rect 524426 525818 524662 526054
rect 524746 525818 524982 526054
rect 524426 525498 524662 525734
rect 524746 525498 524982 525734
rect 531866 711322 532102 711558
rect 532186 711322 532422 711558
rect 531866 711002 532102 711238
rect 532186 711002 532422 711238
rect 528146 673538 528382 673774
rect 528466 673538 528702 673774
rect 528146 673218 528382 673454
rect 528466 673218 528702 673454
rect 528146 637538 528382 637774
rect 528466 637538 528702 637774
rect 528146 637218 528382 637454
rect 528466 637218 528702 637454
rect 528146 601538 528382 601774
rect 528466 601538 528702 601774
rect 528146 601218 528382 601454
rect 528466 601218 528702 601454
rect 528146 565538 528382 565774
rect 528466 565538 528702 565774
rect 528146 565218 528382 565454
rect 528466 565218 528702 565454
rect 528146 529538 528382 529774
rect 528466 529538 528702 529774
rect 528146 529218 528382 529454
rect 528466 529218 528702 529454
rect 524426 489818 524662 490054
rect 524746 489818 524982 490054
rect 524426 489498 524662 489734
rect 524746 489498 524982 489734
rect 524426 453818 524662 454054
rect 524746 453818 524982 454054
rect 524426 453498 524662 453734
rect 524746 453498 524982 453734
rect 528146 493538 528382 493774
rect 528466 493538 528702 493774
rect 528146 493218 528382 493454
rect 528466 493218 528702 493454
rect 528146 457538 528382 457774
rect 528466 457538 528702 457774
rect 528146 457218 528382 457454
rect 528466 457218 528702 457454
rect 525206 435218 525442 435454
rect 525206 434898 525442 435134
rect 524426 417818 524662 418054
rect 524746 417818 524982 418054
rect 524426 417498 524662 417734
rect 524746 417498 524982 417734
rect 524426 381818 524662 382054
rect 524746 381818 524982 382054
rect 524426 381498 524662 381734
rect 524746 381498 524982 381734
rect 524426 345818 524662 346054
rect 524746 345818 524982 346054
rect 524426 345498 524662 345734
rect 524746 345498 524982 345734
rect 524426 309818 524662 310054
rect 524746 309818 524982 310054
rect 524426 309498 524662 309734
rect 524746 309498 524982 309734
rect 524426 273818 524662 274054
rect 524746 273818 524982 274054
rect 524426 273498 524662 273734
rect 524746 273498 524982 273734
rect 529426 438938 529662 439174
rect 529426 438618 529662 438854
rect 528146 421538 528382 421774
rect 528466 421538 528702 421774
rect 528146 421218 528382 421454
rect 528466 421218 528702 421454
rect 528146 385538 528382 385774
rect 528466 385538 528702 385774
rect 528146 385218 528382 385454
rect 528466 385218 528702 385454
rect 528146 349538 528382 349774
rect 528466 349538 528702 349774
rect 528146 349218 528382 349454
rect 528466 349218 528702 349454
rect 531866 677258 532102 677494
rect 532186 677258 532422 677494
rect 531866 676938 532102 677174
rect 532186 676938 532422 677174
rect 531866 641258 532102 641494
rect 532186 641258 532422 641494
rect 531866 640938 532102 641174
rect 532186 640938 532422 641174
rect 531866 605258 532102 605494
rect 532186 605258 532422 605494
rect 531866 604938 532102 605174
rect 532186 604938 532422 605174
rect 531866 569258 532102 569494
rect 532186 569258 532422 569494
rect 531866 568938 532102 569174
rect 532186 568938 532422 569174
rect 531866 533258 532102 533494
rect 532186 533258 532422 533494
rect 531866 532938 532102 533174
rect 532186 532938 532422 533174
rect 531866 497258 532102 497494
rect 532186 497258 532422 497494
rect 531866 496938 532102 497174
rect 532186 496938 532422 497174
rect 531866 461258 532102 461494
rect 532186 461258 532422 461494
rect 531866 460938 532102 461174
rect 532186 460938 532422 461174
rect 541826 704602 542062 704838
rect 542146 704602 542382 704838
rect 541826 704282 542062 704518
rect 542146 704282 542382 704518
rect 541826 687218 542062 687454
rect 542146 687218 542382 687454
rect 541826 686898 542062 687134
rect 542146 686898 542382 687134
rect 541826 651218 542062 651454
rect 542146 651218 542382 651454
rect 541826 650898 542062 651134
rect 542146 650898 542382 651134
rect 541826 615218 542062 615454
rect 542146 615218 542382 615454
rect 541826 614898 542062 615134
rect 542146 614898 542382 615134
rect 541826 579218 542062 579454
rect 542146 579218 542382 579454
rect 541826 578898 542062 579134
rect 542146 578898 542382 579134
rect 541826 543218 542062 543454
rect 542146 543218 542382 543454
rect 541826 542898 542062 543134
rect 542146 542898 542382 543134
rect 541826 507218 542062 507454
rect 542146 507218 542382 507454
rect 541826 506898 542062 507134
rect 542146 506898 542382 507134
rect 541826 471218 542062 471454
rect 542146 471218 542382 471454
rect 541826 470898 542062 471134
rect 542146 470898 542382 471134
rect 545546 705562 545782 705798
rect 545866 705562 546102 705798
rect 545546 705242 545782 705478
rect 545866 705242 546102 705478
rect 545546 690938 545782 691174
rect 545866 690938 546102 691174
rect 545546 690618 545782 690854
rect 545866 690618 546102 690854
rect 545546 654938 545782 655174
rect 545866 654938 546102 655174
rect 545546 654618 545782 654854
rect 545866 654618 546102 654854
rect 545546 618938 545782 619174
rect 545866 618938 546102 619174
rect 545546 618618 545782 618854
rect 545866 618618 546102 618854
rect 545546 582938 545782 583174
rect 545866 582938 546102 583174
rect 545546 582618 545782 582854
rect 545866 582618 546102 582854
rect 545546 546938 545782 547174
rect 545866 546938 546102 547174
rect 545546 546618 545782 546854
rect 545866 546618 546102 546854
rect 545546 510938 545782 511174
rect 545866 510938 546102 511174
rect 545546 510618 545782 510854
rect 545866 510618 546102 510854
rect 545546 474938 545782 475174
rect 545866 474938 546102 475174
rect 545546 474618 545782 474854
rect 545866 474618 546102 474854
rect 537867 438938 538103 439174
rect 537867 438618 538103 438854
rect 549266 706522 549502 706758
rect 549586 706522 549822 706758
rect 549266 706202 549502 706438
rect 549586 706202 549822 706438
rect 549266 694658 549502 694894
rect 549586 694658 549822 694894
rect 549266 694338 549502 694574
rect 549586 694338 549822 694574
rect 549266 658658 549502 658894
rect 549586 658658 549822 658894
rect 549266 658338 549502 658574
rect 549586 658338 549822 658574
rect 549266 622658 549502 622894
rect 549586 622658 549822 622894
rect 549266 622338 549502 622574
rect 549586 622338 549822 622574
rect 549266 586658 549502 586894
rect 549586 586658 549822 586894
rect 549266 586338 549502 586574
rect 549586 586338 549822 586574
rect 549266 550658 549502 550894
rect 549586 550658 549822 550894
rect 549266 550338 549502 550574
rect 549586 550338 549822 550574
rect 549266 514658 549502 514894
rect 549586 514658 549822 514894
rect 549266 514338 549502 514574
rect 549586 514338 549822 514574
rect 549266 478658 549502 478894
rect 549586 478658 549822 478894
rect 549266 478338 549502 478574
rect 549586 478338 549822 478574
rect 549266 442658 549502 442894
rect 549586 442658 549822 442894
rect 549266 442338 549502 442574
rect 549586 442338 549822 442574
rect 545546 438938 545782 439174
rect 545866 438938 546102 439174
rect 545546 438618 545782 438854
rect 545866 438618 546102 438854
rect 533647 435218 533883 435454
rect 533647 434898 533883 435134
rect 542088 435218 542324 435454
rect 542088 434898 542324 435134
rect 531866 425258 532102 425494
rect 532186 425258 532422 425494
rect 531866 424938 532102 425174
rect 532186 424938 532422 425174
rect 531866 389258 532102 389494
rect 532186 389258 532422 389494
rect 531866 388938 532102 389174
rect 532186 388938 532422 389174
rect 531866 353258 532102 353494
rect 532186 353258 532422 353494
rect 531866 352938 532102 353174
rect 532186 352938 532422 353174
rect 528146 313538 528382 313774
rect 528466 313538 528702 313774
rect 528146 313218 528382 313454
rect 528466 313218 528702 313454
rect 528146 277538 528382 277774
rect 528466 277538 528702 277774
rect 528146 277218 528382 277454
rect 528466 277218 528702 277454
rect 531866 317258 532102 317494
rect 532186 317258 532422 317494
rect 531866 316938 532102 317174
rect 532186 316938 532422 317174
rect 531866 281258 532102 281494
rect 532186 281258 532422 281494
rect 531866 280938 532102 281174
rect 532186 280938 532422 281174
rect 479610 258938 479846 259174
rect 479610 258618 479846 258854
rect 510330 258938 510566 259174
rect 510330 258618 510566 258854
rect 464250 255218 464486 255454
rect 464250 254898 464486 255134
rect 494970 255218 495206 255454
rect 494970 254898 495206 255134
rect 525690 255218 525926 255454
rect 525690 254898 525926 255134
rect 459866 245258 460102 245494
rect 460186 245258 460422 245494
rect 459866 244938 460102 245174
rect 460186 244938 460422 245174
rect 541826 399218 542062 399454
rect 542146 399218 542382 399454
rect 541826 398898 542062 399134
rect 542146 398898 542382 399134
rect 541826 363218 542062 363454
rect 542146 363218 542382 363454
rect 541826 362898 542062 363134
rect 542146 362898 542382 363134
rect 541826 327218 542062 327454
rect 542146 327218 542382 327454
rect 541826 326898 542062 327134
rect 542146 326898 542382 327134
rect 546308 438938 546544 439174
rect 546308 438618 546544 438854
rect 545546 402938 545782 403174
rect 545866 402938 546102 403174
rect 545546 402618 545782 402854
rect 545866 402618 546102 402854
rect 545546 366938 545782 367174
rect 545866 366938 546102 367174
rect 545546 366618 545782 366854
rect 545866 366618 546102 366854
rect 545546 330938 545782 331174
rect 545866 330938 546102 331174
rect 545546 330618 545782 330854
rect 545866 330618 546102 330854
rect 541826 291218 542062 291454
rect 542146 291218 542382 291454
rect 541826 290898 542062 291134
rect 542146 290898 542382 291134
rect 531866 245258 532102 245494
rect 532186 245258 532422 245494
rect 531866 244938 532102 245174
rect 532186 244938 532422 245174
rect 479610 222938 479846 223174
rect 479610 222618 479846 222854
rect 510330 222938 510566 223174
rect 510330 222618 510566 222854
rect 464250 219218 464486 219454
rect 464250 218898 464486 219134
rect 494970 219218 495206 219454
rect 494970 218898 495206 219134
rect 525690 219218 525926 219454
rect 525690 218898 525926 219134
rect 459866 209258 460102 209494
rect 460186 209258 460422 209494
rect 459866 208938 460102 209174
rect 460186 208938 460422 209174
rect 531866 209258 532102 209494
rect 532186 209258 532422 209494
rect 531866 208938 532102 209174
rect 532186 208938 532422 209174
rect 459866 173258 460102 173494
rect 460186 173258 460422 173494
rect 459866 172938 460102 173174
rect 460186 172938 460422 173174
rect 459866 137258 460102 137494
rect 460186 137258 460422 137494
rect 459866 136938 460102 137174
rect 460186 136938 460422 137174
rect 459866 101258 460102 101494
rect 460186 101258 460422 101494
rect 459866 100938 460102 101174
rect 460186 100938 460422 101174
rect 459866 65258 460102 65494
rect 460186 65258 460422 65494
rect 459866 64938 460102 65174
rect 460186 64938 460422 65174
rect 459866 29258 460102 29494
rect 460186 29258 460422 29494
rect 459866 28938 460102 29174
rect 460186 28938 460422 29174
rect 456146 -6342 456382 -6106
rect 456466 -6342 456702 -6106
rect 456146 -6662 456382 -6426
rect 456466 -6662 456702 -6426
rect 459866 -7302 460102 -7066
rect 460186 -7302 460422 -7066
rect 459866 -7622 460102 -7386
rect 460186 -7622 460422 -7386
rect 469826 183218 470062 183454
rect 470146 183218 470382 183454
rect 469826 182898 470062 183134
rect 470146 182898 470382 183134
rect 469826 147218 470062 147454
rect 470146 147218 470382 147454
rect 469826 146898 470062 147134
rect 470146 146898 470382 147134
rect 469826 111218 470062 111454
rect 470146 111218 470382 111454
rect 469826 110898 470062 111134
rect 470146 110898 470382 111134
rect 469826 75218 470062 75454
rect 470146 75218 470382 75454
rect 469826 74898 470062 75134
rect 470146 74898 470382 75134
rect 469826 39218 470062 39454
rect 470146 39218 470382 39454
rect 469826 38898 470062 39134
rect 470146 38898 470382 39134
rect 469826 3218 470062 3454
rect 470146 3218 470382 3454
rect 469826 2898 470062 3134
rect 470146 2898 470382 3134
rect 469826 -582 470062 -346
rect 470146 -582 470382 -346
rect 469826 -902 470062 -666
rect 470146 -902 470382 -666
rect 473546 186938 473782 187174
rect 473866 186938 474102 187174
rect 473546 186618 473782 186854
rect 473866 186618 474102 186854
rect 473546 150938 473782 151174
rect 473866 150938 474102 151174
rect 473546 150618 473782 150854
rect 473866 150618 474102 150854
rect 473546 114938 473782 115174
rect 473866 114938 474102 115174
rect 473546 114618 473782 114854
rect 473866 114618 474102 114854
rect 473546 78938 473782 79174
rect 473866 78938 474102 79174
rect 473546 78618 473782 78854
rect 473866 78618 474102 78854
rect 473546 42938 473782 43174
rect 473866 42938 474102 43174
rect 473546 42618 473782 42854
rect 473866 42618 474102 42854
rect 473546 6938 473782 7174
rect 473866 6938 474102 7174
rect 473546 6618 473782 6854
rect 473866 6618 474102 6854
rect 473546 -1542 473782 -1306
rect 473866 -1542 474102 -1306
rect 473546 -1862 473782 -1626
rect 473866 -1862 474102 -1626
rect 477266 190658 477502 190894
rect 477586 190658 477822 190894
rect 477266 190338 477502 190574
rect 477586 190338 477822 190574
rect 477266 154658 477502 154894
rect 477586 154658 477822 154894
rect 477266 154338 477502 154574
rect 477586 154338 477822 154574
rect 477266 118658 477502 118894
rect 477586 118658 477822 118894
rect 477266 118338 477502 118574
rect 477586 118338 477822 118574
rect 477266 82658 477502 82894
rect 477586 82658 477822 82894
rect 477266 82338 477502 82574
rect 477586 82338 477822 82574
rect 477266 46658 477502 46894
rect 477586 46658 477822 46894
rect 477266 46338 477502 46574
rect 477586 46338 477822 46574
rect 477266 10658 477502 10894
rect 477586 10658 477822 10894
rect 477266 10338 477502 10574
rect 477586 10338 477822 10574
rect 477266 -2502 477502 -2266
rect 477586 -2502 477822 -2266
rect 477266 -2822 477502 -2586
rect 477586 -2822 477822 -2586
rect 480986 194378 481222 194614
rect 481306 194378 481542 194614
rect 480986 194058 481222 194294
rect 481306 194058 481542 194294
rect 480986 158378 481222 158614
rect 481306 158378 481542 158614
rect 480986 158058 481222 158294
rect 481306 158058 481542 158294
rect 480986 122378 481222 122614
rect 481306 122378 481542 122614
rect 480986 122058 481222 122294
rect 481306 122058 481542 122294
rect 484706 198098 484942 198334
rect 485026 198098 485262 198334
rect 484706 197778 484942 198014
rect 485026 197778 485262 198014
rect 484706 162098 484942 162334
rect 485026 162098 485262 162334
rect 484706 161778 484942 162014
rect 485026 161778 485262 162014
rect 488426 165818 488662 166054
rect 488746 165818 488982 166054
rect 488426 165498 488662 165734
rect 488746 165498 488982 165734
rect 505826 183218 506062 183454
rect 506146 183218 506382 183454
rect 505826 182898 506062 183134
rect 506146 182898 506382 183134
rect 505826 147218 506062 147454
rect 506146 147218 506382 147454
rect 505826 146898 506062 147134
rect 506146 146898 506382 147134
rect 509546 186938 509782 187174
rect 509866 186938 510102 187174
rect 509546 186618 509782 186854
rect 509866 186618 510102 186854
rect 509546 150938 509782 151174
rect 509866 150938 510102 151174
rect 509546 150618 509782 150854
rect 509866 150618 510102 150854
rect 513266 190658 513502 190894
rect 513586 190658 513822 190894
rect 513266 190338 513502 190574
rect 513586 190338 513822 190574
rect 513266 154658 513502 154894
rect 513586 154658 513822 154894
rect 513266 154338 513502 154574
rect 513586 154338 513822 154574
rect 516986 194378 517222 194614
rect 517306 194378 517542 194614
rect 516986 194058 517222 194294
rect 517306 194058 517542 194294
rect 516986 158378 517222 158614
rect 517306 158378 517542 158614
rect 516986 158058 517222 158294
rect 517306 158058 517542 158294
rect 520706 198098 520942 198334
rect 521026 198098 521262 198334
rect 520706 197778 520942 198014
rect 521026 197778 521262 198014
rect 520706 162098 520942 162334
rect 521026 162098 521262 162334
rect 520706 161778 520942 162014
rect 521026 161778 521262 162014
rect 524426 165818 524662 166054
rect 524746 165818 524982 166054
rect 524426 165498 524662 165734
rect 524746 165498 524982 165734
rect 531866 173258 532102 173494
rect 532186 173258 532422 173494
rect 531866 172938 532102 173174
rect 532186 172938 532422 173174
rect 541826 255218 542062 255454
rect 542146 255218 542382 255454
rect 541826 254898 542062 255134
rect 542146 254898 542382 255134
rect 541826 219218 542062 219454
rect 542146 219218 542382 219454
rect 541826 218898 542062 219134
rect 542146 218898 542382 219134
rect 541826 183218 542062 183454
rect 542146 183218 542382 183454
rect 541826 182898 542062 183134
rect 542146 182898 542382 183134
rect 541826 147218 542062 147454
rect 542146 147218 542382 147454
rect 541826 146898 542062 147134
rect 542146 146898 542382 147134
rect 484706 126098 484942 126334
rect 485026 126098 485262 126334
rect 484706 125778 484942 126014
rect 485026 125778 485262 126014
rect 484250 111218 484486 111454
rect 484250 110898 484486 111134
rect 480986 86378 481222 86614
rect 481306 86378 481542 86614
rect 480986 86058 481222 86294
rect 481306 86058 481542 86294
rect 480986 50378 481222 50614
rect 481306 50378 481542 50614
rect 480986 50058 481222 50294
rect 481306 50058 481542 50294
rect 480986 14378 481222 14614
rect 481306 14378 481542 14614
rect 480986 14058 481222 14294
rect 481306 14058 481542 14294
rect 480986 -3462 481222 -3226
rect 481306 -3462 481542 -3226
rect 480986 -3782 481222 -3546
rect 481306 -3782 481542 -3546
rect 499610 114938 499846 115174
rect 499610 114618 499846 114854
rect 530330 114938 530566 115174
rect 530330 114618 530566 114854
rect 514970 111218 515206 111454
rect 514970 110898 515206 111134
rect 541826 111218 542062 111454
rect 542146 111218 542382 111454
rect 541826 110898 542062 111134
rect 542146 110898 542382 111134
rect 484706 90098 484942 90334
rect 485026 90098 485262 90334
rect 484706 89778 484942 90014
rect 485026 89778 485262 90014
rect 484706 54098 484942 54334
rect 485026 54098 485262 54334
rect 484706 53778 484942 54014
rect 485026 53778 485262 54014
rect 484706 18098 484942 18334
rect 485026 18098 485262 18334
rect 484706 17778 484942 18014
rect 485026 17778 485262 18014
rect 484706 -4422 484942 -4186
rect 485026 -4422 485262 -4186
rect 484706 -4742 484942 -4506
rect 485026 -4742 485262 -4506
rect 488426 57818 488662 58054
rect 488746 57818 488982 58054
rect 488426 57498 488662 57734
rect 488746 57498 488982 57734
rect 488426 21818 488662 22054
rect 488746 21818 488982 22054
rect 488426 21498 488662 21734
rect 488746 21498 488982 21734
rect 488426 -5382 488662 -5146
rect 488746 -5382 488982 -5146
rect 488426 -5702 488662 -5466
rect 488746 -5702 488982 -5466
rect 492146 61538 492382 61774
rect 492466 61538 492702 61774
rect 492146 61218 492382 61454
rect 492466 61218 492702 61454
rect 492146 25538 492382 25774
rect 492466 25538 492702 25774
rect 492146 25218 492382 25454
rect 492466 25218 492702 25454
rect 492146 -6342 492382 -6106
rect 492466 -6342 492702 -6106
rect 492146 -6662 492382 -6426
rect 492466 -6662 492702 -6426
rect 495866 65258 496102 65494
rect 496186 65258 496422 65494
rect 495866 64938 496102 65174
rect 496186 64938 496422 65174
rect 495866 29258 496102 29494
rect 496186 29258 496422 29494
rect 495866 28938 496102 29174
rect 496186 28938 496422 29174
rect 495866 -7302 496102 -7066
rect 496186 -7302 496422 -7066
rect 495866 -7622 496102 -7386
rect 496186 -7622 496422 -7386
rect 505826 75218 506062 75454
rect 506146 75218 506382 75454
rect 505826 74898 506062 75134
rect 506146 74898 506382 75134
rect 505826 39218 506062 39454
rect 506146 39218 506382 39454
rect 505826 38898 506062 39134
rect 506146 38898 506382 39134
rect 505826 3218 506062 3454
rect 506146 3218 506382 3454
rect 505826 2898 506062 3134
rect 506146 2898 506382 3134
rect 505826 -582 506062 -346
rect 506146 -582 506382 -346
rect 505826 -902 506062 -666
rect 506146 -902 506382 -666
rect 509546 78938 509782 79174
rect 509866 78938 510102 79174
rect 509546 78618 509782 78854
rect 509866 78618 510102 78854
rect 509546 42938 509782 43174
rect 509866 42938 510102 43174
rect 509546 42618 509782 42854
rect 509866 42618 510102 42854
rect 509546 6938 509782 7174
rect 509866 6938 510102 7174
rect 509546 6618 509782 6854
rect 509866 6618 510102 6854
rect 509546 -1542 509782 -1306
rect 509866 -1542 510102 -1306
rect 509546 -1862 509782 -1626
rect 509866 -1862 510102 -1626
rect 513266 46658 513502 46894
rect 513586 46658 513822 46894
rect 513266 46338 513502 46574
rect 513586 46338 513822 46574
rect 513266 10658 513502 10894
rect 513586 10658 513822 10894
rect 513266 10338 513502 10574
rect 513586 10338 513822 10574
rect 513266 -2502 513502 -2266
rect 513586 -2502 513822 -2266
rect 513266 -2822 513502 -2586
rect 513586 -2822 513822 -2586
rect 516986 50378 517222 50614
rect 517306 50378 517542 50614
rect 516986 50058 517222 50294
rect 517306 50058 517542 50294
rect 516986 14378 517222 14614
rect 517306 14378 517542 14614
rect 516986 14058 517222 14294
rect 517306 14058 517542 14294
rect 516986 -3462 517222 -3226
rect 517306 -3462 517542 -3226
rect 516986 -3782 517222 -3546
rect 517306 -3782 517542 -3546
rect 520706 54098 520942 54334
rect 521026 54098 521262 54334
rect 520706 53778 520942 54014
rect 521026 53778 521262 54014
rect 520706 18098 520942 18334
rect 521026 18098 521262 18334
rect 520706 17778 520942 18014
rect 521026 17778 521262 18014
rect 520706 -4422 520942 -4186
rect 521026 -4422 521262 -4186
rect 520706 -4742 520942 -4506
rect 521026 -4742 521262 -4506
rect 524426 57818 524662 58054
rect 524746 57818 524982 58054
rect 524426 57498 524662 57734
rect 524746 57498 524982 57734
rect 524426 21818 524662 22054
rect 524746 21818 524982 22054
rect 524426 21498 524662 21734
rect 524746 21498 524982 21734
rect 524426 -5382 524662 -5146
rect 524746 -5382 524982 -5146
rect 524426 -5702 524662 -5466
rect 524746 -5702 524982 -5466
rect 528146 61538 528382 61774
rect 528466 61538 528702 61774
rect 528146 61218 528382 61454
rect 528466 61218 528702 61454
rect 528146 25538 528382 25774
rect 528466 25538 528702 25774
rect 528146 25218 528382 25454
rect 528466 25218 528702 25454
rect 528146 -6342 528382 -6106
rect 528466 -6342 528702 -6106
rect 528146 -6662 528382 -6426
rect 528466 -6662 528702 -6426
rect 531866 65258 532102 65494
rect 532186 65258 532422 65494
rect 531866 64938 532102 65174
rect 532186 64938 532422 65174
rect 531866 29258 532102 29494
rect 532186 29258 532422 29494
rect 531866 28938 532102 29174
rect 532186 28938 532422 29174
rect 531866 -7302 532102 -7066
rect 532186 -7302 532422 -7066
rect 531866 -7622 532102 -7386
rect 532186 -7622 532422 -7386
rect 545546 294938 545782 295174
rect 545866 294938 546102 295174
rect 545546 294618 545782 294854
rect 545866 294618 546102 294854
rect 545546 258938 545782 259174
rect 545866 258938 546102 259174
rect 545546 258618 545782 258854
rect 545866 258618 546102 258854
rect 545546 222938 545782 223174
rect 545866 222938 546102 223174
rect 545546 222618 545782 222854
rect 545866 222618 546102 222854
rect 545546 186938 545782 187174
rect 545866 186938 546102 187174
rect 545546 186618 545782 186854
rect 545866 186618 546102 186854
rect 545546 150938 545782 151174
rect 545866 150938 546102 151174
rect 545546 150618 545782 150854
rect 545866 150618 546102 150854
rect 545546 114938 545782 115174
rect 545866 114938 546102 115174
rect 545546 114618 545782 114854
rect 545866 114618 546102 114854
rect 541826 75218 542062 75454
rect 542146 75218 542382 75454
rect 541826 74898 542062 75134
rect 542146 74898 542382 75134
rect 545546 78938 545782 79174
rect 545866 78938 546102 79174
rect 545546 78618 545782 78854
rect 545866 78618 546102 78854
rect 552986 707482 553222 707718
rect 553306 707482 553542 707718
rect 552986 707162 553222 707398
rect 553306 707162 553542 707398
rect 552986 698378 553222 698614
rect 553306 698378 553542 698614
rect 552986 698058 553222 698294
rect 553306 698058 553542 698294
rect 552986 662378 553222 662614
rect 553306 662378 553542 662614
rect 552986 662058 553222 662294
rect 553306 662058 553542 662294
rect 552986 626378 553222 626614
rect 553306 626378 553542 626614
rect 552986 626058 553222 626294
rect 553306 626058 553542 626294
rect 552986 590378 553222 590614
rect 553306 590378 553542 590614
rect 552986 590058 553222 590294
rect 553306 590058 553542 590294
rect 552986 554378 553222 554614
rect 553306 554378 553542 554614
rect 552986 554058 553222 554294
rect 553306 554058 553542 554294
rect 552986 518378 553222 518614
rect 553306 518378 553542 518614
rect 552986 518058 553222 518294
rect 553306 518058 553542 518294
rect 552986 482378 553222 482614
rect 553306 482378 553542 482614
rect 552986 482058 553222 482294
rect 553306 482058 553542 482294
rect 552986 446378 553222 446614
rect 553306 446378 553542 446614
rect 552986 446058 553222 446294
rect 553306 446058 553542 446294
rect 550529 435218 550765 435454
rect 550529 434898 550765 435134
rect 549266 406658 549502 406894
rect 549586 406658 549822 406894
rect 549266 406338 549502 406574
rect 549586 406338 549822 406574
rect 556706 708442 556942 708678
rect 557026 708442 557262 708678
rect 556706 708122 556942 708358
rect 557026 708122 557262 708358
rect 560426 709402 560662 709638
rect 560746 709402 560982 709638
rect 560426 709082 560662 709318
rect 560746 709082 560982 709318
rect 556706 666098 556942 666334
rect 557026 666098 557262 666334
rect 556706 665778 556942 666014
rect 557026 665778 557262 666014
rect 556706 630098 556942 630334
rect 557026 630098 557262 630334
rect 556706 629778 556942 630014
rect 557026 629778 557262 630014
rect 556706 594098 556942 594334
rect 557026 594098 557262 594334
rect 556706 593778 556942 594014
rect 557026 593778 557262 594014
rect 556706 558098 556942 558334
rect 557026 558098 557262 558334
rect 556706 557778 556942 558014
rect 557026 557778 557262 558014
rect 556706 522098 556942 522334
rect 557026 522098 557262 522334
rect 556706 521778 556942 522014
rect 557026 521778 557262 522014
rect 556706 486098 556942 486334
rect 557026 486098 557262 486334
rect 556706 485778 556942 486014
rect 557026 485778 557262 486014
rect 556706 450098 556942 450334
rect 557026 450098 557262 450334
rect 556706 449778 556942 450014
rect 557026 449778 557262 450014
rect 554749 438938 554985 439174
rect 554749 438618 554985 438854
rect 552986 410378 553222 410614
rect 553306 410378 553542 410614
rect 552986 410058 553222 410294
rect 553306 410058 553542 410294
rect 556706 414098 556942 414334
rect 557026 414098 557262 414334
rect 556706 413778 556942 414014
rect 557026 413778 557262 414014
rect 556706 378007 556942 378243
rect 557026 378007 557262 378243
rect 549266 370658 549502 370894
rect 549586 370658 549822 370894
rect 549266 370338 549502 370574
rect 549586 370338 549822 370574
rect 554918 366938 555154 367174
rect 554918 366618 555154 366854
rect 552952 363218 553188 363454
rect 552952 362898 553188 363134
rect 556885 363218 557121 363454
rect 556885 362898 557121 363134
rect 549266 334658 549502 334894
rect 549586 334658 549822 334894
rect 549266 334338 549502 334574
rect 549586 334338 549822 334574
rect 549266 298658 549502 298894
rect 549586 298658 549822 298894
rect 549266 298338 549502 298574
rect 549586 298338 549822 298574
rect 549266 262658 549502 262894
rect 549586 262658 549822 262894
rect 549266 262338 549502 262574
rect 549586 262338 549822 262574
rect 549266 226658 549502 226894
rect 549586 226658 549822 226894
rect 549266 226338 549502 226574
rect 549586 226338 549822 226574
rect 549266 190658 549502 190894
rect 549586 190658 549822 190894
rect 549266 190338 549502 190574
rect 549586 190338 549822 190574
rect 549266 154658 549502 154894
rect 549586 154658 549822 154894
rect 549266 154338 549502 154574
rect 549586 154338 549822 154574
rect 549266 118658 549502 118894
rect 549586 118658 549822 118894
rect 549266 118338 549502 118574
rect 549586 118338 549822 118574
rect 549266 82658 549502 82894
rect 549586 82658 549822 82894
rect 549266 82338 549502 82574
rect 549586 82338 549822 82574
rect 552986 338378 553222 338614
rect 553306 338378 553542 338614
rect 552986 338058 553222 338294
rect 553306 338058 553542 338294
rect 552986 302378 553222 302614
rect 553306 302378 553542 302614
rect 552986 302058 553222 302294
rect 553306 302058 553542 302294
rect 552986 266378 553222 266614
rect 553306 266378 553542 266614
rect 552986 266058 553222 266294
rect 553306 266058 553542 266294
rect 552986 230378 553222 230614
rect 553306 230378 553542 230614
rect 552986 230058 553222 230294
rect 553306 230058 553542 230294
rect 552986 194378 553222 194614
rect 553306 194378 553542 194614
rect 552986 194058 553222 194294
rect 553306 194058 553542 194294
rect 552986 158378 553222 158614
rect 553306 158378 553542 158614
rect 552986 158058 553222 158294
rect 553306 158058 553542 158294
rect 552986 122378 553222 122614
rect 553306 122378 553542 122614
rect 552986 122058 553222 122294
rect 553306 122058 553542 122294
rect 552986 86378 553222 86614
rect 553306 86378 553542 86614
rect 552986 86058 553222 86294
rect 553306 86058 553542 86294
rect 556706 342098 556942 342334
rect 557026 342098 557262 342334
rect 556706 341778 556942 342014
rect 557026 341778 557262 342014
rect 560426 669818 560662 670054
rect 560746 669818 560982 670054
rect 560426 669498 560662 669734
rect 560746 669498 560982 669734
rect 560426 633818 560662 634054
rect 560746 633818 560982 634054
rect 560426 633498 560662 633734
rect 560746 633498 560982 633734
rect 560426 597818 560662 598054
rect 560746 597818 560982 598054
rect 560426 597498 560662 597734
rect 560746 597498 560982 597734
rect 560426 561818 560662 562054
rect 560746 561818 560982 562054
rect 560426 561498 560662 561734
rect 560746 561498 560982 561734
rect 560426 525818 560662 526054
rect 560746 525818 560982 526054
rect 560426 525498 560662 525734
rect 560746 525498 560982 525734
rect 560426 489818 560662 490054
rect 560746 489818 560982 490054
rect 560426 489498 560662 489734
rect 560746 489498 560982 489734
rect 560426 453818 560662 454054
rect 560746 453818 560982 454054
rect 560426 453498 560662 453734
rect 560746 453498 560982 453734
rect 560426 417818 560662 418054
rect 560746 417818 560982 418054
rect 560426 417498 560662 417734
rect 560746 417498 560982 417734
rect 560426 381818 560662 382054
rect 560746 381818 560982 382054
rect 560426 381498 560662 381734
rect 560746 381498 560982 381734
rect 564146 710362 564382 710598
rect 564466 710362 564702 710598
rect 564146 710042 564382 710278
rect 564466 710042 564702 710278
rect 564146 673538 564382 673774
rect 564466 673538 564702 673774
rect 564146 673218 564382 673454
rect 564466 673218 564702 673454
rect 564146 637538 564382 637774
rect 564466 637538 564702 637774
rect 564146 637218 564382 637454
rect 564466 637218 564702 637454
rect 564146 601538 564382 601774
rect 564466 601538 564702 601774
rect 564146 601218 564382 601454
rect 564466 601218 564702 601454
rect 564146 565538 564382 565774
rect 564466 565538 564702 565774
rect 564146 565218 564382 565454
rect 564466 565218 564702 565454
rect 564146 529538 564382 529774
rect 564466 529538 564702 529774
rect 564146 529218 564382 529454
rect 564466 529218 564702 529454
rect 564146 493538 564382 493774
rect 564466 493538 564702 493774
rect 564146 493218 564382 493454
rect 564466 493218 564702 493454
rect 564146 457538 564382 457774
rect 564466 457538 564702 457774
rect 564146 457218 564382 457454
rect 564466 457218 564702 457454
rect 564146 421538 564382 421774
rect 564466 421538 564702 421774
rect 564146 421218 564382 421454
rect 564466 421218 564702 421454
rect 564146 385538 564382 385774
rect 564466 385538 564702 385774
rect 564146 385218 564382 385454
rect 564466 385218 564702 385454
rect 567866 711322 568102 711558
rect 568186 711322 568422 711558
rect 567866 711002 568102 711238
rect 568186 711002 568422 711238
rect 567866 677258 568102 677494
rect 568186 677258 568422 677494
rect 567866 676938 568102 677174
rect 568186 676938 568422 677174
rect 567866 641258 568102 641494
rect 568186 641258 568422 641494
rect 567866 640938 568102 641174
rect 568186 640938 568422 641174
rect 567866 605258 568102 605494
rect 568186 605258 568422 605494
rect 567866 604938 568102 605174
rect 568186 604938 568422 605174
rect 567866 569258 568102 569494
rect 568186 569258 568422 569494
rect 567866 568938 568102 569174
rect 568186 568938 568422 569174
rect 567866 533258 568102 533494
rect 568186 533258 568422 533494
rect 567866 532938 568102 533174
rect 568186 532938 568422 533174
rect 567866 497258 568102 497494
rect 568186 497258 568422 497494
rect 567866 496938 568102 497174
rect 568186 496938 568422 497174
rect 567866 461258 568102 461494
rect 568186 461258 568422 461494
rect 567866 460938 568102 461174
rect 568186 460938 568422 461174
rect 567866 425258 568102 425494
rect 568186 425258 568422 425494
rect 567866 424938 568102 425174
rect 568186 424938 568422 425174
rect 567866 389258 568102 389494
rect 568186 389258 568422 389494
rect 567866 388938 568102 389174
rect 568186 388938 568422 389174
rect 558851 366938 559087 367174
rect 558851 366618 559087 366854
rect 562784 366938 563020 367174
rect 562784 366618 563020 366854
rect 566717 366938 566953 367174
rect 566717 366618 566953 366854
rect 560818 363218 561054 363454
rect 560818 362898 561054 363134
rect 564751 363218 564987 363454
rect 564751 362898 564987 363134
rect 560426 345818 560662 346054
rect 560746 345818 560982 346054
rect 560426 345498 560662 345734
rect 560746 345498 560982 345734
rect 556706 306098 556942 306334
rect 557026 306098 557262 306334
rect 556706 305778 556942 306014
rect 557026 305778 557262 306014
rect 556706 270098 556942 270334
rect 557026 270098 557262 270334
rect 556706 269778 556942 270014
rect 557026 269778 557262 270014
rect 556706 234098 556942 234334
rect 557026 234098 557262 234334
rect 556706 233778 556942 234014
rect 557026 233778 557262 234014
rect 556706 198098 556942 198334
rect 557026 198098 557262 198334
rect 556706 197778 556942 198014
rect 557026 197778 557262 198014
rect 556706 162098 556942 162334
rect 557026 162098 557262 162334
rect 556706 161778 556942 162014
rect 557026 161778 557262 162014
rect 556706 126098 556942 126334
rect 557026 126098 557262 126334
rect 556706 125778 556942 126014
rect 557026 125778 557262 126014
rect 556706 90098 556942 90334
rect 557026 90098 557262 90334
rect 556706 89778 556942 90014
rect 557026 89778 557262 90014
rect 556706 54098 556942 54334
rect 557026 54098 557262 54334
rect 556706 53778 556942 54014
rect 557026 53778 557262 54014
rect 549266 46658 549502 46894
rect 549586 46658 549822 46894
rect 549266 46338 549502 46574
rect 549586 46338 549822 46574
rect 545930 42938 546166 43174
rect 545930 42618 546166 42854
rect 541826 39218 542062 39454
rect 542146 39218 542382 39454
rect 541826 38898 542062 39134
rect 542146 38898 542382 39134
rect 543458 39218 543694 39454
rect 543458 38898 543694 39134
rect 548403 39218 548639 39454
rect 548403 38898 548639 39134
rect 541826 3218 542062 3454
rect 542146 3218 542382 3454
rect 541826 2898 542062 3134
rect 542146 2898 542382 3134
rect 541826 -582 542062 -346
rect 542146 -582 542382 -346
rect 541826 -902 542062 -666
rect 542146 -902 542382 -666
rect 545546 6938 545782 7174
rect 545866 6938 546102 7174
rect 545546 6618 545782 6854
rect 545866 6618 546102 6854
rect 545546 -1542 545782 -1306
rect 545866 -1542 546102 -1306
rect 545546 -1862 545782 -1626
rect 545866 -1862 546102 -1626
rect 550875 42938 551111 43174
rect 550875 42618 551111 42854
rect 555820 42938 556056 43174
rect 555820 42618 556056 42854
rect 553348 39218 553584 39454
rect 553348 38898 553584 39134
rect 549266 10658 549502 10894
rect 549586 10658 549822 10894
rect 549266 10338 549502 10574
rect 549586 10338 549822 10574
rect 549266 -2502 549502 -2266
rect 549586 -2502 549822 -2266
rect 549266 -2822 549502 -2586
rect 549586 -2822 549822 -2586
rect 552986 14378 553222 14614
rect 553306 14378 553542 14614
rect 552986 14058 553222 14294
rect 553306 14058 553542 14294
rect 552986 -3462 553222 -3226
rect 553306 -3462 553542 -3226
rect 552986 -3782 553222 -3546
rect 553306 -3782 553542 -3546
rect 560426 309818 560662 310054
rect 560746 309818 560982 310054
rect 560426 309498 560662 309734
rect 560746 309498 560982 309734
rect 560426 273818 560662 274054
rect 560746 273818 560982 274054
rect 560426 273498 560662 273734
rect 560746 273498 560982 273734
rect 560426 237818 560662 238054
rect 560746 237818 560982 238054
rect 560426 237498 560662 237734
rect 560746 237498 560982 237734
rect 560426 201818 560662 202054
rect 560746 201818 560982 202054
rect 560426 201498 560662 201734
rect 560746 201498 560982 201734
rect 560426 165818 560662 166054
rect 560746 165818 560982 166054
rect 560426 165498 560662 165734
rect 560746 165498 560982 165734
rect 560426 129818 560662 130054
rect 560746 129818 560982 130054
rect 560426 129498 560662 129734
rect 560746 129498 560982 129734
rect 560426 93818 560662 94054
rect 560746 93818 560982 94054
rect 560426 93498 560662 93734
rect 560746 93498 560982 93734
rect 560426 57818 560662 58054
rect 560746 57818 560982 58054
rect 560426 57498 560662 57734
rect 560746 57498 560982 57734
rect 564146 349538 564382 349774
rect 564466 349538 564702 349774
rect 564146 349218 564382 349454
rect 564466 349218 564702 349454
rect 564146 313538 564382 313774
rect 564466 313538 564702 313774
rect 564146 313218 564382 313454
rect 564466 313218 564702 313454
rect 564146 277538 564382 277774
rect 564466 277538 564702 277774
rect 564146 277218 564382 277454
rect 564466 277218 564702 277454
rect 564146 241538 564382 241774
rect 564466 241538 564702 241774
rect 564146 241218 564382 241454
rect 564466 241218 564702 241454
rect 564146 205538 564382 205774
rect 564466 205538 564702 205774
rect 564146 205218 564382 205454
rect 564466 205218 564702 205454
rect 564146 169538 564382 169774
rect 564466 169538 564702 169774
rect 564146 169218 564382 169454
rect 564466 169218 564702 169454
rect 564146 133538 564382 133774
rect 564466 133538 564702 133774
rect 564146 133218 564382 133454
rect 564466 133218 564702 133454
rect 564146 97538 564382 97774
rect 564466 97538 564702 97774
rect 564146 97218 564382 97454
rect 564466 97218 564702 97454
rect 564146 61538 564382 61774
rect 564466 61538 564702 61774
rect 564146 61218 564382 61454
rect 564466 61218 564702 61454
rect 560765 42938 561001 43174
rect 560765 42618 561001 42854
rect 558293 39218 558529 39454
rect 558293 38898 558529 39134
rect 556706 18098 556942 18334
rect 557026 18098 557262 18334
rect 556706 17778 556942 18014
rect 557026 17778 557262 18014
rect 556706 -4422 556942 -4186
rect 557026 -4422 557262 -4186
rect 556706 -4742 556942 -4506
rect 557026 -4742 557262 -4506
rect 560426 21818 560662 22054
rect 560746 21818 560982 22054
rect 560426 21498 560662 21734
rect 560746 21498 560982 21734
rect 560426 -5382 560662 -5146
rect 560746 -5382 560982 -5146
rect 560426 -5702 560662 -5466
rect 560746 -5702 560982 -5466
rect 564146 25538 564382 25774
rect 564466 25538 564702 25774
rect 564146 25218 564382 25454
rect 564466 25218 564702 25454
rect 564146 -6342 564382 -6106
rect 564466 -6342 564702 -6106
rect 564146 -6662 564382 -6426
rect 564466 -6662 564702 -6426
rect 567866 353258 568102 353494
rect 568186 353258 568422 353494
rect 567866 352938 568102 353174
rect 568186 352938 568422 353174
rect 567866 317258 568102 317494
rect 568186 317258 568422 317494
rect 567866 316938 568102 317174
rect 568186 316938 568422 317174
rect 567866 281258 568102 281494
rect 568186 281258 568422 281494
rect 567866 280938 568102 281174
rect 568186 280938 568422 281174
rect 567866 245258 568102 245494
rect 568186 245258 568422 245494
rect 567866 244938 568102 245174
rect 568186 244938 568422 245174
rect 567866 209258 568102 209494
rect 568186 209258 568422 209494
rect 567866 208938 568102 209174
rect 568186 208938 568422 209174
rect 567866 173258 568102 173494
rect 568186 173258 568422 173494
rect 567866 172938 568102 173174
rect 568186 172938 568422 173174
rect 567866 137258 568102 137494
rect 568186 137258 568422 137494
rect 567866 136938 568102 137174
rect 568186 136938 568422 137174
rect 567866 101258 568102 101494
rect 568186 101258 568422 101494
rect 567866 100938 568102 101174
rect 568186 100938 568422 101174
rect 567866 65258 568102 65494
rect 568186 65258 568422 65494
rect 567866 64938 568102 65174
rect 568186 64938 568422 65174
rect 567866 29258 568102 29494
rect 568186 29258 568422 29494
rect 567866 28938 568102 29174
rect 568186 28938 568422 29174
rect 567866 -7302 568102 -7066
rect 568186 -7302 568422 -7066
rect 567866 -7622 568102 -7386
rect 568186 -7622 568422 -7386
rect 577826 704602 578062 704838
rect 578146 704602 578382 704838
rect 577826 704282 578062 704518
rect 578146 704282 578382 704518
rect 577826 687218 578062 687454
rect 578146 687218 578382 687454
rect 577826 686898 578062 687134
rect 578146 686898 578382 687134
rect 577826 651218 578062 651454
rect 578146 651218 578382 651454
rect 577826 650898 578062 651134
rect 578146 650898 578382 651134
rect 577826 615218 578062 615454
rect 578146 615218 578382 615454
rect 577826 614898 578062 615134
rect 578146 614898 578382 615134
rect 577826 579218 578062 579454
rect 578146 579218 578382 579454
rect 577826 578898 578062 579134
rect 578146 578898 578382 579134
rect 577826 543218 578062 543454
rect 578146 543218 578382 543454
rect 577826 542898 578062 543134
rect 578146 542898 578382 543134
rect 577826 507218 578062 507454
rect 578146 507218 578382 507454
rect 577826 506898 578062 507134
rect 578146 506898 578382 507134
rect 577826 471218 578062 471454
rect 578146 471218 578382 471454
rect 577826 470898 578062 471134
rect 578146 470898 578382 471134
rect 577826 435218 578062 435454
rect 578146 435218 578382 435454
rect 577826 434898 578062 435134
rect 578146 434898 578382 435134
rect 577826 399218 578062 399454
rect 578146 399218 578382 399454
rect 577826 398898 578062 399134
rect 578146 398898 578382 399134
rect 577826 363218 578062 363454
rect 578146 363218 578382 363454
rect 577826 362898 578062 363134
rect 578146 362898 578382 363134
rect 577826 327218 578062 327454
rect 578146 327218 578382 327454
rect 577826 326898 578062 327134
rect 578146 326898 578382 327134
rect 577826 291218 578062 291454
rect 578146 291218 578382 291454
rect 577826 290898 578062 291134
rect 578146 290898 578382 291134
rect 577826 255218 578062 255454
rect 578146 255218 578382 255454
rect 577826 254898 578062 255134
rect 578146 254898 578382 255134
rect 577826 219218 578062 219454
rect 578146 219218 578382 219454
rect 577826 218898 578062 219134
rect 578146 218898 578382 219134
rect 577826 183218 578062 183454
rect 578146 183218 578382 183454
rect 577826 182898 578062 183134
rect 578146 182898 578382 183134
rect 577826 147218 578062 147454
rect 578146 147218 578382 147454
rect 577826 146898 578062 147134
rect 578146 146898 578382 147134
rect 577826 111218 578062 111454
rect 578146 111218 578382 111454
rect 577826 110898 578062 111134
rect 578146 110898 578382 111134
rect 577826 75218 578062 75454
rect 578146 75218 578382 75454
rect 577826 74898 578062 75134
rect 578146 74898 578382 75134
rect 577826 39218 578062 39454
rect 578146 39218 578382 39454
rect 577826 38898 578062 39134
rect 578146 38898 578382 39134
rect 577826 3218 578062 3454
rect 578146 3218 578382 3454
rect 577826 2898 578062 3134
rect 578146 2898 578382 3134
rect 577826 -582 578062 -346
rect 578146 -582 578382 -346
rect 577826 -902 578062 -666
rect 578146 -902 578382 -666
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 581546 705562 581782 705798
rect 581866 705562 582102 705798
rect 581546 705242 581782 705478
rect 581866 705242 582102 705478
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 581546 690938 581782 691174
rect 581866 690938 582102 691174
rect 581546 690618 581782 690854
rect 581866 690618 582102 690854
rect 581546 654938 581782 655174
rect 581866 654938 582102 655174
rect 581546 654618 581782 654854
rect 581866 654618 582102 654854
rect 581546 618938 581782 619174
rect 581866 618938 582102 619174
rect 581546 618618 581782 618854
rect 581866 618618 582102 618854
rect 581546 582938 581782 583174
rect 581866 582938 582102 583174
rect 581546 582618 581782 582854
rect 581866 582618 582102 582854
rect 581546 546938 581782 547174
rect 581866 546938 582102 547174
rect 581546 546618 581782 546854
rect 581866 546618 582102 546854
rect 581546 510938 581782 511174
rect 581866 510938 582102 511174
rect 581546 510618 581782 510854
rect 581866 510618 582102 510854
rect 581546 474938 581782 475174
rect 581866 474938 582102 475174
rect 581546 474618 581782 474854
rect 581866 474618 582102 474854
rect 581546 438938 581782 439174
rect 581866 438938 582102 439174
rect 581546 438618 581782 438854
rect 581866 438618 582102 438854
rect 581546 402938 581782 403174
rect 581866 402938 582102 403174
rect 581546 402618 581782 402854
rect 581866 402618 582102 402854
rect 581546 366938 581782 367174
rect 581866 366938 582102 367174
rect 581546 366618 581782 366854
rect 581866 366618 582102 366854
rect 581546 330938 581782 331174
rect 581866 330938 582102 331174
rect 581546 330618 581782 330854
rect 581866 330618 582102 330854
rect 581546 294938 581782 295174
rect 581866 294938 582102 295174
rect 581546 294618 581782 294854
rect 581866 294618 582102 294854
rect 581546 258938 581782 259174
rect 581866 258938 582102 259174
rect 581546 258618 581782 258854
rect 581866 258618 582102 258854
rect 581546 222938 581782 223174
rect 581866 222938 582102 223174
rect 581546 222618 581782 222854
rect 581866 222618 582102 222854
rect 581546 186938 581782 187174
rect 581866 186938 582102 187174
rect 581546 186618 581782 186854
rect 581866 186618 582102 186854
rect 581546 150938 581782 151174
rect 581866 150938 582102 151174
rect 581546 150618 581782 150854
rect 581866 150618 582102 150854
rect 581546 114938 581782 115174
rect 581866 114938 582102 115174
rect 581546 114618 581782 114854
rect 581866 114618 582102 114854
rect 581546 78938 581782 79174
rect 581866 78938 582102 79174
rect 581546 78618 581782 78854
rect 581866 78618 582102 78854
rect 581546 42938 581782 43174
rect 581866 42938 582102 43174
rect 581546 42618 581782 42854
rect 581866 42618 582102 42854
rect 581546 6938 581782 7174
rect 581866 6938 582102 7174
rect 581546 6618 581782 6854
rect 581866 6618 582102 6854
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 687218 585578 687454
rect 585662 687218 585898 687454
rect 585342 686898 585578 687134
rect 585662 686898 585898 687134
rect 585342 651218 585578 651454
rect 585662 651218 585898 651454
rect 585342 650898 585578 651134
rect 585662 650898 585898 651134
rect 585342 615218 585578 615454
rect 585662 615218 585898 615454
rect 585342 614898 585578 615134
rect 585662 614898 585898 615134
rect 585342 579218 585578 579454
rect 585662 579218 585898 579454
rect 585342 578898 585578 579134
rect 585662 578898 585898 579134
rect 585342 543218 585578 543454
rect 585662 543218 585898 543454
rect 585342 542898 585578 543134
rect 585662 542898 585898 543134
rect 585342 507218 585578 507454
rect 585662 507218 585898 507454
rect 585342 506898 585578 507134
rect 585662 506898 585898 507134
rect 585342 471218 585578 471454
rect 585662 471218 585898 471454
rect 585342 470898 585578 471134
rect 585662 470898 585898 471134
rect 585342 435218 585578 435454
rect 585662 435218 585898 435454
rect 585342 434898 585578 435134
rect 585662 434898 585898 435134
rect 585342 399218 585578 399454
rect 585662 399218 585898 399454
rect 585342 398898 585578 399134
rect 585662 398898 585898 399134
rect 585342 363218 585578 363454
rect 585662 363218 585898 363454
rect 585342 362898 585578 363134
rect 585662 362898 585898 363134
rect 585342 327218 585578 327454
rect 585662 327218 585898 327454
rect 585342 326898 585578 327134
rect 585662 326898 585898 327134
rect 585342 291218 585578 291454
rect 585662 291218 585898 291454
rect 585342 290898 585578 291134
rect 585662 290898 585898 291134
rect 585342 255218 585578 255454
rect 585662 255218 585898 255454
rect 585342 254898 585578 255134
rect 585662 254898 585898 255134
rect 585342 219218 585578 219454
rect 585662 219218 585898 219454
rect 585342 218898 585578 219134
rect 585662 218898 585898 219134
rect 585342 183218 585578 183454
rect 585662 183218 585898 183454
rect 585342 182898 585578 183134
rect 585662 182898 585898 183134
rect 585342 147218 585578 147454
rect 585662 147218 585898 147454
rect 585342 146898 585578 147134
rect 585662 146898 585898 147134
rect 585342 111218 585578 111454
rect 585662 111218 585898 111454
rect 585342 110898 585578 111134
rect 585662 110898 585898 111134
rect 585342 75218 585578 75454
rect 585662 75218 585898 75454
rect 585342 74898 585578 75134
rect 585662 74898 585898 75134
rect 585342 39218 585578 39454
rect 585662 39218 585898 39454
rect 585342 38898 585578 39134
rect 585662 38898 585898 39134
rect 585342 3218 585578 3454
rect 585662 3218 585898 3454
rect 585342 2898 585578 3134
rect 585662 2898 585898 3134
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 690938 586538 691174
rect 586622 690938 586858 691174
rect 586302 690618 586538 690854
rect 586622 690618 586858 690854
rect 586302 654938 586538 655174
rect 586622 654938 586858 655174
rect 586302 654618 586538 654854
rect 586622 654618 586858 654854
rect 586302 618938 586538 619174
rect 586622 618938 586858 619174
rect 586302 618618 586538 618854
rect 586622 618618 586858 618854
rect 586302 582938 586538 583174
rect 586622 582938 586858 583174
rect 586302 582618 586538 582854
rect 586622 582618 586858 582854
rect 586302 546938 586538 547174
rect 586622 546938 586858 547174
rect 586302 546618 586538 546854
rect 586622 546618 586858 546854
rect 586302 510938 586538 511174
rect 586622 510938 586858 511174
rect 586302 510618 586538 510854
rect 586622 510618 586858 510854
rect 586302 474938 586538 475174
rect 586622 474938 586858 475174
rect 586302 474618 586538 474854
rect 586622 474618 586858 474854
rect 586302 438938 586538 439174
rect 586622 438938 586858 439174
rect 586302 438618 586538 438854
rect 586622 438618 586858 438854
rect 586302 402938 586538 403174
rect 586622 402938 586858 403174
rect 586302 402618 586538 402854
rect 586622 402618 586858 402854
rect 586302 366938 586538 367174
rect 586622 366938 586858 367174
rect 586302 366618 586538 366854
rect 586622 366618 586858 366854
rect 586302 330938 586538 331174
rect 586622 330938 586858 331174
rect 586302 330618 586538 330854
rect 586622 330618 586858 330854
rect 586302 294938 586538 295174
rect 586622 294938 586858 295174
rect 586302 294618 586538 294854
rect 586622 294618 586858 294854
rect 586302 258938 586538 259174
rect 586622 258938 586858 259174
rect 586302 258618 586538 258854
rect 586622 258618 586858 258854
rect 586302 222938 586538 223174
rect 586622 222938 586858 223174
rect 586302 222618 586538 222854
rect 586622 222618 586858 222854
rect 586302 186938 586538 187174
rect 586622 186938 586858 187174
rect 586302 186618 586538 186854
rect 586622 186618 586858 186854
rect 586302 150938 586538 151174
rect 586622 150938 586858 151174
rect 586302 150618 586538 150854
rect 586622 150618 586858 150854
rect 586302 114938 586538 115174
rect 586622 114938 586858 115174
rect 586302 114618 586538 114854
rect 586622 114618 586858 114854
rect 586302 78938 586538 79174
rect 586622 78938 586858 79174
rect 586302 78618 586538 78854
rect 586622 78618 586858 78854
rect 586302 42938 586538 43174
rect 586622 42938 586858 43174
rect 586302 42618 586538 42854
rect 586622 42618 586858 42854
rect 586302 6938 586538 7174
rect 586622 6938 586858 7174
rect 586302 6618 586538 6854
rect 586622 6618 586858 6854
rect 581546 -1542 581782 -1306
rect 581866 -1542 582102 -1306
rect 581546 -1862 581782 -1626
rect 581866 -1862 582102 -1626
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 694658 587498 694894
rect 587582 694658 587818 694894
rect 587262 694338 587498 694574
rect 587582 694338 587818 694574
rect 587262 658658 587498 658894
rect 587582 658658 587818 658894
rect 587262 658338 587498 658574
rect 587582 658338 587818 658574
rect 587262 622658 587498 622894
rect 587582 622658 587818 622894
rect 587262 622338 587498 622574
rect 587582 622338 587818 622574
rect 587262 586658 587498 586894
rect 587582 586658 587818 586894
rect 587262 586338 587498 586574
rect 587582 586338 587818 586574
rect 587262 550658 587498 550894
rect 587582 550658 587818 550894
rect 587262 550338 587498 550574
rect 587582 550338 587818 550574
rect 587262 514658 587498 514894
rect 587582 514658 587818 514894
rect 587262 514338 587498 514574
rect 587582 514338 587818 514574
rect 587262 478658 587498 478894
rect 587582 478658 587818 478894
rect 587262 478338 587498 478574
rect 587582 478338 587818 478574
rect 587262 442658 587498 442894
rect 587582 442658 587818 442894
rect 587262 442338 587498 442574
rect 587582 442338 587818 442574
rect 587262 406658 587498 406894
rect 587582 406658 587818 406894
rect 587262 406338 587498 406574
rect 587582 406338 587818 406574
rect 587262 370658 587498 370894
rect 587582 370658 587818 370894
rect 587262 370338 587498 370574
rect 587582 370338 587818 370574
rect 587262 334658 587498 334894
rect 587582 334658 587818 334894
rect 587262 334338 587498 334574
rect 587582 334338 587818 334574
rect 587262 298658 587498 298894
rect 587582 298658 587818 298894
rect 587262 298338 587498 298574
rect 587582 298338 587818 298574
rect 587262 262658 587498 262894
rect 587582 262658 587818 262894
rect 587262 262338 587498 262574
rect 587582 262338 587818 262574
rect 587262 226658 587498 226894
rect 587582 226658 587818 226894
rect 587262 226338 587498 226574
rect 587582 226338 587818 226574
rect 587262 190658 587498 190894
rect 587582 190658 587818 190894
rect 587262 190338 587498 190574
rect 587582 190338 587818 190574
rect 587262 154658 587498 154894
rect 587582 154658 587818 154894
rect 587262 154338 587498 154574
rect 587582 154338 587818 154574
rect 587262 118658 587498 118894
rect 587582 118658 587818 118894
rect 587262 118338 587498 118574
rect 587582 118338 587818 118574
rect 587262 82658 587498 82894
rect 587582 82658 587818 82894
rect 587262 82338 587498 82574
rect 587582 82338 587818 82574
rect 587262 46658 587498 46894
rect 587582 46658 587818 46894
rect 587262 46338 587498 46574
rect 587582 46338 587818 46574
rect 587262 10658 587498 10894
rect 587582 10658 587818 10894
rect 587262 10338 587498 10574
rect 587582 10338 587818 10574
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 698378 588458 698614
rect 588542 698378 588778 698614
rect 588222 698058 588458 698294
rect 588542 698058 588778 698294
rect 588222 662378 588458 662614
rect 588542 662378 588778 662614
rect 588222 662058 588458 662294
rect 588542 662058 588778 662294
rect 588222 626378 588458 626614
rect 588542 626378 588778 626614
rect 588222 626058 588458 626294
rect 588542 626058 588778 626294
rect 588222 590378 588458 590614
rect 588542 590378 588778 590614
rect 588222 590058 588458 590294
rect 588542 590058 588778 590294
rect 588222 554378 588458 554614
rect 588542 554378 588778 554614
rect 588222 554058 588458 554294
rect 588542 554058 588778 554294
rect 588222 518378 588458 518614
rect 588542 518378 588778 518614
rect 588222 518058 588458 518294
rect 588542 518058 588778 518294
rect 588222 482378 588458 482614
rect 588542 482378 588778 482614
rect 588222 482058 588458 482294
rect 588542 482058 588778 482294
rect 588222 446378 588458 446614
rect 588542 446378 588778 446614
rect 588222 446058 588458 446294
rect 588542 446058 588778 446294
rect 588222 410378 588458 410614
rect 588542 410378 588778 410614
rect 588222 410058 588458 410294
rect 588542 410058 588778 410294
rect 588222 374378 588458 374614
rect 588542 374378 588778 374614
rect 588222 374058 588458 374294
rect 588542 374058 588778 374294
rect 588222 338378 588458 338614
rect 588542 338378 588778 338614
rect 588222 338058 588458 338294
rect 588542 338058 588778 338294
rect 588222 302378 588458 302614
rect 588542 302378 588778 302614
rect 588222 302058 588458 302294
rect 588542 302058 588778 302294
rect 588222 266378 588458 266614
rect 588542 266378 588778 266614
rect 588222 266058 588458 266294
rect 588542 266058 588778 266294
rect 588222 230378 588458 230614
rect 588542 230378 588778 230614
rect 588222 230058 588458 230294
rect 588542 230058 588778 230294
rect 588222 194378 588458 194614
rect 588542 194378 588778 194614
rect 588222 194058 588458 194294
rect 588542 194058 588778 194294
rect 588222 158378 588458 158614
rect 588542 158378 588778 158614
rect 588222 158058 588458 158294
rect 588542 158058 588778 158294
rect 588222 122378 588458 122614
rect 588542 122378 588778 122614
rect 588222 122058 588458 122294
rect 588542 122058 588778 122294
rect 588222 86378 588458 86614
rect 588542 86378 588778 86614
rect 588222 86058 588458 86294
rect 588542 86058 588778 86294
rect 588222 50378 588458 50614
rect 588542 50378 588778 50614
rect 588222 50058 588458 50294
rect 588542 50058 588778 50294
rect 588222 14378 588458 14614
rect 588542 14378 588778 14614
rect 588222 14058 588458 14294
rect 588542 14058 588778 14294
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 666098 589418 666334
rect 589502 666098 589738 666334
rect 589182 665778 589418 666014
rect 589502 665778 589738 666014
rect 589182 630098 589418 630334
rect 589502 630098 589738 630334
rect 589182 629778 589418 630014
rect 589502 629778 589738 630014
rect 589182 594098 589418 594334
rect 589502 594098 589738 594334
rect 589182 593778 589418 594014
rect 589502 593778 589738 594014
rect 589182 558098 589418 558334
rect 589502 558098 589738 558334
rect 589182 557778 589418 558014
rect 589502 557778 589738 558014
rect 589182 522098 589418 522334
rect 589502 522098 589738 522334
rect 589182 521778 589418 522014
rect 589502 521778 589738 522014
rect 589182 486098 589418 486334
rect 589502 486098 589738 486334
rect 589182 485778 589418 486014
rect 589502 485778 589738 486014
rect 589182 450098 589418 450334
rect 589502 450098 589738 450334
rect 589182 449778 589418 450014
rect 589502 449778 589738 450014
rect 589182 414098 589418 414334
rect 589502 414098 589738 414334
rect 589182 413778 589418 414014
rect 589502 413778 589738 414014
rect 589182 378098 589418 378334
rect 589502 378098 589738 378334
rect 589182 377778 589418 378014
rect 589502 377778 589738 378014
rect 589182 342098 589418 342334
rect 589502 342098 589738 342334
rect 589182 341778 589418 342014
rect 589502 341778 589738 342014
rect 589182 306098 589418 306334
rect 589502 306098 589738 306334
rect 589182 305778 589418 306014
rect 589502 305778 589738 306014
rect 589182 270098 589418 270334
rect 589502 270098 589738 270334
rect 589182 269778 589418 270014
rect 589502 269778 589738 270014
rect 589182 234098 589418 234334
rect 589502 234098 589738 234334
rect 589182 233778 589418 234014
rect 589502 233778 589738 234014
rect 589182 198098 589418 198334
rect 589502 198098 589738 198334
rect 589182 197778 589418 198014
rect 589502 197778 589738 198014
rect 589182 162098 589418 162334
rect 589502 162098 589738 162334
rect 589182 161778 589418 162014
rect 589502 161778 589738 162014
rect 589182 126098 589418 126334
rect 589502 126098 589738 126334
rect 589182 125778 589418 126014
rect 589502 125778 589738 126014
rect 589182 90098 589418 90334
rect 589502 90098 589738 90334
rect 589182 89778 589418 90014
rect 589502 89778 589738 90014
rect 589182 54098 589418 54334
rect 589502 54098 589738 54334
rect 589182 53778 589418 54014
rect 589502 53778 589738 54014
rect 589182 18098 589418 18334
rect 589502 18098 589738 18334
rect 589182 17778 589418 18014
rect 589502 17778 589738 18014
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 669818 590378 670054
rect 590462 669818 590698 670054
rect 590142 669498 590378 669734
rect 590462 669498 590698 669734
rect 590142 633818 590378 634054
rect 590462 633818 590698 634054
rect 590142 633498 590378 633734
rect 590462 633498 590698 633734
rect 590142 597818 590378 598054
rect 590462 597818 590698 598054
rect 590142 597498 590378 597734
rect 590462 597498 590698 597734
rect 590142 561818 590378 562054
rect 590462 561818 590698 562054
rect 590142 561498 590378 561734
rect 590462 561498 590698 561734
rect 590142 525818 590378 526054
rect 590462 525818 590698 526054
rect 590142 525498 590378 525734
rect 590462 525498 590698 525734
rect 590142 489818 590378 490054
rect 590462 489818 590698 490054
rect 590142 489498 590378 489734
rect 590462 489498 590698 489734
rect 590142 453818 590378 454054
rect 590462 453818 590698 454054
rect 590142 453498 590378 453734
rect 590462 453498 590698 453734
rect 590142 417818 590378 418054
rect 590462 417818 590698 418054
rect 590142 417498 590378 417734
rect 590462 417498 590698 417734
rect 590142 381818 590378 382054
rect 590462 381818 590698 382054
rect 590142 381498 590378 381734
rect 590462 381498 590698 381734
rect 590142 345818 590378 346054
rect 590462 345818 590698 346054
rect 590142 345498 590378 345734
rect 590462 345498 590698 345734
rect 590142 309818 590378 310054
rect 590462 309818 590698 310054
rect 590142 309498 590378 309734
rect 590462 309498 590698 309734
rect 590142 273818 590378 274054
rect 590462 273818 590698 274054
rect 590142 273498 590378 273734
rect 590462 273498 590698 273734
rect 590142 237818 590378 238054
rect 590462 237818 590698 238054
rect 590142 237498 590378 237734
rect 590462 237498 590698 237734
rect 590142 201818 590378 202054
rect 590462 201818 590698 202054
rect 590142 201498 590378 201734
rect 590462 201498 590698 201734
rect 590142 165818 590378 166054
rect 590462 165818 590698 166054
rect 590142 165498 590378 165734
rect 590462 165498 590698 165734
rect 590142 129818 590378 130054
rect 590462 129818 590698 130054
rect 590142 129498 590378 129734
rect 590462 129498 590698 129734
rect 590142 93818 590378 94054
rect 590462 93818 590698 94054
rect 590142 93498 590378 93734
rect 590462 93498 590698 93734
rect 590142 57818 590378 58054
rect 590462 57818 590698 58054
rect 590142 57498 590378 57734
rect 590462 57498 590698 57734
rect 590142 21818 590378 22054
rect 590462 21818 590698 22054
rect 590142 21498 590378 21734
rect 590462 21498 590698 21734
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 673538 591338 673774
rect 591422 673538 591658 673774
rect 591102 673218 591338 673454
rect 591422 673218 591658 673454
rect 591102 637538 591338 637774
rect 591422 637538 591658 637774
rect 591102 637218 591338 637454
rect 591422 637218 591658 637454
rect 591102 601538 591338 601774
rect 591422 601538 591658 601774
rect 591102 601218 591338 601454
rect 591422 601218 591658 601454
rect 591102 565538 591338 565774
rect 591422 565538 591658 565774
rect 591102 565218 591338 565454
rect 591422 565218 591658 565454
rect 591102 529538 591338 529774
rect 591422 529538 591658 529774
rect 591102 529218 591338 529454
rect 591422 529218 591658 529454
rect 591102 493538 591338 493774
rect 591422 493538 591658 493774
rect 591102 493218 591338 493454
rect 591422 493218 591658 493454
rect 591102 457538 591338 457774
rect 591422 457538 591658 457774
rect 591102 457218 591338 457454
rect 591422 457218 591658 457454
rect 591102 421538 591338 421774
rect 591422 421538 591658 421774
rect 591102 421218 591338 421454
rect 591422 421218 591658 421454
rect 591102 385538 591338 385774
rect 591422 385538 591658 385774
rect 591102 385218 591338 385454
rect 591422 385218 591658 385454
rect 591102 349538 591338 349774
rect 591422 349538 591658 349774
rect 591102 349218 591338 349454
rect 591422 349218 591658 349454
rect 591102 313538 591338 313774
rect 591422 313538 591658 313774
rect 591102 313218 591338 313454
rect 591422 313218 591658 313454
rect 591102 277538 591338 277774
rect 591422 277538 591658 277774
rect 591102 277218 591338 277454
rect 591422 277218 591658 277454
rect 591102 241538 591338 241774
rect 591422 241538 591658 241774
rect 591102 241218 591338 241454
rect 591422 241218 591658 241454
rect 591102 205538 591338 205774
rect 591422 205538 591658 205774
rect 591102 205218 591338 205454
rect 591422 205218 591658 205454
rect 591102 169538 591338 169774
rect 591422 169538 591658 169774
rect 591102 169218 591338 169454
rect 591422 169218 591658 169454
rect 591102 133538 591338 133774
rect 591422 133538 591658 133774
rect 591102 133218 591338 133454
rect 591422 133218 591658 133454
rect 591102 97538 591338 97774
rect 591422 97538 591658 97774
rect 591102 97218 591338 97454
rect 591422 97218 591658 97454
rect 591102 61538 591338 61774
rect 591422 61538 591658 61774
rect 591102 61218 591338 61454
rect 591422 61218 591658 61454
rect 591102 25538 591338 25774
rect 591422 25538 591658 25774
rect 591102 25218 591338 25454
rect 591422 25218 591658 25454
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 677258 592298 677494
rect 592382 677258 592618 677494
rect 592062 676938 592298 677174
rect 592382 676938 592618 677174
rect 592062 641258 592298 641494
rect 592382 641258 592618 641494
rect 592062 640938 592298 641174
rect 592382 640938 592618 641174
rect 592062 605258 592298 605494
rect 592382 605258 592618 605494
rect 592062 604938 592298 605174
rect 592382 604938 592618 605174
rect 592062 569258 592298 569494
rect 592382 569258 592618 569494
rect 592062 568938 592298 569174
rect 592382 568938 592618 569174
rect 592062 533258 592298 533494
rect 592382 533258 592618 533494
rect 592062 532938 592298 533174
rect 592382 532938 592618 533174
rect 592062 497258 592298 497494
rect 592382 497258 592618 497494
rect 592062 496938 592298 497174
rect 592382 496938 592618 497174
rect 592062 461258 592298 461494
rect 592382 461258 592618 461494
rect 592062 460938 592298 461174
rect 592382 460938 592618 461174
rect 592062 425258 592298 425494
rect 592382 425258 592618 425494
rect 592062 424938 592298 425174
rect 592382 424938 592618 425174
rect 592062 389258 592298 389494
rect 592382 389258 592618 389494
rect 592062 388938 592298 389174
rect 592382 388938 592618 389174
rect 592062 353258 592298 353494
rect 592382 353258 592618 353494
rect 592062 352938 592298 353174
rect 592382 352938 592618 353174
rect 592062 317258 592298 317494
rect 592382 317258 592618 317494
rect 592062 316938 592298 317174
rect 592382 316938 592618 317174
rect 592062 281258 592298 281494
rect 592382 281258 592618 281494
rect 592062 280938 592298 281174
rect 592382 280938 592618 281174
rect 592062 245258 592298 245494
rect 592382 245258 592618 245494
rect 592062 244938 592298 245174
rect 592382 244938 592618 245174
rect 592062 209258 592298 209494
rect 592382 209258 592618 209494
rect 592062 208938 592298 209174
rect 592382 208938 592618 209174
rect 592062 173258 592298 173494
rect 592382 173258 592618 173494
rect 592062 172938 592298 173174
rect 592382 172938 592618 173174
rect 592062 137258 592298 137494
rect 592382 137258 592618 137494
rect 592062 136938 592298 137174
rect 592382 136938 592618 137174
rect 592062 101258 592298 101494
rect 592382 101258 592618 101494
rect 592062 100938 592298 101174
rect 592382 100938 592618 101174
rect 592062 65258 592298 65494
rect 592382 65258 592618 65494
rect 592062 64938 592298 65174
rect 592382 64938 592618 65174
rect 592062 29258 592298 29494
rect 592382 29258 592618 29494
rect 592062 28938 592298 29174
rect 592382 28938 592618 29174
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 27866 711558
rect 28102 711322 28186 711558
rect 28422 711322 63866 711558
rect 64102 711322 64186 711558
rect 64422 711322 99866 711558
rect 100102 711322 100186 711558
rect 100422 711322 135866 711558
rect 136102 711322 136186 711558
rect 136422 711322 171866 711558
rect 172102 711322 172186 711558
rect 172422 711322 207866 711558
rect 208102 711322 208186 711558
rect 208422 711322 243866 711558
rect 244102 711322 244186 711558
rect 244422 711322 279866 711558
rect 280102 711322 280186 711558
rect 280422 711322 351866 711558
rect 352102 711322 352186 711558
rect 352422 711322 387866 711558
rect 388102 711322 388186 711558
rect 388422 711322 423866 711558
rect 424102 711322 424186 711558
rect 424422 711322 459866 711558
rect 460102 711322 460186 711558
rect 460422 711322 495866 711558
rect 496102 711322 496186 711558
rect 496422 711322 531866 711558
rect 532102 711322 532186 711558
rect 532422 711322 567866 711558
rect 568102 711322 568186 711558
rect 568422 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 27866 711238
rect 28102 711002 28186 711238
rect 28422 711002 63866 711238
rect 64102 711002 64186 711238
rect 64422 711002 99866 711238
rect 100102 711002 100186 711238
rect 100422 711002 135866 711238
rect 136102 711002 136186 711238
rect 136422 711002 171866 711238
rect 172102 711002 172186 711238
rect 172422 711002 207866 711238
rect 208102 711002 208186 711238
rect 208422 711002 243866 711238
rect 244102 711002 244186 711238
rect 244422 711002 279866 711238
rect 280102 711002 280186 711238
rect 280422 711002 351866 711238
rect 352102 711002 352186 711238
rect 352422 711002 387866 711238
rect 388102 711002 388186 711238
rect 388422 711002 423866 711238
rect 424102 711002 424186 711238
rect 424422 711002 459866 711238
rect 460102 711002 460186 711238
rect 460422 711002 495866 711238
rect 496102 711002 496186 711238
rect 496422 711002 531866 711238
rect 532102 711002 532186 711238
rect 532422 711002 567866 711238
rect 568102 711002 568186 711238
rect 568422 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 384146 710598
rect 384382 710362 384466 710598
rect 384702 710362 420146 710598
rect 420382 710362 420466 710598
rect 420702 710362 456146 710598
rect 456382 710362 456466 710598
rect 456702 710362 492146 710598
rect 492382 710362 492466 710598
rect 492702 710362 528146 710598
rect 528382 710362 528466 710598
rect 528702 710362 564146 710598
rect 564382 710362 564466 710598
rect 564702 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 384146 710278
rect 384382 710042 384466 710278
rect 384702 710042 420146 710278
rect 420382 710042 420466 710278
rect 420702 710042 456146 710278
rect 456382 710042 456466 710278
rect 456702 710042 492146 710278
rect 492382 710042 492466 710278
rect 492702 710042 528146 710278
rect 528382 710042 528466 710278
rect 528702 710042 564146 710278
rect 564382 710042 564466 710278
rect 564702 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 20426 709638
rect 20662 709402 20746 709638
rect 20982 709402 380426 709638
rect 380662 709402 380746 709638
rect 380982 709402 416426 709638
rect 416662 709402 416746 709638
rect 416982 709402 452426 709638
rect 452662 709402 452746 709638
rect 452982 709402 488426 709638
rect 488662 709402 488746 709638
rect 488982 709402 524426 709638
rect 524662 709402 524746 709638
rect 524982 709402 560426 709638
rect 560662 709402 560746 709638
rect 560982 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 20426 709318
rect 20662 709082 20746 709318
rect 20982 709082 380426 709318
rect 380662 709082 380746 709318
rect 380982 709082 416426 709318
rect 416662 709082 416746 709318
rect 416982 709082 452426 709318
rect 452662 709082 452746 709318
rect 452982 709082 488426 709318
rect 488662 709082 488746 709318
rect 488982 709082 524426 709318
rect 524662 709082 524746 709318
rect 524982 709082 560426 709318
rect 560662 709082 560746 709318
rect 560982 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 16706 708678
rect 16942 708442 17026 708678
rect 17262 708442 376706 708678
rect 376942 708442 377026 708678
rect 377262 708442 412706 708678
rect 412942 708442 413026 708678
rect 413262 708442 448706 708678
rect 448942 708442 449026 708678
rect 449262 708442 520706 708678
rect 520942 708442 521026 708678
rect 521262 708442 556706 708678
rect 556942 708442 557026 708678
rect 557262 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 16706 708358
rect 16942 708122 17026 708358
rect 17262 708122 376706 708358
rect 376942 708122 377026 708358
rect 377262 708122 412706 708358
rect 412942 708122 413026 708358
rect 413262 708122 448706 708358
rect 448942 708122 449026 708358
rect 449262 708122 520706 708358
rect 520942 708122 521026 708358
rect 521262 708122 556706 708358
rect 556942 708122 557026 708358
rect 557262 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 12986 707718
rect 13222 707482 13306 707718
rect 13542 707482 48986 707718
rect 49222 707482 49306 707718
rect 49542 707482 84986 707718
rect 85222 707482 85306 707718
rect 85542 707482 120986 707718
rect 121222 707482 121306 707718
rect 121542 707482 156986 707718
rect 157222 707482 157306 707718
rect 157542 707482 192986 707718
rect 193222 707482 193306 707718
rect 193542 707482 228986 707718
rect 229222 707482 229306 707718
rect 229542 707482 264986 707718
rect 265222 707482 265306 707718
rect 265542 707482 300986 707718
rect 301222 707482 301306 707718
rect 301542 707482 336986 707718
rect 337222 707482 337306 707718
rect 337542 707482 372986 707718
rect 373222 707482 373306 707718
rect 373542 707482 408986 707718
rect 409222 707482 409306 707718
rect 409542 707482 444986 707718
rect 445222 707482 445306 707718
rect 445542 707482 480986 707718
rect 481222 707482 481306 707718
rect 481542 707482 516986 707718
rect 517222 707482 517306 707718
rect 517542 707482 552986 707718
rect 553222 707482 553306 707718
rect 553542 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 12986 707398
rect 13222 707162 13306 707398
rect 13542 707162 48986 707398
rect 49222 707162 49306 707398
rect 49542 707162 84986 707398
rect 85222 707162 85306 707398
rect 85542 707162 120986 707398
rect 121222 707162 121306 707398
rect 121542 707162 156986 707398
rect 157222 707162 157306 707398
rect 157542 707162 192986 707398
rect 193222 707162 193306 707398
rect 193542 707162 228986 707398
rect 229222 707162 229306 707398
rect 229542 707162 264986 707398
rect 265222 707162 265306 707398
rect 265542 707162 300986 707398
rect 301222 707162 301306 707398
rect 301542 707162 336986 707398
rect 337222 707162 337306 707398
rect 337542 707162 372986 707398
rect 373222 707162 373306 707398
rect 373542 707162 408986 707398
rect 409222 707162 409306 707398
rect 409542 707162 444986 707398
rect 445222 707162 445306 707398
rect 445542 707162 480986 707398
rect 481222 707162 481306 707398
rect 481542 707162 516986 707398
rect 517222 707162 517306 707398
rect 517542 707162 552986 707398
rect 553222 707162 553306 707398
rect 553542 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 9266 706758
rect 9502 706522 9586 706758
rect 9822 706522 45266 706758
rect 45502 706522 45586 706758
rect 45822 706522 81266 706758
rect 81502 706522 81586 706758
rect 81822 706522 117266 706758
rect 117502 706522 117586 706758
rect 117822 706522 153266 706758
rect 153502 706522 153586 706758
rect 153822 706522 189266 706758
rect 189502 706522 189586 706758
rect 189822 706522 225266 706758
rect 225502 706522 225586 706758
rect 225822 706522 261266 706758
rect 261502 706522 261586 706758
rect 261822 706522 297266 706758
rect 297502 706522 297586 706758
rect 297822 706522 333266 706758
rect 333502 706522 333586 706758
rect 333822 706522 369266 706758
rect 369502 706522 369586 706758
rect 369822 706522 405266 706758
rect 405502 706522 405586 706758
rect 405822 706522 441266 706758
rect 441502 706522 441586 706758
rect 441822 706522 477266 706758
rect 477502 706522 477586 706758
rect 477822 706522 513266 706758
rect 513502 706522 513586 706758
rect 513822 706522 549266 706758
rect 549502 706522 549586 706758
rect 549822 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 9266 706438
rect 9502 706202 9586 706438
rect 9822 706202 45266 706438
rect 45502 706202 45586 706438
rect 45822 706202 81266 706438
rect 81502 706202 81586 706438
rect 81822 706202 117266 706438
rect 117502 706202 117586 706438
rect 117822 706202 153266 706438
rect 153502 706202 153586 706438
rect 153822 706202 189266 706438
rect 189502 706202 189586 706438
rect 189822 706202 225266 706438
rect 225502 706202 225586 706438
rect 225822 706202 261266 706438
rect 261502 706202 261586 706438
rect 261822 706202 297266 706438
rect 297502 706202 297586 706438
rect 297822 706202 333266 706438
rect 333502 706202 333586 706438
rect 333822 706202 369266 706438
rect 369502 706202 369586 706438
rect 369822 706202 405266 706438
rect 405502 706202 405586 706438
rect 405822 706202 441266 706438
rect 441502 706202 441586 706438
rect 441822 706202 477266 706438
rect 477502 706202 477586 706438
rect 477822 706202 513266 706438
rect 513502 706202 513586 706438
rect 513822 706202 549266 706438
rect 549502 706202 549586 706438
rect 549822 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 5546 705798
rect 5782 705562 5866 705798
rect 6102 705562 41546 705798
rect 41782 705562 41866 705798
rect 42102 705562 77546 705798
rect 77782 705562 77866 705798
rect 78102 705562 113546 705798
rect 113782 705562 113866 705798
rect 114102 705562 149546 705798
rect 149782 705562 149866 705798
rect 150102 705562 185546 705798
rect 185782 705562 185866 705798
rect 186102 705562 221546 705798
rect 221782 705562 221866 705798
rect 222102 705562 257546 705798
rect 257782 705562 257866 705798
rect 258102 705562 293546 705798
rect 293782 705562 293866 705798
rect 294102 705562 329546 705798
rect 329782 705562 329866 705798
rect 330102 705562 365546 705798
rect 365782 705562 365866 705798
rect 366102 705562 401546 705798
rect 401782 705562 401866 705798
rect 402102 705562 437546 705798
rect 437782 705562 437866 705798
rect 438102 705562 473546 705798
rect 473782 705562 473866 705798
rect 474102 705562 509546 705798
rect 509782 705562 509866 705798
rect 510102 705562 545546 705798
rect 545782 705562 545866 705798
rect 546102 705562 581546 705798
rect 581782 705562 581866 705798
rect 582102 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 5546 705478
rect 5782 705242 5866 705478
rect 6102 705242 41546 705478
rect 41782 705242 41866 705478
rect 42102 705242 77546 705478
rect 77782 705242 77866 705478
rect 78102 705242 113546 705478
rect 113782 705242 113866 705478
rect 114102 705242 149546 705478
rect 149782 705242 149866 705478
rect 150102 705242 185546 705478
rect 185782 705242 185866 705478
rect 186102 705242 221546 705478
rect 221782 705242 221866 705478
rect 222102 705242 257546 705478
rect 257782 705242 257866 705478
rect 258102 705242 293546 705478
rect 293782 705242 293866 705478
rect 294102 705242 329546 705478
rect 329782 705242 329866 705478
rect 330102 705242 365546 705478
rect 365782 705242 365866 705478
rect 366102 705242 401546 705478
rect 401782 705242 401866 705478
rect 402102 705242 437546 705478
rect 437782 705242 437866 705478
rect 438102 705242 473546 705478
rect 473782 705242 473866 705478
rect 474102 705242 509546 705478
rect 509782 705242 509866 705478
rect 510102 705242 545546 705478
rect 545782 705242 545866 705478
rect 546102 705242 581546 705478
rect 581782 705242 581866 705478
rect 582102 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 698614 592650 698646
rect -8726 698378 -4854 698614
rect -4618 698378 -4534 698614
rect -4298 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 588222 698614
rect 588458 698378 588542 698614
rect 588778 698378 592650 698614
rect -8726 698294 592650 698378
rect -8726 698058 -4854 698294
rect -4618 698058 -4534 698294
rect -4298 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 588222 698294
rect 588458 698058 588542 698294
rect 588778 698058 592650 698294
rect -8726 698026 592650 698058
rect -8726 694894 592650 694926
rect -8726 694658 -3894 694894
rect -3658 694658 -3574 694894
rect -3338 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 587262 694894
rect 587498 694658 587582 694894
rect 587818 694658 592650 694894
rect -8726 694574 592650 694658
rect -8726 694338 -3894 694574
rect -3658 694338 -3574 694574
rect -3338 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 587262 694574
rect 587498 694338 587582 694574
rect 587818 694338 592650 694574
rect -8726 694306 592650 694338
rect -8726 691174 592650 691206
rect -8726 690938 -2934 691174
rect -2698 690938 -2614 691174
rect -2378 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 586302 691174
rect 586538 690938 586622 691174
rect 586858 690938 592650 691174
rect -8726 690854 592650 690938
rect -8726 690618 -2934 690854
rect -2698 690618 -2614 690854
rect -2378 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 586302 690854
rect 586538 690618 586622 690854
rect 586858 690618 592650 690854
rect -8726 690586 592650 690618
rect -8726 687454 592650 687486
rect -8726 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 592650 687454
rect -8726 687134 592650 687218
rect -8726 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 592650 687134
rect -8726 686866 592650 686898
rect -8726 677494 592650 677526
rect -8726 677258 -8694 677494
rect -8458 677258 -8374 677494
rect -8138 677258 27866 677494
rect 28102 677258 28186 677494
rect 28422 677258 63866 677494
rect 64102 677258 64186 677494
rect 64422 677258 99866 677494
rect 100102 677258 100186 677494
rect 100422 677258 135866 677494
rect 136102 677258 136186 677494
rect 136422 677258 171866 677494
rect 172102 677258 172186 677494
rect 172422 677258 207866 677494
rect 208102 677258 208186 677494
rect 208422 677258 243866 677494
rect 244102 677258 244186 677494
rect 244422 677258 279866 677494
rect 280102 677258 280186 677494
rect 280422 677258 351866 677494
rect 352102 677258 352186 677494
rect 352422 677258 387866 677494
rect 388102 677258 388186 677494
rect 388422 677258 423866 677494
rect 424102 677258 424186 677494
rect 424422 677258 459866 677494
rect 460102 677258 460186 677494
rect 460422 677258 495866 677494
rect 496102 677258 496186 677494
rect 496422 677258 531866 677494
rect 532102 677258 532186 677494
rect 532422 677258 567866 677494
rect 568102 677258 568186 677494
rect 568422 677258 592062 677494
rect 592298 677258 592382 677494
rect 592618 677258 592650 677494
rect -8726 677174 592650 677258
rect -8726 676938 -8694 677174
rect -8458 676938 -8374 677174
rect -8138 676938 27866 677174
rect 28102 676938 28186 677174
rect 28422 676938 63866 677174
rect 64102 676938 64186 677174
rect 64422 676938 99866 677174
rect 100102 676938 100186 677174
rect 100422 676938 135866 677174
rect 136102 676938 136186 677174
rect 136422 676938 171866 677174
rect 172102 676938 172186 677174
rect 172422 676938 207866 677174
rect 208102 676938 208186 677174
rect 208422 676938 243866 677174
rect 244102 676938 244186 677174
rect 244422 676938 279866 677174
rect 280102 676938 280186 677174
rect 280422 676938 351866 677174
rect 352102 676938 352186 677174
rect 352422 676938 387866 677174
rect 388102 676938 388186 677174
rect 388422 676938 423866 677174
rect 424102 676938 424186 677174
rect 424422 676938 459866 677174
rect 460102 676938 460186 677174
rect 460422 676938 495866 677174
rect 496102 676938 496186 677174
rect 496422 676938 531866 677174
rect 532102 676938 532186 677174
rect 532422 676938 567866 677174
rect 568102 676938 568186 677174
rect 568422 676938 592062 677174
rect 592298 676938 592382 677174
rect 592618 676938 592650 677174
rect -8726 676906 592650 676938
rect -8726 673774 592650 673806
rect -8726 673538 -7734 673774
rect -7498 673538 -7414 673774
rect -7178 673538 384146 673774
rect 384382 673538 384466 673774
rect 384702 673538 420146 673774
rect 420382 673538 420466 673774
rect 420702 673538 456146 673774
rect 456382 673538 456466 673774
rect 456702 673538 492146 673774
rect 492382 673538 492466 673774
rect 492702 673538 528146 673774
rect 528382 673538 528466 673774
rect 528702 673538 564146 673774
rect 564382 673538 564466 673774
rect 564702 673538 591102 673774
rect 591338 673538 591422 673774
rect 591658 673538 592650 673774
rect -8726 673454 592650 673538
rect -8726 673218 -7734 673454
rect -7498 673218 -7414 673454
rect -7178 673218 384146 673454
rect 384382 673218 384466 673454
rect 384702 673218 420146 673454
rect 420382 673218 420466 673454
rect 420702 673218 456146 673454
rect 456382 673218 456466 673454
rect 456702 673218 492146 673454
rect 492382 673218 492466 673454
rect 492702 673218 528146 673454
rect 528382 673218 528466 673454
rect 528702 673218 564146 673454
rect 564382 673218 564466 673454
rect 564702 673218 591102 673454
rect 591338 673218 591422 673454
rect 591658 673218 592650 673454
rect -8726 673186 592650 673218
rect -8726 670054 592650 670086
rect -8726 669818 -6774 670054
rect -6538 669818 -6454 670054
rect -6218 669818 20426 670054
rect 20662 669818 20746 670054
rect 20982 669818 380426 670054
rect 380662 669818 380746 670054
rect 380982 669818 416426 670054
rect 416662 669818 416746 670054
rect 416982 669818 452426 670054
rect 452662 669818 452746 670054
rect 452982 669818 488426 670054
rect 488662 669818 488746 670054
rect 488982 669818 524426 670054
rect 524662 669818 524746 670054
rect 524982 669818 560426 670054
rect 560662 669818 560746 670054
rect 560982 669818 590142 670054
rect 590378 669818 590462 670054
rect 590698 669818 592650 670054
rect -8726 669734 592650 669818
rect -8726 669498 -6774 669734
rect -6538 669498 -6454 669734
rect -6218 669498 20426 669734
rect 20662 669498 20746 669734
rect 20982 669498 380426 669734
rect 380662 669498 380746 669734
rect 380982 669498 416426 669734
rect 416662 669498 416746 669734
rect 416982 669498 452426 669734
rect 452662 669498 452746 669734
rect 452982 669498 488426 669734
rect 488662 669498 488746 669734
rect 488982 669498 524426 669734
rect 524662 669498 524746 669734
rect 524982 669498 560426 669734
rect 560662 669498 560746 669734
rect 560982 669498 590142 669734
rect 590378 669498 590462 669734
rect 590698 669498 592650 669734
rect -8726 669466 592650 669498
rect -8726 666334 592650 666366
rect -8726 666098 -5814 666334
rect -5578 666098 -5494 666334
rect -5258 666098 16706 666334
rect 16942 666098 17026 666334
rect 17262 666098 376706 666334
rect 376942 666098 377026 666334
rect 377262 666098 412706 666334
rect 412942 666098 413026 666334
rect 413262 666098 448706 666334
rect 448942 666098 449026 666334
rect 449262 666098 520706 666334
rect 520942 666098 521026 666334
rect 521262 666098 556706 666334
rect 556942 666098 557026 666334
rect 557262 666098 589182 666334
rect 589418 666098 589502 666334
rect 589738 666098 592650 666334
rect -8726 666014 592650 666098
rect -8726 665778 -5814 666014
rect -5578 665778 -5494 666014
rect -5258 665778 16706 666014
rect 16942 665778 17026 666014
rect 17262 665778 376706 666014
rect 376942 665778 377026 666014
rect 377262 665778 412706 666014
rect 412942 665778 413026 666014
rect 413262 665778 448706 666014
rect 448942 665778 449026 666014
rect 449262 665778 520706 666014
rect 520942 665778 521026 666014
rect 521262 665778 556706 666014
rect 556942 665778 557026 666014
rect 557262 665778 589182 666014
rect 589418 665778 589502 666014
rect 589738 665778 592650 666014
rect -8726 665746 592650 665778
rect -8726 662614 592650 662646
rect -8726 662378 -4854 662614
rect -4618 662378 -4534 662614
rect -4298 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 588222 662614
rect 588458 662378 588542 662614
rect 588778 662378 592650 662614
rect -8726 662294 592650 662378
rect -8726 662058 -4854 662294
rect -4618 662058 -4534 662294
rect -4298 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 588222 662294
rect 588458 662058 588542 662294
rect 588778 662058 592650 662294
rect -8726 662026 592650 662058
rect -8726 658894 592650 658926
rect -8726 658658 -3894 658894
rect -3658 658658 -3574 658894
rect -3338 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 587262 658894
rect 587498 658658 587582 658894
rect 587818 658658 592650 658894
rect -8726 658574 592650 658658
rect -8726 658338 -3894 658574
rect -3658 658338 -3574 658574
rect -3338 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 587262 658574
rect 587498 658338 587582 658574
rect 587818 658338 592650 658574
rect -8726 658306 592650 658338
rect -8726 655174 592650 655206
rect -8726 654938 -2934 655174
rect -2698 654938 -2614 655174
rect -2378 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 39610 655174
rect 39846 654938 70330 655174
rect 70566 654938 101050 655174
rect 101286 654938 131770 655174
rect 132006 654938 162490 655174
rect 162726 654938 193210 655174
rect 193446 654938 223930 655174
rect 224166 654938 254650 655174
rect 254886 654938 285370 655174
rect 285606 654938 316090 655174
rect 316326 654938 346810 655174
rect 347046 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 479610 655174
rect 479846 654938 510330 655174
rect 510566 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 586302 655174
rect 586538 654938 586622 655174
rect 586858 654938 592650 655174
rect -8726 654854 592650 654938
rect -8726 654618 -2934 654854
rect -2698 654618 -2614 654854
rect -2378 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 39610 654854
rect 39846 654618 70330 654854
rect 70566 654618 101050 654854
rect 101286 654618 131770 654854
rect 132006 654618 162490 654854
rect 162726 654618 193210 654854
rect 193446 654618 223930 654854
rect 224166 654618 254650 654854
rect 254886 654618 285370 654854
rect 285606 654618 316090 654854
rect 316326 654618 346810 654854
rect 347046 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 479610 654854
rect 479846 654618 510330 654854
rect 510566 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 586302 654854
rect 586538 654618 586622 654854
rect 586858 654618 592650 654854
rect -8726 654586 592650 654618
rect -8726 651454 592650 651486
rect -8726 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 24250 651454
rect 24486 651218 54970 651454
rect 55206 651218 85690 651454
rect 85926 651218 116410 651454
rect 116646 651218 147130 651454
rect 147366 651218 177850 651454
rect 178086 651218 208570 651454
rect 208806 651218 239290 651454
rect 239526 651218 270010 651454
rect 270246 651218 300730 651454
rect 300966 651218 331450 651454
rect 331686 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 464250 651454
rect 464486 651218 494970 651454
rect 495206 651218 525690 651454
rect 525926 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 592650 651454
rect -8726 651134 592650 651218
rect -8726 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 24250 651134
rect 24486 650898 54970 651134
rect 55206 650898 85690 651134
rect 85926 650898 116410 651134
rect 116646 650898 147130 651134
rect 147366 650898 177850 651134
rect 178086 650898 208570 651134
rect 208806 650898 239290 651134
rect 239526 650898 270010 651134
rect 270246 650898 300730 651134
rect 300966 650898 331450 651134
rect 331686 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 464250 651134
rect 464486 650898 494970 651134
rect 495206 650898 525690 651134
rect 525926 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 592650 651134
rect -8726 650866 592650 650898
rect -8726 641494 592650 641526
rect -8726 641258 -8694 641494
rect -8458 641258 -8374 641494
rect -8138 641258 27866 641494
rect 28102 641258 28186 641494
rect 28422 641258 387866 641494
rect 388102 641258 388186 641494
rect 388422 641258 423866 641494
rect 424102 641258 424186 641494
rect 424422 641258 531866 641494
rect 532102 641258 532186 641494
rect 532422 641258 567866 641494
rect 568102 641258 568186 641494
rect 568422 641258 592062 641494
rect 592298 641258 592382 641494
rect 592618 641258 592650 641494
rect -8726 641174 592650 641258
rect -8726 640938 -8694 641174
rect -8458 640938 -8374 641174
rect -8138 640938 27866 641174
rect 28102 640938 28186 641174
rect 28422 640938 387866 641174
rect 388102 640938 388186 641174
rect 388422 640938 423866 641174
rect 424102 640938 424186 641174
rect 424422 640938 531866 641174
rect 532102 640938 532186 641174
rect 532422 640938 567866 641174
rect 568102 640938 568186 641174
rect 568422 640938 592062 641174
rect 592298 640938 592382 641174
rect 592618 640938 592650 641174
rect -8726 640906 592650 640938
rect -8726 637774 592650 637806
rect -8726 637538 -7734 637774
rect -7498 637538 -7414 637774
rect -7178 637538 384146 637774
rect 384382 637538 384466 637774
rect 384702 637538 420146 637774
rect 420382 637538 420466 637774
rect 420702 637538 456146 637774
rect 456382 637538 456466 637774
rect 456702 637538 528146 637774
rect 528382 637538 528466 637774
rect 528702 637538 564146 637774
rect 564382 637538 564466 637774
rect 564702 637538 591102 637774
rect 591338 637538 591422 637774
rect 591658 637538 592650 637774
rect -8726 637454 592650 637538
rect -8726 637218 -7734 637454
rect -7498 637218 -7414 637454
rect -7178 637218 384146 637454
rect 384382 637218 384466 637454
rect 384702 637218 420146 637454
rect 420382 637218 420466 637454
rect 420702 637218 456146 637454
rect 456382 637218 456466 637454
rect 456702 637218 528146 637454
rect 528382 637218 528466 637454
rect 528702 637218 564146 637454
rect 564382 637218 564466 637454
rect 564702 637218 591102 637454
rect 591338 637218 591422 637454
rect 591658 637218 592650 637454
rect -8726 637186 592650 637218
rect -8726 634054 592650 634086
rect -8726 633818 -6774 634054
rect -6538 633818 -6454 634054
rect -6218 633818 20426 634054
rect 20662 633818 20746 634054
rect 20982 633818 380426 634054
rect 380662 633818 380746 634054
rect 380982 633818 416426 634054
rect 416662 633818 416746 634054
rect 416982 633818 452426 634054
rect 452662 633818 452746 634054
rect 452982 633818 524426 634054
rect 524662 633818 524746 634054
rect 524982 633818 560426 634054
rect 560662 633818 560746 634054
rect 560982 633818 590142 634054
rect 590378 633818 590462 634054
rect 590698 633818 592650 634054
rect -8726 633734 592650 633818
rect -8726 633498 -6774 633734
rect -6538 633498 -6454 633734
rect -6218 633498 20426 633734
rect 20662 633498 20746 633734
rect 20982 633498 380426 633734
rect 380662 633498 380746 633734
rect 380982 633498 416426 633734
rect 416662 633498 416746 633734
rect 416982 633498 452426 633734
rect 452662 633498 452746 633734
rect 452982 633498 524426 633734
rect 524662 633498 524746 633734
rect 524982 633498 560426 633734
rect 560662 633498 560746 633734
rect 560982 633498 590142 633734
rect 590378 633498 590462 633734
rect 590698 633498 592650 633734
rect -8726 633466 592650 633498
rect -8726 630334 592650 630366
rect -8726 630098 -5814 630334
rect -5578 630098 -5494 630334
rect -5258 630098 16706 630334
rect 16942 630098 17026 630334
rect 17262 630098 376706 630334
rect 376942 630098 377026 630334
rect 377262 630098 412706 630334
rect 412942 630098 413026 630334
rect 413262 630098 448706 630334
rect 448942 630098 449026 630334
rect 449262 630098 520706 630334
rect 520942 630098 521026 630334
rect 521262 630098 556706 630334
rect 556942 630098 557026 630334
rect 557262 630098 589182 630334
rect 589418 630098 589502 630334
rect 589738 630098 592650 630334
rect -8726 630014 592650 630098
rect -8726 629778 -5814 630014
rect -5578 629778 -5494 630014
rect -5258 629778 16706 630014
rect 16942 629778 17026 630014
rect 17262 629778 376706 630014
rect 376942 629778 377026 630014
rect 377262 629778 412706 630014
rect 412942 629778 413026 630014
rect 413262 629778 448706 630014
rect 448942 629778 449026 630014
rect 449262 629778 520706 630014
rect 520942 629778 521026 630014
rect 521262 629778 556706 630014
rect 556942 629778 557026 630014
rect 557262 629778 589182 630014
rect 589418 629778 589502 630014
rect 589738 629778 592650 630014
rect -8726 629746 592650 629778
rect -8726 626614 592650 626646
rect -8726 626378 -4854 626614
rect -4618 626378 -4534 626614
rect -4298 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 372986 626614
rect 373222 626378 373306 626614
rect 373542 626378 408986 626614
rect 409222 626378 409306 626614
rect 409542 626378 444986 626614
rect 445222 626378 445306 626614
rect 445542 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 588222 626614
rect 588458 626378 588542 626614
rect 588778 626378 592650 626614
rect -8726 626294 592650 626378
rect -8726 626058 -4854 626294
rect -4618 626058 -4534 626294
rect -4298 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 372986 626294
rect 373222 626058 373306 626294
rect 373542 626058 408986 626294
rect 409222 626058 409306 626294
rect 409542 626058 444986 626294
rect 445222 626058 445306 626294
rect 445542 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 588222 626294
rect 588458 626058 588542 626294
rect 588778 626058 592650 626294
rect -8726 626026 592650 626058
rect -8726 622894 592650 622926
rect -8726 622658 -3894 622894
rect -3658 622658 -3574 622894
rect -3338 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 369266 622894
rect 369502 622658 369586 622894
rect 369822 622658 405266 622894
rect 405502 622658 405586 622894
rect 405822 622658 441266 622894
rect 441502 622658 441586 622894
rect 441822 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 587262 622894
rect 587498 622658 587582 622894
rect 587818 622658 592650 622894
rect -8726 622574 592650 622658
rect -8726 622338 -3894 622574
rect -3658 622338 -3574 622574
rect -3338 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 369266 622574
rect 369502 622338 369586 622574
rect 369822 622338 405266 622574
rect 405502 622338 405586 622574
rect 405822 622338 441266 622574
rect 441502 622338 441586 622574
rect 441822 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 587262 622574
rect 587498 622338 587582 622574
rect 587818 622338 592650 622574
rect -8726 622306 592650 622338
rect -8726 619174 592650 619206
rect -8726 618938 -2934 619174
rect -2698 618938 -2614 619174
rect -2378 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 39610 619174
rect 39846 618938 70330 619174
rect 70566 618938 101050 619174
rect 101286 618938 131770 619174
rect 132006 618938 162490 619174
rect 162726 618938 193210 619174
rect 193446 618938 223930 619174
rect 224166 618938 254650 619174
rect 254886 618938 285370 619174
rect 285606 618938 316090 619174
rect 316326 618938 346810 619174
rect 347046 618938 365546 619174
rect 365782 618938 365866 619174
rect 366102 618938 401546 619174
rect 401782 618938 401866 619174
rect 402102 618938 437546 619174
rect 437782 618938 437866 619174
rect 438102 618938 479610 619174
rect 479846 618938 510330 619174
rect 510566 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 586302 619174
rect 586538 618938 586622 619174
rect 586858 618938 592650 619174
rect -8726 618854 592650 618938
rect -8726 618618 -2934 618854
rect -2698 618618 -2614 618854
rect -2378 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 39610 618854
rect 39846 618618 70330 618854
rect 70566 618618 101050 618854
rect 101286 618618 131770 618854
rect 132006 618618 162490 618854
rect 162726 618618 193210 618854
rect 193446 618618 223930 618854
rect 224166 618618 254650 618854
rect 254886 618618 285370 618854
rect 285606 618618 316090 618854
rect 316326 618618 346810 618854
rect 347046 618618 365546 618854
rect 365782 618618 365866 618854
rect 366102 618618 401546 618854
rect 401782 618618 401866 618854
rect 402102 618618 437546 618854
rect 437782 618618 437866 618854
rect 438102 618618 479610 618854
rect 479846 618618 510330 618854
rect 510566 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 586302 618854
rect 586538 618618 586622 618854
rect 586858 618618 592650 618854
rect -8726 618586 592650 618618
rect -8726 615454 592650 615486
rect -8726 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 24250 615454
rect 24486 615218 54970 615454
rect 55206 615218 85690 615454
rect 85926 615218 116410 615454
rect 116646 615218 147130 615454
rect 147366 615218 177850 615454
rect 178086 615218 208570 615454
rect 208806 615218 239290 615454
rect 239526 615218 270010 615454
rect 270246 615218 300730 615454
rect 300966 615218 331450 615454
rect 331686 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 464250 615454
rect 464486 615218 494970 615454
rect 495206 615218 525690 615454
rect 525926 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 592650 615454
rect -8726 615134 592650 615218
rect -8726 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 24250 615134
rect 24486 614898 54970 615134
rect 55206 614898 85690 615134
rect 85926 614898 116410 615134
rect 116646 614898 147130 615134
rect 147366 614898 177850 615134
rect 178086 614898 208570 615134
rect 208806 614898 239290 615134
rect 239526 614898 270010 615134
rect 270246 614898 300730 615134
rect 300966 614898 331450 615134
rect 331686 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 464250 615134
rect 464486 614898 494970 615134
rect 495206 614898 525690 615134
rect 525926 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 592650 615134
rect -8726 614866 592650 614898
rect -8726 605494 592650 605526
rect -8726 605258 -8694 605494
rect -8458 605258 -8374 605494
rect -8138 605258 27866 605494
rect 28102 605258 28186 605494
rect 28422 605258 387866 605494
rect 388102 605258 388186 605494
rect 388422 605258 423866 605494
rect 424102 605258 424186 605494
rect 424422 605258 531866 605494
rect 532102 605258 532186 605494
rect 532422 605258 567866 605494
rect 568102 605258 568186 605494
rect 568422 605258 592062 605494
rect 592298 605258 592382 605494
rect 592618 605258 592650 605494
rect -8726 605174 592650 605258
rect -8726 604938 -8694 605174
rect -8458 604938 -8374 605174
rect -8138 604938 27866 605174
rect 28102 604938 28186 605174
rect 28422 604938 387866 605174
rect 388102 604938 388186 605174
rect 388422 604938 423866 605174
rect 424102 604938 424186 605174
rect 424422 604938 531866 605174
rect 532102 604938 532186 605174
rect 532422 604938 567866 605174
rect 568102 604938 568186 605174
rect 568422 604938 592062 605174
rect 592298 604938 592382 605174
rect 592618 604938 592650 605174
rect -8726 604906 592650 604938
rect -8726 601774 592650 601806
rect -8726 601538 -7734 601774
rect -7498 601538 -7414 601774
rect -7178 601538 384146 601774
rect 384382 601538 384466 601774
rect 384702 601538 420146 601774
rect 420382 601538 420466 601774
rect 420702 601538 456146 601774
rect 456382 601538 456466 601774
rect 456702 601538 528146 601774
rect 528382 601538 528466 601774
rect 528702 601538 564146 601774
rect 564382 601538 564466 601774
rect 564702 601538 591102 601774
rect 591338 601538 591422 601774
rect 591658 601538 592650 601774
rect -8726 601454 592650 601538
rect -8726 601218 -7734 601454
rect -7498 601218 -7414 601454
rect -7178 601218 384146 601454
rect 384382 601218 384466 601454
rect 384702 601218 420146 601454
rect 420382 601218 420466 601454
rect 420702 601218 456146 601454
rect 456382 601218 456466 601454
rect 456702 601218 528146 601454
rect 528382 601218 528466 601454
rect 528702 601218 564146 601454
rect 564382 601218 564466 601454
rect 564702 601218 591102 601454
rect 591338 601218 591422 601454
rect 591658 601218 592650 601454
rect -8726 601186 592650 601218
rect -8726 598054 592650 598086
rect -8726 597818 -6774 598054
rect -6538 597818 -6454 598054
rect -6218 597818 20426 598054
rect 20662 597818 20746 598054
rect 20982 597818 380426 598054
rect 380662 597818 380746 598054
rect 380982 597818 416426 598054
rect 416662 597818 416746 598054
rect 416982 597818 452426 598054
rect 452662 597818 452746 598054
rect 452982 597818 488426 598054
rect 488662 597818 488746 598054
rect 488982 597818 524426 598054
rect 524662 597818 524746 598054
rect 524982 597818 560426 598054
rect 560662 597818 560746 598054
rect 560982 597818 590142 598054
rect 590378 597818 590462 598054
rect 590698 597818 592650 598054
rect -8726 597734 592650 597818
rect -8726 597498 -6774 597734
rect -6538 597498 -6454 597734
rect -6218 597498 20426 597734
rect 20662 597498 20746 597734
rect 20982 597498 380426 597734
rect 380662 597498 380746 597734
rect 380982 597498 416426 597734
rect 416662 597498 416746 597734
rect 416982 597498 452426 597734
rect 452662 597498 452746 597734
rect 452982 597498 488426 597734
rect 488662 597498 488746 597734
rect 488982 597498 524426 597734
rect 524662 597498 524746 597734
rect 524982 597498 560426 597734
rect 560662 597498 560746 597734
rect 560982 597498 590142 597734
rect 590378 597498 590462 597734
rect 590698 597498 592650 597734
rect -8726 597466 592650 597498
rect -8726 594334 592650 594366
rect -8726 594098 -5814 594334
rect -5578 594098 -5494 594334
rect -5258 594098 16706 594334
rect 16942 594098 17026 594334
rect 17262 594098 376706 594334
rect 376942 594098 377026 594334
rect 377262 594098 412706 594334
rect 412942 594098 413026 594334
rect 413262 594098 448706 594334
rect 448942 594098 449026 594334
rect 449262 594098 484706 594334
rect 484942 594098 485026 594334
rect 485262 594098 520706 594334
rect 520942 594098 521026 594334
rect 521262 594098 556706 594334
rect 556942 594098 557026 594334
rect 557262 594098 589182 594334
rect 589418 594098 589502 594334
rect 589738 594098 592650 594334
rect -8726 594014 592650 594098
rect -8726 593778 -5814 594014
rect -5578 593778 -5494 594014
rect -5258 593778 16706 594014
rect 16942 593778 17026 594014
rect 17262 593778 376706 594014
rect 376942 593778 377026 594014
rect 377262 593778 412706 594014
rect 412942 593778 413026 594014
rect 413262 593778 448706 594014
rect 448942 593778 449026 594014
rect 449262 593778 484706 594014
rect 484942 593778 485026 594014
rect 485262 593778 520706 594014
rect 520942 593778 521026 594014
rect 521262 593778 556706 594014
rect 556942 593778 557026 594014
rect 557262 593778 589182 594014
rect 589418 593778 589502 594014
rect 589738 593778 592650 594014
rect -8726 593746 592650 593778
rect -8726 590614 592650 590646
rect -8726 590378 -4854 590614
rect -4618 590378 -4534 590614
rect -4298 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 372986 590614
rect 373222 590378 373306 590614
rect 373542 590378 408986 590614
rect 409222 590378 409306 590614
rect 409542 590378 444986 590614
rect 445222 590378 445306 590614
rect 445542 590378 480986 590614
rect 481222 590378 481306 590614
rect 481542 590378 516986 590614
rect 517222 590378 517306 590614
rect 517542 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 588222 590614
rect 588458 590378 588542 590614
rect 588778 590378 592650 590614
rect -8726 590294 592650 590378
rect -8726 590058 -4854 590294
rect -4618 590058 -4534 590294
rect -4298 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 372986 590294
rect 373222 590058 373306 590294
rect 373542 590058 408986 590294
rect 409222 590058 409306 590294
rect 409542 590058 444986 590294
rect 445222 590058 445306 590294
rect 445542 590058 480986 590294
rect 481222 590058 481306 590294
rect 481542 590058 516986 590294
rect 517222 590058 517306 590294
rect 517542 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 588222 590294
rect 588458 590058 588542 590294
rect 588778 590058 592650 590294
rect -8726 590026 592650 590058
rect -8726 586894 592650 586926
rect -8726 586658 -3894 586894
rect -3658 586658 -3574 586894
rect -3338 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 369266 586894
rect 369502 586658 369586 586894
rect 369822 586658 405266 586894
rect 405502 586658 405586 586894
rect 405822 586658 441266 586894
rect 441502 586658 441586 586894
rect 441822 586658 477266 586894
rect 477502 586658 477586 586894
rect 477822 586658 513266 586894
rect 513502 586658 513586 586894
rect 513822 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 587262 586894
rect 587498 586658 587582 586894
rect 587818 586658 592650 586894
rect -8726 586574 592650 586658
rect -8726 586338 -3894 586574
rect -3658 586338 -3574 586574
rect -3338 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 369266 586574
rect 369502 586338 369586 586574
rect 369822 586338 405266 586574
rect 405502 586338 405586 586574
rect 405822 586338 441266 586574
rect 441502 586338 441586 586574
rect 441822 586338 477266 586574
rect 477502 586338 477586 586574
rect 477822 586338 513266 586574
rect 513502 586338 513586 586574
rect 513822 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 587262 586574
rect 587498 586338 587582 586574
rect 587818 586338 592650 586574
rect -8726 586306 592650 586338
rect -8726 583174 592650 583206
rect -8726 582938 -2934 583174
rect -2698 582938 -2614 583174
rect -2378 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 39610 583174
rect 39846 582938 70330 583174
rect 70566 582938 101050 583174
rect 101286 582938 131770 583174
rect 132006 582938 162490 583174
rect 162726 582938 193210 583174
rect 193446 582938 223930 583174
rect 224166 582938 254650 583174
rect 254886 582938 285370 583174
rect 285606 582938 316090 583174
rect 316326 582938 346810 583174
rect 347046 582938 365546 583174
rect 365782 582938 365866 583174
rect 366102 582938 401546 583174
rect 401782 582938 401866 583174
rect 402102 582938 437546 583174
rect 437782 582938 437866 583174
rect 438102 582938 473546 583174
rect 473782 582938 473866 583174
rect 474102 582938 509546 583174
rect 509782 582938 509866 583174
rect 510102 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 586302 583174
rect 586538 582938 586622 583174
rect 586858 582938 592650 583174
rect -8726 582854 592650 582938
rect -8726 582618 -2934 582854
rect -2698 582618 -2614 582854
rect -2378 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 39610 582854
rect 39846 582618 70330 582854
rect 70566 582618 101050 582854
rect 101286 582618 131770 582854
rect 132006 582618 162490 582854
rect 162726 582618 193210 582854
rect 193446 582618 223930 582854
rect 224166 582618 254650 582854
rect 254886 582618 285370 582854
rect 285606 582618 316090 582854
rect 316326 582618 346810 582854
rect 347046 582618 365546 582854
rect 365782 582618 365866 582854
rect 366102 582618 401546 582854
rect 401782 582618 401866 582854
rect 402102 582618 437546 582854
rect 437782 582618 437866 582854
rect 438102 582618 473546 582854
rect 473782 582618 473866 582854
rect 474102 582618 509546 582854
rect 509782 582618 509866 582854
rect 510102 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 586302 582854
rect 586538 582618 586622 582854
rect 586858 582618 592650 582854
rect -8726 582586 592650 582618
rect -8726 579454 592650 579486
rect -8726 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 24250 579454
rect 24486 579218 54970 579454
rect 55206 579218 85690 579454
rect 85926 579218 116410 579454
rect 116646 579218 147130 579454
rect 147366 579218 177850 579454
rect 178086 579218 208570 579454
rect 208806 579218 239290 579454
rect 239526 579218 270010 579454
rect 270246 579218 300730 579454
rect 300966 579218 331450 579454
rect 331686 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 592650 579454
rect -8726 579134 592650 579218
rect -8726 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 24250 579134
rect 24486 578898 54970 579134
rect 55206 578898 85690 579134
rect 85926 578898 116410 579134
rect 116646 578898 147130 579134
rect 147366 578898 177850 579134
rect 178086 578898 208570 579134
rect 208806 578898 239290 579134
rect 239526 578898 270010 579134
rect 270246 578898 300730 579134
rect 300966 578898 331450 579134
rect 331686 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 592650 579134
rect -8726 578866 592650 578898
rect -8726 569494 592650 569526
rect -8726 569258 -8694 569494
rect -8458 569258 -8374 569494
rect -8138 569258 27866 569494
rect 28102 569258 28186 569494
rect 28422 569258 387866 569494
rect 388102 569258 388186 569494
rect 388422 569258 423866 569494
rect 424102 569258 424186 569494
rect 424422 569258 459866 569494
rect 460102 569258 460186 569494
rect 460422 569258 495866 569494
rect 496102 569258 496186 569494
rect 496422 569258 531866 569494
rect 532102 569258 532186 569494
rect 532422 569258 567866 569494
rect 568102 569258 568186 569494
rect 568422 569258 592062 569494
rect 592298 569258 592382 569494
rect 592618 569258 592650 569494
rect -8726 569174 592650 569258
rect -8726 568938 -8694 569174
rect -8458 568938 -8374 569174
rect -8138 568938 27866 569174
rect 28102 568938 28186 569174
rect 28422 568938 387866 569174
rect 388102 568938 388186 569174
rect 388422 568938 423866 569174
rect 424102 568938 424186 569174
rect 424422 568938 459866 569174
rect 460102 568938 460186 569174
rect 460422 568938 495866 569174
rect 496102 568938 496186 569174
rect 496422 568938 531866 569174
rect 532102 568938 532186 569174
rect 532422 568938 567866 569174
rect 568102 568938 568186 569174
rect 568422 568938 592062 569174
rect 592298 568938 592382 569174
rect 592618 568938 592650 569174
rect -8726 568906 592650 568938
rect -8726 565774 592650 565806
rect -8726 565538 -7734 565774
rect -7498 565538 -7414 565774
rect -7178 565538 384146 565774
rect 384382 565538 384466 565774
rect 384702 565538 420146 565774
rect 420382 565538 420466 565774
rect 420702 565538 456146 565774
rect 456382 565538 456466 565774
rect 456702 565538 492146 565774
rect 492382 565538 492466 565774
rect 492702 565538 528146 565774
rect 528382 565538 528466 565774
rect 528702 565538 564146 565774
rect 564382 565538 564466 565774
rect 564702 565538 591102 565774
rect 591338 565538 591422 565774
rect 591658 565538 592650 565774
rect -8726 565454 592650 565538
rect -8726 565218 -7734 565454
rect -7498 565218 -7414 565454
rect -7178 565218 384146 565454
rect 384382 565218 384466 565454
rect 384702 565218 420146 565454
rect 420382 565218 420466 565454
rect 420702 565218 456146 565454
rect 456382 565218 456466 565454
rect 456702 565218 492146 565454
rect 492382 565218 492466 565454
rect 492702 565218 528146 565454
rect 528382 565218 528466 565454
rect 528702 565218 564146 565454
rect 564382 565218 564466 565454
rect 564702 565218 591102 565454
rect 591338 565218 591422 565454
rect 591658 565218 592650 565454
rect -8726 565186 592650 565218
rect -8726 562054 592650 562086
rect -8726 561818 -6774 562054
rect -6538 561818 -6454 562054
rect -6218 561818 20426 562054
rect 20662 561818 20746 562054
rect 20982 561818 380426 562054
rect 380662 561818 380746 562054
rect 380982 561818 416426 562054
rect 416662 561818 416746 562054
rect 416982 561818 452426 562054
rect 452662 561818 452746 562054
rect 452982 561818 488426 562054
rect 488662 561818 488746 562054
rect 488982 561818 524426 562054
rect 524662 561818 524746 562054
rect 524982 561818 560426 562054
rect 560662 561818 560746 562054
rect 560982 561818 590142 562054
rect 590378 561818 590462 562054
rect 590698 561818 592650 562054
rect -8726 561734 592650 561818
rect -8726 561498 -6774 561734
rect -6538 561498 -6454 561734
rect -6218 561498 20426 561734
rect 20662 561498 20746 561734
rect 20982 561498 380426 561734
rect 380662 561498 380746 561734
rect 380982 561498 416426 561734
rect 416662 561498 416746 561734
rect 416982 561498 452426 561734
rect 452662 561498 452746 561734
rect 452982 561498 488426 561734
rect 488662 561498 488746 561734
rect 488982 561498 524426 561734
rect 524662 561498 524746 561734
rect 524982 561498 560426 561734
rect 560662 561498 560746 561734
rect 560982 561498 590142 561734
rect 590378 561498 590462 561734
rect 590698 561498 592650 561734
rect -8726 561466 592650 561498
rect -8726 558334 592650 558366
rect -8726 558098 -5814 558334
rect -5578 558098 -5494 558334
rect -5258 558098 16706 558334
rect 16942 558098 17026 558334
rect 17262 558098 376706 558334
rect 376942 558098 377026 558334
rect 377262 558098 412706 558334
rect 412942 558098 413026 558334
rect 413262 558098 448706 558334
rect 448942 558098 449026 558334
rect 449262 558098 484706 558334
rect 484942 558098 485026 558334
rect 485262 558098 520706 558334
rect 520942 558098 521026 558334
rect 521262 558098 556706 558334
rect 556942 558098 557026 558334
rect 557262 558098 589182 558334
rect 589418 558098 589502 558334
rect 589738 558098 592650 558334
rect -8726 558014 592650 558098
rect -8726 557778 -5814 558014
rect -5578 557778 -5494 558014
rect -5258 557778 16706 558014
rect 16942 557778 17026 558014
rect 17262 557778 376706 558014
rect 376942 557778 377026 558014
rect 377262 557778 412706 558014
rect 412942 557778 413026 558014
rect 413262 557778 448706 558014
rect 448942 557778 449026 558014
rect 449262 557778 484706 558014
rect 484942 557778 485026 558014
rect 485262 557778 520706 558014
rect 520942 557778 521026 558014
rect 521262 557778 556706 558014
rect 556942 557778 557026 558014
rect 557262 557778 589182 558014
rect 589418 557778 589502 558014
rect 589738 557778 592650 558014
rect -8726 557746 592650 557778
rect -8726 554614 592650 554646
rect -8726 554378 -4854 554614
rect -4618 554378 -4534 554614
rect -4298 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 372986 554614
rect 373222 554378 373306 554614
rect 373542 554378 408986 554614
rect 409222 554378 409306 554614
rect 409542 554378 444986 554614
rect 445222 554378 445306 554614
rect 445542 554378 480986 554614
rect 481222 554378 481306 554614
rect 481542 554378 516986 554614
rect 517222 554378 517306 554614
rect 517542 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 588222 554614
rect 588458 554378 588542 554614
rect 588778 554378 592650 554614
rect -8726 554294 592650 554378
rect -8726 554058 -4854 554294
rect -4618 554058 -4534 554294
rect -4298 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 372986 554294
rect 373222 554058 373306 554294
rect 373542 554058 408986 554294
rect 409222 554058 409306 554294
rect 409542 554058 444986 554294
rect 445222 554058 445306 554294
rect 445542 554058 480986 554294
rect 481222 554058 481306 554294
rect 481542 554058 516986 554294
rect 517222 554058 517306 554294
rect 517542 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 588222 554294
rect 588458 554058 588542 554294
rect 588778 554058 592650 554294
rect -8726 554026 592650 554058
rect -8726 550894 592650 550926
rect -8726 550658 -3894 550894
rect -3658 550658 -3574 550894
rect -3338 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 369266 550894
rect 369502 550658 369586 550894
rect 369822 550658 405266 550894
rect 405502 550658 405586 550894
rect 405822 550658 441266 550894
rect 441502 550658 441586 550894
rect 441822 550658 477266 550894
rect 477502 550658 477586 550894
rect 477822 550658 513266 550894
rect 513502 550658 513586 550894
rect 513822 550658 549266 550894
rect 549502 550658 549586 550894
rect 549822 550658 587262 550894
rect 587498 550658 587582 550894
rect 587818 550658 592650 550894
rect -8726 550574 592650 550658
rect -8726 550338 -3894 550574
rect -3658 550338 -3574 550574
rect -3338 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 369266 550574
rect 369502 550338 369586 550574
rect 369822 550338 405266 550574
rect 405502 550338 405586 550574
rect 405822 550338 441266 550574
rect 441502 550338 441586 550574
rect 441822 550338 477266 550574
rect 477502 550338 477586 550574
rect 477822 550338 513266 550574
rect 513502 550338 513586 550574
rect 513822 550338 549266 550574
rect 549502 550338 549586 550574
rect 549822 550338 587262 550574
rect 587498 550338 587582 550574
rect 587818 550338 592650 550574
rect -8726 550306 592650 550338
rect -8726 547174 592650 547206
rect -8726 546938 -2934 547174
rect -2698 546938 -2614 547174
rect -2378 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 39610 547174
rect 39846 546938 70330 547174
rect 70566 546938 101050 547174
rect 101286 546938 131770 547174
rect 132006 546938 162490 547174
rect 162726 546938 193210 547174
rect 193446 546938 223930 547174
rect 224166 546938 254650 547174
rect 254886 546938 285370 547174
rect 285606 546938 316090 547174
rect 316326 546938 346810 547174
rect 347046 546938 365546 547174
rect 365782 546938 365866 547174
rect 366102 546938 401546 547174
rect 401782 546938 401866 547174
rect 402102 546938 437546 547174
rect 437782 546938 437866 547174
rect 438102 546938 473546 547174
rect 473782 546938 473866 547174
rect 474102 546938 509546 547174
rect 509782 546938 509866 547174
rect 510102 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 586302 547174
rect 586538 546938 586622 547174
rect 586858 546938 592650 547174
rect -8726 546854 592650 546938
rect -8726 546618 -2934 546854
rect -2698 546618 -2614 546854
rect -2378 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 39610 546854
rect 39846 546618 70330 546854
rect 70566 546618 101050 546854
rect 101286 546618 131770 546854
rect 132006 546618 162490 546854
rect 162726 546618 193210 546854
rect 193446 546618 223930 546854
rect 224166 546618 254650 546854
rect 254886 546618 285370 546854
rect 285606 546618 316090 546854
rect 316326 546618 346810 546854
rect 347046 546618 365546 546854
rect 365782 546618 365866 546854
rect 366102 546618 401546 546854
rect 401782 546618 401866 546854
rect 402102 546618 437546 546854
rect 437782 546618 437866 546854
rect 438102 546618 473546 546854
rect 473782 546618 473866 546854
rect 474102 546618 509546 546854
rect 509782 546618 509866 546854
rect 510102 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 586302 546854
rect 586538 546618 586622 546854
rect 586858 546618 592650 546854
rect -8726 546586 592650 546618
rect -8726 543454 592650 543486
rect -8726 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 24250 543454
rect 24486 543218 54970 543454
rect 55206 543218 85690 543454
rect 85926 543218 116410 543454
rect 116646 543218 147130 543454
rect 147366 543218 177850 543454
rect 178086 543218 208570 543454
rect 208806 543218 239290 543454
rect 239526 543218 270010 543454
rect 270246 543218 300730 543454
rect 300966 543218 331450 543454
rect 331686 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 592650 543454
rect -8726 543134 592650 543218
rect -8726 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 24250 543134
rect 24486 542898 54970 543134
rect 55206 542898 85690 543134
rect 85926 542898 116410 543134
rect 116646 542898 147130 543134
rect 147366 542898 177850 543134
rect 178086 542898 208570 543134
rect 208806 542898 239290 543134
rect 239526 542898 270010 543134
rect 270246 542898 300730 543134
rect 300966 542898 331450 543134
rect 331686 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 592650 543134
rect -8726 542866 592650 542898
rect -8726 533494 592650 533526
rect -8726 533258 -8694 533494
rect -8458 533258 -8374 533494
rect -8138 533258 27866 533494
rect 28102 533258 28186 533494
rect 28422 533258 387866 533494
rect 388102 533258 388186 533494
rect 388422 533258 423866 533494
rect 424102 533258 424186 533494
rect 424422 533258 459866 533494
rect 460102 533258 460186 533494
rect 460422 533258 495866 533494
rect 496102 533258 496186 533494
rect 496422 533258 531866 533494
rect 532102 533258 532186 533494
rect 532422 533258 567866 533494
rect 568102 533258 568186 533494
rect 568422 533258 592062 533494
rect 592298 533258 592382 533494
rect 592618 533258 592650 533494
rect -8726 533174 592650 533258
rect -8726 532938 -8694 533174
rect -8458 532938 -8374 533174
rect -8138 532938 27866 533174
rect 28102 532938 28186 533174
rect 28422 532938 387866 533174
rect 388102 532938 388186 533174
rect 388422 532938 423866 533174
rect 424102 532938 424186 533174
rect 424422 532938 459866 533174
rect 460102 532938 460186 533174
rect 460422 532938 495866 533174
rect 496102 532938 496186 533174
rect 496422 532938 531866 533174
rect 532102 532938 532186 533174
rect 532422 532938 567866 533174
rect 568102 532938 568186 533174
rect 568422 532938 592062 533174
rect 592298 532938 592382 533174
rect 592618 532938 592650 533174
rect -8726 532906 592650 532938
rect -8726 529774 592650 529806
rect -8726 529538 -7734 529774
rect -7498 529538 -7414 529774
rect -7178 529538 384146 529774
rect 384382 529538 384466 529774
rect 384702 529538 420146 529774
rect 420382 529538 420466 529774
rect 420702 529538 456146 529774
rect 456382 529538 456466 529774
rect 456702 529538 492146 529774
rect 492382 529538 492466 529774
rect 492702 529538 528146 529774
rect 528382 529538 528466 529774
rect 528702 529538 564146 529774
rect 564382 529538 564466 529774
rect 564702 529538 591102 529774
rect 591338 529538 591422 529774
rect 591658 529538 592650 529774
rect -8726 529454 592650 529538
rect -8726 529218 -7734 529454
rect -7498 529218 -7414 529454
rect -7178 529218 384146 529454
rect 384382 529218 384466 529454
rect 384702 529218 420146 529454
rect 420382 529218 420466 529454
rect 420702 529218 456146 529454
rect 456382 529218 456466 529454
rect 456702 529218 492146 529454
rect 492382 529218 492466 529454
rect 492702 529218 528146 529454
rect 528382 529218 528466 529454
rect 528702 529218 564146 529454
rect 564382 529218 564466 529454
rect 564702 529218 591102 529454
rect 591338 529218 591422 529454
rect 591658 529218 592650 529454
rect -8726 529186 592650 529218
rect -8726 526054 592650 526086
rect -8726 525818 -6774 526054
rect -6538 525818 -6454 526054
rect -6218 525818 20426 526054
rect 20662 525818 20746 526054
rect 20982 525818 380426 526054
rect 380662 525818 380746 526054
rect 380982 525818 416426 526054
rect 416662 525818 416746 526054
rect 416982 525818 452426 526054
rect 452662 525818 452746 526054
rect 452982 525818 488426 526054
rect 488662 525818 488746 526054
rect 488982 525818 524426 526054
rect 524662 525818 524746 526054
rect 524982 525818 560426 526054
rect 560662 525818 560746 526054
rect 560982 525818 590142 526054
rect 590378 525818 590462 526054
rect 590698 525818 592650 526054
rect -8726 525734 592650 525818
rect -8726 525498 -6774 525734
rect -6538 525498 -6454 525734
rect -6218 525498 20426 525734
rect 20662 525498 20746 525734
rect 20982 525498 380426 525734
rect 380662 525498 380746 525734
rect 380982 525498 416426 525734
rect 416662 525498 416746 525734
rect 416982 525498 452426 525734
rect 452662 525498 452746 525734
rect 452982 525498 488426 525734
rect 488662 525498 488746 525734
rect 488982 525498 524426 525734
rect 524662 525498 524746 525734
rect 524982 525498 560426 525734
rect 560662 525498 560746 525734
rect 560982 525498 590142 525734
rect 590378 525498 590462 525734
rect 590698 525498 592650 525734
rect -8726 525466 592650 525498
rect -8726 522334 592650 522366
rect -8726 522098 -5814 522334
rect -5578 522098 -5494 522334
rect -5258 522098 16706 522334
rect 16942 522098 17026 522334
rect 17262 522098 376706 522334
rect 376942 522098 377026 522334
rect 377262 522098 412706 522334
rect 412942 522098 413026 522334
rect 413262 522098 448706 522334
rect 448942 522098 449026 522334
rect 449262 522098 484706 522334
rect 484942 522098 485026 522334
rect 485262 522098 520706 522334
rect 520942 522098 521026 522334
rect 521262 522098 556706 522334
rect 556942 522098 557026 522334
rect 557262 522098 589182 522334
rect 589418 522098 589502 522334
rect 589738 522098 592650 522334
rect -8726 522014 592650 522098
rect -8726 521778 -5814 522014
rect -5578 521778 -5494 522014
rect -5258 521778 16706 522014
rect 16942 521778 17026 522014
rect 17262 521778 376706 522014
rect 376942 521778 377026 522014
rect 377262 521778 412706 522014
rect 412942 521778 413026 522014
rect 413262 521778 448706 522014
rect 448942 521778 449026 522014
rect 449262 521778 484706 522014
rect 484942 521778 485026 522014
rect 485262 521778 520706 522014
rect 520942 521778 521026 522014
rect 521262 521778 556706 522014
rect 556942 521778 557026 522014
rect 557262 521778 589182 522014
rect 589418 521778 589502 522014
rect 589738 521778 592650 522014
rect -8726 521746 592650 521778
rect -8726 518614 592650 518646
rect -8726 518378 -4854 518614
rect -4618 518378 -4534 518614
rect -4298 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 372986 518614
rect 373222 518378 373306 518614
rect 373542 518378 408986 518614
rect 409222 518378 409306 518614
rect 409542 518378 444986 518614
rect 445222 518378 445306 518614
rect 445542 518378 480986 518614
rect 481222 518378 481306 518614
rect 481542 518378 516986 518614
rect 517222 518378 517306 518614
rect 517542 518378 552986 518614
rect 553222 518378 553306 518614
rect 553542 518378 588222 518614
rect 588458 518378 588542 518614
rect 588778 518378 592650 518614
rect -8726 518294 592650 518378
rect -8726 518058 -4854 518294
rect -4618 518058 -4534 518294
rect -4298 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 372986 518294
rect 373222 518058 373306 518294
rect 373542 518058 408986 518294
rect 409222 518058 409306 518294
rect 409542 518058 444986 518294
rect 445222 518058 445306 518294
rect 445542 518058 480986 518294
rect 481222 518058 481306 518294
rect 481542 518058 516986 518294
rect 517222 518058 517306 518294
rect 517542 518058 552986 518294
rect 553222 518058 553306 518294
rect 553542 518058 588222 518294
rect 588458 518058 588542 518294
rect 588778 518058 592650 518294
rect -8726 518026 592650 518058
rect -8726 514894 592650 514926
rect -8726 514658 -3894 514894
rect -3658 514658 -3574 514894
rect -3338 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 369266 514894
rect 369502 514658 369586 514894
rect 369822 514658 405266 514894
rect 405502 514658 405586 514894
rect 405822 514658 441266 514894
rect 441502 514658 441586 514894
rect 441822 514658 477266 514894
rect 477502 514658 477586 514894
rect 477822 514658 513266 514894
rect 513502 514658 513586 514894
rect 513822 514658 549266 514894
rect 549502 514658 549586 514894
rect 549822 514658 587262 514894
rect 587498 514658 587582 514894
rect 587818 514658 592650 514894
rect -8726 514574 592650 514658
rect -8726 514338 -3894 514574
rect -3658 514338 -3574 514574
rect -3338 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 369266 514574
rect 369502 514338 369586 514574
rect 369822 514338 405266 514574
rect 405502 514338 405586 514574
rect 405822 514338 441266 514574
rect 441502 514338 441586 514574
rect 441822 514338 477266 514574
rect 477502 514338 477586 514574
rect 477822 514338 513266 514574
rect 513502 514338 513586 514574
rect 513822 514338 549266 514574
rect 549502 514338 549586 514574
rect 549822 514338 587262 514574
rect 587498 514338 587582 514574
rect 587818 514338 592650 514574
rect -8726 514306 592650 514338
rect -8726 511174 592650 511206
rect -8726 510938 -2934 511174
rect -2698 510938 -2614 511174
rect -2378 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 39610 511174
rect 39846 510938 70330 511174
rect 70566 510938 101050 511174
rect 101286 510938 131770 511174
rect 132006 510938 162490 511174
rect 162726 510938 193210 511174
rect 193446 510938 223930 511174
rect 224166 510938 254650 511174
rect 254886 510938 285370 511174
rect 285606 510938 316090 511174
rect 316326 510938 346810 511174
rect 347046 510938 365546 511174
rect 365782 510938 365866 511174
rect 366102 510938 401546 511174
rect 401782 510938 401866 511174
rect 402102 510938 437546 511174
rect 437782 510938 437866 511174
rect 438102 510938 453424 511174
rect 453660 510938 455862 511174
rect 456098 510938 458300 511174
rect 458536 510938 460738 511174
rect 460974 510938 473546 511174
rect 473782 510938 473866 511174
rect 474102 510938 483424 511174
rect 483660 510938 485862 511174
rect 486098 510938 488300 511174
rect 488536 510938 490738 511174
rect 490974 510938 509546 511174
rect 509782 510938 509866 511174
rect 510102 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 586302 511174
rect 586538 510938 586622 511174
rect 586858 510938 592650 511174
rect -8726 510854 592650 510938
rect -8726 510618 -2934 510854
rect -2698 510618 -2614 510854
rect -2378 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 39610 510854
rect 39846 510618 70330 510854
rect 70566 510618 101050 510854
rect 101286 510618 131770 510854
rect 132006 510618 162490 510854
rect 162726 510618 193210 510854
rect 193446 510618 223930 510854
rect 224166 510618 254650 510854
rect 254886 510618 285370 510854
rect 285606 510618 316090 510854
rect 316326 510618 346810 510854
rect 347046 510618 365546 510854
rect 365782 510618 365866 510854
rect 366102 510618 401546 510854
rect 401782 510618 401866 510854
rect 402102 510618 437546 510854
rect 437782 510618 437866 510854
rect 438102 510618 453424 510854
rect 453660 510618 455862 510854
rect 456098 510618 458300 510854
rect 458536 510618 460738 510854
rect 460974 510618 473546 510854
rect 473782 510618 473866 510854
rect 474102 510618 483424 510854
rect 483660 510618 485862 510854
rect 486098 510618 488300 510854
rect 488536 510618 490738 510854
rect 490974 510618 509546 510854
rect 509782 510618 509866 510854
rect 510102 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 586302 510854
rect 586538 510618 586622 510854
rect 586858 510618 592650 510854
rect -8726 510586 592650 510618
rect -8726 507454 592650 507486
rect -8726 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 24250 507454
rect 24486 507218 54970 507454
rect 55206 507218 85690 507454
rect 85926 507218 116410 507454
rect 116646 507218 147130 507454
rect 147366 507218 177850 507454
rect 178086 507218 208570 507454
rect 208806 507218 239290 507454
rect 239526 507218 270010 507454
rect 270246 507218 300730 507454
rect 300966 507218 331450 507454
rect 331686 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 452205 507454
rect 452441 507218 454643 507454
rect 454879 507218 457081 507454
rect 457317 507218 459519 507454
rect 459755 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 482205 507454
rect 482441 507218 484643 507454
rect 484879 507218 487081 507454
rect 487317 507218 489519 507454
rect 489755 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 592650 507454
rect -8726 507134 592650 507218
rect -8726 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 24250 507134
rect 24486 506898 54970 507134
rect 55206 506898 85690 507134
rect 85926 506898 116410 507134
rect 116646 506898 147130 507134
rect 147366 506898 177850 507134
rect 178086 506898 208570 507134
rect 208806 506898 239290 507134
rect 239526 506898 270010 507134
rect 270246 506898 300730 507134
rect 300966 506898 331450 507134
rect 331686 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 452205 507134
rect 452441 506898 454643 507134
rect 454879 506898 457081 507134
rect 457317 506898 459519 507134
rect 459755 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 482205 507134
rect 482441 506898 484643 507134
rect 484879 506898 487081 507134
rect 487317 506898 489519 507134
rect 489755 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 592650 507134
rect -8726 506866 592650 506898
rect -8726 497494 592650 497526
rect -8726 497258 -8694 497494
rect -8458 497258 -8374 497494
rect -8138 497258 27866 497494
rect 28102 497258 28186 497494
rect 28422 497258 387866 497494
rect 388102 497258 388186 497494
rect 388422 497258 423866 497494
rect 424102 497258 424186 497494
rect 424422 497258 459866 497494
rect 460102 497258 460186 497494
rect 460422 497258 495866 497494
rect 496102 497258 496186 497494
rect 496422 497258 531866 497494
rect 532102 497258 532186 497494
rect 532422 497258 567866 497494
rect 568102 497258 568186 497494
rect 568422 497258 592062 497494
rect 592298 497258 592382 497494
rect 592618 497258 592650 497494
rect -8726 497174 592650 497258
rect -8726 496938 -8694 497174
rect -8458 496938 -8374 497174
rect -8138 496938 27866 497174
rect 28102 496938 28186 497174
rect 28422 496938 387866 497174
rect 388102 496938 388186 497174
rect 388422 496938 423866 497174
rect 424102 496938 424186 497174
rect 424422 496938 459866 497174
rect 460102 496938 460186 497174
rect 460422 496938 495866 497174
rect 496102 496938 496186 497174
rect 496422 496938 531866 497174
rect 532102 496938 532186 497174
rect 532422 496938 567866 497174
rect 568102 496938 568186 497174
rect 568422 496938 592062 497174
rect 592298 496938 592382 497174
rect 592618 496938 592650 497174
rect -8726 496906 592650 496938
rect -8726 493774 592650 493806
rect -8726 493538 -7734 493774
rect -7498 493538 -7414 493774
rect -7178 493538 384146 493774
rect 384382 493538 384466 493774
rect 384702 493538 420146 493774
rect 420382 493538 420466 493774
rect 420702 493538 456146 493774
rect 456382 493538 456466 493774
rect 456702 493538 492146 493774
rect 492382 493538 492466 493774
rect 492702 493538 528146 493774
rect 528382 493538 528466 493774
rect 528702 493538 564146 493774
rect 564382 493538 564466 493774
rect 564702 493538 591102 493774
rect 591338 493538 591422 493774
rect 591658 493538 592650 493774
rect -8726 493454 592650 493538
rect -8726 493218 -7734 493454
rect -7498 493218 -7414 493454
rect -7178 493218 384146 493454
rect 384382 493218 384466 493454
rect 384702 493218 420146 493454
rect 420382 493218 420466 493454
rect 420702 493218 456146 493454
rect 456382 493218 456466 493454
rect 456702 493218 492146 493454
rect 492382 493218 492466 493454
rect 492702 493218 528146 493454
rect 528382 493218 528466 493454
rect 528702 493218 564146 493454
rect 564382 493218 564466 493454
rect 564702 493218 591102 493454
rect 591338 493218 591422 493454
rect 591658 493218 592650 493454
rect -8726 493186 592650 493218
rect -8726 490054 592650 490086
rect -8726 489818 -6774 490054
rect -6538 489818 -6454 490054
rect -6218 489818 20426 490054
rect 20662 489818 20746 490054
rect 20982 489818 380426 490054
rect 380662 489818 380746 490054
rect 380982 489818 416426 490054
rect 416662 489818 416746 490054
rect 416982 489818 452426 490054
rect 452662 489818 452746 490054
rect 452982 489818 488426 490054
rect 488662 489818 488746 490054
rect 488982 489818 524426 490054
rect 524662 489818 524746 490054
rect 524982 489818 560426 490054
rect 560662 489818 560746 490054
rect 560982 489818 590142 490054
rect 590378 489818 590462 490054
rect 590698 489818 592650 490054
rect -8726 489734 592650 489818
rect -8726 489498 -6774 489734
rect -6538 489498 -6454 489734
rect -6218 489498 20426 489734
rect 20662 489498 20746 489734
rect 20982 489498 380426 489734
rect 380662 489498 380746 489734
rect 380982 489498 416426 489734
rect 416662 489498 416746 489734
rect 416982 489498 452426 489734
rect 452662 489498 452746 489734
rect 452982 489498 488426 489734
rect 488662 489498 488746 489734
rect 488982 489498 524426 489734
rect 524662 489498 524746 489734
rect 524982 489498 560426 489734
rect 560662 489498 560746 489734
rect 560982 489498 590142 489734
rect 590378 489498 590462 489734
rect 590698 489498 592650 489734
rect -8726 489466 592650 489498
rect -8726 486334 592650 486366
rect -8726 486098 -5814 486334
rect -5578 486098 -5494 486334
rect -5258 486098 16706 486334
rect 16942 486098 17026 486334
rect 17262 486098 376706 486334
rect 376942 486098 377026 486334
rect 377262 486098 412706 486334
rect 412942 486098 413026 486334
rect 413262 486098 448706 486334
rect 448942 486098 449026 486334
rect 449262 486098 484706 486334
rect 484942 486098 485026 486334
rect 485262 486098 520706 486334
rect 520942 486098 521026 486334
rect 521262 486098 556706 486334
rect 556942 486098 557026 486334
rect 557262 486098 589182 486334
rect 589418 486098 589502 486334
rect 589738 486098 592650 486334
rect -8726 486014 592650 486098
rect -8726 485778 -5814 486014
rect -5578 485778 -5494 486014
rect -5258 485778 16706 486014
rect 16942 485778 17026 486014
rect 17262 485778 376706 486014
rect 376942 485778 377026 486014
rect 377262 485778 412706 486014
rect 412942 485778 413026 486014
rect 413262 485778 448706 486014
rect 448942 485778 449026 486014
rect 449262 485778 484706 486014
rect 484942 485778 485026 486014
rect 485262 485778 520706 486014
rect 520942 485778 521026 486014
rect 521262 485778 556706 486014
rect 556942 485778 557026 486014
rect 557262 485778 589182 486014
rect 589418 485778 589502 486014
rect 589738 485778 592650 486014
rect -8726 485746 592650 485778
rect -8726 482614 592650 482646
rect -8726 482378 -4854 482614
rect -4618 482378 -4534 482614
rect -4298 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 372986 482614
rect 373222 482378 373306 482614
rect 373542 482378 408986 482614
rect 409222 482378 409306 482614
rect 409542 482378 444986 482614
rect 445222 482378 445306 482614
rect 445542 482378 480986 482614
rect 481222 482378 481306 482614
rect 481542 482378 516986 482614
rect 517222 482378 517306 482614
rect 517542 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 588222 482614
rect 588458 482378 588542 482614
rect 588778 482378 592650 482614
rect -8726 482294 592650 482378
rect -8726 482058 -4854 482294
rect -4618 482058 -4534 482294
rect -4298 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 372986 482294
rect 373222 482058 373306 482294
rect 373542 482058 408986 482294
rect 409222 482058 409306 482294
rect 409542 482058 444986 482294
rect 445222 482058 445306 482294
rect 445542 482058 480986 482294
rect 481222 482058 481306 482294
rect 481542 482058 516986 482294
rect 517222 482058 517306 482294
rect 517542 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 588222 482294
rect 588458 482058 588542 482294
rect 588778 482058 592650 482294
rect -8726 482026 592650 482058
rect -8726 478894 592650 478926
rect -8726 478658 -3894 478894
rect -3658 478658 -3574 478894
rect -3338 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 369266 478894
rect 369502 478658 369586 478894
rect 369822 478658 405266 478894
rect 405502 478658 405586 478894
rect 405822 478658 441266 478894
rect 441502 478658 441586 478894
rect 441822 478658 477266 478894
rect 477502 478658 477586 478894
rect 477822 478658 513266 478894
rect 513502 478658 513586 478894
rect 513822 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 587262 478894
rect 587498 478658 587582 478894
rect 587818 478658 592650 478894
rect -8726 478574 592650 478658
rect -8726 478338 -3894 478574
rect -3658 478338 -3574 478574
rect -3338 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 369266 478574
rect 369502 478338 369586 478574
rect 369822 478338 405266 478574
rect 405502 478338 405586 478574
rect 405822 478338 441266 478574
rect 441502 478338 441586 478574
rect 441822 478338 477266 478574
rect 477502 478338 477586 478574
rect 477822 478338 513266 478574
rect 513502 478338 513586 478574
rect 513822 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 587262 478574
rect 587498 478338 587582 478574
rect 587818 478338 592650 478574
rect -8726 478306 592650 478338
rect -8726 475174 592650 475206
rect -8726 474938 -2934 475174
rect -2698 474938 -2614 475174
rect -2378 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 39610 475174
rect 39846 474938 70330 475174
rect 70566 474938 101050 475174
rect 101286 474938 131770 475174
rect 132006 474938 162490 475174
rect 162726 474938 193210 475174
rect 193446 474938 223930 475174
rect 224166 474938 254650 475174
rect 254886 474938 285370 475174
rect 285606 474938 316090 475174
rect 316326 474938 346810 475174
rect 347046 474938 365546 475174
rect 365782 474938 365866 475174
rect 366102 474938 401546 475174
rect 401782 474938 401866 475174
rect 402102 474938 437546 475174
rect 437782 474938 437866 475174
rect 438102 474938 473546 475174
rect 473782 474938 473866 475174
rect 474102 474938 509546 475174
rect 509782 474938 509866 475174
rect 510102 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 586302 475174
rect 586538 474938 586622 475174
rect 586858 474938 592650 475174
rect -8726 474854 592650 474938
rect -8726 474618 -2934 474854
rect -2698 474618 -2614 474854
rect -2378 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 39610 474854
rect 39846 474618 70330 474854
rect 70566 474618 101050 474854
rect 101286 474618 131770 474854
rect 132006 474618 162490 474854
rect 162726 474618 193210 474854
rect 193446 474618 223930 474854
rect 224166 474618 254650 474854
rect 254886 474618 285370 474854
rect 285606 474618 316090 474854
rect 316326 474618 346810 474854
rect 347046 474618 365546 474854
rect 365782 474618 365866 474854
rect 366102 474618 401546 474854
rect 401782 474618 401866 474854
rect 402102 474618 437546 474854
rect 437782 474618 437866 474854
rect 438102 474618 473546 474854
rect 473782 474618 473866 474854
rect 474102 474618 509546 474854
rect 509782 474618 509866 474854
rect 510102 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 586302 474854
rect 586538 474618 586622 474854
rect 586858 474618 592650 474854
rect -8726 474586 592650 474618
rect -8726 471454 592650 471486
rect -8726 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 24250 471454
rect 24486 471218 54970 471454
rect 55206 471218 85690 471454
rect 85926 471218 116410 471454
rect 116646 471218 147130 471454
rect 147366 471218 177850 471454
rect 178086 471218 208570 471454
rect 208806 471218 239290 471454
rect 239526 471218 270010 471454
rect 270246 471218 300730 471454
rect 300966 471218 331450 471454
rect 331686 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 592650 471454
rect -8726 471134 592650 471218
rect -8726 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 24250 471134
rect 24486 470898 54970 471134
rect 55206 470898 85690 471134
rect 85926 470898 116410 471134
rect 116646 470898 147130 471134
rect 147366 470898 177850 471134
rect 178086 470898 208570 471134
rect 208806 470898 239290 471134
rect 239526 470898 270010 471134
rect 270246 470898 300730 471134
rect 300966 470898 331450 471134
rect 331686 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 592650 471134
rect -8726 470866 592650 470898
rect -8726 461494 592650 461526
rect -8726 461258 -8694 461494
rect -8458 461258 -8374 461494
rect -8138 461258 27866 461494
rect 28102 461258 28186 461494
rect 28422 461258 387866 461494
rect 388102 461258 388186 461494
rect 388422 461258 423866 461494
rect 424102 461258 424186 461494
rect 424422 461258 459866 461494
rect 460102 461258 460186 461494
rect 460422 461258 495866 461494
rect 496102 461258 496186 461494
rect 496422 461258 531866 461494
rect 532102 461258 532186 461494
rect 532422 461258 567866 461494
rect 568102 461258 568186 461494
rect 568422 461258 592062 461494
rect 592298 461258 592382 461494
rect 592618 461258 592650 461494
rect -8726 461174 592650 461258
rect -8726 460938 -8694 461174
rect -8458 460938 -8374 461174
rect -8138 460938 27866 461174
rect 28102 460938 28186 461174
rect 28422 460938 387866 461174
rect 388102 460938 388186 461174
rect 388422 460938 423866 461174
rect 424102 460938 424186 461174
rect 424422 460938 459866 461174
rect 460102 460938 460186 461174
rect 460422 460938 495866 461174
rect 496102 460938 496186 461174
rect 496422 460938 531866 461174
rect 532102 460938 532186 461174
rect 532422 460938 567866 461174
rect 568102 460938 568186 461174
rect 568422 460938 592062 461174
rect 592298 460938 592382 461174
rect 592618 460938 592650 461174
rect -8726 460906 592650 460938
rect -8726 457774 592650 457806
rect -8726 457538 -7734 457774
rect -7498 457538 -7414 457774
rect -7178 457538 384146 457774
rect 384382 457538 384466 457774
rect 384702 457538 420146 457774
rect 420382 457538 420466 457774
rect 420702 457538 456146 457774
rect 456382 457538 456466 457774
rect 456702 457538 492146 457774
rect 492382 457538 492466 457774
rect 492702 457538 528146 457774
rect 528382 457538 528466 457774
rect 528702 457538 564146 457774
rect 564382 457538 564466 457774
rect 564702 457538 591102 457774
rect 591338 457538 591422 457774
rect 591658 457538 592650 457774
rect -8726 457454 592650 457538
rect -8726 457218 -7734 457454
rect -7498 457218 -7414 457454
rect -7178 457218 384146 457454
rect 384382 457218 384466 457454
rect 384702 457218 420146 457454
rect 420382 457218 420466 457454
rect 420702 457218 456146 457454
rect 456382 457218 456466 457454
rect 456702 457218 492146 457454
rect 492382 457218 492466 457454
rect 492702 457218 528146 457454
rect 528382 457218 528466 457454
rect 528702 457218 564146 457454
rect 564382 457218 564466 457454
rect 564702 457218 591102 457454
rect 591338 457218 591422 457454
rect 591658 457218 592650 457454
rect -8726 457186 592650 457218
rect -8726 454054 592650 454086
rect -8726 453818 -6774 454054
rect -6538 453818 -6454 454054
rect -6218 453818 20426 454054
rect 20662 453818 20746 454054
rect 20982 453818 380426 454054
rect 380662 453818 380746 454054
rect 380982 453818 416426 454054
rect 416662 453818 416746 454054
rect 416982 453818 452426 454054
rect 452662 453818 452746 454054
rect 452982 454007 524426 454054
rect 452982 453818 488426 454007
rect -8726 453771 488426 453818
rect 488662 453771 488746 454007
rect 488982 453818 524426 454007
rect 524662 453818 524746 454054
rect 524982 453818 560426 454054
rect 560662 453818 560746 454054
rect 560982 453818 590142 454054
rect 590378 453818 590462 454054
rect 590698 453818 592650 454054
rect 488982 453771 592650 453818
rect -8726 453734 592650 453771
rect -8726 453498 -6774 453734
rect -6538 453498 -6454 453734
rect -6218 453498 20426 453734
rect 20662 453498 20746 453734
rect 20982 453498 380426 453734
rect 380662 453498 380746 453734
rect 380982 453498 416426 453734
rect 416662 453498 416746 453734
rect 416982 453498 452426 453734
rect 452662 453498 452746 453734
rect 452982 453498 524426 453734
rect 524662 453498 524746 453734
rect 524982 453498 560426 453734
rect 560662 453498 560746 453734
rect 560982 453498 590142 453734
rect 590378 453498 590462 453734
rect 590698 453498 592650 453734
rect -8726 453466 592650 453498
rect -8726 450334 592650 450366
rect -8726 450098 -5814 450334
rect -5578 450098 -5494 450334
rect -5258 450098 16706 450334
rect 16942 450098 17026 450334
rect 17262 450098 376706 450334
rect 376942 450098 377026 450334
rect 377262 450098 412706 450334
rect 412942 450098 413026 450334
rect 413262 450098 448706 450334
rect 448942 450098 449026 450334
rect 449262 450098 484706 450334
rect 484942 450098 485026 450334
rect 485262 450098 520706 450334
rect 520942 450098 521026 450334
rect 521262 450098 556706 450334
rect 556942 450098 557026 450334
rect 557262 450098 589182 450334
rect 589418 450098 589502 450334
rect 589738 450098 592650 450334
rect -8726 450014 592650 450098
rect -8726 449778 -5814 450014
rect -5578 449778 -5494 450014
rect -5258 449778 16706 450014
rect 16942 449778 17026 450014
rect 17262 449778 376706 450014
rect 376942 449778 377026 450014
rect 377262 449778 412706 450014
rect 412942 449778 413026 450014
rect 413262 449778 448706 450014
rect 448942 449778 449026 450014
rect 449262 449778 484706 450014
rect 484942 449778 485026 450014
rect 485262 449778 520706 450014
rect 520942 449778 521026 450014
rect 521262 449778 556706 450014
rect 556942 449778 557026 450014
rect 557262 449778 589182 450014
rect 589418 449778 589502 450014
rect 589738 449778 592650 450014
rect -8726 449746 592650 449778
rect -8726 446614 592650 446646
rect -8726 446378 -4854 446614
rect -4618 446378 -4534 446614
rect -4298 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 372986 446614
rect 373222 446378 373306 446614
rect 373542 446378 408986 446614
rect 409222 446378 409306 446614
rect 409542 446378 444986 446614
rect 445222 446378 445306 446614
rect 445542 446378 516986 446614
rect 517222 446378 517306 446614
rect 517542 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 588222 446614
rect 588458 446378 588542 446614
rect 588778 446378 592650 446614
rect -8726 446294 592650 446378
rect -8726 446058 -4854 446294
rect -4618 446058 -4534 446294
rect -4298 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 372986 446294
rect 373222 446058 373306 446294
rect 373542 446058 408986 446294
rect 409222 446058 409306 446294
rect 409542 446058 444986 446294
rect 445222 446058 445306 446294
rect 445542 446058 516986 446294
rect 517222 446058 517306 446294
rect 517542 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 588222 446294
rect 588458 446058 588542 446294
rect 588778 446058 592650 446294
rect -8726 446026 592650 446058
rect -8726 442894 592650 442926
rect -8726 442658 -3894 442894
rect -3658 442658 -3574 442894
rect -3338 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 369266 442894
rect 369502 442658 369586 442894
rect 369822 442658 405266 442894
rect 405502 442658 405586 442894
rect 405822 442658 477266 442894
rect 477502 442658 477586 442894
rect 477822 442658 513266 442894
rect 513502 442658 513586 442894
rect 513822 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 587262 442894
rect 587498 442658 587582 442894
rect 587818 442658 592650 442894
rect -8726 442574 592650 442658
rect -8726 442338 -3894 442574
rect -3658 442338 -3574 442574
rect -3338 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 369266 442574
rect 369502 442338 369586 442574
rect 369822 442338 405266 442574
rect 405502 442338 405586 442574
rect 405822 442338 477266 442574
rect 477502 442338 477586 442574
rect 477822 442338 513266 442574
rect 513502 442338 513586 442574
rect 513822 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 587262 442574
rect 587498 442338 587582 442574
rect 587818 442338 592650 442574
rect -8726 442306 592650 442338
rect -8726 439174 592650 439206
rect -8726 438938 -2934 439174
rect -2698 438938 -2614 439174
rect -2378 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 39610 439174
rect 39846 438938 70330 439174
rect 70566 438938 101050 439174
rect 101286 438938 131770 439174
rect 132006 438938 162490 439174
rect 162726 438938 193210 439174
rect 193446 438938 223930 439174
rect 224166 438938 254650 439174
rect 254886 438938 285370 439174
rect 285606 438938 316090 439174
rect 316326 438938 346810 439174
rect 347046 438938 365546 439174
rect 365782 438938 365866 439174
rect 366102 438938 401546 439174
rect 401782 438938 401866 439174
rect 402102 438938 426666 439174
rect 426902 438938 432347 439174
rect 432583 438938 438028 439174
rect 438264 438938 443709 439174
rect 443945 438938 475930 439174
rect 476166 438938 480875 439174
rect 481111 438938 485820 439174
rect 486056 438938 490765 439174
rect 491001 438938 509546 439174
rect 509782 438938 509866 439174
rect 510102 438938 529426 439174
rect 529662 438938 537867 439174
rect 538103 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 546308 439174
rect 546544 438938 554749 439174
rect 554985 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 586302 439174
rect 586538 438938 586622 439174
rect 586858 438938 592650 439174
rect -8726 438854 592650 438938
rect -8726 438618 -2934 438854
rect -2698 438618 -2614 438854
rect -2378 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 39610 438854
rect 39846 438618 70330 438854
rect 70566 438618 101050 438854
rect 101286 438618 131770 438854
rect 132006 438618 162490 438854
rect 162726 438618 193210 438854
rect 193446 438618 223930 438854
rect 224166 438618 254650 438854
rect 254886 438618 285370 438854
rect 285606 438618 316090 438854
rect 316326 438618 346810 438854
rect 347046 438618 365546 438854
rect 365782 438618 365866 438854
rect 366102 438618 401546 438854
rect 401782 438618 401866 438854
rect 402102 438618 426666 438854
rect 426902 438618 432347 438854
rect 432583 438618 438028 438854
rect 438264 438618 443709 438854
rect 443945 438618 475930 438854
rect 476166 438618 480875 438854
rect 481111 438618 485820 438854
rect 486056 438618 490765 438854
rect 491001 438618 509546 438854
rect 509782 438618 509866 438854
rect 510102 438618 529426 438854
rect 529662 438618 537867 438854
rect 538103 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 546308 438854
rect 546544 438618 554749 438854
rect 554985 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 586302 438854
rect 586538 438618 586622 438854
rect 586858 438618 592650 438854
rect -8726 438586 592650 438618
rect -8726 435454 592650 435486
rect -8726 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 24250 435454
rect 24486 435218 54970 435454
rect 55206 435218 85690 435454
rect 85926 435218 116410 435454
rect 116646 435218 147130 435454
rect 147366 435218 177850 435454
rect 178086 435218 208570 435454
rect 208806 435218 239290 435454
rect 239526 435218 270010 435454
rect 270246 435218 300730 435454
rect 300966 435218 331450 435454
rect 331686 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 423826 435454
rect 424062 435218 429507 435454
rect 429743 435218 435188 435454
rect 435424 435218 440869 435454
rect 441105 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 473458 435454
rect 473694 435218 478403 435454
rect 478639 435218 483348 435454
rect 483584 435218 488293 435454
rect 488529 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 525206 435454
rect 525442 435218 533647 435454
rect 533883 435218 542088 435454
rect 542324 435218 550529 435454
rect 550765 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 592650 435454
rect -8726 435134 592650 435218
rect -8726 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 24250 435134
rect 24486 434898 54970 435134
rect 55206 434898 85690 435134
rect 85926 434898 116410 435134
rect 116646 434898 147130 435134
rect 147366 434898 177850 435134
rect 178086 434898 208570 435134
rect 208806 434898 239290 435134
rect 239526 434898 270010 435134
rect 270246 434898 300730 435134
rect 300966 434898 331450 435134
rect 331686 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 423826 435134
rect 424062 434898 429507 435134
rect 429743 434898 435188 435134
rect 435424 434898 440869 435134
rect 441105 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 473458 435134
rect 473694 434898 478403 435134
rect 478639 434898 483348 435134
rect 483584 434898 488293 435134
rect 488529 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 525206 435134
rect 525442 434898 533647 435134
rect 533883 434898 542088 435134
rect 542324 434898 550529 435134
rect 550765 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 592650 435134
rect -8726 434866 592650 434898
rect -8726 425494 592650 425526
rect -8726 425258 -8694 425494
rect -8458 425258 -8374 425494
rect -8138 425258 27866 425494
rect 28102 425258 28186 425494
rect 28422 425258 387866 425494
rect 388102 425258 388186 425494
rect 388422 425258 459866 425494
rect 460102 425258 460186 425494
rect 460422 425258 495866 425494
rect 496102 425258 496186 425494
rect 496422 425258 531866 425494
rect 532102 425258 532186 425494
rect 532422 425258 567866 425494
rect 568102 425258 568186 425494
rect 568422 425258 592062 425494
rect 592298 425258 592382 425494
rect 592618 425258 592650 425494
rect -8726 425174 592650 425258
rect -8726 424938 -8694 425174
rect -8458 424938 -8374 425174
rect -8138 424938 27866 425174
rect 28102 424938 28186 425174
rect 28422 424938 387866 425174
rect 388102 424938 388186 425174
rect 388422 424938 459866 425174
rect 460102 424938 460186 425174
rect 460422 424938 495866 425174
rect 496102 424938 496186 425174
rect 496422 424938 531866 425174
rect 532102 424938 532186 425174
rect 532422 424938 567866 425174
rect 568102 424938 568186 425174
rect 568422 424938 592062 425174
rect 592298 424938 592382 425174
rect 592618 424938 592650 425174
rect -8726 424906 592650 424938
rect -8726 421774 592650 421806
rect -8726 421538 -7734 421774
rect -7498 421538 -7414 421774
rect -7178 421538 384146 421774
rect 384382 421538 384466 421774
rect 384702 421538 420146 421774
rect 420382 421538 420466 421774
rect 420702 421538 456146 421774
rect 456382 421538 456466 421774
rect 456702 421538 492146 421774
rect 492382 421538 492466 421774
rect 492702 421538 528146 421774
rect 528382 421538 528466 421774
rect 528702 421538 564146 421774
rect 564382 421538 564466 421774
rect 564702 421538 591102 421774
rect 591338 421538 591422 421774
rect 591658 421538 592650 421774
rect -8726 421454 592650 421538
rect -8726 421218 -7734 421454
rect -7498 421218 -7414 421454
rect -7178 421218 384146 421454
rect 384382 421218 384466 421454
rect 384702 421218 420146 421454
rect 420382 421218 420466 421454
rect 420702 421218 456146 421454
rect 456382 421218 456466 421454
rect 456702 421218 492146 421454
rect 492382 421218 492466 421454
rect 492702 421218 528146 421454
rect 528382 421218 528466 421454
rect 528702 421218 564146 421454
rect 564382 421218 564466 421454
rect 564702 421218 591102 421454
rect 591338 421218 591422 421454
rect 591658 421218 592650 421454
rect -8726 421186 592650 421218
rect -8726 418054 592650 418086
rect -8726 417818 -6774 418054
rect -6538 417818 -6454 418054
rect -6218 417818 20426 418054
rect 20662 417818 20746 418054
rect 20982 417818 380426 418054
rect 380662 417818 380746 418054
rect 380982 417818 416426 418054
rect 416662 417818 416746 418054
rect 416982 417818 452426 418054
rect 452662 417818 452746 418054
rect 452982 417818 524426 418054
rect 524662 417818 524746 418054
rect 524982 417818 560426 418054
rect 560662 417818 560746 418054
rect 560982 417818 590142 418054
rect 590378 417818 590462 418054
rect 590698 417818 592650 418054
rect -8726 417734 592650 417818
rect -8726 417498 -6774 417734
rect -6538 417498 -6454 417734
rect -6218 417498 20426 417734
rect 20662 417498 20746 417734
rect 20982 417498 380426 417734
rect 380662 417498 380746 417734
rect 380982 417498 416426 417734
rect 416662 417498 416746 417734
rect 416982 417498 452426 417734
rect 452662 417498 452746 417734
rect 452982 417498 524426 417734
rect 524662 417498 524746 417734
rect 524982 417498 560426 417734
rect 560662 417498 560746 417734
rect 560982 417498 590142 417734
rect 590378 417498 590462 417734
rect 590698 417498 592650 417734
rect -8726 417466 592650 417498
rect -8726 414334 592650 414366
rect -8726 414098 -5814 414334
rect -5578 414098 -5494 414334
rect -5258 414098 16706 414334
rect 16942 414098 17026 414334
rect 17262 414098 376706 414334
rect 376942 414098 377026 414334
rect 377262 414098 412706 414334
rect 412942 414098 413026 414334
rect 413262 414098 448706 414334
rect 448942 414098 449026 414334
rect 449262 414098 484706 414334
rect 484942 414098 485026 414334
rect 485262 414098 520706 414334
rect 520942 414098 521026 414334
rect 521262 414098 556706 414334
rect 556942 414098 557026 414334
rect 557262 414098 589182 414334
rect 589418 414098 589502 414334
rect 589738 414098 592650 414334
rect -8726 414014 592650 414098
rect -8726 413778 -5814 414014
rect -5578 413778 -5494 414014
rect -5258 413778 16706 414014
rect 16942 413778 17026 414014
rect 17262 413778 376706 414014
rect 376942 413778 377026 414014
rect 377262 413778 412706 414014
rect 412942 413778 413026 414014
rect 413262 413778 448706 414014
rect 448942 413778 449026 414014
rect 449262 413778 484706 414014
rect 484942 413778 485026 414014
rect 485262 413778 520706 414014
rect 520942 413778 521026 414014
rect 521262 413778 556706 414014
rect 556942 413778 557026 414014
rect 557262 413778 589182 414014
rect 589418 413778 589502 414014
rect 589738 413778 592650 414014
rect -8726 413746 592650 413778
rect -8726 410614 592650 410646
rect -8726 410378 -4854 410614
rect -4618 410378 -4534 410614
rect -4298 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 372986 410614
rect 373222 410378 373306 410614
rect 373542 410378 408986 410614
rect 409222 410378 409306 410614
rect 409542 410378 444986 410614
rect 445222 410378 445306 410614
rect 445542 410378 516986 410614
rect 517222 410378 517306 410614
rect 517542 410378 552986 410614
rect 553222 410378 553306 410614
rect 553542 410378 588222 410614
rect 588458 410378 588542 410614
rect 588778 410378 592650 410614
rect -8726 410294 592650 410378
rect -8726 410058 -4854 410294
rect -4618 410058 -4534 410294
rect -4298 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 372986 410294
rect 373222 410058 373306 410294
rect 373542 410058 408986 410294
rect 409222 410058 409306 410294
rect 409542 410058 444986 410294
rect 445222 410058 445306 410294
rect 445542 410058 516986 410294
rect 517222 410058 517306 410294
rect 517542 410058 552986 410294
rect 553222 410058 553306 410294
rect 553542 410058 588222 410294
rect 588458 410058 588542 410294
rect 588778 410058 592650 410294
rect -8726 410026 592650 410058
rect -8726 406894 592650 406926
rect -8726 406658 -3894 406894
rect -3658 406658 -3574 406894
rect -3338 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 369266 406894
rect 369502 406658 369586 406894
rect 369822 406658 405266 406894
rect 405502 406658 405586 406894
rect 405822 406658 441266 406894
rect 441502 406658 441586 406894
rect 441822 406658 477266 406894
rect 477502 406658 477586 406894
rect 477822 406658 513266 406894
rect 513502 406658 513586 406894
rect 513822 406658 549266 406894
rect 549502 406658 549586 406894
rect 549822 406658 587262 406894
rect 587498 406658 587582 406894
rect 587818 406658 592650 406894
rect -8726 406574 592650 406658
rect -8726 406338 -3894 406574
rect -3658 406338 -3574 406574
rect -3338 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 369266 406574
rect 369502 406338 369586 406574
rect 369822 406338 405266 406574
rect 405502 406338 405586 406574
rect 405822 406338 441266 406574
rect 441502 406338 441586 406574
rect 441822 406338 477266 406574
rect 477502 406338 477586 406574
rect 477822 406338 513266 406574
rect 513502 406338 513586 406574
rect 513822 406338 549266 406574
rect 549502 406338 549586 406574
rect 549822 406338 587262 406574
rect 587498 406338 587582 406574
rect 587818 406338 592650 406574
rect -8726 406306 592650 406338
rect -8726 403174 592650 403206
rect -8726 402938 -2934 403174
rect -2698 402938 -2614 403174
rect -2378 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 39610 403174
rect 39846 402938 70330 403174
rect 70566 402938 101050 403174
rect 101286 402938 131770 403174
rect 132006 402938 162490 403174
rect 162726 402938 193210 403174
rect 193446 402938 223930 403174
rect 224166 402938 254650 403174
rect 254886 402938 285370 403174
rect 285606 402938 316090 403174
rect 316326 402938 346810 403174
rect 347046 402938 365546 403174
rect 365782 402938 365866 403174
rect 366102 402938 401546 403174
rect 401782 402938 401866 403174
rect 402102 402938 437546 403174
rect 437782 402938 437866 403174
rect 438102 402938 509546 403174
rect 509782 402938 509866 403174
rect 510102 402938 545546 403174
rect 545782 402938 545866 403174
rect 546102 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 586302 403174
rect 586538 402938 586622 403174
rect 586858 402938 592650 403174
rect -8726 402854 592650 402938
rect -8726 402618 -2934 402854
rect -2698 402618 -2614 402854
rect -2378 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 39610 402854
rect 39846 402618 70330 402854
rect 70566 402618 101050 402854
rect 101286 402618 131770 402854
rect 132006 402618 162490 402854
rect 162726 402618 193210 402854
rect 193446 402618 223930 402854
rect 224166 402618 254650 402854
rect 254886 402618 285370 402854
rect 285606 402618 316090 402854
rect 316326 402618 346810 402854
rect 347046 402618 365546 402854
rect 365782 402618 365866 402854
rect 366102 402618 401546 402854
rect 401782 402618 401866 402854
rect 402102 402618 437546 402854
rect 437782 402618 437866 402854
rect 438102 402618 509546 402854
rect 509782 402618 509866 402854
rect 510102 402618 545546 402854
rect 545782 402618 545866 402854
rect 546102 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 586302 402854
rect 586538 402618 586622 402854
rect 586858 402618 592650 402854
rect -8726 402586 592650 402618
rect -8726 399454 592650 399486
rect -8726 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 24250 399454
rect 24486 399218 54970 399454
rect 55206 399218 85690 399454
rect 85926 399218 116410 399454
rect 116646 399218 147130 399454
rect 147366 399218 177850 399454
rect 178086 399218 208570 399454
rect 208806 399218 239290 399454
rect 239526 399218 270010 399454
rect 270246 399218 300730 399454
rect 300966 399218 331450 399454
rect 331686 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 592650 399454
rect -8726 399134 592650 399218
rect -8726 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 24250 399134
rect 24486 398898 54970 399134
rect 55206 398898 85690 399134
rect 85926 398898 116410 399134
rect 116646 398898 147130 399134
rect 147366 398898 177850 399134
rect 178086 398898 208570 399134
rect 208806 398898 239290 399134
rect 239526 398898 270010 399134
rect 270246 398898 300730 399134
rect 300966 398898 331450 399134
rect 331686 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 592650 399134
rect -8726 398866 592650 398898
rect -8726 389494 592650 389526
rect -8726 389258 -8694 389494
rect -8458 389258 -8374 389494
rect -8138 389258 27866 389494
rect 28102 389258 28186 389494
rect 28422 389258 387866 389494
rect 388102 389258 388186 389494
rect 388422 389258 423866 389494
rect 424102 389258 424186 389494
rect 424422 389258 459866 389494
rect 460102 389258 460186 389494
rect 460422 389258 495866 389494
rect 496102 389258 496186 389494
rect 496422 389258 531866 389494
rect 532102 389258 532186 389494
rect 532422 389258 567866 389494
rect 568102 389258 568186 389494
rect 568422 389258 592062 389494
rect 592298 389258 592382 389494
rect 592618 389258 592650 389494
rect -8726 389174 592650 389258
rect -8726 388938 -8694 389174
rect -8458 388938 -8374 389174
rect -8138 388938 27866 389174
rect 28102 388938 28186 389174
rect 28422 388938 387866 389174
rect 388102 388938 388186 389174
rect 388422 388938 423866 389174
rect 424102 388938 424186 389174
rect 424422 388938 459866 389174
rect 460102 388938 460186 389174
rect 460422 388938 495866 389174
rect 496102 388938 496186 389174
rect 496422 388938 531866 389174
rect 532102 388938 532186 389174
rect 532422 388938 567866 389174
rect 568102 388938 568186 389174
rect 568422 388938 592062 389174
rect 592298 388938 592382 389174
rect 592618 388938 592650 389174
rect -8726 388906 592650 388938
rect -8726 385774 592650 385806
rect -8726 385538 -7734 385774
rect -7498 385538 -7414 385774
rect -7178 385538 384146 385774
rect 384382 385538 384466 385774
rect 384702 385538 420146 385774
rect 420382 385538 420466 385774
rect 420702 385538 456146 385774
rect 456382 385538 456466 385774
rect 456702 385538 528146 385774
rect 528382 385538 528466 385774
rect 528702 385538 564146 385774
rect 564382 385538 564466 385774
rect 564702 385538 591102 385774
rect 591338 385538 591422 385774
rect 591658 385538 592650 385774
rect -8726 385454 592650 385538
rect -8726 385218 -7734 385454
rect -7498 385218 -7414 385454
rect -7178 385218 384146 385454
rect 384382 385218 384466 385454
rect 384702 385218 420146 385454
rect 420382 385218 420466 385454
rect 420702 385218 456146 385454
rect 456382 385218 456466 385454
rect 456702 385218 528146 385454
rect 528382 385218 528466 385454
rect 528702 385218 564146 385454
rect 564382 385218 564466 385454
rect 564702 385218 591102 385454
rect 591338 385218 591422 385454
rect 591658 385218 592650 385454
rect -8726 385186 592650 385218
rect -8726 382054 592650 382086
rect -8726 381818 -6774 382054
rect -6538 381818 -6454 382054
rect -6218 381818 20426 382054
rect 20662 381818 20746 382054
rect 20982 381818 380426 382054
rect 380662 381818 380746 382054
rect 380982 381818 416426 382054
rect 416662 381818 416746 382054
rect 416982 381818 452426 382054
rect 452662 381818 452746 382054
rect 452982 381818 524426 382054
rect 524662 381818 524746 382054
rect 524982 381818 560426 382054
rect 560662 381818 560746 382054
rect 560982 381818 590142 382054
rect 590378 381818 590462 382054
rect 590698 381818 592650 382054
rect -8726 381734 592650 381818
rect -8726 381498 -6774 381734
rect -6538 381498 -6454 381734
rect -6218 381498 20426 381734
rect 20662 381498 20746 381734
rect 20982 381498 380426 381734
rect 380662 381498 380746 381734
rect 380982 381498 416426 381734
rect 416662 381498 416746 381734
rect 416982 381498 452426 381734
rect 452662 381498 452746 381734
rect 452982 381498 524426 381734
rect 524662 381498 524746 381734
rect 524982 381498 560426 381734
rect 560662 381498 560746 381734
rect 560982 381498 590142 381734
rect 590378 381498 590462 381734
rect 590698 381498 592650 381734
rect -8726 381466 592650 381498
rect -8726 378334 592650 378366
rect -8726 378098 -5814 378334
rect -5578 378098 -5494 378334
rect -5258 378098 16706 378334
rect 16942 378098 17026 378334
rect 17262 378098 376706 378334
rect 376942 378098 377026 378334
rect 377262 378098 412706 378334
rect 412942 378098 413026 378334
rect 413262 378098 448706 378334
rect 448942 378098 449026 378334
rect 449262 378098 520706 378334
rect 520942 378098 521026 378334
rect 521262 378243 589182 378334
rect 521262 378098 556706 378243
rect -8726 378014 556706 378098
rect -8726 377778 -5814 378014
rect -5578 377778 -5494 378014
rect -5258 377778 16706 378014
rect 16942 377778 17026 378014
rect 17262 377778 376706 378014
rect 376942 377778 377026 378014
rect 377262 377778 412706 378014
rect 412942 377778 413026 378014
rect 413262 377778 448706 378014
rect 448942 377778 449026 378014
rect 449262 377778 520706 378014
rect 520942 377778 521026 378014
rect 521262 378007 556706 378014
rect 556942 378007 557026 378243
rect 557262 378098 589182 378243
rect 589418 378098 589502 378334
rect 589738 378098 592650 378334
rect 557262 378014 592650 378098
rect 557262 378007 589182 378014
rect 521262 377778 589182 378007
rect 589418 377778 589502 378014
rect 589738 377778 592650 378014
rect -8726 377746 592650 377778
rect -8726 374614 592650 374646
rect -8726 374378 -4854 374614
rect -4618 374378 -4534 374614
rect -4298 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 372986 374614
rect 373222 374378 373306 374614
rect 373542 374378 408986 374614
rect 409222 374378 409306 374614
rect 409542 374378 444986 374614
rect 445222 374378 445306 374614
rect 445542 374378 516986 374614
rect 517222 374378 517306 374614
rect 517542 374378 588222 374614
rect 588458 374378 588542 374614
rect 588778 374378 592650 374614
rect -8726 374294 592650 374378
rect -8726 374058 -4854 374294
rect -4618 374058 -4534 374294
rect -4298 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 372986 374294
rect 373222 374058 373306 374294
rect 373542 374058 408986 374294
rect 409222 374058 409306 374294
rect 409542 374058 444986 374294
rect 445222 374058 445306 374294
rect 445542 374058 516986 374294
rect 517222 374058 517306 374294
rect 517542 374058 588222 374294
rect 588458 374058 588542 374294
rect 588778 374058 592650 374294
rect -8726 374026 592650 374058
rect -8726 370894 592650 370926
rect -8726 370658 -3894 370894
rect -3658 370658 -3574 370894
rect -3338 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 369266 370894
rect 369502 370658 369586 370894
rect 369822 370658 405266 370894
rect 405502 370658 405586 370894
rect 405822 370658 441266 370894
rect 441502 370658 441586 370894
rect 441822 370658 513266 370894
rect 513502 370658 513586 370894
rect 513822 370658 549266 370894
rect 549502 370658 549586 370894
rect 549822 370658 587262 370894
rect 587498 370658 587582 370894
rect 587818 370658 592650 370894
rect -8726 370574 592650 370658
rect -8726 370338 -3894 370574
rect -3658 370338 -3574 370574
rect -3338 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 369266 370574
rect 369502 370338 369586 370574
rect 369822 370338 405266 370574
rect 405502 370338 405586 370574
rect 405822 370338 441266 370574
rect 441502 370338 441586 370574
rect 441822 370338 513266 370574
rect 513502 370338 513586 370574
rect 513822 370338 549266 370574
rect 549502 370338 549586 370574
rect 549822 370338 587262 370574
rect 587498 370338 587582 370574
rect 587818 370338 592650 370574
rect -8726 370306 592650 370338
rect -8726 367174 592650 367206
rect -8726 366938 -2934 367174
rect -2698 366938 -2614 367174
rect -2378 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 39610 367174
rect 39846 366938 70330 367174
rect 70566 366938 101050 367174
rect 101286 366938 131770 367174
rect 132006 366938 162490 367174
rect 162726 366938 193210 367174
rect 193446 366938 223930 367174
rect 224166 366938 254650 367174
rect 254886 366938 285370 367174
rect 285606 366938 316090 367174
rect 316326 366938 346810 367174
rect 347046 366938 365546 367174
rect 365782 366938 365866 367174
rect 366102 366938 401546 367174
rect 401782 366938 401866 367174
rect 402102 366938 437546 367174
rect 437782 366938 437866 367174
rect 438102 366938 469610 367174
rect 469846 366938 500330 367174
rect 500566 366938 509546 367174
rect 509782 366938 509866 367174
rect 510102 366938 545546 367174
rect 545782 366938 545866 367174
rect 546102 366938 554918 367174
rect 555154 366938 558851 367174
rect 559087 366938 562784 367174
rect 563020 366938 566717 367174
rect 566953 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 586302 367174
rect 586538 366938 586622 367174
rect 586858 366938 592650 367174
rect -8726 366854 592650 366938
rect -8726 366618 -2934 366854
rect -2698 366618 -2614 366854
rect -2378 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 39610 366854
rect 39846 366618 70330 366854
rect 70566 366618 101050 366854
rect 101286 366618 131770 366854
rect 132006 366618 162490 366854
rect 162726 366618 193210 366854
rect 193446 366618 223930 366854
rect 224166 366618 254650 366854
rect 254886 366618 285370 366854
rect 285606 366618 316090 366854
rect 316326 366618 346810 366854
rect 347046 366618 365546 366854
rect 365782 366618 365866 366854
rect 366102 366618 401546 366854
rect 401782 366618 401866 366854
rect 402102 366618 437546 366854
rect 437782 366618 437866 366854
rect 438102 366618 469610 366854
rect 469846 366618 500330 366854
rect 500566 366618 509546 366854
rect 509782 366618 509866 366854
rect 510102 366618 545546 366854
rect 545782 366618 545866 366854
rect 546102 366618 554918 366854
rect 555154 366618 558851 366854
rect 559087 366618 562784 366854
rect 563020 366618 566717 366854
rect 566953 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 586302 366854
rect 586538 366618 586622 366854
rect 586858 366618 592650 366854
rect -8726 366586 592650 366618
rect -8726 363454 592650 363486
rect -8726 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 24250 363454
rect 24486 363218 54970 363454
rect 55206 363218 85690 363454
rect 85926 363218 116410 363454
rect 116646 363218 147130 363454
rect 147366 363218 177850 363454
rect 178086 363218 208570 363454
rect 208806 363218 239290 363454
rect 239526 363218 270010 363454
rect 270246 363218 300730 363454
rect 300966 363218 331450 363454
rect 331686 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 454250 363454
rect 454486 363218 484970 363454
rect 485206 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 552952 363454
rect 553188 363218 556885 363454
rect 557121 363218 560818 363454
rect 561054 363218 564751 363454
rect 564987 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 592650 363454
rect -8726 363134 592650 363218
rect -8726 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 24250 363134
rect 24486 362898 54970 363134
rect 55206 362898 85690 363134
rect 85926 362898 116410 363134
rect 116646 362898 147130 363134
rect 147366 362898 177850 363134
rect 178086 362898 208570 363134
rect 208806 362898 239290 363134
rect 239526 362898 270010 363134
rect 270246 362898 300730 363134
rect 300966 362898 331450 363134
rect 331686 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 454250 363134
rect 454486 362898 484970 363134
rect 485206 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 552952 363134
rect 553188 362898 556885 363134
rect 557121 362898 560818 363134
rect 561054 362898 564751 363134
rect 564987 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 592650 363134
rect -8726 362866 592650 362898
rect -8726 353494 592650 353526
rect -8726 353258 -8694 353494
rect -8458 353258 -8374 353494
rect -8138 353258 27866 353494
rect 28102 353258 28186 353494
rect 28422 353258 387866 353494
rect 388102 353258 388186 353494
rect 388422 353258 423866 353494
rect 424102 353258 424186 353494
rect 424422 353258 459866 353494
rect 460102 353258 460186 353494
rect 460422 353258 495866 353494
rect 496102 353258 496186 353494
rect 496422 353258 531866 353494
rect 532102 353258 532186 353494
rect 532422 353258 567866 353494
rect 568102 353258 568186 353494
rect 568422 353258 592062 353494
rect 592298 353258 592382 353494
rect 592618 353258 592650 353494
rect -8726 353174 592650 353258
rect -8726 352938 -8694 353174
rect -8458 352938 -8374 353174
rect -8138 352938 27866 353174
rect 28102 352938 28186 353174
rect 28422 352938 387866 353174
rect 388102 352938 388186 353174
rect 388422 352938 423866 353174
rect 424102 352938 424186 353174
rect 424422 352938 459866 353174
rect 460102 352938 460186 353174
rect 460422 352938 495866 353174
rect 496102 352938 496186 353174
rect 496422 352938 531866 353174
rect 532102 352938 532186 353174
rect 532422 352938 567866 353174
rect 568102 352938 568186 353174
rect 568422 352938 592062 353174
rect 592298 352938 592382 353174
rect 592618 352938 592650 353174
rect -8726 352906 592650 352938
rect -8726 349774 592650 349806
rect -8726 349538 -7734 349774
rect -7498 349538 -7414 349774
rect -7178 349538 384146 349774
rect 384382 349538 384466 349774
rect 384702 349538 420146 349774
rect 420382 349538 420466 349774
rect 420702 349538 456146 349774
rect 456382 349538 456466 349774
rect 456702 349538 528146 349774
rect 528382 349538 528466 349774
rect 528702 349538 564146 349774
rect 564382 349538 564466 349774
rect 564702 349538 591102 349774
rect 591338 349538 591422 349774
rect 591658 349538 592650 349774
rect -8726 349454 592650 349538
rect -8726 349218 -7734 349454
rect -7498 349218 -7414 349454
rect -7178 349218 384146 349454
rect 384382 349218 384466 349454
rect 384702 349218 420146 349454
rect 420382 349218 420466 349454
rect 420702 349218 456146 349454
rect 456382 349218 456466 349454
rect 456702 349218 528146 349454
rect 528382 349218 528466 349454
rect 528702 349218 564146 349454
rect 564382 349218 564466 349454
rect 564702 349218 591102 349454
rect 591338 349218 591422 349454
rect 591658 349218 592650 349454
rect -8726 349186 592650 349218
rect -8726 346054 592650 346086
rect -8726 345818 -6774 346054
rect -6538 345818 -6454 346054
rect -6218 345818 20426 346054
rect 20662 345818 20746 346054
rect 20982 345818 380426 346054
rect 380662 345818 380746 346054
rect 380982 345818 416426 346054
rect 416662 345818 416746 346054
rect 416982 345818 452426 346054
rect 452662 345818 452746 346054
rect 452982 345818 524426 346054
rect 524662 345818 524746 346054
rect 524982 345818 560426 346054
rect 560662 345818 560746 346054
rect 560982 345818 590142 346054
rect 590378 345818 590462 346054
rect 590698 345818 592650 346054
rect -8726 345734 592650 345818
rect -8726 345498 -6774 345734
rect -6538 345498 -6454 345734
rect -6218 345498 20426 345734
rect 20662 345498 20746 345734
rect 20982 345498 380426 345734
rect 380662 345498 380746 345734
rect 380982 345498 416426 345734
rect 416662 345498 416746 345734
rect 416982 345498 452426 345734
rect 452662 345498 452746 345734
rect 452982 345498 524426 345734
rect 524662 345498 524746 345734
rect 524982 345498 560426 345734
rect 560662 345498 560746 345734
rect 560982 345498 590142 345734
rect 590378 345498 590462 345734
rect 590698 345498 592650 345734
rect -8726 345466 592650 345498
rect -8726 342334 592650 342366
rect -8726 342098 -5814 342334
rect -5578 342098 -5494 342334
rect -5258 342098 16706 342334
rect 16942 342098 17026 342334
rect 17262 342098 376706 342334
rect 376942 342098 377026 342334
rect 377262 342098 412706 342334
rect 412942 342098 413026 342334
rect 413262 342098 448706 342334
rect 448942 342098 449026 342334
rect 449262 342098 520706 342334
rect 520942 342098 521026 342334
rect 521262 342098 556706 342334
rect 556942 342098 557026 342334
rect 557262 342098 589182 342334
rect 589418 342098 589502 342334
rect 589738 342098 592650 342334
rect -8726 342014 592650 342098
rect -8726 341778 -5814 342014
rect -5578 341778 -5494 342014
rect -5258 341778 16706 342014
rect 16942 341778 17026 342014
rect 17262 341778 376706 342014
rect 376942 341778 377026 342014
rect 377262 341778 412706 342014
rect 412942 341778 413026 342014
rect 413262 341778 448706 342014
rect 448942 341778 449026 342014
rect 449262 341778 520706 342014
rect 520942 341778 521026 342014
rect 521262 341778 556706 342014
rect 556942 341778 557026 342014
rect 557262 341778 589182 342014
rect 589418 341778 589502 342014
rect 589738 341778 592650 342014
rect -8726 341746 592650 341778
rect -8726 338614 592650 338646
rect -8726 338378 -4854 338614
rect -4618 338378 -4534 338614
rect -4298 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 372986 338614
rect 373222 338378 373306 338614
rect 373542 338378 408986 338614
rect 409222 338378 409306 338614
rect 409542 338378 444986 338614
rect 445222 338378 445306 338614
rect 445542 338378 516986 338614
rect 517222 338378 517306 338614
rect 517542 338378 552986 338614
rect 553222 338378 553306 338614
rect 553542 338378 588222 338614
rect 588458 338378 588542 338614
rect 588778 338378 592650 338614
rect -8726 338294 592650 338378
rect -8726 338058 -4854 338294
rect -4618 338058 -4534 338294
rect -4298 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 372986 338294
rect 373222 338058 373306 338294
rect 373542 338058 408986 338294
rect 409222 338058 409306 338294
rect 409542 338058 444986 338294
rect 445222 338058 445306 338294
rect 445542 338058 516986 338294
rect 517222 338058 517306 338294
rect 517542 338058 552986 338294
rect 553222 338058 553306 338294
rect 553542 338058 588222 338294
rect 588458 338058 588542 338294
rect 588778 338058 592650 338294
rect -8726 338026 592650 338058
rect -8726 334894 592650 334926
rect -8726 334658 -3894 334894
rect -3658 334658 -3574 334894
rect -3338 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 369266 334894
rect 369502 334658 369586 334894
rect 369822 334658 405266 334894
rect 405502 334658 405586 334894
rect 405822 334658 441266 334894
rect 441502 334658 441586 334894
rect 441822 334658 513266 334894
rect 513502 334658 513586 334894
rect 513822 334658 549266 334894
rect 549502 334658 549586 334894
rect 549822 334658 587262 334894
rect 587498 334658 587582 334894
rect 587818 334658 592650 334894
rect -8726 334574 592650 334658
rect -8726 334338 -3894 334574
rect -3658 334338 -3574 334574
rect -3338 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 369266 334574
rect 369502 334338 369586 334574
rect 369822 334338 405266 334574
rect 405502 334338 405586 334574
rect 405822 334338 441266 334574
rect 441502 334338 441586 334574
rect 441822 334338 513266 334574
rect 513502 334338 513586 334574
rect 513822 334338 549266 334574
rect 549502 334338 549586 334574
rect 549822 334338 587262 334574
rect 587498 334338 587582 334574
rect 587818 334338 592650 334574
rect -8726 334306 592650 334338
rect -8726 331174 592650 331206
rect -8726 330938 -2934 331174
rect -2698 330938 -2614 331174
rect -2378 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 39610 331174
rect 39846 330938 70330 331174
rect 70566 330938 101050 331174
rect 101286 330938 131770 331174
rect 132006 330938 162490 331174
rect 162726 330938 193210 331174
rect 193446 330938 223930 331174
rect 224166 330938 254650 331174
rect 254886 330938 285370 331174
rect 285606 330938 316090 331174
rect 316326 330938 346810 331174
rect 347046 330938 365546 331174
rect 365782 330938 365866 331174
rect 366102 330938 401546 331174
rect 401782 330938 401866 331174
rect 402102 330938 407932 331174
rect 408168 330938 414878 331174
rect 415114 330938 421824 331174
rect 422060 330938 428770 331174
rect 429006 330938 437546 331174
rect 437782 330938 437866 331174
rect 438102 330938 469610 331174
rect 469846 330938 500330 331174
rect 500566 330938 509546 331174
rect 509782 330938 509866 331174
rect 510102 330938 545546 331174
rect 545782 330938 545866 331174
rect 546102 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 586302 331174
rect 586538 330938 586622 331174
rect 586858 330938 592650 331174
rect -8726 330854 592650 330938
rect -8726 330618 -2934 330854
rect -2698 330618 -2614 330854
rect -2378 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 39610 330854
rect 39846 330618 70330 330854
rect 70566 330618 101050 330854
rect 101286 330618 131770 330854
rect 132006 330618 162490 330854
rect 162726 330618 193210 330854
rect 193446 330618 223930 330854
rect 224166 330618 254650 330854
rect 254886 330618 285370 330854
rect 285606 330618 316090 330854
rect 316326 330618 346810 330854
rect 347046 330618 365546 330854
rect 365782 330618 365866 330854
rect 366102 330618 401546 330854
rect 401782 330618 401866 330854
rect 402102 330618 407932 330854
rect 408168 330618 414878 330854
rect 415114 330618 421824 330854
rect 422060 330618 428770 330854
rect 429006 330618 437546 330854
rect 437782 330618 437866 330854
rect 438102 330618 469610 330854
rect 469846 330618 500330 330854
rect 500566 330618 509546 330854
rect 509782 330618 509866 330854
rect 510102 330618 545546 330854
rect 545782 330618 545866 330854
rect 546102 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 586302 330854
rect 586538 330618 586622 330854
rect 586858 330618 592650 330854
rect -8726 330586 592650 330618
rect -8726 327454 592650 327486
rect -8726 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 24250 327454
rect 24486 327218 54970 327454
rect 55206 327218 85690 327454
rect 85926 327218 116410 327454
rect 116646 327218 147130 327454
rect 147366 327218 177850 327454
rect 178086 327218 208570 327454
rect 208806 327218 239290 327454
rect 239526 327218 270010 327454
rect 270246 327218 300730 327454
rect 300966 327218 331450 327454
rect 331686 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 404459 327454
rect 404695 327218 411405 327454
rect 411641 327218 418351 327454
rect 418587 327218 425297 327454
rect 425533 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 454250 327454
rect 454486 327218 484970 327454
rect 485206 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 592650 327454
rect -8726 327134 592650 327218
rect -8726 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 24250 327134
rect 24486 326898 54970 327134
rect 55206 326898 85690 327134
rect 85926 326898 116410 327134
rect 116646 326898 147130 327134
rect 147366 326898 177850 327134
rect 178086 326898 208570 327134
rect 208806 326898 239290 327134
rect 239526 326898 270010 327134
rect 270246 326898 300730 327134
rect 300966 326898 331450 327134
rect 331686 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 404459 327134
rect 404695 326898 411405 327134
rect 411641 326898 418351 327134
rect 418587 326898 425297 327134
rect 425533 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 454250 327134
rect 454486 326898 484970 327134
rect 485206 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 592650 327134
rect -8726 326866 592650 326898
rect -8726 317494 592650 317526
rect -8726 317258 -8694 317494
rect -8458 317258 -8374 317494
rect -8138 317258 27866 317494
rect 28102 317258 28186 317494
rect 28422 317258 387866 317494
rect 388102 317258 388186 317494
rect 388422 317258 423866 317494
rect 424102 317258 424186 317494
rect 424422 317258 459866 317494
rect 460102 317258 460186 317494
rect 460422 317258 495866 317494
rect 496102 317258 496186 317494
rect 496422 317258 531866 317494
rect 532102 317258 532186 317494
rect 532422 317258 567866 317494
rect 568102 317258 568186 317494
rect 568422 317258 592062 317494
rect 592298 317258 592382 317494
rect 592618 317258 592650 317494
rect -8726 317174 592650 317258
rect -8726 316938 -8694 317174
rect -8458 316938 -8374 317174
rect -8138 316938 27866 317174
rect 28102 316938 28186 317174
rect 28422 316938 387866 317174
rect 388102 316938 388186 317174
rect 388422 316938 423866 317174
rect 424102 316938 424186 317174
rect 424422 316938 459866 317174
rect 460102 316938 460186 317174
rect 460422 316938 495866 317174
rect 496102 316938 496186 317174
rect 496422 316938 531866 317174
rect 532102 316938 532186 317174
rect 532422 316938 567866 317174
rect 568102 316938 568186 317174
rect 568422 316938 592062 317174
rect 592298 316938 592382 317174
rect 592618 316938 592650 317174
rect -8726 316906 592650 316938
rect -8726 313774 592650 313806
rect -8726 313538 -7734 313774
rect -7498 313538 -7414 313774
rect -7178 313538 384146 313774
rect 384382 313538 384466 313774
rect 384702 313538 420146 313774
rect 420382 313538 420466 313774
rect 420702 313538 456146 313774
rect 456382 313538 456466 313774
rect 456702 313538 492146 313774
rect 492382 313538 492466 313774
rect 492702 313538 528146 313774
rect 528382 313538 528466 313774
rect 528702 313538 564146 313774
rect 564382 313538 564466 313774
rect 564702 313538 591102 313774
rect 591338 313538 591422 313774
rect 591658 313538 592650 313774
rect -8726 313454 592650 313538
rect -8726 313218 -7734 313454
rect -7498 313218 -7414 313454
rect -7178 313218 384146 313454
rect 384382 313218 384466 313454
rect 384702 313218 420146 313454
rect 420382 313218 420466 313454
rect 420702 313218 456146 313454
rect 456382 313218 456466 313454
rect 456702 313218 492146 313454
rect 492382 313218 492466 313454
rect 492702 313218 528146 313454
rect 528382 313218 528466 313454
rect 528702 313218 564146 313454
rect 564382 313218 564466 313454
rect 564702 313218 591102 313454
rect 591338 313218 591422 313454
rect 591658 313218 592650 313454
rect -8726 313186 592650 313218
rect -8726 310054 592650 310086
rect -8726 309818 -6774 310054
rect -6538 309818 -6454 310054
rect -6218 309818 20426 310054
rect 20662 309818 20746 310054
rect 20982 309818 380426 310054
rect 380662 309818 380746 310054
rect 380982 309818 416426 310054
rect 416662 309818 416746 310054
rect 416982 309818 452426 310054
rect 452662 309818 452746 310054
rect 452982 309818 488426 310054
rect 488662 309818 488746 310054
rect 488982 309818 524426 310054
rect 524662 309818 524746 310054
rect 524982 309818 560426 310054
rect 560662 309818 560746 310054
rect 560982 309818 590142 310054
rect 590378 309818 590462 310054
rect 590698 309818 592650 310054
rect -8726 309734 592650 309818
rect -8726 309498 -6774 309734
rect -6538 309498 -6454 309734
rect -6218 309498 20426 309734
rect 20662 309498 20746 309734
rect 20982 309498 380426 309734
rect 380662 309498 380746 309734
rect 380982 309498 416426 309734
rect 416662 309498 416746 309734
rect 416982 309498 452426 309734
rect 452662 309498 452746 309734
rect 452982 309498 488426 309734
rect 488662 309498 488746 309734
rect 488982 309498 524426 309734
rect 524662 309498 524746 309734
rect 524982 309498 560426 309734
rect 560662 309498 560746 309734
rect 560982 309498 590142 309734
rect 590378 309498 590462 309734
rect 590698 309498 592650 309734
rect -8726 309466 592650 309498
rect -8726 306334 592650 306366
rect -8726 306098 -5814 306334
rect -5578 306098 -5494 306334
rect -5258 306098 16706 306334
rect 16942 306098 17026 306334
rect 17262 306098 376706 306334
rect 376942 306098 377026 306334
rect 377262 306098 412706 306334
rect 412942 306098 413026 306334
rect 413262 306098 448706 306334
rect 448942 306098 449026 306334
rect 449262 306098 484706 306334
rect 484942 306098 485026 306334
rect 485262 306098 520706 306334
rect 520942 306098 521026 306334
rect 521262 306098 556706 306334
rect 556942 306098 557026 306334
rect 557262 306098 589182 306334
rect 589418 306098 589502 306334
rect 589738 306098 592650 306334
rect -8726 306014 592650 306098
rect -8726 305778 -5814 306014
rect -5578 305778 -5494 306014
rect -5258 305778 16706 306014
rect 16942 305778 17026 306014
rect 17262 305778 376706 306014
rect 376942 305778 377026 306014
rect 377262 305778 412706 306014
rect 412942 305778 413026 306014
rect 413262 305778 448706 306014
rect 448942 305778 449026 306014
rect 449262 305778 484706 306014
rect 484942 305778 485026 306014
rect 485262 305778 520706 306014
rect 520942 305778 521026 306014
rect 521262 305778 556706 306014
rect 556942 305778 557026 306014
rect 557262 305778 589182 306014
rect 589418 305778 589502 306014
rect 589738 305778 592650 306014
rect -8726 305746 592650 305778
rect -8726 302614 592650 302646
rect -8726 302378 -4854 302614
rect -4618 302378 -4534 302614
rect -4298 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 372986 302614
rect 373222 302378 373306 302614
rect 373542 302378 408986 302614
rect 409222 302378 409306 302614
rect 409542 302378 444986 302614
rect 445222 302378 445306 302614
rect 445542 302378 480986 302614
rect 481222 302378 481306 302614
rect 481542 302378 516986 302614
rect 517222 302378 517306 302614
rect 517542 302378 552986 302614
rect 553222 302378 553306 302614
rect 553542 302378 588222 302614
rect 588458 302378 588542 302614
rect 588778 302378 592650 302614
rect -8726 302294 592650 302378
rect -8726 302058 -4854 302294
rect -4618 302058 -4534 302294
rect -4298 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 372986 302294
rect 373222 302058 373306 302294
rect 373542 302058 408986 302294
rect 409222 302058 409306 302294
rect 409542 302058 444986 302294
rect 445222 302058 445306 302294
rect 445542 302058 480986 302294
rect 481222 302058 481306 302294
rect 481542 302058 516986 302294
rect 517222 302058 517306 302294
rect 517542 302058 552986 302294
rect 553222 302058 553306 302294
rect 553542 302058 588222 302294
rect 588458 302058 588542 302294
rect 588778 302058 592650 302294
rect -8726 302026 592650 302058
rect -8726 298894 592650 298926
rect -8726 298658 -3894 298894
rect -3658 298658 -3574 298894
rect -3338 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 369266 298894
rect 369502 298658 369586 298894
rect 369822 298658 405266 298894
rect 405502 298658 405586 298894
rect 405822 298658 441266 298894
rect 441502 298658 441586 298894
rect 441822 298658 477266 298894
rect 477502 298658 477586 298894
rect 477822 298658 513266 298894
rect 513502 298658 513586 298894
rect 513822 298658 549266 298894
rect 549502 298658 549586 298894
rect 549822 298658 587262 298894
rect 587498 298658 587582 298894
rect 587818 298658 592650 298894
rect -8726 298574 592650 298658
rect -8726 298338 -3894 298574
rect -3658 298338 -3574 298574
rect -3338 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 369266 298574
rect 369502 298338 369586 298574
rect 369822 298338 405266 298574
rect 405502 298338 405586 298574
rect 405822 298338 441266 298574
rect 441502 298338 441586 298574
rect 441822 298338 477266 298574
rect 477502 298338 477586 298574
rect 477822 298338 513266 298574
rect 513502 298338 513586 298574
rect 513822 298338 549266 298574
rect 549502 298338 549586 298574
rect 549822 298338 587262 298574
rect 587498 298338 587582 298574
rect 587818 298338 592650 298574
rect -8726 298306 592650 298338
rect -8726 295174 592650 295206
rect -8726 294938 -2934 295174
rect -2698 294938 -2614 295174
rect -2378 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 39610 295174
rect 39846 294938 70330 295174
rect 70566 294938 101050 295174
rect 101286 294938 131770 295174
rect 132006 294938 162490 295174
rect 162726 294938 193210 295174
rect 193446 294938 223930 295174
rect 224166 294938 254650 295174
rect 254886 294938 285370 295174
rect 285606 294938 316090 295174
rect 316326 294938 346810 295174
rect 347046 294938 365546 295174
rect 365782 294938 365866 295174
rect 366102 294938 401546 295174
rect 401782 294938 401866 295174
rect 402102 294938 437546 295174
rect 437782 294938 437866 295174
rect 438102 294938 509546 295174
rect 509782 294938 509866 295174
rect 510102 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 586302 295174
rect 586538 294938 586622 295174
rect 586858 294938 592650 295174
rect -8726 294854 592650 294938
rect -8726 294618 -2934 294854
rect -2698 294618 -2614 294854
rect -2378 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 39610 294854
rect 39846 294618 70330 294854
rect 70566 294618 101050 294854
rect 101286 294618 131770 294854
rect 132006 294618 162490 294854
rect 162726 294618 193210 294854
rect 193446 294618 223930 294854
rect 224166 294618 254650 294854
rect 254886 294618 285370 294854
rect 285606 294618 316090 294854
rect 316326 294618 346810 294854
rect 347046 294618 365546 294854
rect 365782 294618 365866 294854
rect 366102 294618 401546 294854
rect 401782 294618 401866 294854
rect 402102 294618 437546 294854
rect 437782 294618 437866 294854
rect 438102 294618 509546 294854
rect 509782 294618 509866 294854
rect 510102 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 586302 294854
rect 586538 294618 586622 294854
rect 586858 294618 592650 294854
rect -8726 294586 592650 294618
rect -8726 291454 592650 291486
rect -8726 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 24250 291454
rect 24486 291218 54970 291454
rect 55206 291218 85690 291454
rect 85926 291218 116410 291454
rect 116646 291218 147130 291454
rect 147366 291218 177850 291454
rect 178086 291218 208570 291454
rect 208806 291218 239290 291454
rect 239526 291218 270010 291454
rect 270246 291218 300730 291454
rect 300966 291218 331450 291454
rect 331686 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 592650 291454
rect -8726 291134 592650 291218
rect -8726 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 24250 291134
rect 24486 290898 54970 291134
rect 55206 290898 85690 291134
rect 85926 290898 116410 291134
rect 116646 290898 147130 291134
rect 147366 290898 177850 291134
rect 178086 290898 208570 291134
rect 208806 290898 239290 291134
rect 239526 290898 270010 291134
rect 270246 290898 300730 291134
rect 300966 290898 331450 291134
rect 331686 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 592650 291134
rect -8726 290866 592650 290898
rect -8726 281494 592650 281526
rect -8726 281258 -8694 281494
rect -8458 281258 -8374 281494
rect -8138 281258 27866 281494
rect 28102 281258 28186 281494
rect 28422 281258 387866 281494
rect 388102 281258 388186 281494
rect 388422 281258 423866 281494
rect 424102 281258 424186 281494
rect 424422 281258 459866 281494
rect 460102 281258 460186 281494
rect 460422 281258 495866 281494
rect 496102 281258 496186 281494
rect 496422 281258 531866 281494
rect 532102 281258 532186 281494
rect 532422 281258 567866 281494
rect 568102 281258 568186 281494
rect 568422 281258 592062 281494
rect 592298 281258 592382 281494
rect 592618 281258 592650 281494
rect -8726 281174 592650 281258
rect -8726 280938 -8694 281174
rect -8458 280938 -8374 281174
rect -8138 280938 27866 281174
rect 28102 280938 28186 281174
rect 28422 280938 387866 281174
rect 388102 280938 388186 281174
rect 388422 280938 423866 281174
rect 424102 280938 424186 281174
rect 424422 280938 459866 281174
rect 460102 280938 460186 281174
rect 460422 280938 495866 281174
rect 496102 280938 496186 281174
rect 496422 280938 531866 281174
rect 532102 280938 532186 281174
rect 532422 280938 567866 281174
rect 568102 280938 568186 281174
rect 568422 280938 592062 281174
rect 592298 280938 592382 281174
rect 592618 280938 592650 281174
rect -8726 280906 592650 280938
rect -8726 277774 592650 277806
rect -8726 277538 -7734 277774
rect -7498 277538 -7414 277774
rect -7178 277538 384146 277774
rect 384382 277538 384466 277774
rect 384702 277538 420146 277774
rect 420382 277538 420466 277774
rect 420702 277538 456146 277774
rect 456382 277538 456466 277774
rect 456702 277538 492146 277774
rect 492382 277538 492466 277774
rect 492702 277538 528146 277774
rect 528382 277538 528466 277774
rect 528702 277538 564146 277774
rect 564382 277538 564466 277774
rect 564702 277538 591102 277774
rect 591338 277538 591422 277774
rect 591658 277538 592650 277774
rect -8726 277454 592650 277538
rect -8726 277218 -7734 277454
rect -7498 277218 -7414 277454
rect -7178 277218 384146 277454
rect 384382 277218 384466 277454
rect 384702 277218 420146 277454
rect 420382 277218 420466 277454
rect 420702 277218 456146 277454
rect 456382 277218 456466 277454
rect 456702 277218 492146 277454
rect 492382 277218 492466 277454
rect 492702 277218 528146 277454
rect 528382 277218 528466 277454
rect 528702 277218 564146 277454
rect 564382 277218 564466 277454
rect 564702 277218 591102 277454
rect 591338 277218 591422 277454
rect 591658 277218 592650 277454
rect -8726 277186 592650 277218
rect -8726 274054 592650 274086
rect -8726 273818 -6774 274054
rect -6538 273818 -6454 274054
rect -6218 273818 20426 274054
rect 20662 273818 20746 274054
rect 20982 273818 380426 274054
rect 380662 273818 380746 274054
rect 380982 273818 416426 274054
rect 416662 273818 416746 274054
rect 416982 273818 452426 274054
rect 452662 273818 452746 274054
rect 452982 273818 488426 274054
rect 488662 273818 488746 274054
rect 488982 273818 524426 274054
rect 524662 273818 524746 274054
rect 524982 273818 560426 274054
rect 560662 273818 560746 274054
rect 560982 273818 590142 274054
rect 590378 273818 590462 274054
rect 590698 273818 592650 274054
rect -8726 273734 592650 273818
rect -8726 273498 -6774 273734
rect -6538 273498 -6454 273734
rect -6218 273498 20426 273734
rect 20662 273498 20746 273734
rect 20982 273498 380426 273734
rect 380662 273498 380746 273734
rect 380982 273498 416426 273734
rect 416662 273498 416746 273734
rect 416982 273498 452426 273734
rect 452662 273498 452746 273734
rect 452982 273498 488426 273734
rect 488662 273498 488746 273734
rect 488982 273498 524426 273734
rect 524662 273498 524746 273734
rect 524982 273498 560426 273734
rect 560662 273498 560746 273734
rect 560982 273498 590142 273734
rect 590378 273498 590462 273734
rect 590698 273498 592650 273734
rect -8726 273466 592650 273498
rect -8726 270334 592650 270366
rect -8726 270098 -5814 270334
rect -5578 270098 -5494 270334
rect -5258 270098 16706 270334
rect 16942 270098 17026 270334
rect 17262 270098 376706 270334
rect 376942 270098 377026 270334
rect 377262 270098 412706 270334
rect 412942 270098 413026 270334
rect 413262 270098 448706 270334
rect 448942 270098 449026 270334
rect 449262 270098 484706 270334
rect 484942 270098 485026 270334
rect 485262 270098 520706 270334
rect 520942 270098 521026 270334
rect 521262 270098 556706 270334
rect 556942 270098 557026 270334
rect 557262 270098 589182 270334
rect 589418 270098 589502 270334
rect 589738 270098 592650 270334
rect -8726 270014 592650 270098
rect -8726 269778 -5814 270014
rect -5578 269778 -5494 270014
rect -5258 269778 16706 270014
rect 16942 269778 17026 270014
rect 17262 269778 376706 270014
rect 376942 269778 377026 270014
rect 377262 269778 412706 270014
rect 412942 269778 413026 270014
rect 413262 269778 448706 270014
rect 448942 269778 449026 270014
rect 449262 269778 484706 270014
rect 484942 269778 485026 270014
rect 485262 269778 520706 270014
rect 520942 269778 521026 270014
rect 521262 269778 556706 270014
rect 556942 269778 557026 270014
rect 557262 269778 589182 270014
rect 589418 269778 589502 270014
rect 589738 269778 592650 270014
rect -8726 269746 592650 269778
rect -8726 266614 592650 266646
rect -8726 266378 -4854 266614
rect -4618 266378 -4534 266614
rect -4298 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 372986 266614
rect 373222 266378 373306 266614
rect 373542 266378 408986 266614
rect 409222 266378 409306 266614
rect 409542 266378 444986 266614
rect 445222 266378 445306 266614
rect 445542 266378 480986 266614
rect 481222 266378 481306 266614
rect 481542 266378 516986 266614
rect 517222 266378 517306 266614
rect 517542 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 588222 266614
rect 588458 266378 588542 266614
rect 588778 266378 592650 266614
rect -8726 266294 592650 266378
rect -8726 266058 -4854 266294
rect -4618 266058 -4534 266294
rect -4298 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 372986 266294
rect 373222 266058 373306 266294
rect 373542 266058 408986 266294
rect 409222 266058 409306 266294
rect 409542 266058 444986 266294
rect 445222 266058 445306 266294
rect 445542 266058 480986 266294
rect 481222 266058 481306 266294
rect 481542 266058 516986 266294
rect 517222 266058 517306 266294
rect 517542 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 588222 266294
rect 588458 266058 588542 266294
rect 588778 266058 592650 266294
rect -8726 266026 592650 266058
rect -8726 262894 592650 262926
rect -8726 262658 -3894 262894
rect -3658 262658 -3574 262894
rect -3338 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 369266 262894
rect 369502 262658 369586 262894
rect 369822 262658 405266 262894
rect 405502 262658 405586 262894
rect 405822 262658 441266 262894
rect 441502 262658 441586 262894
rect 441822 262658 477266 262894
rect 477502 262658 477586 262894
rect 477822 262658 513266 262894
rect 513502 262658 513586 262894
rect 513822 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 587262 262894
rect 587498 262658 587582 262894
rect 587818 262658 592650 262894
rect -8726 262574 592650 262658
rect -8726 262338 -3894 262574
rect -3658 262338 -3574 262574
rect -3338 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 369266 262574
rect 369502 262338 369586 262574
rect 369822 262338 405266 262574
rect 405502 262338 405586 262574
rect 405822 262338 441266 262574
rect 441502 262338 441586 262574
rect 441822 262338 477266 262574
rect 477502 262338 477586 262574
rect 477822 262338 513266 262574
rect 513502 262338 513586 262574
rect 513822 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 587262 262574
rect 587498 262338 587582 262574
rect 587818 262338 592650 262574
rect -8726 262306 592650 262338
rect -8726 259174 592650 259206
rect -8726 258938 -2934 259174
rect -2698 258938 -2614 259174
rect -2378 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 39610 259174
rect 39846 258938 70330 259174
rect 70566 258938 101050 259174
rect 101286 258938 131770 259174
rect 132006 258938 162490 259174
rect 162726 258938 193210 259174
rect 193446 258938 223930 259174
rect 224166 258938 254650 259174
rect 254886 258938 285370 259174
rect 285606 258938 316090 259174
rect 316326 258938 346810 259174
rect 347046 258938 365546 259174
rect 365782 258938 365866 259174
rect 366102 258938 401546 259174
rect 401782 258938 401866 259174
rect 402102 258938 437546 259174
rect 437782 258938 437866 259174
rect 438102 258938 479610 259174
rect 479846 258938 510330 259174
rect 510566 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 586302 259174
rect 586538 258938 586622 259174
rect 586858 258938 592650 259174
rect -8726 258854 592650 258938
rect -8726 258618 -2934 258854
rect -2698 258618 -2614 258854
rect -2378 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 39610 258854
rect 39846 258618 70330 258854
rect 70566 258618 101050 258854
rect 101286 258618 131770 258854
rect 132006 258618 162490 258854
rect 162726 258618 193210 258854
rect 193446 258618 223930 258854
rect 224166 258618 254650 258854
rect 254886 258618 285370 258854
rect 285606 258618 316090 258854
rect 316326 258618 346810 258854
rect 347046 258618 365546 258854
rect 365782 258618 365866 258854
rect 366102 258618 401546 258854
rect 401782 258618 401866 258854
rect 402102 258618 437546 258854
rect 437782 258618 437866 258854
rect 438102 258618 479610 258854
rect 479846 258618 510330 258854
rect 510566 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 586302 258854
rect 586538 258618 586622 258854
rect 586858 258618 592650 258854
rect -8726 258586 592650 258618
rect -8726 255454 592650 255486
rect -8726 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 24250 255454
rect 24486 255218 54970 255454
rect 55206 255218 85690 255454
rect 85926 255218 116410 255454
rect 116646 255218 147130 255454
rect 147366 255218 177850 255454
rect 178086 255218 208570 255454
rect 208806 255218 239290 255454
rect 239526 255218 270010 255454
rect 270246 255218 300730 255454
rect 300966 255218 331450 255454
rect 331686 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 464250 255454
rect 464486 255218 494970 255454
rect 495206 255218 525690 255454
rect 525926 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 592650 255454
rect -8726 255134 592650 255218
rect -8726 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 24250 255134
rect 24486 254898 54970 255134
rect 55206 254898 85690 255134
rect 85926 254898 116410 255134
rect 116646 254898 147130 255134
rect 147366 254898 177850 255134
rect 178086 254898 208570 255134
rect 208806 254898 239290 255134
rect 239526 254898 270010 255134
rect 270246 254898 300730 255134
rect 300966 254898 331450 255134
rect 331686 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 464250 255134
rect 464486 254898 494970 255134
rect 495206 254898 525690 255134
rect 525926 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 592650 255134
rect -8726 254866 592650 254898
rect -8726 245494 592650 245526
rect -8726 245258 -8694 245494
rect -8458 245258 -8374 245494
rect -8138 245258 27866 245494
rect 28102 245258 28186 245494
rect 28422 245258 387866 245494
rect 388102 245258 388186 245494
rect 388422 245258 423866 245494
rect 424102 245258 424186 245494
rect 424422 245258 459866 245494
rect 460102 245258 460186 245494
rect 460422 245258 531866 245494
rect 532102 245258 532186 245494
rect 532422 245258 567866 245494
rect 568102 245258 568186 245494
rect 568422 245258 592062 245494
rect 592298 245258 592382 245494
rect 592618 245258 592650 245494
rect -8726 245174 592650 245258
rect -8726 244938 -8694 245174
rect -8458 244938 -8374 245174
rect -8138 244938 27866 245174
rect 28102 244938 28186 245174
rect 28422 244938 387866 245174
rect 388102 244938 388186 245174
rect 388422 244938 423866 245174
rect 424102 244938 424186 245174
rect 424422 244938 459866 245174
rect 460102 244938 460186 245174
rect 460422 244938 531866 245174
rect 532102 244938 532186 245174
rect 532422 244938 567866 245174
rect 568102 244938 568186 245174
rect 568422 244938 592062 245174
rect 592298 244938 592382 245174
rect 592618 244938 592650 245174
rect -8726 244906 592650 244938
rect -8726 241774 592650 241806
rect -8726 241538 -7734 241774
rect -7498 241538 -7414 241774
rect -7178 241538 384146 241774
rect 384382 241538 384466 241774
rect 384702 241538 420146 241774
rect 420382 241538 420466 241774
rect 420702 241538 456146 241774
rect 456382 241538 456466 241774
rect 456702 241538 564146 241774
rect 564382 241538 564466 241774
rect 564702 241538 591102 241774
rect 591338 241538 591422 241774
rect 591658 241538 592650 241774
rect -8726 241454 592650 241538
rect -8726 241218 -7734 241454
rect -7498 241218 -7414 241454
rect -7178 241218 384146 241454
rect 384382 241218 384466 241454
rect 384702 241218 420146 241454
rect 420382 241218 420466 241454
rect 420702 241218 456146 241454
rect 456382 241218 456466 241454
rect 456702 241218 564146 241454
rect 564382 241218 564466 241454
rect 564702 241218 591102 241454
rect 591338 241218 591422 241454
rect 591658 241218 592650 241454
rect -8726 241186 592650 241218
rect -8726 238054 592650 238086
rect -8726 237818 -6774 238054
rect -6538 237818 -6454 238054
rect -6218 237818 20426 238054
rect 20662 237818 20746 238054
rect 20982 237818 380426 238054
rect 380662 237818 380746 238054
rect 380982 237818 416426 238054
rect 416662 237818 416746 238054
rect 416982 237818 452426 238054
rect 452662 237818 452746 238054
rect 452982 237818 560426 238054
rect 560662 237818 560746 238054
rect 560982 237818 590142 238054
rect 590378 237818 590462 238054
rect 590698 237818 592650 238054
rect -8726 237734 592650 237818
rect -8726 237498 -6774 237734
rect -6538 237498 -6454 237734
rect -6218 237498 20426 237734
rect 20662 237498 20746 237734
rect 20982 237498 380426 237734
rect 380662 237498 380746 237734
rect 380982 237498 416426 237734
rect 416662 237498 416746 237734
rect 416982 237498 452426 237734
rect 452662 237498 452746 237734
rect 452982 237498 560426 237734
rect 560662 237498 560746 237734
rect 560982 237498 590142 237734
rect 590378 237498 590462 237734
rect 590698 237498 592650 237734
rect -8726 237466 592650 237498
rect -8726 234334 592650 234366
rect -8726 234098 -5814 234334
rect -5578 234098 -5494 234334
rect -5258 234098 16706 234334
rect 16942 234098 17026 234334
rect 17262 234098 376706 234334
rect 376942 234098 377026 234334
rect 377262 234098 412706 234334
rect 412942 234098 413026 234334
rect 413262 234098 448706 234334
rect 448942 234098 449026 234334
rect 449262 234098 556706 234334
rect 556942 234098 557026 234334
rect 557262 234098 589182 234334
rect 589418 234098 589502 234334
rect 589738 234098 592650 234334
rect -8726 234014 592650 234098
rect -8726 233778 -5814 234014
rect -5578 233778 -5494 234014
rect -5258 233778 16706 234014
rect 16942 233778 17026 234014
rect 17262 233778 376706 234014
rect 376942 233778 377026 234014
rect 377262 233778 412706 234014
rect 412942 233778 413026 234014
rect 413262 233778 448706 234014
rect 448942 233778 449026 234014
rect 449262 233778 556706 234014
rect 556942 233778 557026 234014
rect 557262 233778 589182 234014
rect 589418 233778 589502 234014
rect 589738 233778 592650 234014
rect -8726 233746 592650 233778
rect -8726 230614 592650 230646
rect -8726 230378 -4854 230614
rect -4618 230378 -4534 230614
rect -4298 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 372986 230614
rect 373222 230378 373306 230614
rect 373542 230378 408986 230614
rect 409222 230378 409306 230614
rect 409542 230378 444986 230614
rect 445222 230378 445306 230614
rect 445542 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 588222 230614
rect 588458 230378 588542 230614
rect 588778 230378 592650 230614
rect -8726 230294 592650 230378
rect -8726 230058 -4854 230294
rect -4618 230058 -4534 230294
rect -4298 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 372986 230294
rect 373222 230058 373306 230294
rect 373542 230058 408986 230294
rect 409222 230058 409306 230294
rect 409542 230058 444986 230294
rect 445222 230058 445306 230294
rect 445542 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 588222 230294
rect 588458 230058 588542 230294
rect 588778 230058 592650 230294
rect -8726 230026 592650 230058
rect -8726 226894 592650 226926
rect -8726 226658 -3894 226894
rect -3658 226658 -3574 226894
rect -3338 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 369266 226894
rect 369502 226658 369586 226894
rect 369822 226658 405266 226894
rect 405502 226658 405586 226894
rect 405822 226658 441266 226894
rect 441502 226658 441586 226894
rect 441822 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 587262 226894
rect 587498 226658 587582 226894
rect 587818 226658 592650 226894
rect -8726 226574 592650 226658
rect -8726 226338 -3894 226574
rect -3658 226338 -3574 226574
rect -3338 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 369266 226574
rect 369502 226338 369586 226574
rect 369822 226338 405266 226574
rect 405502 226338 405586 226574
rect 405822 226338 441266 226574
rect 441502 226338 441586 226574
rect 441822 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 587262 226574
rect 587498 226338 587582 226574
rect 587818 226338 592650 226574
rect -8726 226306 592650 226338
rect -8726 223174 592650 223206
rect -8726 222938 -2934 223174
rect -2698 222938 -2614 223174
rect -2378 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 39610 223174
rect 39846 222938 70330 223174
rect 70566 222938 101050 223174
rect 101286 222938 131770 223174
rect 132006 222938 162490 223174
rect 162726 222938 193210 223174
rect 193446 222938 223930 223174
rect 224166 222938 254650 223174
rect 254886 222938 285370 223174
rect 285606 222938 316090 223174
rect 316326 222938 346810 223174
rect 347046 222938 365546 223174
rect 365782 222938 365866 223174
rect 366102 222938 401546 223174
rect 401782 222938 401866 223174
rect 402102 222938 437546 223174
rect 437782 222938 437866 223174
rect 438102 222938 479610 223174
rect 479846 222938 510330 223174
rect 510566 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 586302 223174
rect 586538 222938 586622 223174
rect 586858 222938 592650 223174
rect -8726 222854 592650 222938
rect -8726 222618 -2934 222854
rect -2698 222618 -2614 222854
rect -2378 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 39610 222854
rect 39846 222618 70330 222854
rect 70566 222618 101050 222854
rect 101286 222618 131770 222854
rect 132006 222618 162490 222854
rect 162726 222618 193210 222854
rect 193446 222618 223930 222854
rect 224166 222618 254650 222854
rect 254886 222618 285370 222854
rect 285606 222618 316090 222854
rect 316326 222618 346810 222854
rect 347046 222618 365546 222854
rect 365782 222618 365866 222854
rect 366102 222618 401546 222854
rect 401782 222618 401866 222854
rect 402102 222618 437546 222854
rect 437782 222618 437866 222854
rect 438102 222618 479610 222854
rect 479846 222618 510330 222854
rect 510566 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 586302 222854
rect 586538 222618 586622 222854
rect 586858 222618 592650 222854
rect -8726 222586 592650 222618
rect -8726 219454 592650 219486
rect -8726 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 24250 219454
rect 24486 219218 54970 219454
rect 55206 219218 85690 219454
rect 85926 219218 116410 219454
rect 116646 219218 147130 219454
rect 147366 219218 177850 219454
rect 178086 219218 208570 219454
rect 208806 219218 239290 219454
rect 239526 219218 270010 219454
rect 270246 219218 300730 219454
rect 300966 219218 331450 219454
rect 331686 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 464250 219454
rect 464486 219218 494970 219454
rect 495206 219218 525690 219454
rect 525926 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 592650 219454
rect -8726 219134 592650 219218
rect -8726 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 24250 219134
rect 24486 218898 54970 219134
rect 55206 218898 85690 219134
rect 85926 218898 116410 219134
rect 116646 218898 147130 219134
rect 147366 218898 177850 219134
rect 178086 218898 208570 219134
rect 208806 218898 239290 219134
rect 239526 218898 270010 219134
rect 270246 218898 300730 219134
rect 300966 218898 331450 219134
rect 331686 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 464250 219134
rect 464486 218898 494970 219134
rect 495206 218898 525690 219134
rect 525926 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 592650 219134
rect -8726 218866 592650 218898
rect -8726 209494 592650 209526
rect -8726 209258 -8694 209494
rect -8458 209258 -8374 209494
rect -8138 209258 27866 209494
rect 28102 209258 28186 209494
rect 28422 209258 387866 209494
rect 388102 209258 388186 209494
rect 388422 209258 423866 209494
rect 424102 209258 424186 209494
rect 424422 209258 459866 209494
rect 460102 209258 460186 209494
rect 460422 209258 531866 209494
rect 532102 209258 532186 209494
rect 532422 209258 567866 209494
rect 568102 209258 568186 209494
rect 568422 209258 592062 209494
rect 592298 209258 592382 209494
rect 592618 209258 592650 209494
rect -8726 209174 592650 209258
rect -8726 208938 -8694 209174
rect -8458 208938 -8374 209174
rect -8138 208938 27866 209174
rect 28102 208938 28186 209174
rect 28422 208938 387866 209174
rect 388102 208938 388186 209174
rect 388422 208938 423866 209174
rect 424102 208938 424186 209174
rect 424422 208938 459866 209174
rect 460102 208938 460186 209174
rect 460422 208938 531866 209174
rect 532102 208938 532186 209174
rect 532422 208938 567866 209174
rect 568102 208938 568186 209174
rect 568422 208938 592062 209174
rect 592298 208938 592382 209174
rect 592618 208938 592650 209174
rect -8726 208906 592650 208938
rect -8726 205774 592650 205806
rect -8726 205538 -7734 205774
rect -7498 205538 -7414 205774
rect -7178 205538 384146 205774
rect 384382 205538 384466 205774
rect 384702 205538 420146 205774
rect 420382 205538 420466 205774
rect 420702 205538 456146 205774
rect 456382 205538 456466 205774
rect 456702 205538 564146 205774
rect 564382 205538 564466 205774
rect 564702 205538 591102 205774
rect 591338 205538 591422 205774
rect 591658 205538 592650 205774
rect -8726 205454 592650 205538
rect -8726 205218 -7734 205454
rect -7498 205218 -7414 205454
rect -7178 205218 384146 205454
rect 384382 205218 384466 205454
rect 384702 205218 420146 205454
rect 420382 205218 420466 205454
rect 420702 205218 456146 205454
rect 456382 205218 456466 205454
rect 456702 205218 564146 205454
rect 564382 205218 564466 205454
rect 564702 205218 591102 205454
rect 591338 205218 591422 205454
rect 591658 205218 592650 205454
rect -8726 205186 592650 205218
rect -8726 202054 592650 202086
rect -8726 201818 -6774 202054
rect -6538 201818 -6454 202054
rect -6218 201818 20426 202054
rect 20662 201818 20746 202054
rect 20982 201818 380426 202054
rect 380662 201818 380746 202054
rect 380982 201818 416426 202054
rect 416662 201818 416746 202054
rect 416982 201818 452426 202054
rect 452662 201818 452746 202054
rect 452982 201818 560426 202054
rect 560662 201818 560746 202054
rect 560982 201818 590142 202054
rect 590378 201818 590462 202054
rect 590698 201818 592650 202054
rect -8726 201734 592650 201818
rect -8726 201498 -6774 201734
rect -6538 201498 -6454 201734
rect -6218 201498 20426 201734
rect 20662 201498 20746 201734
rect 20982 201498 380426 201734
rect 380662 201498 380746 201734
rect 380982 201498 416426 201734
rect 416662 201498 416746 201734
rect 416982 201498 452426 201734
rect 452662 201498 452746 201734
rect 452982 201498 560426 201734
rect 560662 201498 560746 201734
rect 560982 201498 590142 201734
rect 590378 201498 590462 201734
rect 590698 201498 592650 201734
rect -8726 201466 592650 201498
rect -8726 198334 592650 198366
rect -8726 198098 -5814 198334
rect -5578 198098 -5494 198334
rect -5258 198098 16706 198334
rect 16942 198098 17026 198334
rect 17262 198098 376706 198334
rect 376942 198098 377026 198334
rect 377262 198098 412706 198334
rect 412942 198098 413026 198334
rect 413262 198098 448706 198334
rect 448942 198098 449026 198334
rect 449262 198098 484706 198334
rect 484942 198098 485026 198334
rect 485262 198098 520706 198334
rect 520942 198098 521026 198334
rect 521262 198098 556706 198334
rect 556942 198098 557026 198334
rect 557262 198098 589182 198334
rect 589418 198098 589502 198334
rect 589738 198098 592650 198334
rect -8726 198014 592650 198098
rect -8726 197778 -5814 198014
rect -5578 197778 -5494 198014
rect -5258 197778 16706 198014
rect 16942 197778 17026 198014
rect 17262 197778 376706 198014
rect 376942 197778 377026 198014
rect 377262 197778 412706 198014
rect 412942 197778 413026 198014
rect 413262 197778 448706 198014
rect 448942 197778 449026 198014
rect 449262 197778 484706 198014
rect 484942 197778 485026 198014
rect 485262 197778 520706 198014
rect 520942 197778 521026 198014
rect 521262 197778 556706 198014
rect 556942 197778 557026 198014
rect 557262 197778 589182 198014
rect 589418 197778 589502 198014
rect 589738 197778 592650 198014
rect -8726 197746 592650 197778
rect -8726 194614 592650 194646
rect -8726 194378 -4854 194614
rect -4618 194378 -4534 194614
rect -4298 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 372986 194614
rect 373222 194378 373306 194614
rect 373542 194378 408986 194614
rect 409222 194378 409306 194614
rect 409542 194378 444986 194614
rect 445222 194378 445306 194614
rect 445542 194378 480986 194614
rect 481222 194378 481306 194614
rect 481542 194378 516986 194614
rect 517222 194378 517306 194614
rect 517542 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 588222 194614
rect 588458 194378 588542 194614
rect 588778 194378 592650 194614
rect -8726 194294 592650 194378
rect -8726 194058 -4854 194294
rect -4618 194058 -4534 194294
rect -4298 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 372986 194294
rect 373222 194058 373306 194294
rect 373542 194058 408986 194294
rect 409222 194058 409306 194294
rect 409542 194058 444986 194294
rect 445222 194058 445306 194294
rect 445542 194058 480986 194294
rect 481222 194058 481306 194294
rect 481542 194058 516986 194294
rect 517222 194058 517306 194294
rect 517542 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 588222 194294
rect 588458 194058 588542 194294
rect 588778 194058 592650 194294
rect -8726 194026 592650 194058
rect -8726 190894 592650 190926
rect -8726 190658 -3894 190894
rect -3658 190658 -3574 190894
rect -3338 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 369266 190894
rect 369502 190658 369586 190894
rect 369822 190658 405266 190894
rect 405502 190658 405586 190894
rect 405822 190658 441266 190894
rect 441502 190658 441586 190894
rect 441822 190658 477266 190894
rect 477502 190658 477586 190894
rect 477822 190658 513266 190894
rect 513502 190658 513586 190894
rect 513822 190658 549266 190894
rect 549502 190658 549586 190894
rect 549822 190658 587262 190894
rect 587498 190658 587582 190894
rect 587818 190658 592650 190894
rect -8726 190574 592650 190658
rect -8726 190338 -3894 190574
rect -3658 190338 -3574 190574
rect -3338 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 369266 190574
rect 369502 190338 369586 190574
rect 369822 190338 405266 190574
rect 405502 190338 405586 190574
rect 405822 190338 441266 190574
rect 441502 190338 441586 190574
rect 441822 190338 477266 190574
rect 477502 190338 477586 190574
rect 477822 190338 513266 190574
rect 513502 190338 513586 190574
rect 513822 190338 549266 190574
rect 549502 190338 549586 190574
rect 549822 190338 587262 190574
rect 587498 190338 587582 190574
rect 587818 190338 592650 190574
rect -8726 190306 592650 190338
rect -8726 187174 592650 187206
rect -8726 186938 -2934 187174
rect -2698 186938 -2614 187174
rect -2378 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 39610 187174
rect 39846 186938 70330 187174
rect 70566 186938 101050 187174
rect 101286 186938 131770 187174
rect 132006 186938 162490 187174
rect 162726 186938 193210 187174
rect 193446 186938 223930 187174
rect 224166 186938 254650 187174
rect 254886 186938 285370 187174
rect 285606 186938 316090 187174
rect 316326 186938 346810 187174
rect 347046 186938 365546 187174
rect 365782 186938 365866 187174
rect 366102 186938 401546 187174
rect 401782 186938 401866 187174
rect 402102 186938 437546 187174
rect 437782 186938 437866 187174
rect 438102 186938 473546 187174
rect 473782 186938 473866 187174
rect 474102 186938 509546 187174
rect 509782 186938 509866 187174
rect 510102 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 586302 187174
rect 586538 186938 586622 187174
rect 586858 186938 592650 187174
rect -8726 186854 592650 186938
rect -8726 186618 -2934 186854
rect -2698 186618 -2614 186854
rect -2378 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 39610 186854
rect 39846 186618 70330 186854
rect 70566 186618 101050 186854
rect 101286 186618 131770 186854
rect 132006 186618 162490 186854
rect 162726 186618 193210 186854
rect 193446 186618 223930 186854
rect 224166 186618 254650 186854
rect 254886 186618 285370 186854
rect 285606 186618 316090 186854
rect 316326 186618 346810 186854
rect 347046 186618 365546 186854
rect 365782 186618 365866 186854
rect 366102 186618 401546 186854
rect 401782 186618 401866 186854
rect 402102 186618 437546 186854
rect 437782 186618 437866 186854
rect 438102 186618 473546 186854
rect 473782 186618 473866 186854
rect 474102 186618 509546 186854
rect 509782 186618 509866 186854
rect 510102 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 586302 186854
rect 586538 186618 586622 186854
rect 586858 186618 592650 186854
rect -8726 186586 592650 186618
rect -8726 183454 592650 183486
rect -8726 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 24250 183454
rect 24486 183218 54970 183454
rect 55206 183218 85690 183454
rect 85926 183218 116410 183454
rect 116646 183218 147130 183454
rect 147366 183218 177850 183454
rect 178086 183218 208570 183454
rect 208806 183218 239290 183454
rect 239526 183218 270010 183454
rect 270246 183218 300730 183454
rect 300966 183218 331450 183454
rect 331686 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 592650 183454
rect -8726 183134 592650 183218
rect -8726 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 24250 183134
rect 24486 182898 54970 183134
rect 55206 182898 85690 183134
rect 85926 182898 116410 183134
rect 116646 182898 147130 183134
rect 147366 182898 177850 183134
rect 178086 182898 208570 183134
rect 208806 182898 239290 183134
rect 239526 182898 270010 183134
rect 270246 182898 300730 183134
rect 300966 182898 331450 183134
rect 331686 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 592650 183134
rect -8726 182866 592650 182898
rect -8726 173494 592650 173526
rect -8726 173258 -8694 173494
rect -8458 173258 -8374 173494
rect -8138 173258 27866 173494
rect 28102 173258 28186 173494
rect 28422 173258 387866 173494
rect 388102 173258 388186 173494
rect 388422 173258 423866 173494
rect 424102 173258 424186 173494
rect 424422 173258 459866 173494
rect 460102 173258 460186 173494
rect 460422 173258 531866 173494
rect 532102 173258 532186 173494
rect 532422 173258 567866 173494
rect 568102 173258 568186 173494
rect 568422 173258 592062 173494
rect 592298 173258 592382 173494
rect 592618 173258 592650 173494
rect -8726 173174 592650 173258
rect -8726 172938 -8694 173174
rect -8458 172938 -8374 173174
rect -8138 172938 27866 173174
rect 28102 172938 28186 173174
rect 28422 172938 387866 173174
rect 388102 172938 388186 173174
rect 388422 172938 423866 173174
rect 424102 172938 424186 173174
rect 424422 172938 459866 173174
rect 460102 172938 460186 173174
rect 460422 172938 531866 173174
rect 532102 172938 532186 173174
rect 532422 172938 567866 173174
rect 568102 172938 568186 173174
rect 568422 172938 592062 173174
rect 592298 172938 592382 173174
rect 592618 172938 592650 173174
rect -8726 172906 592650 172938
rect -8726 169774 592650 169806
rect -8726 169538 -7734 169774
rect -7498 169538 -7414 169774
rect -7178 169538 384146 169774
rect 384382 169538 384466 169774
rect 384702 169538 420146 169774
rect 420382 169538 420466 169774
rect 420702 169538 456146 169774
rect 456382 169538 456466 169774
rect 456702 169538 564146 169774
rect 564382 169538 564466 169774
rect 564702 169538 591102 169774
rect 591338 169538 591422 169774
rect 591658 169538 592650 169774
rect -8726 169454 592650 169538
rect -8726 169218 -7734 169454
rect -7498 169218 -7414 169454
rect -7178 169218 384146 169454
rect 384382 169218 384466 169454
rect 384702 169218 420146 169454
rect 420382 169218 420466 169454
rect 420702 169218 456146 169454
rect 456382 169218 456466 169454
rect 456702 169218 564146 169454
rect 564382 169218 564466 169454
rect 564702 169218 591102 169454
rect 591338 169218 591422 169454
rect 591658 169218 592650 169454
rect -8726 169186 592650 169218
rect -8726 166054 592650 166086
rect -8726 165818 -6774 166054
rect -6538 165818 -6454 166054
rect -6218 165818 20426 166054
rect 20662 165818 20746 166054
rect 20982 165818 380426 166054
rect 380662 165818 380746 166054
rect 380982 165818 416426 166054
rect 416662 165818 416746 166054
rect 416982 165818 452426 166054
rect 452662 165818 452746 166054
rect 452982 165818 488426 166054
rect 488662 165818 488746 166054
rect 488982 165818 524426 166054
rect 524662 165818 524746 166054
rect 524982 165818 560426 166054
rect 560662 165818 560746 166054
rect 560982 165818 590142 166054
rect 590378 165818 590462 166054
rect 590698 165818 592650 166054
rect -8726 165734 592650 165818
rect -8726 165498 -6774 165734
rect -6538 165498 -6454 165734
rect -6218 165498 20426 165734
rect 20662 165498 20746 165734
rect 20982 165498 380426 165734
rect 380662 165498 380746 165734
rect 380982 165498 416426 165734
rect 416662 165498 416746 165734
rect 416982 165498 452426 165734
rect 452662 165498 452746 165734
rect 452982 165498 488426 165734
rect 488662 165498 488746 165734
rect 488982 165498 524426 165734
rect 524662 165498 524746 165734
rect 524982 165498 560426 165734
rect 560662 165498 560746 165734
rect 560982 165498 590142 165734
rect 590378 165498 590462 165734
rect 590698 165498 592650 165734
rect -8726 165466 592650 165498
rect -8726 162334 592650 162366
rect -8726 162098 -5814 162334
rect -5578 162098 -5494 162334
rect -5258 162098 16706 162334
rect 16942 162098 17026 162334
rect 17262 162098 376706 162334
rect 376942 162098 377026 162334
rect 377262 162098 412706 162334
rect 412942 162098 413026 162334
rect 413262 162098 448706 162334
rect 448942 162098 449026 162334
rect 449262 162098 484706 162334
rect 484942 162098 485026 162334
rect 485262 162098 520706 162334
rect 520942 162098 521026 162334
rect 521262 162098 556706 162334
rect 556942 162098 557026 162334
rect 557262 162098 589182 162334
rect 589418 162098 589502 162334
rect 589738 162098 592650 162334
rect -8726 162014 592650 162098
rect -8726 161778 -5814 162014
rect -5578 161778 -5494 162014
rect -5258 161778 16706 162014
rect 16942 161778 17026 162014
rect 17262 161778 376706 162014
rect 376942 161778 377026 162014
rect 377262 161778 412706 162014
rect 412942 161778 413026 162014
rect 413262 161778 448706 162014
rect 448942 161778 449026 162014
rect 449262 161778 484706 162014
rect 484942 161778 485026 162014
rect 485262 161778 520706 162014
rect 520942 161778 521026 162014
rect 521262 161778 556706 162014
rect 556942 161778 557026 162014
rect 557262 161778 589182 162014
rect 589418 161778 589502 162014
rect 589738 161778 592650 162014
rect -8726 161746 592650 161778
rect -8726 158614 592650 158646
rect -8726 158378 -4854 158614
rect -4618 158378 -4534 158614
rect -4298 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 372986 158614
rect 373222 158378 373306 158614
rect 373542 158378 408986 158614
rect 409222 158378 409306 158614
rect 409542 158378 480986 158614
rect 481222 158378 481306 158614
rect 481542 158378 516986 158614
rect 517222 158378 517306 158614
rect 517542 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 588222 158614
rect 588458 158378 588542 158614
rect 588778 158378 592650 158614
rect -8726 158294 592650 158378
rect -8726 158058 -4854 158294
rect -4618 158058 -4534 158294
rect -4298 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 372986 158294
rect 373222 158058 373306 158294
rect 373542 158058 408986 158294
rect 409222 158058 409306 158294
rect 409542 158058 480986 158294
rect 481222 158058 481306 158294
rect 481542 158058 516986 158294
rect 517222 158058 517306 158294
rect 517542 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 588222 158294
rect 588458 158058 588542 158294
rect 588778 158058 592650 158294
rect -8726 158026 592650 158058
rect -8726 154894 592650 154926
rect -8726 154658 -3894 154894
rect -3658 154658 -3574 154894
rect -3338 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 369266 154894
rect 369502 154658 369586 154894
rect 369822 154658 405266 154894
rect 405502 154658 405586 154894
rect 405822 154658 477266 154894
rect 477502 154658 477586 154894
rect 477822 154658 513266 154894
rect 513502 154658 513586 154894
rect 513822 154658 549266 154894
rect 549502 154658 549586 154894
rect 549822 154658 587262 154894
rect 587498 154658 587582 154894
rect 587818 154658 592650 154894
rect -8726 154574 592650 154658
rect -8726 154338 -3894 154574
rect -3658 154338 -3574 154574
rect -3338 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 369266 154574
rect 369502 154338 369586 154574
rect 369822 154338 405266 154574
rect 405502 154338 405586 154574
rect 405822 154338 477266 154574
rect 477502 154338 477586 154574
rect 477822 154338 513266 154574
rect 513502 154338 513586 154574
rect 513822 154338 549266 154574
rect 549502 154338 549586 154574
rect 549822 154338 587262 154574
rect 587498 154338 587582 154574
rect 587818 154338 592650 154574
rect -8726 154306 592650 154338
rect -8726 151174 592650 151206
rect -8726 150938 -2934 151174
rect -2698 150938 -2614 151174
rect -2378 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 39610 151174
rect 39846 150938 70330 151174
rect 70566 150938 101050 151174
rect 101286 150938 131770 151174
rect 132006 150938 162490 151174
rect 162726 150938 193210 151174
rect 193446 150938 223930 151174
rect 224166 150938 254650 151174
rect 254886 150938 285370 151174
rect 285606 150938 316090 151174
rect 316326 150938 346810 151174
rect 347046 150938 365546 151174
rect 365782 150938 365866 151174
rect 366102 150938 401546 151174
rect 401782 150938 401866 151174
rect 402102 150938 429610 151174
rect 429846 150938 473546 151174
rect 473782 150938 473866 151174
rect 474102 150938 509546 151174
rect 509782 150938 509866 151174
rect 510102 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 586302 151174
rect 586538 150938 586622 151174
rect 586858 150938 592650 151174
rect -8726 150854 592650 150938
rect -8726 150618 -2934 150854
rect -2698 150618 -2614 150854
rect -2378 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 39610 150854
rect 39846 150618 70330 150854
rect 70566 150618 101050 150854
rect 101286 150618 131770 150854
rect 132006 150618 162490 150854
rect 162726 150618 193210 150854
rect 193446 150618 223930 150854
rect 224166 150618 254650 150854
rect 254886 150618 285370 150854
rect 285606 150618 316090 150854
rect 316326 150618 346810 150854
rect 347046 150618 365546 150854
rect 365782 150618 365866 150854
rect 366102 150618 401546 150854
rect 401782 150618 401866 150854
rect 402102 150618 429610 150854
rect 429846 150618 473546 150854
rect 473782 150618 473866 150854
rect 474102 150618 509546 150854
rect 509782 150618 509866 150854
rect 510102 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 586302 150854
rect 586538 150618 586622 150854
rect 586858 150618 592650 150854
rect -8726 150586 592650 150618
rect -8726 147454 592650 147486
rect -8726 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 24250 147454
rect 24486 147218 54970 147454
rect 55206 147218 85690 147454
rect 85926 147218 116410 147454
rect 116646 147218 147130 147454
rect 147366 147218 177850 147454
rect 178086 147218 208570 147454
rect 208806 147218 239290 147454
rect 239526 147218 270010 147454
rect 270246 147218 300730 147454
rect 300966 147218 331450 147454
rect 331686 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 414250 147454
rect 414486 147218 444970 147454
rect 445206 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 592650 147454
rect -8726 147134 592650 147218
rect -8726 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 24250 147134
rect 24486 146898 54970 147134
rect 55206 146898 85690 147134
rect 85926 146898 116410 147134
rect 116646 146898 147130 147134
rect 147366 146898 177850 147134
rect 178086 146898 208570 147134
rect 208806 146898 239290 147134
rect 239526 146898 270010 147134
rect 270246 146898 300730 147134
rect 300966 146898 331450 147134
rect 331686 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 414250 147134
rect 414486 146898 444970 147134
rect 445206 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 592650 147134
rect -8726 146866 592650 146898
rect -8726 137494 592650 137526
rect -8726 137258 -8694 137494
rect -8458 137258 -8374 137494
rect -8138 137258 27866 137494
rect 28102 137258 28186 137494
rect 28422 137258 387866 137494
rect 388102 137258 388186 137494
rect 388422 137258 459866 137494
rect 460102 137258 460186 137494
rect 460422 137258 567866 137494
rect 568102 137258 568186 137494
rect 568422 137258 592062 137494
rect 592298 137258 592382 137494
rect 592618 137258 592650 137494
rect -8726 137174 592650 137258
rect -8726 136938 -8694 137174
rect -8458 136938 -8374 137174
rect -8138 136938 27866 137174
rect 28102 136938 28186 137174
rect 28422 136938 387866 137174
rect 388102 136938 388186 137174
rect 388422 136938 459866 137174
rect 460102 136938 460186 137174
rect 460422 136938 567866 137174
rect 568102 136938 568186 137174
rect 568422 136938 592062 137174
rect 592298 136938 592382 137174
rect 592618 136938 592650 137174
rect -8726 136906 592650 136938
rect -8726 133774 592650 133806
rect -8726 133538 -7734 133774
rect -7498 133538 -7414 133774
rect -7178 133538 384146 133774
rect 384382 133538 384466 133774
rect 384702 133538 456146 133774
rect 456382 133538 456466 133774
rect 456702 133538 564146 133774
rect 564382 133538 564466 133774
rect 564702 133538 591102 133774
rect 591338 133538 591422 133774
rect 591658 133538 592650 133774
rect -8726 133454 592650 133538
rect -8726 133218 -7734 133454
rect -7498 133218 -7414 133454
rect -7178 133218 384146 133454
rect 384382 133218 384466 133454
rect 384702 133218 456146 133454
rect 456382 133218 456466 133454
rect 456702 133218 564146 133454
rect 564382 133218 564466 133454
rect 564702 133218 591102 133454
rect 591338 133218 591422 133454
rect 591658 133218 592650 133454
rect -8726 133186 592650 133218
rect -8726 130054 592650 130086
rect -8726 129818 -6774 130054
rect -6538 129818 -6454 130054
rect -6218 129818 20426 130054
rect 20662 129818 20746 130054
rect 20982 129818 380426 130054
rect 380662 129818 380746 130054
rect 380982 129818 452426 130054
rect 452662 129818 452746 130054
rect 452982 129818 560426 130054
rect 560662 129818 560746 130054
rect 560982 129818 590142 130054
rect 590378 129818 590462 130054
rect 590698 129818 592650 130054
rect -8726 129734 592650 129818
rect -8726 129498 -6774 129734
rect -6538 129498 -6454 129734
rect -6218 129498 20426 129734
rect 20662 129498 20746 129734
rect 20982 129498 380426 129734
rect 380662 129498 380746 129734
rect 380982 129498 452426 129734
rect 452662 129498 452746 129734
rect 452982 129498 560426 129734
rect 560662 129498 560746 129734
rect 560982 129498 590142 129734
rect 590378 129498 590462 129734
rect 590698 129498 592650 129734
rect -8726 129466 592650 129498
rect -8726 126334 592650 126366
rect -8726 126098 -5814 126334
rect -5578 126098 -5494 126334
rect -5258 126098 16706 126334
rect 16942 126098 17026 126334
rect 17262 126098 376706 126334
rect 376942 126098 377026 126334
rect 377262 126098 412706 126334
rect 412942 126098 413026 126334
rect 413262 126098 448706 126334
rect 448942 126098 449026 126334
rect 449262 126098 484706 126334
rect 484942 126098 485026 126334
rect 485262 126098 556706 126334
rect 556942 126098 557026 126334
rect 557262 126098 589182 126334
rect 589418 126098 589502 126334
rect 589738 126098 592650 126334
rect -8726 126014 592650 126098
rect -8726 125778 -5814 126014
rect -5578 125778 -5494 126014
rect -5258 125778 16706 126014
rect 16942 125778 17026 126014
rect 17262 125778 376706 126014
rect 376942 125778 377026 126014
rect 377262 125778 412706 126014
rect 412942 125778 413026 126014
rect 413262 125778 448706 126014
rect 448942 125778 449026 126014
rect 449262 125778 484706 126014
rect 484942 125778 485026 126014
rect 485262 125778 556706 126014
rect 556942 125778 557026 126014
rect 557262 125778 589182 126014
rect 589418 125778 589502 126014
rect 589738 125778 592650 126014
rect -8726 125746 592650 125778
rect -8726 122614 592650 122646
rect -8726 122378 -4854 122614
rect -4618 122378 -4534 122614
rect -4298 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 372986 122614
rect 373222 122378 373306 122614
rect 373542 122378 408986 122614
rect 409222 122378 409306 122614
rect 409542 122378 480986 122614
rect 481222 122378 481306 122614
rect 481542 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 588222 122614
rect 588458 122378 588542 122614
rect 588778 122378 592650 122614
rect -8726 122294 592650 122378
rect -8726 122058 -4854 122294
rect -4618 122058 -4534 122294
rect -4298 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 372986 122294
rect 373222 122058 373306 122294
rect 373542 122058 408986 122294
rect 409222 122058 409306 122294
rect 409542 122058 480986 122294
rect 481222 122058 481306 122294
rect 481542 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 588222 122294
rect 588458 122058 588542 122294
rect 588778 122058 592650 122294
rect -8726 122026 592650 122058
rect -8726 118894 592650 118926
rect -8726 118658 -3894 118894
rect -3658 118658 -3574 118894
rect -3338 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 369266 118894
rect 369502 118658 369586 118894
rect 369822 118658 405266 118894
rect 405502 118658 405586 118894
rect 405822 118658 441266 118894
rect 441502 118658 441586 118894
rect 441822 118658 477266 118894
rect 477502 118658 477586 118894
rect 477822 118658 549266 118894
rect 549502 118658 549586 118894
rect 549822 118658 587262 118894
rect 587498 118658 587582 118894
rect 587818 118658 592650 118894
rect -8726 118574 592650 118658
rect -8726 118338 -3894 118574
rect -3658 118338 -3574 118574
rect -3338 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 369266 118574
rect 369502 118338 369586 118574
rect 369822 118338 405266 118574
rect 405502 118338 405586 118574
rect 405822 118338 441266 118574
rect 441502 118338 441586 118574
rect 441822 118338 477266 118574
rect 477502 118338 477586 118574
rect 477822 118338 549266 118574
rect 549502 118338 549586 118574
rect 549822 118338 587262 118574
rect 587498 118338 587582 118574
rect 587818 118338 592650 118574
rect -8726 118306 592650 118338
rect -8726 115174 592650 115206
rect -8726 114938 -2934 115174
rect -2698 114938 -2614 115174
rect -2378 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 39610 115174
rect 39846 114938 70330 115174
rect 70566 114938 101050 115174
rect 101286 114938 131770 115174
rect 132006 114938 162490 115174
rect 162726 114938 193210 115174
rect 193446 114938 223930 115174
rect 224166 114938 254650 115174
rect 254886 114938 285370 115174
rect 285606 114938 316090 115174
rect 316326 114938 346810 115174
rect 347046 114938 365546 115174
rect 365782 114938 365866 115174
rect 366102 114938 401546 115174
rect 401782 114938 401866 115174
rect 402102 114938 437546 115174
rect 437782 114938 437866 115174
rect 438102 114938 473546 115174
rect 473782 114938 473866 115174
rect 474102 114938 499610 115174
rect 499846 114938 530330 115174
rect 530566 114938 545546 115174
rect 545782 114938 545866 115174
rect 546102 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 586302 115174
rect 586538 114938 586622 115174
rect 586858 114938 592650 115174
rect -8726 114854 592650 114938
rect -8726 114618 -2934 114854
rect -2698 114618 -2614 114854
rect -2378 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 39610 114854
rect 39846 114618 70330 114854
rect 70566 114618 101050 114854
rect 101286 114618 131770 114854
rect 132006 114618 162490 114854
rect 162726 114618 193210 114854
rect 193446 114618 223930 114854
rect 224166 114618 254650 114854
rect 254886 114618 285370 114854
rect 285606 114618 316090 114854
rect 316326 114618 346810 114854
rect 347046 114618 365546 114854
rect 365782 114618 365866 114854
rect 366102 114618 401546 114854
rect 401782 114618 401866 114854
rect 402102 114618 437546 114854
rect 437782 114618 437866 114854
rect 438102 114618 473546 114854
rect 473782 114618 473866 114854
rect 474102 114618 499610 114854
rect 499846 114618 530330 114854
rect 530566 114618 545546 114854
rect 545782 114618 545866 114854
rect 546102 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 586302 114854
rect 586538 114618 586622 114854
rect 586858 114618 592650 114854
rect -8726 114586 592650 114618
rect -8726 111454 592650 111486
rect -8726 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 24250 111454
rect 24486 111218 54970 111454
rect 55206 111218 85690 111454
rect 85926 111218 116410 111454
rect 116646 111218 147130 111454
rect 147366 111218 177850 111454
rect 178086 111218 208570 111454
rect 208806 111218 239290 111454
rect 239526 111218 270010 111454
rect 270246 111218 300730 111454
rect 300966 111218 331450 111454
rect 331686 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 484250 111454
rect 484486 111218 514970 111454
rect 515206 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 592650 111454
rect -8726 111134 592650 111218
rect -8726 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 24250 111134
rect 24486 110898 54970 111134
rect 55206 110898 85690 111134
rect 85926 110898 116410 111134
rect 116646 110898 147130 111134
rect 147366 110898 177850 111134
rect 178086 110898 208570 111134
rect 208806 110898 239290 111134
rect 239526 110898 270010 111134
rect 270246 110898 300730 111134
rect 300966 110898 331450 111134
rect 331686 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 484250 111134
rect 484486 110898 514970 111134
rect 515206 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 592650 111134
rect -8726 110866 592650 110898
rect -8726 101494 592650 101526
rect -8726 101258 -8694 101494
rect -8458 101258 -8374 101494
rect -8138 101258 27866 101494
rect 28102 101258 28186 101494
rect 28422 101258 387866 101494
rect 388102 101258 388186 101494
rect 388422 101258 423866 101494
rect 424102 101258 424186 101494
rect 424422 101258 459866 101494
rect 460102 101258 460186 101494
rect 460422 101258 567866 101494
rect 568102 101258 568186 101494
rect 568422 101258 592062 101494
rect 592298 101258 592382 101494
rect 592618 101258 592650 101494
rect -8726 101174 592650 101258
rect -8726 100938 -8694 101174
rect -8458 100938 -8374 101174
rect -8138 100938 27866 101174
rect 28102 100938 28186 101174
rect 28422 100938 387866 101174
rect 388102 100938 388186 101174
rect 388422 100938 423866 101174
rect 424102 100938 424186 101174
rect 424422 100938 459866 101174
rect 460102 100938 460186 101174
rect 460422 100938 567866 101174
rect 568102 100938 568186 101174
rect 568422 100938 592062 101174
rect 592298 100938 592382 101174
rect 592618 100938 592650 101174
rect -8726 100906 592650 100938
rect -8726 97774 592650 97806
rect -8726 97538 -7734 97774
rect -7498 97538 -7414 97774
rect -7178 97538 384146 97774
rect 384382 97538 384466 97774
rect 384702 97538 420146 97774
rect 420382 97538 420466 97774
rect 420702 97538 456146 97774
rect 456382 97538 456466 97774
rect 456702 97538 564146 97774
rect 564382 97538 564466 97774
rect 564702 97538 591102 97774
rect 591338 97538 591422 97774
rect 591658 97538 592650 97774
rect -8726 97454 592650 97538
rect -8726 97218 -7734 97454
rect -7498 97218 -7414 97454
rect -7178 97218 384146 97454
rect 384382 97218 384466 97454
rect 384702 97218 420146 97454
rect 420382 97218 420466 97454
rect 420702 97218 456146 97454
rect 456382 97218 456466 97454
rect 456702 97218 564146 97454
rect 564382 97218 564466 97454
rect 564702 97218 591102 97454
rect 591338 97218 591422 97454
rect 591658 97218 592650 97454
rect -8726 97186 592650 97218
rect -8726 94054 592650 94086
rect -8726 93818 -6774 94054
rect -6538 93818 -6454 94054
rect -6218 93818 20426 94054
rect 20662 93818 20746 94054
rect 20982 93818 380426 94054
rect 380662 93818 380746 94054
rect 380982 93818 416426 94054
rect 416662 93818 416746 94054
rect 416982 93818 452426 94054
rect 452662 93818 452746 94054
rect 452982 93818 560426 94054
rect 560662 93818 560746 94054
rect 560982 93818 590142 94054
rect 590378 93818 590462 94054
rect 590698 93818 592650 94054
rect -8726 93734 592650 93818
rect -8726 93498 -6774 93734
rect -6538 93498 -6454 93734
rect -6218 93498 20426 93734
rect 20662 93498 20746 93734
rect 20982 93498 380426 93734
rect 380662 93498 380746 93734
rect 380982 93498 416426 93734
rect 416662 93498 416746 93734
rect 416982 93498 452426 93734
rect 452662 93498 452746 93734
rect 452982 93498 560426 93734
rect 560662 93498 560746 93734
rect 560982 93498 590142 93734
rect 590378 93498 590462 93734
rect 590698 93498 592650 93734
rect -8726 93466 592650 93498
rect -8726 90334 592650 90366
rect -8726 90098 -5814 90334
rect -5578 90098 -5494 90334
rect -5258 90098 16706 90334
rect 16942 90098 17026 90334
rect 17262 90098 376706 90334
rect 376942 90098 377026 90334
rect 377262 90098 412706 90334
rect 412942 90098 413026 90334
rect 413262 90098 448706 90334
rect 448942 90098 449026 90334
rect 449262 90098 484706 90334
rect 484942 90098 485026 90334
rect 485262 90098 556706 90334
rect 556942 90098 557026 90334
rect 557262 90098 589182 90334
rect 589418 90098 589502 90334
rect 589738 90098 592650 90334
rect -8726 90014 592650 90098
rect -8726 89778 -5814 90014
rect -5578 89778 -5494 90014
rect -5258 89778 16706 90014
rect 16942 89778 17026 90014
rect 17262 89778 376706 90014
rect 376942 89778 377026 90014
rect 377262 89778 412706 90014
rect 412942 89778 413026 90014
rect 413262 89778 448706 90014
rect 448942 89778 449026 90014
rect 449262 89778 484706 90014
rect 484942 89778 485026 90014
rect 485262 89778 556706 90014
rect 556942 89778 557026 90014
rect 557262 89778 589182 90014
rect 589418 89778 589502 90014
rect 589738 89778 592650 90014
rect -8726 89746 592650 89778
rect -8726 86614 592650 86646
rect -8726 86378 -4854 86614
rect -4618 86378 -4534 86614
rect -4298 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 372986 86614
rect 373222 86378 373306 86614
rect 373542 86378 408986 86614
rect 409222 86378 409306 86614
rect 409542 86378 444986 86614
rect 445222 86378 445306 86614
rect 445542 86378 480986 86614
rect 481222 86378 481306 86614
rect 481542 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 588222 86614
rect 588458 86378 588542 86614
rect 588778 86378 592650 86614
rect -8726 86294 592650 86378
rect -8726 86058 -4854 86294
rect -4618 86058 -4534 86294
rect -4298 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 372986 86294
rect 373222 86058 373306 86294
rect 373542 86058 408986 86294
rect 409222 86058 409306 86294
rect 409542 86058 444986 86294
rect 445222 86058 445306 86294
rect 445542 86058 480986 86294
rect 481222 86058 481306 86294
rect 481542 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 588222 86294
rect 588458 86058 588542 86294
rect 588778 86058 592650 86294
rect -8726 86026 592650 86058
rect -8726 82894 592650 82926
rect -8726 82658 -3894 82894
rect -3658 82658 -3574 82894
rect -3338 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 369266 82894
rect 369502 82658 369586 82894
rect 369822 82658 405266 82894
rect 405502 82658 405586 82894
rect 405822 82658 441266 82894
rect 441502 82658 441586 82894
rect 441822 82658 477266 82894
rect 477502 82658 477586 82894
rect 477822 82658 549266 82894
rect 549502 82658 549586 82894
rect 549822 82658 587262 82894
rect 587498 82658 587582 82894
rect 587818 82658 592650 82894
rect -8726 82574 592650 82658
rect -8726 82338 -3894 82574
rect -3658 82338 -3574 82574
rect -3338 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 369266 82574
rect 369502 82338 369586 82574
rect 369822 82338 405266 82574
rect 405502 82338 405586 82574
rect 405822 82338 441266 82574
rect 441502 82338 441586 82574
rect 441822 82338 477266 82574
rect 477502 82338 477586 82574
rect 477822 82338 549266 82574
rect 549502 82338 549586 82574
rect 549822 82338 587262 82574
rect 587498 82338 587582 82574
rect 587818 82338 592650 82574
rect -8726 82306 592650 82338
rect -8726 79174 592650 79206
rect -8726 78938 -2934 79174
rect -2698 78938 -2614 79174
rect -2378 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 39610 79174
rect 39846 78938 70330 79174
rect 70566 78938 101050 79174
rect 101286 78938 131770 79174
rect 132006 78938 162490 79174
rect 162726 78938 193210 79174
rect 193446 78938 223930 79174
rect 224166 78938 254650 79174
rect 254886 78938 285370 79174
rect 285606 78938 316090 79174
rect 316326 78938 346810 79174
rect 347046 78938 365546 79174
rect 365782 78938 365866 79174
rect 366102 78938 401546 79174
rect 401782 78938 401866 79174
rect 402102 78938 437546 79174
rect 437782 78938 437866 79174
rect 438102 78938 473546 79174
rect 473782 78938 473866 79174
rect 474102 78938 509546 79174
rect 509782 78938 509866 79174
rect 510102 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 586302 79174
rect 586538 78938 586622 79174
rect 586858 78938 592650 79174
rect -8726 78854 592650 78938
rect -8726 78618 -2934 78854
rect -2698 78618 -2614 78854
rect -2378 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 39610 78854
rect 39846 78618 70330 78854
rect 70566 78618 101050 78854
rect 101286 78618 131770 78854
rect 132006 78618 162490 78854
rect 162726 78618 193210 78854
rect 193446 78618 223930 78854
rect 224166 78618 254650 78854
rect 254886 78618 285370 78854
rect 285606 78618 316090 78854
rect 316326 78618 346810 78854
rect 347046 78618 365546 78854
rect 365782 78618 365866 78854
rect 366102 78618 401546 78854
rect 401782 78618 401866 78854
rect 402102 78618 437546 78854
rect 437782 78618 437866 78854
rect 438102 78618 473546 78854
rect 473782 78618 473866 78854
rect 474102 78618 509546 78854
rect 509782 78618 509866 78854
rect 510102 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 586302 78854
rect 586538 78618 586622 78854
rect 586858 78618 592650 78854
rect -8726 78586 592650 78618
rect -8726 75454 592650 75486
rect -8726 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 24250 75454
rect 24486 75218 54970 75454
rect 55206 75218 85690 75454
rect 85926 75218 116410 75454
rect 116646 75218 147130 75454
rect 147366 75218 177850 75454
rect 178086 75218 208570 75454
rect 208806 75218 239290 75454
rect 239526 75218 270010 75454
rect 270246 75218 300730 75454
rect 300966 75218 331450 75454
rect 331686 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 592650 75454
rect -8726 75134 592650 75218
rect -8726 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 24250 75134
rect 24486 74898 54970 75134
rect 55206 74898 85690 75134
rect 85926 74898 116410 75134
rect 116646 74898 147130 75134
rect 147366 74898 177850 75134
rect 178086 74898 208570 75134
rect 208806 74898 239290 75134
rect 239526 74898 270010 75134
rect 270246 74898 300730 75134
rect 300966 74898 331450 75134
rect 331686 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 592650 75134
rect -8726 74866 592650 74898
rect -8726 65494 592650 65526
rect -8726 65258 -8694 65494
rect -8458 65258 -8374 65494
rect -8138 65258 27866 65494
rect 28102 65258 28186 65494
rect 28422 65258 387866 65494
rect 388102 65258 388186 65494
rect 388422 65258 423866 65494
rect 424102 65258 424186 65494
rect 424422 65258 459866 65494
rect 460102 65258 460186 65494
rect 460422 65258 495866 65494
rect 496102 65258 496186 65494
rect 496422 65258 531866 65494
rect 532102 65258 532186 65494
rect 532422 65258 567866 65494
rect 568102 65258 568186 65494
rect 568422 65258 592062 65494
rect 592298 65258 592382 65494
rect 592618 65258 592650 65494
rect -8726 65174 592650 65258
rect -8726 64938 -8694 65174
rect -8458 64938 -8374 65174
rect -8138 64938 27866 65174
rect 28102 64938 28186 65174
rect 28422 64938 387866 65174
rect 388102 64938 388186 65174
rect 388422 64938 423866 65174
rect 424102 64938 424186 65174
rect 424422 64938 459866 65174
rect 460102 64938 460186 65174
rect 460422 64938 495866 65174
rect 496102 64938 496186 65174
rect 496422 64938 531866 65174
rect 532102 64938 532186 65174
rect 532422 64938 567866 65174
rect 568102 64938 568186 65174
rect 568422 64938 592062 65174
rect 592298 64938 592382 65174
rect 592618 64938 592650 65174
rect -8726 64906 592650 64938
rect -8726 61774 592650 61806
rect -8726 61538 -7734 61774
rect -7498 61538 -7414 61774
rect -7178 61538 384146 61774
rect 384382 61538 384466 61774
rect 384702 61538 420146 61774
rect 420382 61538 420466 61774
rect 420702 61538 456146 61774
rect 456382 61538 456466 61774
rect 456702 61538 492146 61774
rect 492382 61538 492466 61774
rect 492702 61538 528146 61774
rect 528382 61538 528466 61774
rect 528702 61538 564146 61774
rect 564382 61538 564466 61774
rect 564702 61538 591102 61774
rect 591338 61538 591422 61774
rect 591658 61538 592650 61774
rect -8726 61454 592650 61538
rect -8726 61218 -7734 61454
rect -7498 61218 -7414 61454
rect -7178 61218 384146 61454
rect 384382 61218 384466 61454
rect 384702 61218 420146 61454
rect 420382 61218 420466 61454
rect 420702 61218 456146 61454
rect 456382 61218 456466 61454
rect 456702 61218 492146 61454
rect 492382 61218 492466 61454
rect 492702 61218 528146 61454
rect 528382 61218 528466 61454
rect 528702 61218 564146 61454
rect 564382 61218 564466 61454
rect 564702 61218 591102 61454
rect 591338 61218 591422 61454
rect 591658 61218 592650 61454
rect -8726 61186 592650 61218
rect -8726 58054 592650 58086
rect -8726 57818 -6774 58054
rect -6538 57818 -6454 58054
rect -6218 57818 20426 58054
rect 20662 57818 20746 58054
rect 20982 57818 380426 58054
rect 380662 57818 380746 58054
rect 380982 57818 416426 58054
rect 416662 57818 416746 58054
rect 416982 57818 452426 58054
rect 452662 57818 452746 58054
rect 452982 57818 488426 58054
rect 488662 57818 488746 58054
rect 488982 57818 524426 58054
rect 524662 57818 524746 58054
rect 524982 57818 560426 58054
rect 560662 57818 560746 58054
rect 560982 57818 590142 58054
rect 590378 57818 590462 58054
rect 590698 57818 592650 58054
rect -8726 57734 592650 57818
rect -8726 57498 -6774 57734
rect -6538 57498 -6454 57734
rect -6218 57498 20426 57734
rect 20662 57498 20746 57734
rect 20982 57498 380426 57734
rect 380662 57498 380746 57734
rect 380982 57498 416426 57734
rect 416662 57498 416746 57734
rect 416982 57498 452426 57734
rect 452662 57498 452746 57734
rect 452982 57498 488426 57734
rect 488662 57498 488746 57734
rect 488982 57498 524426 57734
rect 524662 57498 524746 57734
rect 524982 57498 560426 57734
rect 560662 57498 560746 57734
rect 560982 57498 590142 57734
rect 590378 57498 590462 57734
rect 590698 57498 592650 57734
rect -8726 57466 592650 57498
rect -8726 54334 592650 54366
rect -8726 54098 -5814 54334
rect -5578 54098 -5494 54334
rect -5258 54098 16706 54334
rect 16942 54098 17026 54334
rect 17262 54098 376706 54334
rect 376942 54098 377026 54334
rect 377262 54098 412706 54334
rect 412942 54098 413026 54334
rect 413262 54098 448706 54334
rect 448942 54098 449026 54334
rect 449262 54098 484706 54334
rect 484942 54098 485026 54334
rect 485262 54098 520706 54334
rect 520942 54098 521026 54334
rect 521262 54098 556706 54334
rect 556942 54098 557026 54334
rect 557262 54098 589182 54334
rect 589418 54098 589502 54334
rect 589738 54098 592650 54334
rect -8726 54014 592650 54098
rect -8726 53778 -5814 54014
rect -5578 53778 -5494 54014
rect -5258 53778 16706 54014
rect 16942 53778 17026 54014
rect 17262 53778 376706 54014
rect 376942 53778 377026 54014
rect 377262 53778 412706 54014
rect 412942 53778 413026 54014
rect 413262 53778 448706 54014
rect 448942 53778 449026 54014
rect 449262 53778 484706 54014
rect 484942 53778 485026 54014
rect 485262 53778 520706 54014
rect 520942 53778 521026 54014
rect 521262 53778 556706 54014
rect 556942 53778 557026 54014
rect 557262 53778 589182 54014
rect 589418 53778 589502 54014
rect 589738 53778 592650 54014
rect -8726 53746 592650 53778
rect -8726 50614 592650 50646
rect -8726 50378 -4854 50614
rect -4618 50378 -4534 50614
rect -4298 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 372986 50614
rect 373222 50378 373306 50614
rect 373542 50378 408986 50614
rect 409222 50378 409306 50614
rect 409542 50378 444986 50614
rect 445222 50378 445306 50614
rect 445542 50378 480986 50614
rect 481222 50378 481306 50614
rect 481542 50378 516986 50614
rect 517222 50378 517306 50614
rect 517542 50378 588222 50614
rect 588458 50378 588542 50614
rect 588778 50378 592650 50614
rect -8726 50294 592650 50378
rect -8726 50058 -4854 50294
rect -4618 50058 -4534 50294
rect -4298 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 372986 50294
rect 373222 50058 373306 50294
rect 373542 50058 408986 50294
rect 409222 50058 409306 50294
rect 409542 50058 444986 50294
rect 445222 50058 445306 50294
rect 445542 50058 480986 50294
rect 481222 50058 481306 50294
rect 481542 50058 516986 50294
rect 517222 50058 517306 50294
rect 517542 50058 588222 50294
rect 588458 50058 588542 50294
rect 588778 50058 592650 50294
rect -8726 50026 592650 50058
rect -8726 46894 592650 46926
rect -8726 46658 -3894 46894
rect -3658 46658 -3574 46894
rect -3338 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 45266 46894
rect 45502 46658 45586 46894
rect 45822 46658 81266 46894
rect 81502 46658 81586 46894
rect 81822 46658 117266 46894
rect 117502 46658 117586 46894
rect 117822 46658 153266 46894
rect 153502 46658 153586 46894
rect 153822 46658 189266 46894
rect 189502 46658 189586 46894
rect 189822 46658 225266 46894
rect 225502 46658 225586 46894
rect 225822 46658 261266 46894
rect 261502 46658 261586 46894
rect 261822 46658 297266 46894
rect 297502 46658 297586 46894
rect 297822 46658 333266 46894
rect 333502 46658 333586 46894
rect 333822 46658 369266 46894
rect 369502 46658 369586 46894
rect 369822 46658 405266 46894
rect 405502 46658 405586 46894
rect 405822 46658 441266 46894
rect 441502 46658 441586 46894
rect 441822 46658 477266 46894
rect 477502 46658 477586 46894
rect 477822 46658 513266 46894
rect 513502 46658 513586 46894
rect 513822 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 587262 46894
rect 587498 46658 587582 46894
rect 587818 46658 592650 46894
rect -8726 46574 592650 46658
rect -8726 46338 -3894 46574
rect -3658 46338 -3574 46574
rect -3338 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 45266 46574
rect 45502 46338 45586 46574
rect 45822 46338 81266 46574
rect 81502 46338 81586 46574
rect 81822 46338 117266 46574
rect 117502 46338 117586 46574
rect 117822 46338 153266 46574
rect 153502 46338 153586 46574
rect 153822 46338 189266 46574
rect 189502 46338 189586 46574
rect 189822 46338 225266 46574
rect 225502 46338 225586 46574
rect 225822 46338 261266 46574
rect 261502 46338 261586 46574
rect 261822 46338 297266 46574
rect 297502 46338 297586 46574
rect 297822 46338 333266 46574
rect 333502 46338 333586 46574
rect 333822 46338 369266 46574
rect 369502 46338 369586 46574
rect 369822 46338 405266 46574
rect 405502 46338 405586 46574
rect 405822 46338 441266 46574
rect 441502 46338 441586 46574
rect 441822 46338 477266 46574
rect 477502 46338 477586 46574
rect 477822 46338 513266 46574
rect 513502 46338 513586 46574
rect 513822 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 587262 46574
rect 587498 46338 587582 46574
rect 587818 46338 592650 46574
rect -8726 46306 592650 46338
rect -8726 43174 592650 43206
rect -8726 42938 -2934 43174
rect -2698 42938 -2614 43174
rect -2378 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 77546 43174
rect 77782 42938 77866 43174
rect 78102 42938 113546 43174
rect 113782 42938 113866 43174
rect 114102 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 221546 43174
rect 221782 42938 221866 43174
rect 222102 42938 257546 43174
rect 257782 42938 257866 43174
rect 258102 42938 293546 43174
rect 293782 42938 293866 43174
rect 294102 42938 329546 43174
rect 329782 42938 329866 43174
rect 330102 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 401546 43174
rect 401782 42938 401866 43174
rect 402102 42938 437546 43174
rect 437782 42938 437866 43174
rect 438102 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 545930 43174
rect 546166 42938 550875 43174
rect 551111 42938 555820 43174
rect 556056 42938 560765 43174
rect 561001 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 586302 43174
rect 586538 42938 586622 43174
rect 586858 42938 592650 43174
rect -8726 42854 592650 42938
rect -8726 42618 -2934 42854
rect -2698 42618 -2614 42854
rect -2378 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 77546 42854
rect 77782 42618 77866 42854
rect 78102 42618 113546 42854
rect 113782 42618 113866 42854
rect 114102 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 221546 42854
rect 221782 42618 221866 42854
rect 222102 42618 257546 42854
rect 257782 42618 257866 42854
rect 258102 42618 293546 42854
rect 293782 42618 293866 42854
rect 294102 42618 329546 42854
rect 329782 42618 329866 42854
rect 330102 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 401546 42854
rect 401782 42618 401866 42854
rect 402102 42618 437546 42854
rect 437782 42618 437866 42854
rect 438102 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 545930 42854
rect 546166 42618 550875 42854
rect 551111 42618 555820 42854
rect 556056 42618 560765 42854
rect 561001 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 586302 42854
rect 586538 42618 586622 42854
rect 586858 42618 592650 42854
rect -8726 42586 592650 42618
rect -8726 39454 592650 39486
rect -8726 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 543458 39454
rect 543694 39218 548403 39454
rect 548639 39218 553348 39454
rect 553584 39218 558293 39454
rect 558529 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 592650 39454
rect -8726 39134 592650 39218
rect -8726 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 543458 39134
rect 543694 38898 548403 39134
rect 548639 38898 553348 39134
rect 553584 38898 558293 39134
rect 558529 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 592650 39134
rect -8726 38866 592650 38898
rect -8726 29494 592650 29526
rect -8726 29258 -8694 29494
rect -8458 29258 -8374 29494
rect -8138 29258 27866 29494
rect 28102 29258 28186 29494
rect 28422 29258 63866 29494
rect 64102 29258 64186 29494
rect 64422 29258 99866 29494
rect 100102 29258 100186 29494
rect 100422 29258 135866 29494
rect 136102 29258 136186 29494
rect 136422 29258 171866 29494
rect 172102 29258 172186 29494
rect 172422 29258 207866 29494
rect 208102 29258 208186 29494
rect 208422 29258 243866 29494
rect 244102 29258 244186 29494
rect 244422 29258 279866 29494
rect 280102 29258 280186 29494
rect 280422 29258 315866 29494
rect 316102 29258 316186 29494
rect 316422 29258 351866 29494
rect 352102 29258 352186 29494
rect 352422 29258 387866 29494
rect 388102 29258 388186 29494
rect 388422 29258 423866 29494
rect 424102 29258 424186 29494
rect 424422 29258 459866 29494
rect 460102 29258 460186 29494
rect 460422 29258 495866 29494
rect 496102 29258 496186 29494
rect 496422 29258 531866 29494
rect 532102 29258 532186 29494
rect 532422 29258 567866 29494
rect 568102 29258 568186 29494
rect 568422 29258 592062 29494
rect 592298 29258 592382 29494
rect 592618 29258 592650 29494
rect -8726 29174 592650 29258
rect -8726 28938 -8694 29174
rect -8458 28938 -8374 29174
rect -8138 28938 27866 29174
rect 28102 28938 28186 29174
rect 28422 28938 63866 29174
rect 64102 28938 64186 29174
rect 64422 28938 99866 29174
rect 100102 28938 100186 29174
rect 100422 28938 135866 29174
rect 136102 28938 136186 29174
rect 136422 28938 171866 29174
rect 172102 28938 172186 29174
rect 172422 28938 207866 29174
rect 208102 28938 208186 29174
rect 208422 28938 243866 29174
rect 244102 28938 244186 29174
rect 244422 28938 279866 29174
rect 280102 28938 280186 29174
rect 280422 28938 315866 29174
rect 316102 28938 316186 29174
rect 316422 28938 351866 29174
rect 352102 28938 352186 29174
rect 352422 28938 387866 29174
rect 388102 28938 388186 29174
rect 388422 28938 423866 29174
rect 424102 28938 424186 29174
rect 424422 28938 459866 29174
rect 460102 28938 460186 29174
rect 460422 28938 495866 29174
rect 496102 28938 496186 29174
rect 496422 28938 531866 29174
rect 532102 28938 532186 29174
rect 532422 28938 567866 29174
rect 568102 28938 568186 29174
rect 568422 28938 592062 29174
rect 592298 28938 592382 29174
rect 592618 28938 592650 29174
rect -8726 28906 592650 28938
rect -8726 25774 592650 25806
rect -8726 25538 -7734 25774
rect -7498 25538 -7414 25774
rect -7178 25538 24146 25774
rect 24382 25538 24466 25774
rect 24702 25538 60146 25774
rect 60382 25538 60466 25774
rect 60702 25538 96146 25774
rect 96382 25538 96466 25774
rect 96702 25538 132146 25774
rect 132382 25538 132466 25774
rect 132702 25538 168146 25774
rect 168382 25538 168466 25774
rect 168702 25538 204146 25774
rect 204382 25538 204466 25774
rect 204702 25538 240146 25774
rect 240382 25538 240466 25774
rect 240702 25538 276146 25774
rect 276382 25538 276466 25774
rect 276702 25538 312146 25774
rect 312382 25538 312466 25774
rect 312702 25538 348146 25774
rect 348382 25538 348466 25774
rect 348702 25538 384146 25774
rect 384382 25538 384466 25774
rect 384702 25538 420146 25774
rect 420382 25538 420466 25774
rect 420702 25538 456146 25774
rect 456382 25538 456466 25774
rect 456702 25538 492146 25774
rect 492382 25538 492466 25774
rect 492702 25538 528146 25774
rect 528382 25538 528466 25774
rect 528702 25538 564146 25774
rect 564382 25538 564466 25774
rect 564702 25538 591102 25774
rect 591338 25538 591422 25774
rect 591658 25538 592650 25774
rect -8726 25454 592650 25538
rect -8726 25218 -7734 25454
rect -7498 25218 -7414 25454
rect -7178 25218 24146 25454
rect 24382 25218 24466 25454
rect 24702 25218 60146 25454
rect 60382 25218 60466 25454
rect 60702 25218 96146 25454
rect 96382 25218 96466 25454
rect 96702 25218 132146 25454
rect 132382 25218 132466 25454
rect 132702 25218 168146 25454
rect 168382 25218 168466 25454
rect 168702 25218 204146 25454
rect 204382 25218 204466 25454
rect 204702 25218 240146 25454
rect 240382 25218 240466 25454
rect 240702 25218 276146 25454
rect 276382 25218 276466 25454
rect 276702 25218 312146 25454
rect 312382 25218 312466 25454
rect 312702 25218 348146 25454
rect 348382 25218 348466 25454
rect 348702 25218 384146 25454
rect 384382 25218 384466 25454
rect 384702 25218 420146 25454
rect 420382 25218 420466 25454
rect 420702 25218 456146 25454
rect 456382 25218 456466 25454
rect 456702 25218 492146 25454
rect 492382 25218 492466 25454
rect 492702 25218 528146 25454
rect 528382 25218 528466 25454
rect 528702 25218 564146 25454
rect 564382 25218 564466 25454
rect 564702 25218 591102 25454
rect 591338 25218 591422 25454
rect 591658 25218 592650 25454
rect -8726 25186 592650 25218
rect -8726 22054 592650 22086
rect -8726 21818 -6774 22054
rect -6538 21818 -6454 22054
rect -6218 21818 20426 22054
rect 20662 21818 20746 22054
rect 20982 21818 56426 22054
rect 56662 21818 56746 22054
rect 56982 21818 92426 22054
rect 92662 21818 92746 22054
rect 92982 21818 128426 22054
rect 128662 21818 128746 22054
rect 128982 21818 164426 22054
rect 164662 21818 164746 22054
rect 164982 21818 200426 22054
rect 200662 21818 200746 22054
rect 200982 21818 236426 22054
rect 236662 21818 236746 22054
rect 236982 21818 272426 22054
rect 272662 21818 272746 22054
rect 272982 21818 308426 22054
rect 308662 21818 308746 22054
rect 308982 21818 344426 22054
rect 344662 21818 344746 22054
rect 344982 21818 380426 22054
rect 380662 21818 380746 22054
rect 380982 21818 416426 22054
rect 416662 21818 416746 22054
rect 416982 21818 452426 22054
rect 452662 21818 452746 22054
rect 452982 21818 488426 22054
rect 488662 21818 488746 22054
rect 488982 21818 524426 22054
rect 524662 21818 524746 22054
rect 524982 21818 560426 22054
rect 560662 21818 560746 22054
rect 560982 21818 590142 22054
rect 590378 21818 590462 22054
rect 590698 21818 592650 22054
rect -8726 21734 592650 21818
rect -8726 21498 -6774 21734
rect -6538 21498 -6454 21734
rect -6218 21498 20426 21734
rect 20662 21498 20746 21734
rect 20982 21498 56426 21734
rect 56662 21498 56746 21734
rect 56982 21498 92426 21734
rect 92662 21498 92746 21734
rect 92982 21498 128426 21734
rect 128662 21498 128746 21734
rect 128982 21498 164426 21734
rect 164662 21498 164746 21734
rect 164982 21498 200426 21734
rect 200662 21498 200746 21734
rect 200982 21498 236426 21734
rect 236662 21498 236746 21734
rect 236982 21498 272426 21734
rect 272662 21498 272746 21734
rect 272982 21498 308426 21734
rect 308662 21498 308746 21734
rect 308982 21498 344426 21734
rect 344662 21498 344746 21734
rect 344982 21498 380426 21734
rect 380662 21498 380746 21734
rect 380982 21498 416426 21734
rect 416662 21498 416746 21734
rect 416982 21498 452426 21734
rect 452662 21498 452746 21734
rect 452982 21498 488426 21734
rect 488662 21498 488746 21734
rect 488982 21498 524426 21734
rect 524662 21498 524746 21734
rect 524982 21498 560426 21734
rect 560662 21498 560746 21734
rect 560982 21498 590142 21734
rect 590378 21498 590462 21734
rect 590698 21498 592650 21734
rect -8726 21466 592650 21498
rect -8726 18334 592650 18366
rect -8726 18098 -5814 18334
rect -5578 18098 -5494 18334
rect -5258 18098 16706 18334
rect 16942 18098 17026 18334
rect 17262 18098 52706 18334
rect 52942 18098 53026 18334
rect 53262 18098 88706 18334
rect 88942 18098 89026 18334
rect 89262 18098 124706 18334
rect 124942 18098 125026 18334
rect 125262 18098 160706 18334
rect 160942 18098 161026 18334
rect 161262 18098 196706 18334
rect 196942 18098 197026 18334
rect 197262 18098 232706 18334
rect 232942 18098 233026 18334
rect 233262 18098 268706 18334
rect 268942 18098 269026 18334
rect 269262 18098 304706 18334
rect 304942 18098 305026 18334
rect 305262 18098 340706 18334
rect 340942 18098 341026 18334
rect 341262 18098 376706 18334
rect 376942 18098 377026 18334
rect 377262 18098 412706 18334
rect 412942 18098 413026 18334
rect 413262 18098 448706 18334
rect 448942 18098 449026 18334
rect 449262 18098 484706 18334
rect 484942 18098 485026 18334
rect 485262 18098 520706 18334
rect 520942 18098 521026 18334
rect 521262 18098 556706 18334
rect 556942 18098 557026 18334
rect 557262 18098 589182 18334
rect 589418 18098 589502 18334
rect 589738 18098 592650 18334
rect -8726 18014 592650 18098
rect -8726 17778 -5814 18014
rect -5578 17778 -5494 18014
rect -5258 17778 16706 18014
rect 16942 17778 17026 18014
rect 17262 17778 52706 18014
rect 52942 17778 53026 18014
rect 53262 17778 88706 18014
rect 88942 17778 89026 18014
rect 89262 17778 124706 18014
rect 124942 17778 125026 18014
rect 125262 17778 160706 18014
rect 160942 17778 161026 18014
rect 161262 17778 196706 18014
rect 196942 17778 197026 18014
rect 197262 17778 232706 18014
rect 232942 17778 233026 18014
rect 233262 17778 268706 18014
rect 268942 17778 269026 18014
rect 269262 17778 304706 18014
rect 304942 17778 305026 18014
rect 305262 17778 340706 18014
rect 340942 17778 341026 18014
rect 341262 17778 376706 18014
rect 376942 17778 377026 18014
rect 377262 17778 412706 18014
rect 412942 17778 413026 18014
rect 413262 17778 448706 18014
rect 448942 17778 449026 18014
rect 449262 17778 484706 18014
rect 484942 17778 485026 18014
rect 485262 17778 520706 18014
rect 520942 17778 521026 18014
rect 521262 17778 556706 18014
rect 556942 17778 557026 18014
rect 557262 17778 589182 18014
rect 589418 17778 589502 18014
rect 589738 17778 592650 18014
rect -8726 17746 592650 17778
rect -8726 14614 592650 14646
rect -8726 14378 -4854 14614
rect -4618 14378 -4534 14614
rect -4298 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 588222 14614
rect 588458 14378 588542 14614
rect 588778 14378 592650 14614
rect -8726 14294 592650 14378
rect -8726 14058 -4854 14294
rect -4618 14058 -4534 14294
rect -4298 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 588222 14294
rect 588458 14058 588542 14294
rect 588778 14058 592650 14294
rect -8726 14026 592650 14058
rect -8726 10894 592650 10926
rect -8726 10658 -3894 10894
rect -3658 10658 -3574 10894
rect -3338 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 587262 10894
rect 587498 10658 587582 10894
rect 587818 10658 592650 10894
rect -8726 10574 592650 10658
rect -8726 10338 -3894 10574
rect -3658 10338 -3574 10574
rect -3338 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 587262 10574
rect 587498 10338 587582 10574
rect 587818 10338 592650 10574
rect -8726 10306 592650 10338
rect -8726 7174 592650 7206
rect -8726 6938 -2934 7174
rect -2698 6938 -2614 7174
rect -2378 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 586302 7174
rect 586538 6938 586622 7174
rect 586858 6938 592650 7174
rect -8726 6854 592650 6938
rect -8726 6618 -2934 6854
rect -2698 6618 -2614 6854
rect -2378 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 586302 6854
rect 586538 6618 586622 6854
rect 586858 6618 592650 6854
rect -8726 6586 592650 6618
rect -8726 3454 592650 3486
rect -8726 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 592650 3454
rect -8726 3134 592650 3218
rect -8726 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 592650 3134
rect -8726 2866 592650 2898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 5546 -1306
rect 5782 -1542 5866 -1306
rect 6102 -1542 41546 -1306
rect 41782 -1542 41866 -1306
rect 42102 -1542 77546 -1306
rect 77782 -1542 77866 -1306
rect 78102 -1542 113546 -1306
rect 113782 -1542 113866 -1306
rect 114102 -1542 149546 -1306
rect 149782 -1542 149866 -1306
rect 150102 -1542 185546 -1306
rect 185782 -1542 185866 -1306
rect 186102 -1542 221546 -1306
rect 221782 -1542 221866 -1306
rect 222102 -1542 257546 -1306
rect 257782 -1542 257866 -1306
rect 258102 -1542 293546 -1306
rect 293782 -1542 293866 -1306
rect 294102 -1542 329546 -1306
rect 329782 -1542 329866 -1306
rect 330102 -1542 365546 -1306
rect 365782 -1542 365866 -1306
rect 366102 -1542 401546 -1306
rect 401782 -1542 401866 -1306
rect 402102 -1542 437546 -1306
rect 437782 -1542 437866 -1306
rect 438102 -1542 473546 -1306
rect 473782 -1542 473866 -1306
rect 474102 -1542 509546 -1306
rect 509782 -1542 509866 -1306
rect 510102 -1542 545546 -1306
rect 545782 -1542 545866 -1306
rect 546102 -1542 581546 -1306
rect 581782 -1542 581866 -1306
rect 582102 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 5546 -1626
rect 5782 -1862 5866 -1626
rect 6102 -1862 41546 -1626
rect 41782 -1862 41866 -1626
rect 42102 -1862 77546 -1626
rect 77782 -1862 77866 -1626
rect 78102 -1862 113546 -1626
rect 113782 -1862 113866 -1626
rect 114102 -1862 149546 -1626
rect 149782 -1862 149866 -1626
rect 150102 -1862 185546 -1626
rect 185782 -1862 185866 -1626
rect 186102 -1862 221546 -1626
rect 221782 -1862 221866 -1626
rect 222102 -1862 257546 -1626
rect 257782 -1862 257866 -1626
rect 258102 -1862 293546 -1626
rect 293782 -1862 293866 -1626
rect 294102 -1862 329546 -1626
rect 329782 -1862 329866 -1626
rect 330102 -1862 365546 -1626
rect 365782 -1862 365866 -1626
rect 366102 -1862 401546 -1626
rect 401782 -1862 401866 -1626
rect 402102 -1862 437546 -1626
rect 437782 -1862 437866 -1626
rect 438102 -1862 473546 -1626
rect 473782 -1862 473866 -1626
rect 474102 -1862 509546 -1626
rect 509782 -1862 509866 -1626
rect 510102 -1862 545546 -1626
rect 545782 -1862 545866 -1626
rect 546102 -1862 581546 -1626
rect 581782 -1862 581866 -1626
rect 582102 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 9266 -2266
rect 9502 -2502 9586 -2266
rect 9822 -2502 45266 -2266
rect 45502 -2502 45586 -2266
rect 45822 -2502 81266 -2266
rect 81502 -2502 81586 -2266
rect 81822 -2502 117266 -2266
rect 117502 -2502 117586 -2266
rect 117822 -2502 153266 -2266
rect 153502 -2502 153586 -2266
rect 153822 -2502 189266 -2266
rect 189502 -2502 189586 -2266
rect 189822 -2502 225266 -2266
rect 225502 -2502 225586 -2266
rect 225822 -2502 261266 -2266
rect 261502 -2502 261586 -2266
rect 261822 -2502 297266 -2266
rect 297502 -2502 297586 -2266
rect 297822 -2502 333266 -2266
rect 333502 -2502 333586 -2266
rect 333822 -2502 369266 -2266
rect 369502 -2502 369586 -2266
rect 369822 -2502 405266 -2266
rect 405502 -2502 405586 -2266
rect 405822 -2502 441266 -2266
rect 441502 -2502 441586 -2266
rect 441822 -2502 477266 -2266
rect 477502 -2502 477586 -2266
rect 477822 -2502 513266 -2266
rect 513502 -2502 513586 -2266
rect 513822 -2502 549266 -2266
rect 549502 -2502 549586 -2266
rect 549822 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 9266 -2586
rect 9502 -2822 9586 -2586
rect 9822 -2822 45266 -2586
rect 45502 -2822 45586 -2586
rect 45822 -2822 81266 -2586
rect 81502 -2822 81586 -2586
rect 81822 -2822 117266 -2586
rect 117502 -2822 117586 -2586
rect 117822 -2822 153266 -2586
rect 153502 -2822 153586 -2586
rect 153822 -2822 189266 -2586
rect 189502 -2822 189586 -2586
rect 189822 -2822 225266 -2586
rect 225502 -2822 225586 -2586
rect 225822 -2822 261266 -2586
rect 261502 -2822 261586 -2586
rect 261822 -2822 297266 -2586
rect 297502 -2822 297586 -2586
rect 297822 -2822 333266 -2586
rect 333502 -2822 333586 -2586
rect 333822 -2822 369266 -2586
rect 369502 -2822 369586 -2586
rect 369822 -2822 405266 -2586
rect 405502 -2822 405586 -2586
rect 405822 -2822 441266 -2586
rect 441502 -2822 441586 -2586
rect 441822 -2822 477266 -2586
rect 477502 -2822 477586 -2586
rect 477822 -2822 513266 -2586
rect 513502 -2822 513586 -2586
rect 513822 -2822 549266 -2586
rect 549502 -2822 549586 -2586
rect 549822 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 12986 -3226
rect 13222 -3462 13306 -3226
rect 13542 -3462 48986 -3226
rect 49222 -3462 49306 -3226
rect 49542 -3462 84986 -3226
rect 85222 -3462 85306 -3226
rect 85542 -3462 120986 -3226
rect 121222 -3462 121306 -3226
rect 121542 -3462 156986 -3226
rect 157222 -3462 157306 -3226
rect 157542 -3462 192986 -3226
rect 193222 -3462 193306 -3226
rect 193542 -3462 228986 -3226
rect 229222 -3462 229306 -3226
rect 229542 -3462 264986 -3226
rect 265222 -3462 265306 -3226
rect 265542 -3462 300986 -3226
rect 301222 -3462 301306 -3226
rect 301542 -3462 336986 -3226
rect 337222 -3462 337306 -3226
rect 337542 -3462 372986 -3226
rect 373222 -3462 373306 -3226
rect 373542 -3462 408986 -3226
rect 409222 -3462 409306 -3226
rect 409542 -3462 444986 -3226
rect 445222 -3462 445306 -3226
rect 445542 -3462 480986 -3226
rect 481222 -3462 481306 -3226
rect 481542 -3462 516986 -3226
rect 517222 -3462 517306 -3226
rect 517542 -3462 552986 -3226
rect 553222 -3462 553306 -3226
rect 553542 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 12986 -3546
rect 13222 -3782 13306 -3546
rect 13542 -3782 48986 -3546
rect 49222 -3782 49306 -3546
rect 49542 -3782 84986 -3546
rect 85222 -3782 85306 -3546
rect 85542 -3782 120986 -3546
rect 121222 -3782 121306 -3546
rect 121542 -3782 156986 -3546
rect 157222 -3782 157306 -3546
rect 157542 -3782 192986 -3546
rect 193222 -3782 193306 -3546
rect 193542 -3782 228986 -3546
rect 229222 -3782 229306 -3546
rect 229542 -3782 264986 -3546
rect 265222 -3782 265306 -3546
rect 265542 -3782 300986 -3546
rect 301222 -3782 301306 -3546
rect 301542 -3782 336986 -3546
rect 337222 -3782 337306 -3546
rect 337542 -3782 372986 -3546
rect 373222 -3782 373306 -3546
rect 373542 -3782 408986 -3546
rect 409222 -3782 409306 -3546
rect 409542 -3782 444986 -3546
rect 445222 -3782 445306 -3546
rect 445542 -3782 480986 -3546
rect 481222 -3782 481306 -3546
rect 481542 -3782 516986 -3546
rect 517222 -3782 517306 -3546
rect 517542 -3782 552986 -3546
rect 553222 -3782 553306 -3546
rect 553542 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 16706 -4186
rect 16942 -4422 17026 -4186
rect 17262 -4422 52706 -4186
rect 52942 -4422 53026 -4186
rect 53262 -4422 88706 -4186
rect 88942 -4422 89026 -4186
rect 89262 -4422 124706 -4186
rect 124942 -4422 125026 -4186
rect 125262 -4422 160706 -4186
rect 160942 -4422 161026 -4186
rect 161262 -4422 196706 -4186
rect 196942 -4422 197026 -4186
rect 197262 -4422 232706 -4186
rect 232942 -4422 233026 -4186
rect 233262 -4422 268706 -4186
rect 268942 -4422 269026 -4186
rect 269262 -4422 304706 -4186
rect 304942 -4422 305026 -4186
rect 305262 -4422 340706 -4186
rect 340942 -4422 341026 -4186
rect 341262 -4422 376706 -4186
rect 376942 -4422 377026 -4186
rect 377262 -4422 412706 -4186
rect 412942 -4422 413026 -4186
rect 413262 -4422 448706 -4186
rect 448942 -4422 449026 -4186
rect 449262 -4422 484706 -4186
rect 484942 -4422 485026 -4186
rect 485262 -4422 520706 -4186
rect 520942 -4422 521026 -4186
rect 521262 -4422 556706 -4186
rect 556942 -4422 557026 -4186
rect 557262 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 16706 -4506
rect 16942 -4742 17026 -4506
rect 17262 -4742 52706 -4506
rect 52942 -4742 53026 -4506
rect 53262 -4742 88706 -4506
rect 88942 -4742 89026 -4506
rect 89262 -4742 124706 -4506
rect 124942 -4742 125026 -4506
rect 125262 -4742 160706 -4506
rect 160942 -4742 161026 -4506
rect 161262 -4742 196706 -4506
rect 196942 -4742 197026 -4506
rect 197262 -4742 232706 -4506
rect 232942 -4742 233026 -4506
rect 233262 -4742 268706 -4506
rect 268942 -4742 269026 -4506
rect 269262 -4742 304706 -4506
rect 304942 -4742 305026 -4506
rect 305262 -4742 340706 -4506
rect 340942 -4742 341026 -4506
rect 341262 -4742 376706 -4506
rect 376942 -4742 377026 -4506
rect 377262 -4742 412706 -4506
rect 412942 -4742 413026 -4506
rect 413262 -4742 448706 -4506
rect 448942 -4742 449026 -4506
rect 449262 -4742 484706 -4506
rect 484942 -4742 485026 -4506
rect 485262 -4742 520706 -4506
rect 520942 -4742 521026 -4506
rect 521262 -4742 556706 -4506
rect 556942 -4742 557026 -4506
rect 557262 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 20426 -5146
rect 20662 -5382 20746 -5146
rect 20982 -5382 56426 -5146
rect 56662 -5382 56746 -5146
rect 56982 -5382 92426 -5146
rect 92662 -5382 92746 -5146
rect 92982 -5382 128426 -5146
rect 128662 -5382 128746 -5146
rect 128982 -5382 164426 -5146
rect 164662 -5382 164746 -5146
rect 164982 -5382 200426 -5146
rect 200662 -5382 200746 -5146
rect 200982 -5382 236426 -5146
rect 236662 -5382 236746 -5146
rect 236982 -5382 272426 -5146
rect 272662 -5382 272746 -5146
rect 272982 -5382 308426 -5146
rect 308662 -5382 308746 -5146
rect 308982 -5382 344426 -5146
rect 344662 -5382 344746 -5146
rect 344982 -5382 380426 -5146
rect 380662 -5382 380746 -5146
rect 380982 -5382 416426 -5146
rect 416662 -5382 416746 -5146
rect 416982 -5382 452426 -5146
rect 452662 -5382 452746 -5146
rect 452982 -5382 488426 -5146
rect 488662 -5382 488746 -5146
rect 488982 -5382 524426 -5146
rect 524662 -5382 524746 -5146
rect 524982 -5382 560426 -5146
rect 560662 -5382 560746 -5146
rect 560982 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 20426 -5466
rect 20662 -5702 20746 -5466
rect 20982 -5702 56426 -5466
rect 56662 -5702 56746 -5466
rect 56982 -5702 92426 -5466
rect 92662 -5702 92746 -5466
rect 92982 -5702 128426 -5466
rect 128662 -5702 128746 -5466
rect 128982 -5702 164426 -5466
rect 164662 -5702 164746 -5466
rect 164982 -5702 200426 -5466
rect 200662 -5702 200746 -5466
rect 200982 -5702 236426 -5466
rect 236662 -5702 236746 -5466
rect 236982 -5702 272426 -5466
rect 272662 -5702 272746 -5466
rect 272982 -5702 308426 -5466
rect 308662 -5702 308746 -5466
rect 308982 -5702 344426 -5466
rect 344662 -5702 344746 -5466
rect 344982 -5702 380426 -5466
rect 380662 -5702 380746 -5466
rect 380982 -5702 416426 -5466
rect 416662 -5702 416746 -5466
rect 416982 -5702 452426 -5466
rect 452662 -5702 452746 -5466
rect 452982 -5702 488426 -5466
rect 488662 -5702 488746 -5466
rect 488982 -5702 524426 -5466
rect 524662 -5702 524746 -5466
rect 524982 -5702 560426 -5466
rect 560662 -5702 560746 -5466
rect 560982 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 24146 -6106
rect 24382 -6342 24466 -6106
rect 24702 -6342 60146 -6106
rect 60382 -6342 60466 -6106
rect 60702 -6342 96146 -6106
rect 96382 -6342 96466 -6106
rect 96702 -6342 132146 -6106
rect 132382 -6342 132466 -6106
rect 132702 -6342 168146 -6106
rect 168382 -6342 168466 -6106
rect 168702 -6342 204146 -6106
rect 204382 -6342 204466 -6106
rect 204702 -6342 240146 -6106
rect 240382 -6342 240466 -6106
rect 240702 -6342 276146 -6106
rect 276382 -6342 276466 -6106
rect 276702 -6342 312146 -6106
rect 312382 -6342 312466 -6106
rect 312702 -6342 348146 -6106
rect 348382 -6342 348466 -6106
rect 348702 -6342 384146 -6106
rect 384382 -6342 384466 -6106
rect 384702 -6342 420146 -6106
rect 420382 -6342 420466 -6106
rect 420702 -6342 456146 -6106
rect 456382 -6342 456466 -6106
rect 456702 -6342 492146 -6106
rect 492382 -6342 492466 -6106
rect 492702 -6342 528146 -6106
rect 528382 -6342 528466 -6106
rect 528702 -6342 564146 -6106
rect 564382 -6342 564466 -6106
rect 564702 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 24146 -6426
rect 24382 -6662 24466 -6426
rect 24702 -6662 60146 -6426
rect 60382 -6662 60466 -6426
rect 60702 -6662 96146 -6426
rect 96382 -6662 96466 -6426
rect 96702 -6662 132146 -6426
rect 132382 -6662 132466 -6426
rect 132702 -6662 168146 -6426
rect 168382 -6662 168466 -6426
rect 168702 -6662 204146 -6426
rect 204382 -6662 204466 -6426
rect 204702 -6662 240146 -6426
rect 240382 -6662 240466 -6426
rect 240702 -6662 276146 -6426
rect 276382 -6662 276466 -6426
rect 276702 -6662 312146 -6426
rect 312382 -6662 312466 -6426
rect 312702 -6662 348146 -6426
rect 348382 -6662 348466 -6426
rect 348702 -6662 384146 -6426
rect 384382 -6662 384466 -6426
rect 384702 -6662 420146 -6426
rect 420382 -6662 420466 -6426
rect 420702 -6662 456146 -6426
rect 456382 -6662 456466 -6426
rect 456702 -6662 492146 -6426
rect 492382 -6662 492466 -6426
rect 492702 -6662 528146 -6426
rect 528382 -6662 528466 -6426
rect 528702 -6662 564146 -6426
rect 564382 -6662 564466 -6426
rect 564702 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 27866 -7066
rect 28102 -7302 28186 -7066
rect 28422 -7302 63866 -7066
rect 64102 -7302 64186 -7066
rect 64422 -7302 99866 -7066
rect 100102 -7302 100186 -7066
rect 100422 -7302 135866 -7066
rect 136102 -7302 136186 -7066
rect 136422 -7302 171866 -7066
rect 172102 -7302 172186 -7066
rect 172422 -7302 207866 -7066
rect 208102 -7302 208186 -7066
rect 208422 -7302 243866 -7066
rect 244102 -7302 244186 -7066
rect 244422 -7302 279866 -7066
rect 280102 -7302 280186 -7066
rect 280422 -7302 315866 -7066
rect 316102 -7302 316186 -7066
rect 316422 -7302 351866 -7066
rect 352102 -7302 352186 -7066
rect 352422 -7302 387866 -7066
rect 388102 -7302 388186 -7066
rect 388422 -7302 423866 -7066
rect 424102 -7302 424186 -7066
rect 424422 -7302 459866 -7066
rect 460102 -7302 460186 -7066
rect 460422 -7302 495866 -7066
rect 496102 -7302 496186 -7066
rect 496422 -7302 531866 -7066
rect 532102 -7302 532186 -7066
rect 532422 -7302 567866 -7066
rect 568102 -7302 568186 -7066
rect 568422 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 27866 -7386
rect 28102 -7622 28186 -7386
rect 28422 -7622 63866 -7386
rect 64102 -7622 64186 -7386
rect 64422 -7622 99866 -7386
rect 100102 -7622 100186 -7386
rect 100422 -7622 135866 -7386
rect 136102 -7622 136186 -7386
rect 136422 -7622 171866 -7386
rect 172102 -7622 172186 -7386
rect 172422 -7622 207866 -7386
rect 208102 -7622 208186 -7386
rect 208422 -7622 243866 -7386
rect 244102 -7622 244186 -7386
rect 244422 -7622 279866 -7386
rect 280102 -7622 280186 -7386
rect 280422 -7622 315866 -7386
rect 316102 -7622 316186 -7386
rect 316422 -7622 351866 -7386
rect 352102 -7622 352186 -7386
rect 352422 -7622 387866 -7386
rect 388102 -7622 388186 -7386
rect 388422 -7622 423866 -7386
rect 424102 -7622 424186 -7386
rect 424422 -7622 459866 -7386
rect 460102 -7622 460186 -7386
rect 460422 -7622 495866 -7386
rect 496102 -7622 496186 -7386
rect 496422 -7622 531866 -7386
rect 532102 -7622 532186 -7386
rect 532422 -7622 567866 -7386
rect 568102 -7622 568186 -7386
rect 568422 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use posit_unit  posit_unit
timestamp 0
transform 1 0 460000 0 1 200000
box 0 2128 70000 67504
use multiplexer  proj_multiplexer
timestamp 0
transform 1 0 450000 0 1 322000
box 0 0 60000 64000
use tholin_avalonsemi_5401  tholin_avalonsemi_5401
timestamp 0
transform 1 0 520000 0 1 425000
box 1066 0 36000 36000
use tholin_avalonsemi_tbb1143  tholin_avalonsemi_tbb1143
timestamp 0
transform 1 0 400000 0 1 305000
box 1066 2048 30000 30000
use tt2_tholin_diceroll  tt2_tholin_diceroll
timestamp 0
transform 1 0 470000 0 1 432000
box 1066 0 21043 22000
use tt2_tholin_multiplexed_counter  tt2_tholin_multiplexed_counter
timestamp 0
transform 1 0 550000 0 1 360000
box 842 0 17098 18000
use tt2_tholin_multiplier  tt2_tholin_multiplier
timestamp 0
transform 1 0 450000 0 1 500000
box 0 0 11118 16584
use tt2_tholin_namebadge  tt2_tholin_namebadge
timestamp 0
transform 1 0 420000 0 1 420000
box 1066 0 23987 25000
use tune_player  tune_player
timestamp 0
transform 1 0 540000 0 1 30000
box 0 2128 21043 19632
use wrapped_6502  wrapped_6502
timestamp 0
transform 1 0 410000 0 1 120000
box 1066 1504 40000 40000
use wrapped_MC14500  wrapped_MC14500
timestamp 0
transform 1 0 480000 0 1 500000
box 566 0 12000 18000
use wrapped_as1802  wrapped_as1802
timestamp 0
transform 1 0 480000 0 1 80000
box 1066 2128 60000 60000
use wrapped_as2650  wrapped_as2650
timestamp 0
transform 1 0 460000 0 1 600000
box 0 0 68816 67992
use wrapped_as512512512  wrapped_as512512512
timestamp 0
transform 1 0 20000 0 1 45000
box 1066 2128 340000 637616
<< labels >>
flabel metal3 s 583520 285276 584960 285516 0 FreeSans 960 0 0 0 analog_io[0]
port 0 nsew signal bidirectional
flabel metal2 s 446098 703520 446210 704960 0 FreeSans 448 90 0 0 analog_io[10]
port 1 nsew signal bidirectional
flabel metal2 s 381146 703520 381258 704960 0 FreeSans 448 90 0 0 analog_io[11]
port 2 nsew signal bidirectional
flabel metal2 s 316286 703520 316398 704960 0 FreeSans 448 90 0 0 analog_io[12]
port 3 nsew signal bidirectional
flabel metal2 s 251426 703520 251538 704960 0 FreeSans 448 90 0 0 analog_io[13]
port 4 nsew signal bidirectional
flabel metal2 s 186474 703520 186586 704960 0 FreeSans 448 90 0 0 analog_io[14]
port 5 nsew signal bidirectional
flabel metal2 s 121614 703520 121726 704960 0 FreeSans 448 90 0 0 analog_io[15]
port 6 nsew signal bidirectional
flabel metal2 s 56754 703520 56866 704960 0 FreeSans 448 90 0 0 analog_io[16]
port 7 nsew signal bidirectional
flabel metal3 s -960 697220 480 697460 0 FreeSans 960 0 0 0 analog_io[17]
port 8 nsew signal bidirectional
flabel metal3 s -960 644996 480 645236 0 FreeSans 960 0 0 0 analog_io[18]
port 9 nsew signal bidirectional
flabel metal3 s -960 592908 480 593148 0 FreeSans 960 0 0 0 analog_io[19]
port 10 nsew signal bidirectional
flabel metal3 s 583520 338452 584960 338692 0 FreeSans 960 0 0 0 analog_io[1]
port 11 nsew signal bidirectional
flabel metal3 s -960 540684 480 540924 0 FreeSans 960 0 0 0 analog_io[20]
port 12 nsew signal bidirectional
flabel metal3 s -960 488596 480 488836 0 FreeSans 960 0 0 0 analog_io[21]
port 13 nsew signal bidirectional
flabel metal3 s -960 436508 480 436748 0 FreeSans 960 0 0 0 analog_io[22]
port 14 nsew signal bidirectional
flabel metal3 s -960 384284 480 384524 0 FreeSans 960 0 0 0 analog_io[23]
port 15 nsew signal bidirectional
flabel metal3 s -960 332196 480 332436 0 FreeSans 960 0 0 0 analog_io[24]
port 16 nsew signal bidirectional
flabel metal3 s -960 279972 480 280212 0 FreeSans 960 0 0 0 analog_io[25]
port 17 nsew signal bidirectional
flabel metal3 s -960 227884 480 228124 0 FreeSans 960 0 0 0 analog_io[26]
port 18 nsew signal bidirectional
flabel metal3 s -960 175796 480 176036 0 FreeSans 960 0 0 0 analog_io[27]
port 19 nsew signal bidirectional
flabel metal3 s -960 123572 480 123812 0 FreeSans 960 0 0 0 analog_io[28]
port 20 nsew signal bidirectional
flabel metal3 s 583520 391628 584960 391868 0 FreeSans 960 0 0 0 analog_io[2]
port 21 nsew signal bidirectional
flabel metal3 s 583520 444668 584960 444908 0 FreeSans 960 0 0 0 analog_io[3]
port 22 nsew signal bidirectional
flabel metal3 s 583520 497844 584960 498084 0 FreeSans 960 0 0 0 analog_io[4]
port 23 nsew signal bidirectional
flabel metal3 s 583520 551020 584960 551260 0 FreeSans 960 0 0 0 analog_io[5]
port 24 nsew signal bidirectional
flabel metal3 s 583520 604060 584960 604300 0 FreeSans 960 0 0 0 analog_io[6]
port 25 nsew signal bidirectional
flabel metal3 s 583520 657236 584960 657476 0 FreeSans 960 0 0 0 analog_io[7]
port 26 nsew signal bidirectional
flabel metal2 s 575818 703520 575930 704960 0 FreeSans 448 90 0 0 analog_io[8]
port 27 nsew signal bidirectional
flabel metal2 s 510958 703520 511070 704960 0 FreeSans 448 90 0 0 analog_io[9]
port 28 nsew signal bidirectional
flabel metal3 s 583520 6476 584960 6716 0 FreeSans 960 0 0 0 io_in[0]
port 29 nsew signal input
flabel metal3 s 583520 457996 584960 458236 0 FreeSans 960 0 0 0 io_in[10]
port 30 nsew signal input
flabel metal3 s 583520 511172 584960 511412 0 FreeSans 960 0 0 0 io_in[11]
port 31 nsew signal input
flabel metal3 s 583520 564212 584960 564452 0 FreeSans 960 0 0 0 io_in[12]
port 32 nsew signal input
flabel metal3 s 583520 617388 584960 617628 0 FreeSans 960 0 0 0 io_in[13]
port 33 nsew signal input
flabel metal3 s 583520 670564 584960 670804 0 FreeSans 960 0 0 0 io_in[14]
port 34 nsew signal input
flabel metal2 s 559626 703520 559738 704960 0 FreeSans 448 90 0 0 io_in[15]
port 35 nsew signal input
flabel metal2 s 494766 703520 494878 704960 0 FreeSans 448 90 0 0 io_in[16]
port 36 nsew signal input
flabel metal2 s 429814 703520 429926 704960 0 FreeSans 448 90 0 0 io_in[17]
port 37 nsew signal input
flabel metal2 s 364954 703520 365066 704960 0 FreeSans 448 90 0 0 io_in[18]
port 38 nsew signal input
flabel metal2 s 300094 703520 300206 704960 0 FreeSans 448 90 0 0 io_in[19]
port 39 nsew signal input
flabel metal3 s 583520 46188 584960 46428 0 FreeSans 960 0 0 0 io_in[1]
port 40 nsew signal input
flabel metal2 s 235142 703520 235254 704960 0 FreeSans 448 90 0 0 io_in[20]
port 41 nsew signal input
flabel metal2 s 170282 703520 170394 704960 0 FreeSans 448 90 0 0 io_in[21]
port 42 nsew signal input
flabel metal2 s 105422 703520 105534 704960 0 FreeSans 448 90 0 0 io_in[22]
port 43 nsew signal input
flabel metal2 s 40470 703520 40582 704960 0 FreeSans 448 90 0 0 io_in[23]
port 44 nsew signal input
flabel metal3 s -960 684164 480 684404 0 FreeSans 960 0 0 0 io_in[24]
port 45 nsew signal input
flabel metal3 s -960 631940 480 632180 0 FreeSans 960 0 0 0 io_in[25]
port 46 nsew signal input
flabel metal3 s -960 579852 480 580092 0 FreeSans 960 0 0 0 io_in[26]
port 47 nsew signal input
flabel metal3 s -960 527764 480 528004 0 FreeSans 960 0 0 0 io_in[27]
port 48 nsew signal input
flabel metal3 s -960 475540 480 475780 0 FreeSans 960 0 0 0 io_in[28]
port 49 nsew signal input
flabel metal3 s -960 423452 480 423692 0 FreeSans 960 0 0 0 io_in[29]
port 50 nsew signal input
flabel metal3 s 583520 86036 584960 86276 0 FreeSans 960 0 0 0 io_in[2]
port 51 nsew signal input
flabel metal3 s -960 371228 480 371468 0 FreeSans 960 0 0 0 io_in[30]
port 52 nsew signal input
flabel metal3 s -960 319140 480 319380 0 FreeSans 960 0 0 0 io_in[31]
port 53 nsew signal input
flabel metal3 s -960 267052 480 267292 0 FreeSans 960 0 0 0 io_in[32]
port 54 nsew signal input
flabel metal3 s -960 214828 480 215068 0 FreeSans 960 0 0 0 io_in[33]
port 55 nsew signal input
flabel metal3 s -960 162740 480 162980 0 FreeSans 960 0 0 0 io_in[34]
port 56 nsew signal input
flabel metal3 s -960 110516 480 110756 0 FreeSans 960 0 0 0 io_in[35]
port 57 nsew signal input
flabel metal3 s -960 71484 480 71724 0 FreeSans 960 0 0 0 io_in[36]
port 58 nsew signal input
flabel metal3 s -960 32316 480 32556 0 FreeSans 960 0 0 0 io_in[37]
port 59 nsew signal input
flabel metal3 s 583520 125884 584960 126124 0 FreeSans 960 0 0 0 io_in[3]
port 60 nsew signal input
flabel metal3 s 583520 165732 584960 165972 0 FreeSans 960 0 0 0 io_in[4]
port 61 nsew signal input
flabel metal3 s 583520 205580 584960 205820 0 FreeSans 960 0 0 0 io_in[5]
port 62 nsew signal input
flabel metal3 s 583520 245428 584960 245668 0 FreeSans 960 0 0 0 io_in[6]
port 63 nsew signal input
flabel metal3 s 583520 298604 584960 298844 0 FreeSans 960 0 0 0 io_in[7]
port 64 nsew signal input
flabel metal3 s 583520 351780 584960 352020 0 FreeSans 960 0 0 0 io_in[8]
port 65 nsew signal input
flabel metal3 s 583520 404820 584960 405060 0 FreeSans 960 0 0 0 io_in[9]
port 66 nsew signal input
flabel metal3 s 583520 32996 584960 33236 0 FreeSans 960 0 0 0 io_oeb[0]
port 67 nsew signal tristate
flabel metal3 s 583520 484516 584960 484756 0 FreeSans 960 0 0 0 io_oeb[10]
port 68 nsew signal tristate
flabel metal3 s 583520 537692 584960 537932 0 FreeSans 960 0 0 0 io_oeb[11]
port 69 nsew signal tristate
flabel metal3 s 583520 590868 584960 591108 0 FreeSans 960 0 0 0 io_oeb[12]
port 70 nsew signal tristate
flabel metal3 s 583520 643908 584960 644148 0 FreeSans 960 0 0 0 io_oeb[13]
port 71 nsew signal tristate
flabel metal3 s 583520 697084 584960 697324 0 FreeSans 960 0 0 0 io_oeb[14]
port 72 nsew signal tristate
flabel metal2 s 527150 703520 527262 704960 0 FreeSans 448 90 0 0 io_oeb[15]
port 73 nsew signal tristate
flabel metal2 s 462290 703520 462402 704960 0 FreeSans 448 90 0 0 io_oeb[16]
port 74 nsew signal tristate
flabel metal2 s 397430 703520 397542 704960 0 FreeSans 448 90 0 0 io_oeb[17]
port 75 nsew signal tristate
flabel metal2 s 332478 703520 332590 704960 0 FreeSans 448 90 0 0 io_oeb[18]
port 76 nsew signal tristate
flabel metal2 s 267618 703520 267730 704960 0 FreeSans 448 90 0 0 io_oeb[19]
port 77 nsew signal tristate
flabel metal3 s 583520 72844 584960 73084 0 FreeSans 960 0 0 0 io_oeb[1]
port 78 nsew signal tristate
flabel metal2 s 202758 703520 202870 704960 0 FreeSans 448 90 0 0 io_oeb[20]
port 79 nsew signal tristate
flabel metal2 s 137806 703520 137918 704960 0 FreeSans 448 90 0 0 io_oeb[21]
port 80 nsew signal tristate
flabel metal2 s 72946 703520 73058 704960 0 FreeSans 448 90 0 0 io_oeb[22]
port 81 nsew signal tristate
flabel metal2 s 8086 703520 8198 704960 0 FreeSans 448 90 0 0 io_oeb[23]
port 82 nsew signal tristate
flabel metal3 s -960 658052 480 658292 0 FreeSans 960 0 0 0 io_oeb[24]
port 83 nsew signal tristate
flabel metal3 s -960 605964 480 606204 0 FreeSans 960 0 0 0 io_oeb[25]
port 84 nsew signal tristate
flabel metal3 s -960 553740 480 553980 0 FreeSans 960 0 0 0 io_oeb[26]
port 85 nsew signal tristate
flabel metal3 s -960 501652 480 501892 0 FreeSans 960 0 0 0 io_oeb[27]
port 86 nsew signal tristate
flabel metal3 s -960 449428 480 449668 0 FreeSans 960 0 0 0 io_oeb[28]
port 87 nsew signal tristate
flabel metal3 s -960 397340 480 397580 0 FreeSans 960 0 0 0 io_oeb[29]
port 88 nsew signal tristate
flabel metal3 s 583520 112692 584960 112932 0 FreeSans 960 0 0 0 io_oeb[2]
port 89 nsew signal tristate
flabel metal3 s -960 345252 480 345492 0 FreeSans 960 0 0 0 io_oeb[30]
port 90 nsew signal tristate
flabel metal3 s -960 293028 480 293268 0 FreeSans 960 0 0 0 io_oeb[31]
port 91 nsew signal tristate
flabel metal3 s -960 240940 480 241180 0 FreeSans 960 0 0 0 io_oeb[32]
port 92 nsew signal tristate
flabel metal3 s -960 188716 480 188956 0 FreeSans 960 0 0 0 io_oeb[33]
port 93 nsew signal tristate
flabel metal3 s -960 136628 480 136868 0 FreeSans 960 0 0 0 io_oeb[34]
port 94 nsew signal tristate
flabel metal3 s -960 84540 480 84780 0 FreeSans 960 0 0 0 io_oeb[35]
port 95 nsew signal tristate
flabel metal3 s -960 45372 480 45612 0 FreeSans 960 0 0 0 io_oeb[36]
port 96 nsew signal tristate
flabel metal3 s -960 6340 480 6580 0 FreeSans 960 0 0 0 io_oeb[37]
port 97 nsew signal tristate
flabel metal3 s 583520 152540 584960 152780 0 FreeSans 960 0 0 0 io_oeb[3]
port 98 nsew signal tristate
flabel metal3 s 583520 192388 584960 192628 0 FreeSans 960 0 0 0 io_oeb[4]
port 99 nsew signal tristate
flabel metal3 s 583520 232236 584960 232476 0 FreeSans 960 0 0 0 io_oeb[5]
port 100 nsew signal tristate
flabel metal3 s 583520 272084 584960 272324 0 FreeSans 960 0 0 0 io_oeb[6]
port 101 nsew signal tristate
flabel metal3 s 583520 325124 584960 325364 0 FreeSans 960 0 0 0 io_oeb[7]
port 102 nsew signal tristate
flabel metal3 s 583520 378300 584960 378540 0 FreeSans 960 0 0 0 io_oeb[8]
port 103 nsew signal tristate
flabel metal3 s 583520 431476 584960 431716 0 FreeSans 960 0 0 0 io_oeb[9]
port 104 nsew signal tristate
flabel metal3 s 583520 19668 584960 19908 0 FreeSans 960 0 0 0 io_out[0]
port 105 nsew signal tristate
flabel metal3 s 583520 471324 584960 471564 0 FreeSans 960 0 0 0 io_out[10]
port 106 nsew signal tristate
flabel metal3 s 583520 524364 584960 524604 0 FreeSans 960 0 0 0 io_out[11]
port 107 nsew signal tristate
flabel metal3 s 583520 577540 584960 577780 0 FreeSans 960 0 0 0 io_out[12]
port 108 nsew signal tristate
flabel metal3 s 583520 630716 584960 630956 0 FreeSans 960 0 0 0 io_out[13]
port 109 nsew signal tristate
flabel metal3 s 583520 683756 584960 683996 0 FreeSans 960 0 0 0 io_out[14]
port 110 nsew signal tristate
flabel metal2 s 543434 703520 543546 704960 0 FreeSans 448 90 0 0 io_out[15]
port 111 nsew signal tristate
flabel metal2 s 478482 703520 478594 704960 0 FreeSans 448 90 0 0 io_out[16]
port 112 nsew signal tristate
flabel metal2 s 413622 703520 413734 704960 0 FreeSans 448 90 0 0 io_out[17]
port 113 nsew signal tristate
flabel metal2 s 348762 703520 348874 704960 0 FreeSans 448 90 0 0 io_out[18]
port 114 nsew signal tristate
flabel metal2 s 283810 703520 283922 704960 0 FreeSans 448 90 0 0 io_out[19]
port 115 nsew signal tristate
flabel metal3 s 583520 59516 584960 59756 0 FreeSans 960 0 0 0 io_out[1]
port 116 nsew signal tristate
flabel metal2 s 218950 703520 219062 704960 0 FreeSans 448 90 0 0 io_out[20]
port 117 nsew signal tristate
flabel metal2 s 154090 703520 154202 704960 0 FreeSans 448 90 0 0 io_out[21]
port 118 nsew signal tristate
flabel metal2 s 89138 703520 89250 704960 0 FreeSans 448 90 0 0 io_out[22]
port 119 nsew signal tristate
flabel metal2 s 24278 703520 24390 704960 0 FreeSans 448 90 0 0 io_out[23]
port 120 nsew signal tristate
flabel metal3 s -960 671108 480 671348 0 FreeSans 960 0 0 0 io_out[24]
port 121 nsew signal tristate
flabel metal3 s -960 619020 480 619260 0 FreeSans 960 0 0 0 io_out[25]
port 122 nsew signal tristate
flabel metal3 s -960 566796 480 567036 0 FreeSans 960 0 0 0 io_out[26]
port 123 nsew signal tristate
flabel metal3 s -960 514708 480 514948 0 FreeSans 960 0 0 0 io_out[27]
port 124 nsew signal tristate
flabel metal3 s -960 462484 480 462724 0 FreeSans 960 0 0 0 io_out[28]
port 125 nsew signal tristate
flabel metal3 s -960 410396 480 410636 0 FreeSans 960 0 0 0 io_out[29]
port 126 nsew signal tristate
flabel metal3 s 583520 99364 584960 99604 0 FreeSans 960 0 0 0 io_out[2]
port 127 nsew signal tristate
flabel metal3 s -960 358308 480 358548 0 FreeSans 960 0 0 0 io_out[30]
port 128 nsew signal tristate
flabel metal3 s -960 306084 480 306324 0 FreeSans 960 0 0 0 io_out[31]
port 129 nsew signal tristate
flabel metal3 s -960 253996 480 254236 0 FreeSans 960 0 0 0 io_out[32]
port 130 nsew signal tristate
flabel metal3 s -960 201772 480 202012 0 FreeSans 960 0 0 0 io_out[33]
port 131 nsew signal tristate
flabel metal3 s -960 149684 480 149924 0 FreeSans 960 0 0 0 io_out[34]
port 132 nsew signal tristate
flabel metal3 s -960 97460 480 97700 0 FreeSans 960 0 0 0 io_out[35]
port 133 nsew signal tristate
flabel metal3 s -960 58428 480 58668 0 FreeSans 960 0 0 0 io_out[36]
port 134 nsew signal tristate
flabel metal3 s -960 19260 480 19500 0 FreeSans 960 0 0 0 io_out[37]
port 135 nsew signal tristate
flabel metal3 s 583520 139212 584960 139452 0 FreeSans 960 0 0 0 io_out[3]
port 136 nsew signal tristate
flabel metal3 s 583520 179060 584960 179300 0 FreeSans 960 0 0 0 io_out[4]
port 137 nsew signal tristate
flabel metal3 s 583520 218908 584960 219148 0 FreeSans 960 0 0 0 io_out[5]
port 138 nsew signal tristate
flabel metal3 s 583520 258756 584960 258996 0 FreeSans 960 0 0 0 io_out[6]
port 139 nsew signal tristate
flabel metal3 s 583520 311932 584960 312172 0 FreeSans 960 0 0 0 io_out[7]
port 140 nsew signal tristate
flabel metal3 s 583520 364972 584960 365212 0 FreeSans 960 0 0 0 io_out[8]
port 141 nsew signal tristate
flabel metal3 s 583520 418148 584960 418388 0 FreeSans 960 0 0 0 io_out[9]
port 142 nsew signal tristate
flabel metal2 s 125846 -960 125958 480 0 FreeSans 448 90 0 0 la_data_in[0]
port 143 nsew signal input
flabel metal2 s 480506 -960 480618 480 0 FreeSans 448 90 0 0 la_data_in[100]
port 144 nsew signal input
flabel metal2 s 484002 -960 484114 480 0 FreeSans 448 90 0 0 la_data_in[101]
port 145 nsew signal input
flabel metal2 s 487590 -960 487702 480 0 FreeSans 448 90 0 0 la_data_in[102]
port 146 nsew signal input
flabel metal2 s 491086 -960 491198 480 0 FreeSans 448 90 0 0 la_data_in[103]
port 147 nsew signal input
flabel metal2 s 494674 -960 494786 480 0 FreeSans 448 90 0 0 la_data_in[104]
port 148 nsew signal input
flabel metal2 s 498170 -960 498282 480 0 FreeSans 448 90 0 0 la_data_in[105]
port 149 nsew signal input
flabel metal2 s 501758 -960 501870 480 0 FreeSans 448 90 0 0 la_data_in[106]
port 150 nsew signal input
flabel metal2 s 505346 -960 505458 480 0 FreeSans 448 90 0 0 la_data_in[107]
port 151 nsew signal input
flabel metal2 s 508842 -960 508954 480 0 FreeSans 448 90 0 0 la_data_in[108]
port 152 nsew signal input
flabel metal2 s 512430 -960 512542 480 0 FreeSans 448 90 0 0 la_data_in[109]
port 153 nsew signal input
flabel metal2 s 161266 -960 161378 480 0 FreeSans 448 90 0 0 la_data_in[10]
port 154 nsew signal input
flabel metal2 s 515926 -960 516038 480 0 FreeSans 448 90 0 0 la_data_in[110]
port 155 nsew signal input
flabel metal2 s 519514 -960 519626 480 0 FreeSans 448 90 0 0 la_data_in[111]
port 156 nsew signal input
flabel metal2 s 523010 -960 523122 480 0 FreeSans 448 90 0 0 la_data_in[112]
port 157 nsew signal input
flabel metal2 s 526598 -960 526710 480 0 FreeSans 448 90 0 0 la_data_in[113]
port 158 nsew signal input
flabel metal2 s 530094 -960 530206 480 0 FreeSans 448 90 0 0 la_data_in[114]
port 159 nsew signal input
flabel metal2 s 533682 -960 533794 480 0 FreeSans 448 90 0 0 la_data_in[115]
port 160 nsew signal input
flabel metal2 s 537178 -960 537290 480 0 FreeSans 448 90 0 0 la_data_in[116]
port 161 nsew signal input
flabel metal2 s 540766 -960 540878 480 0 FreeSans 448 90 0 0 la_data_in[117]
port 162 nsew signal input
flabel metal2 s 544354 -960 544466 480 0 FreeSans 448 90 0 0 la_data_in[118]
port 163 nsew signal input
flabel metal2 s 547850 -960 547962 480 0 FreeSans 448 90 0 0 la_data_in[119]
port 164 nsew signal input
flabel metal2 s 164854 -960 164966 480 0 FreeSans 448 90 0 0 la_data_in[11]
port 165 nsew signal input
flabel metal2 s 551438 -960 551550 480 0 FreeSans 448 90 0 0 la_data_in[120]
port 166 nsew signal input
flabel metal2 s 554934 -960 555046 480 0 FreeSans 448 90 0 0 la_data_in[121]
port 167 nsew signal input
flabel metal2 s 558522 -960 558634 480 0 FreeSans 448 90 0 0 la_data_in[122]
port 168 nsew signal input
flabel metal2 s 562018 -960 562130 480 0 FreeSans 448 90 0 0 la_data_in[123]
port 169 nsew signal input
flabel metal2 s 565606 -960 565718 480 0 FreeSans 448 90 0 0 la_data_in[124]
port 170 nsew signal input
flabel metal2 s 569102 -960 569214 480 0 FreeSans 448 90 0 0 la_data_in[125]
port 171 nsew signal input
flabel metal2 s 572690 -960 572802 480 0 FreeSans 448 90 0 0 la_data_in[126]
port 172 nsew signal input
flabel metal2 s 576278 -960 576390 480 0 FreeSans 448 90 0 0 la_data_in[127]
port 173 nsew signal input
flabel metal2 s 168350 -960 168462 480 0 FreeSans 448 90 0 0 la_data_in[12]
port 174 nsew signal input
flabel metal2 s 171938 -960 172050 480 0 FreeSans 448 90 0 0 la_data_in[13]
port 175 nsew signal input
flabel metal2 s 175434 -960 175546 480 0 FreeSans 448 90 0 0 la_data_in[14]
port 176 nsew signal input
flabel metal2 s 179022 -960 179134 480 0 FreeSans 448 90 0 0 la_data_in[15]
port 177 nsew signal input
flabel metal2 s 182518 -960 182630 480 0 FreeSans 448 90 0 0 la_data_in[16]
port 178 nsew signal input
flabel metal2 s 186106 -960 186218 480 0 FreeSans 448 90 0 0 la_data_in[17]
port 179 nsew signal input
flabel metal2 s 189694 -960 189806 480 0 FreeSans 448 90 0 0 la_data_in[18]
port 180 nsew signal input
flabel metal2 s 193190 -960 193302 480 0 FreeSans 448 90 0 0 la_data_in[19]
port 181 nsew signal input
flabel metal2 s 129342 -960 129454 480 0 FreeSans 448 90 0 0 la_data_in[1]
port 182 nsew signal input
flabel metal2 s 196778 -960 196890 480 0 FreeSans 448 90 0 0 la_data_in[20]
port 183 nsew signal input
flabel metal2 s 200274 -960 200386 480 0 FreeSans 448 90 0 0 la_data_in[21]
port 184 nsew signal input
flabel metal2 s 203862 -960 203974 480 0 FreeSans 448 90 0 0 la_data_in[22]
port 185 nsew signal input
flabel metal2 s 207358 -960 207470 480 0 FreeSans 448 90 0 0 la_data_in[23]
port 186 nsew signal input
flabel metal2 s 210946 -960 211058 480 0 FreeSans 448 90 0 0 la_data_in[24]
port 187 nsew signal input
flabel metal2 s 214442 -960 214554 480 0 FreeSans 448 90 0 0 la_data_in[25]
port 188 nsew signal input
flabel metal2 s 218030 -960 218142 480 0 FreeSans 448 90 0 0 la_data_in[26]
port 189 nsew signal input
flabel metal2 s 221526 -960 221638 480 0 FreeSans 448 90 0 0 la_data_in[27]
port 190 nsew signal input
flabel metal2 s 225114 -960 225226 480 0 FreeSans 448 90 0 0 la_data_in[28]
port 191 nsew signal input
flabel metal2 s 228702 -960 228814 480 0 FreeSans 448 90 0 0 la_data_in[29]
port 192 nsew signal input
flabel metal2 s 132930 -960 133042 480 0 FreeSans 448 90 0 0 la_data_in[2]
port 193 nsew signal input
flabel metal2 s 232198 -960 232310 480 0 FreeSans 448 90 0 0 la_data_in[30]
port 194 nsew signal input
flabel metal2 s 235786 -960 235898 480 0 FreeSans 448 90 0 0 la_data_in[31]
port 195 nsew signal input
flabel metal2 s 239282 -960 239394 480 0 FreeSans 448 90 0 0 la_data_in[32]
port 196 nsew signal input
flabel metal2 s 242870 -960 242982 480 0 FreeSans 448 90 0 0 la_data_in[33]
port 197 nsew signal input
flabel metal2 s 246366 -960 246478 480 0 FreeSans 448 90 0 0 la_data_in[34]
port 198 nsew signal input
flabel metal2 s 249954 -960 250066 480 0 FreeSans 448 90 0 0 la_data_in[35]
port 199 nsew signal input
flabel metal2 s 253450 -960 253562 480 0 FreeSans 448 90 0 0 la_data_in[36]
port 200 nsew signal input
flabel metal2 s 257038 -960 257150 480 0 FreeSans 448 90 0 0 la_data_in[37]
port 201 nsew signal input
flabel metal2 s 260626 -960 260738 480 0 FreeSans 448 90 0 0 la_data_in[38]
port 202 nsew signal input
flabel metal2 s 264122 -960 264234 480 0 FreeSans 448 90 0 0 la_data_in[39]
port 203 nsew signal input
flabel metal2 s 136426 -960 136538 480 0 FreeSans 448 90 0 0 la_data_in[3]
port 204 nsew signal input
flabel metal2 s 267710 -960 267822 480 0 FreeSans 448 90 0 0 la_data_in[40]
port 205 nsew signal input
flabel metal2 s 271206 -960 271318 480 0 FreeSans 448 90 0 0 la_data_in[41]
port 206 nsew signal input
flabel metal2 s 274794 -960 274906 480 0 FreeSans 448 90 0 0 la_data_in[42]
port 207 nsew signal input
flabel metal2 s 278290 -960 278402 480 0 FreeSans 448 90 0 0 la_data_in[43]
port 208 nsew signal input
flabel metal2 s 281878 -960 281990 480 0 FreeSans 448 90 0 0 la_data_in[44]
port 209 nsew signal input
flabel metal2 s 285374 -960 285486 480 0 FreeSans 448 90 0 0 la_data_in[45]
port 210 nsew signal input
flabel metal2 s 288962 -960 289074 480 0 FreeSans 448 90 0 0 la_data_in[46]
port 211 nsew signal input
flabel metal2 s 292550 -960 292662 480 0 FreeSans 448 90 0 0 la_data_in[47]
port 212 nsew signal input
flabel metal2 s 296046 -960 296158 480 0 FreeSans 448 90 0 0 la_data_in[48]
port 213 nsew signal input
flabel metal2 s 299634 -960 299746 480 0 FreeSans 448 90 0 0 la_data_in[49]
port 214 nsew signal input
flabel metal2 s 140014 -960 140126 480 0 FreeSans 448 90 0 0 la_data_in[4]
port 215 nsew signal input
flabel metal2 s 303130 -960 303242 480 0 FreeSans 448 90 0 0 la_data_in[50]
port 216 nsew signal input
flabel metal2 s 306718 -960 306830 480 0 FreeSans 448 90 0 0 la_data_in[51]
port 217 nsew signal input
flabel metal2 s 310214 -960 310326 480 0 FreeSans 448 90 0 0 la_data_in[52]
port 218 nsew signal input
flabel metal2 s 313802 -960 313914 480 0 FreeSans 448 90 0 0 la_data_in[53]
port 219 nsew signal input
flabel metal2 s 317298 -960 317410 480 0 FreeSans 448 90 0 0 la_data_in[54]
port 220 nsew signal input
flabel metal2 s 320886 -960 320998 480 0 FreeSans 448 90 0 0 la_data_in[55]
port 221 nsew signal input
flabel metal2 s 324382 -960 324494 480 0 FreeSans 448 90 0 0 la_data_in[56]
port 222 nsew signal input
flabel metal2 s 327970 -960 328082 480 0 FreeSans 448 90 0 0 la_data_in[57]
port 223 nsew signal input
flabel metal2 s 331558 -960 331670 480 0 FreeSans 448 90 0 0 la_data_in[58]
port 224 nsew signal input
flabel metal2 s 335054 -960 335166 480 0 FreeSans 448 90 0 0 la_data_in[59]
port 225 nsew signal input
flabel metal2 s 143510 -960 143622 480 0 FreeSans 448 90 0 0 la_data_in[5]
port 226 nsew signal input
flabel metal2 s 338642 -960 338754 480 0 FreeSans 448 90 0 0 la_data_in[60]
port 227 nsew signal input
flabel metal2 s 342138 -960 342250 480 0 FreeSans 448 90 0 0 la_data_in[61]
port 228 nsew signal input
flabel metal2 s 345726 -960 345838 480 0 FreeSans 448 90 0 0 la_data_in[62]
port 229 nsew signal input
flabel metal2 s 349222 -960 349334 480 0 FreeSans 448 90 0 0 la_data_in[63]
port 230 nsew signal input
flabel metal2 s 352810 -960 352922 480 0 FreeSans 448 90 0 0 la_data_in[64]
port 231 nsew signal input
flabel metal2 s 356306 -960 356418 480 0 FreeSans 448 90 0 0 la_data_in[65]
port 232 nsew signal input
flabel metal2 s 359894 -960 360006 480 0 FreeSans 448 90 0 0 la_data_in[66]
port 233 nsew signal input
flabel metal2 s 363482 -960 363594 480 0 FreeSans 448 90 0 0 la_data_in[67]
port 234 nsew signal input
flabel metal2 s 366978 -960 367090 480 0 FreeSans 448 90 0 0 la_data_in[68]
port 235 nsew signal input
flabel metal2 s 370566 -960 370678 480 0 FreeSans 448 90 0 0 la_data_in[69]
port 236 nsew signal input
flabel metal2 s 147098 -960 147210 480 0 FreeSans 448 90 0 0 la_data_in[6]
port 237 nsew signal input
flabel metal2 s 374062 -960 374174 480 0 FreeSans 448 90 0 0 la_data_in[70]
port 238 nsew signal input
flabel metal2 s 377650 -960 377762 480 0 FreeSans 448 90 0 0 la_data_in[71]
port 239 nsew signal input
flabel metal2 s 381146 -960 381258 480 0 FreeSans 448 90 0 0 la_data_in[72]
port 240 nsew signal input
flabel metal2 s 384734 -960 384846 480 0 FreeSans 448 90 0 0 la_data_in[73]
port 241 nsew signal input
flabel metal2 s 388230 -960 388342 480 0 FreeSans 448 90 0 0 la_data_in[74]
port 242 nsew signal input
flabel metal2 s 391818 -960 391930 480 0 FreeSans 448 90 0 0 la_data_in[75]
port 243 nsew signal input
flabel metal2 s 395314 -960 395426 480 0 FreeSans 448 90 0 0 la_data_in[76]
port 244 nsew signal input
flabel metal2 s 398902 -960 399014 480 0 FreeSans 448 90 0 0 la_data_in[77]
port 245 nsew signal input
flabel metal2 s 402490 -960 402602 480 0 FreeSans 448 90 0 0 la_data_in[78]
port 246 nsew signal input
flabel metal2 s 405986 -960 406098 480 0 FreeSans 448 90 0 0 la_data_in[79]
port 247 nsew signal input
flabel metal2 s 150594 -960 150706 480 0 FreeSans 448 90 0 0 la_data_in[7]
port 248 nsew signal input
flabel metal2 s 409574 -960 409686 480 0 FreeSans 448 90 0 0 la_data_in[80]
port 249 nsew signal input
flabel metal2 s 413070 -960 413182 480 0 FreeSans 448 90 0 0 la_data_in[81]
port 250 nsew signal input
flabel metal2 s 416658 -960 416770 480 0 FreeSans 448 90 0 0 la_data_in[82]
port 251 nsew signal input
flabel metal2 s 420154 -960 420266 480 0 FreeSans 448 90 0 0 la_data_in[83]
port 252 nsew signal input
flabel metal2 s 423742 -960 423854 480 0 FreeSans 448 90 0 0 la_data_in[84]
port 253 nsew signal input
flabel metal2 s 427238 -960 427350 480 0 FreeSans 448 90 0 0 la_data_in[85]
port 254 nsew signal input
flabel metal2 s 430826 -960 430938 480 0 FreeSans 448 90 0 0 la_data_in[86]
port 255 nsew signal input
flabel metal2 s 434414 -960 434526 480 0 FreeSans 448 90 0 0 la_data_in[87]
port 256 nsew signal input
flabel metal2 s 437910 -960 438022 480 0 FreeSans 448 90 0 0 la_data_in[88]
port 257 nsew signal input
flabel metal2 s 441498 -960 441610 480 0 FreeSans 448 90 0 0 la_data_in[89]
port 258 nsew signal input
flabel metal2 s 154182 -960 154294 480 0 FreeSans 448 90 0 0 la_data_in[8]
port 259 nsew signal input
flabel metal2 s 444994 -960 445106 480 0 FreeSans 448 90 0 0 la_data_in[90]
port 260 nsew signal input
flabel metal2 s 448582 -960 448694 480 0 FreeSans 448 90 0 0 la_data_in[91]
port 261 nsew signal input
flabel metal2 s 452078 -960 452190 480 0 FreeSans 448 90 0 0 la_data_in[92]
port 262 nsew signal input
flabel metal2 s 455666 -960 455778 480 0 FreeSans 448 90 0 0 la_data_in[93]
port 263 nsew signal input
flabel metal2 s 459162 -960 459274 480 0 FreeSans 448 90 0 0 la_data_in[94]
port 264 nsew signal input
flabel metal2 s 462750 -960 462862 480 0 FreeSans 448 90 0 0 la_data_in[95]
port 265 nsew signal input
flabel metal2 s 466246 -960 466358 480 0 FreeSans 448 90 0 0 la_data_in[96]
port 266 nsew signal input
flabel metal2 s 469834 -960 469946 480 0 FreeSans 448 90 0 0 la_data_in[97]
port 267 nsew signal input
flabel metal2 s 473422 -960 473534 480 0 FreeSans 448 90 0 0 la_data_in[98]
port 268 nsew signal input
flabel metal2 s 476918 -960 477030 480 0 FreeSans 448 90 0 0 la_data_in[99]
port 269 nsew signal input
flabel metal2 s 157770 -960 157882 480 0 FreeSans 448 90 0 0 la_data_in[9]
port 270 nsew signal input
flabel metal2 s 126950 -960 127062 480 0 FreeSans 448 90 0 0 la_data_out[0]
port 271 nsew signal tristate
flabel metal2 s 481702 -960 481814 480 0 FreeSans 448 90 0 0 la_data_out[100]
port 272 nsew signal tristate
flabel metal2 s 485198 -960 485310 480 0 FreeSans 448 90 0 0 la_data_out[101]
port 273 nsew signal tristate
flabel metal2 s 488786 -960 488898 480 0 FreeSans 448 90 0 0 la_data_out[102]
port 274 nsew signal tristate
flabel metal2 s 492282 -960 492394 480 0 FreeSans 448 90 0 0 la_data_out[103]
port 275 nsew signal tristate
flabel metal2 s 495870 -960 495982 480 0 FreeSans 448 90 0 0 la_data_out[104]
port 276 nsew signal tristate
flabel metal2 s 499366 -960 499478 480 0 FreeSans 448 90 0 0 la_data_out[105]
port 277 nsew signal tristate
flabel metal2 s 502954 -960 503066 480 0 FreeSans 448 90 0 0 la_data_out[106]
port 278 nsew signal tristate
flabel metal2 s 506450 -960 506562 480 0 FreeSans 448 90 0 0 la_data_out[107]
port 279 nsew signal tristate
flabel metal2 s 510038 -960 510150 480 0 FreeSans 448 90 0 0 la_data_out[108]
port 280 nsew signal tristate
flabel metal2 s 513534 -960 513646 480 0 FreeSans 448 90 0 0 la_data_out[109]
port 281 nsew signal tristate
flabel metal2 s 162462 -960 162574 480 0 FreeSans 448 90 0 0 la_data_out[10]
port 282 nsew signal tristate
flabel metal2 s 517122 -960 517234 480 0 FreeSans 448 90 0 0 la_data_out[110]
port 283 nsew signal tristate
flabel metal2 s 520710 -960 520822 480 0 FreeSans 448 90 0 0 la_data_out[111]
port 284 nsew signal tristate
flabel metal2 s 524206 -960 524318 480 0 FreeSans 448 90 0 0 la_data_out[112]
port 285 nsew signal tristate
flabel metal2 s 527794 -960 527906 480 0 FreeSans 448 90 0 0 la_data_out[113]
port 286 nsew signal tristate
flabel metal2 s 531290 -960 531402 480 0 FreeSans 448 90 0 0 la_data_out[114]
port 287 nsew signal tristate
flabel metal2 s 534878 -960 534990 480 0 FreeSans 448 90 0 0 la_data_out[115]
port 288 nsew signal tristate
flabel metal2 s 538374 -960 538486 480 0 FreeSans 448 90 0 0 la_data_out[116]
port 289 nsew signal tristate
flabel metal2 s 541962 -960 542074 480 0 FreeSans 448 90 0 0 la_data_out[117]
port 290 nsew signal tristate
flabel metal2 s 545458 -960 545570 480 0 FreeSans 448 90 0 0 la_data_out[118]
port 291 nsew signal tristate
flabel metal2 s 549046 -960 549158 480 0 FreeSans 448 90 0 0 la_data_out[119]
port 292 nsew signal tristate
flabel metal2 s 166050 -960 166162 480 0 FreeSans 448 90 0 0 la_data_out[11]
port 293 nsew signal tristate
flabel metal2 s 552634 -960 552746 480 0 FreeSans 448 90 0 0 la_data_out[120]
port 294 nsew signal tristate
flabel metal2 s 556130 -960 556242 480 0 FreeSans 448 90 0 0 la_data_out[121]
port 295 nsew signal tristate
flabel metal2 s 559718 -960 559830 480 0 FreeSans 448 90 0 0 la_data_out[122]
port 296 nsew signal tristate
flabel metal2 s 563214 -960 563326 480 0 FreeSans 448 90 0 0 la_data_out[123]
port 297 nsew signal tristate
flabel metal2 s 566802 -960 566914 480 0 FreeSans 448 90 0 0 la_data_out[124]
port 298 nsew signal tristate
flabel metal2 s 570298 -960 570410 480 0 FreeSans 448 90 0 0 la_data_out[125]
port 299 nsew signal tristate
flabel metal2 s 573886 -960 573998 480 0 FreeSans 448 90 0 0 la_data_out[126]
port 300 nsew signal tristate
flabel metal2 s 577382 -960 577494 480 0 FreeSans 448 90 0 0 la_data_out[127]
port 301 nsew signal tristate
flabel metal2 s 169546 -960 169658 480 0 FreeSans 448 90 0 0 la_data_out[12]
port 302 nsew signal tristate
flabel metal2 s 173134 -960 173246 480 0 FreeSans 448 90 0 0 la_data_out[13]
port 303 nsew signal tristate
flabel metal2 s 176630 -960 176742 480 0 FreeSans 448 90 0 0 la_data_out[14]
port 304 nsew signal tristate
flabel metal2 s 180218 -960 180330 480 0 FreeSans 448 90 0 0 la_data_out[15]
port 305 nsew signal tristate
flabel metal2 s 183714 -960 183826 480 0 FreeSans 448 90 0 0 la_data_out[16]
port 306 nsew signal tristate
flabel metal2 s 187302 -960 187414 480 0 FreeSans 448 90 0 0 la_data_out[17]
port 307 nsew signal tristate
flabel metal2 s 190798 -960 190910 480 0 FreeSans 448 90 0 0 la_data_out[18]
port 308 nsew signal tristate
flabel metal2 s 194386 -960 194498 480 0 FreeSans 448 90 0 0 la_data_out[19]
port 309 nsew signal tristate
flabel metal2 s 130538 -960 130650 480 0 FreeSans 448 90 0 0 la_data_out[1]
port 310 nsew signal tristate
flabel metal2 s 197882 -960 197994 480 0 FreeSans 448 90 0 0 la_data_out[20]
port 311 nsew signal tristate
flabel metal2 s 201470 -960 201582 480 0 FreeSans 448 90 0 0 la_data_out[21]
port 312 nsew signal tristate
flabel metal2 s 205058 -960 205170 480 0 FreeSans 448 90 0 0 la_data_out[22]
port 313 nsew signal tristate
flabel metal2 s 208554 -960 208666 480 0 FreeSans 448 90 0 0 la_data_out[23]
port 314 nsew signal tristate
flabel metal2 s 212142 -960 212254 480 0 FreeSans 448 90 0 0 la_data_out[24]
port 315 nsew signal tristate
flabel metal2 s 215638 -960 215750 480 0 FreeSans 448 90 0 0 la_data_out[25]
port 316 nsew signal tristate
flabel metal2 s 219226 -960 219338 480 0 FreeSans 448 90 0 0 la_data_out[26]
port 317 nsew signal tristate
flabel metal2 s 222722 -960 222834 480 0 FreeSans 448 90 0 0 la_data_out[27]
port 318 nsew signal tristate
flabel metal2 s 226310 -960 226422 480 0 FreeSans 448 90 0 0 la_data_out[28]
port 319 nsew signal tristate
flabel metal2 s 229806 -960 229918 480 0 FreeSans 448 90 0 0 la_data_out[29]
port 320 nsew signal tristate
flabel metal2 s 134126 -960 134238 480 0 FreeSans 448 90 0 0 la_data_out[2]
port 321 nsew signal tristate
flabel metal2 s 233394 -960 233506 480 0 FreeSans 448 90 0 0 la_data_out[30]
port 322 nsew signal tristate
flabel metal2 s 236982 -960 237094 480 0 FreeSans 448 90 0 0 la_data_out[31]
port 323 nsew signal tristate
flabel metal2 s 240478 -960 240590 480 0 FreeSans 448 90 0 0 la_data_out[32]
port 324 nsew signal tristate
flabel metal2 s 244066 -960 244178 480 0 FreeSans 448 90 0 0 la_data_out[33]
port 325 nsew signal tristate
flabel metal2 s 247562 -960 247674 480 0 FreeSans 448 90 0 0 la_data_out[34]
port 326 nsew signal tristate
flabel metal2 s 251150 -960 251262 480 0 FreeSans 448 90 0 0 la_data_out[35]
port 327 nsew signal tristate
flabel metal2 s 254646 -960 254758 480 0 FreeSans 448 90 0 0 la_data_out[36]
port 328 nsew signal tristate
flabel metal2 s 258234 -960 258346 480 0 FreeSans 448 90 0 0 la_data_out[37]
port 329 nsew signal tristate
flabel metal2 s 261730 -960 261842 480 0 FreeSans 448 90 0 0 la_data_out[38]
port 330 nsew signal tristate
flabel metal2 s 265318 -960 265430 480 0 FreeSans 448 90 0 0 la_data_out[39]
port 331 nsew signal tristate
flabel metal2 s 137622 -960 137734 480 0 FreeSans 448 90 0 0 la_data_out[3]
port 332 nsew signal tristate
flabel metal2 s 268814 -960 268926 480 0 FreeSans 448 90 0 0 la_data_out[40]
port 333 nsew signal tristate
flabel metal2 s 272402 -960 272514 480 0 FreeSans 448 90 0 0 la_data_out[41]
port 334 nsew signal tristate
flabel metal2 s 275990 -960 276102 480 0 FreeSans 448 90 0 0 la_data_out[42]
port 335 nsew signal tristate
flabel metal2 s 279486 -960 279598 480 0 FreeSans 448 90 0 0 la_data_out[43]
port 336 nsew signal tristate
flabel metal2 s 283074 -960 283186 480 0 FreeSans 448 90 0 0 la_data_out[44]
port 337 nsew signal tristate
flabel metal2 s 286570 -960 286682 480 0 FreeSans 448 90 0 0 la_data_out[45]
port 338 nsew signal tristate
flabel metal2 s 290158 -960 290270 480 0 FreeSans 448 90 0 0 la_data_out[46]
port 339 nsew signal tristate
flabel metal2 s 293654 -960 293766 480 0 FreeSans 448 90 0 0 la_data_out[47]
port 340 nsew signal tristate
flabel metal2 s 297242 -960 297354 480 0 FreeSans 448 90 0 0 la_data_out[48]
port 341 nsew signal tristate
flabel metal2 s 300738 -960 300850 480 0 FreeSans 448 90 0 0 la_data_out[49]
port 342 nsew signal tristate
flabel metal2 s 141210 -960 141322 480 0 FreeSans 448 90 0 0 la_data_out[4]
port 343 nsew signal tristate
flabel metal2 s 304326 -960 304438 480 0 FreeSans 448 90 0 0 la_data_out[50]
port 344 nsew signal tristate
flabel metal2 s 307914 -960 308026 480 0 FreeSans 448 90 0 0 la_data_out[51]
port 345 nsew signal tristate
flabel metal2 s 311410 -960 311522 480 0 FreeSans 448 90 0 0 la_data_out[52]
port 346 nsew signal tristate
flabel metal2 s 314998 -960 315110 480 0 FreeSans 448 90 0 0 la_data_out[53]
port 347 nsew signal tristate
flabel metal2 s 318494 -960 318606 480 0 FreeSans 448 90 0 0 la_data_out[54]
port 348 nsew signal tristate
flabel metal2 s 322082 -960 322194 480 0 FreeSans 448 90 0 0 la_data_out[55]
port 349 nsew signal tristate
flabel metal2 s 325578 -960 325690 480 0 FreeSans 448 90 0 0 la_data_out[56]
port 350 nsew signal tristate
flabel metal2 s 329166 -960 329278 480 0 FreeSans 448 90 0 0 la_data_out[57]
port 351 nsew signal tristate
flabel metal2 s 332662 -960 332774 480 0 FreeSans 448 90 0 0 la_data_out[58]
port 352 nsew signal tristate
flabel metal2 s 336250 -960 336362 480 0 FreeSans 448 90 0 0 la_data_out[59]
port 353 nsew signal tristate
flabel metal2 s 144706 -960 144818 480 0 FreeSans 448 90 0 0 la_data_out[5]
port 354 nsew signal tristate
flabel metal2 s 339838 -960 339950 480 0 FreeSans 448 90 0 0 la_data_out[60]
port 355 nsew signal tristate
flabel metal2 s 343334 -960 343446 480 0 FreeSans 448 90 0 0 la_data_out[61]
port 356 nsew signal tristate
flabel metal2 s 346922 -960 347034 480 0 FreeSans 448 90 0 0 la_data_out[62]
port 357 nsew signal tristate
flabel metal2 s 350418 -960 350530 480 0 FreeSans 448 90 0 0 la_data_out[63]
port 358 nsew signal tristate
flabel metal2 s 354006 -960 354118 480 0 FreeSans 448 90 0 0 la_data_out[64]
port 359 nsew signal tristate
flabel metal2 s 357502 -960 357614 480 0 FreeSans 448 90 0 0 la_data_out[65]
port 360 nsew signal tristate
flabel metal2 s 361090 -960 361202 480 0 FreeSans 448 90 0 0 la_data_out[66]
port 361 nsew signal tristate
flabel metal2 s 364586 -960 364698 480 0 FreeSans 448 90 0 0 la_data_out[67]
port 362 nsew signal tristate
flabel metal2 s 368174 -960 368286 480 0 FreeSans 448 90 0 0 la_data_out[68]
port 363 nsew signal tristate
flabel metal2 s 371670 -960 371782 480 0 FreeSans 448 90 0 0 la_data_out[69]
port 364 nsew signal tristate
flabel metal2 s 148294 -960 148406 480 0 FreeSans 448 90 0 0 la_data_out[6]
port 365 nsew signal tristate
flabel metal2 s 375258 -960 375370 480 0 FreeSans 448 90 0 0 la_data_out[70]
port 366 nsew signal tristate
flabel metal2 s 378846 -960 378958 480 0 FreeSans 448 90 0 0 la_data_out[71]
port 367 nsew signal tristate
flabel metal2 s 382342 -960 382454 480 0 FreeSans 448 90 0 0 la_data_out[72]
port 368 nsew signal tristate
flabel metal2 s 385930 -960 386042 480 0 FreeSans 448 90 0 0 la_data_out[73]
port 369 nsew signal tristate
flabel metal2 s 389426 -960 389538 480 0 FreeSans 448 90 0 0 la_data_out[74]
port 370 nsew signal tristate
flabel metal2 s 393014 -960 393126 480 0 FreeSans 448 90 0 0 la_data_out[75]
port 371 nsew signal tristate
flabel metal2 s 396510 -960 396622 480 0 FreeSans 448 90 0 0 la_data_out[76]
port 372 nsew signal tristate
flabel metal2 s 400098 -960 400210 480 0 FreeSans 448 90 0 0 la_data_out[77]
port 373 nsew signal tristate
flabel metal2 s 403594 -960 403706 480 0 FreeSans 448 90 0 0 la_data_out[78]
port 374 nsew signal tristate
flabel metal2 s 407182 -960 407294 480 0 FreeSans 448 90 0 0 la_data_out[79]
port 375 nsew signal tristate
flabel metal2 s 151790 -960 151902 480 0 FreeSans 448 90 0 0 la_data_out[7]
port 376 nsew signal tristate
flabel metal2 s 410770 -960 410882 480 0 FreeSans 448 90 0 0 la_data_out[80]
port 377 nsew signal tristate
flabel metal2 s 414266 -960 414378 480 0 FreeSans 448 90 0 0 la_data_out[81]
port 378 nsew signal tristate
flabel metal2 s 417854 -960 417966 480 0 FreeSans 448 90 0 0 la_data_out[82]
port 379 nsew signal tristate
flabel metal2 s 421350 -960 421462 480 0 FreeSans 448 90 0 0 la_data_out[83]
port 380 nsew signal tristate
flabel metal2 s 424938 -960 425050 480 0 FreeSans 448 90 0 0 la_data_out[84]
port 381 nsew signal tristate
flabel metal2 s 428434 -960 428546 480 0 FreeSans 448 90 0 0 la_data_out[85]
port 382 nsew signal tristate
flabel metal2 s 432022 -960 432134 480 0 FreeSans 448 90 0 0 la_data_out[86]
port 383 nsew signal tristate
flabel metal2 s 435518 -960 435630 480 0 FreeSans 448 90 0 0 la_data_out[87]
port 384 nsew signal tristate
flabel metal2 s 439106 -960 439218 480 0 FreeSans 448 90 0 0 la_data_out[88]
port 385 nsew signal tristate
flabel metal2 s 442602 -960 442714 480 0 FreeSans 448 90 0 0 la_data_out[89]
port 386 nsew signal tristate
flabel metal2 s 155378 -960 155490 480 0 FreeSans 448 90 0 0 la_data_out[8]
port 387 nsew signal tristate
flabel metal2 s 446190 -960 446302 480 0 FreeSans 448 90 0 0 la_data_out[90]
port 388 nsew signal tristate
flabel metal2 s 449778 -960 449890 480 0 FreeSans 448 90 0 0 la_data_out[91]
port 389 nsew signal tristate
flabel metal2 s 453274 -960 453386 480 0 FreeSans 448 90 0 0 la_data_out[92]
port 390 nsew signal tristate
flabel metal2 s 456862 -960 456974 480 0 FreeSans 448 90 0 0 la_data_out[93]
port 391 nsew signal tristate
flabel metal2 s 460358 -960 460470 480 0 FreeSans 448 90 0 0 la_data_out[94]
port 392 nsew signal tristate
flabel metal2 s 463946 -960 464058 480 0 FreeSans 448 90 0 0 la_data_out[95]
port 393 nsew signal tristate
flabel metal2 s 467442 -960 467554 480 0 FreeSans 448 90 0 0 la_data_out[96]
port 394 nsew signal tristate
flabel metal2 s 471030 -960 471142 480 0 FreeSans 448 90 0 0 la_data_out[97]
port 395 nsew signal tristate
flabel metal2 s 474526 -960 474638 480 0 FreeSans 448 90 0 0 la_data_out[98]
port 396 nsew signal tristate
flabel metal2 s 478114 -960 478226 480 0 FreeSans 448 90 0 0 la_data_out[99]
port 397 nsew signal tristate
flabel metal2 s 158874 -960 158986 480 0 FreeSans 448 90 0 0 la_data_out[9]
port 398 nsew signal tristate
flabel metal2 s 128146 -960 128258 480 0 FreeSans 448 90 0 0 la_oenb[0]
port 399 nsew signal input
flabel metal2 s 482806 -960 482918 480 0 FreeSans 448 90 0 0 la_oenb[100]
port 400 nsew signal input
flabel metal2 s 486394 -960 486506 480 0 FreeSans 448 90 0 0 la_oenb[101]
port 401 nsew signal input
flabel metal2 s 489890 -960 490002 480 0 FreeSans 448 90 0 0 la_oenb[102]
port 402 nsew signal input
flabel metal2 s 493478 -960 493590 480 0 FreeSans 448 90 0 0 la_oenb[103]
port 403 nsew signal input
flabel metal2 s 497066 -960 497178 480 0 FreeSans 448 90 0 0 la_oenb[104]
port 404 nsew signal input
flabel metal2 s 500562 -960 500674 480 0 FreeSans 448 90 0 0 la_oenb[105]
port 405 nsew signal input
flabel metal2 s 504150 -960 504262 480 0 FreeSans 448 90 0 0 la_oenb[106]
port 406 nsew signal input
flabel metal2 s 507646 -960 507758 480 0 FreeSans 448 90 0 0 la_oenb[107]
port 407 nsew signal input
flabel metal2 s 511234 -960 511346 480 0 FreeSans 448 90 0 0 la_oenb[108]
port 408 nsew signal input
flabel metal2 s 514730 -960 514842 480 0 FreeSans 448 90 0 0 la_oenb[109]
port 409 nsew signal input
flabel metal2 s 163658 -960 163770 480 0 FreeSans 448 90 0 0 la_oenb[10]
port 410 nsew signal input
flabel metal2 s 518318 -960 518430 480 0 FreeSans 448 90 0 0 la_oenb[110]
port 411 nsew signal input
flabel metal2 s 521814 -960 521926 480 0 FreeSans 448 90 0 0 la_oenb[111]
port 412 nsew signal input
flabel metal2 s 525402 -960 525514 480 0 FreeSans 448 90 0 0 la_oenb[112]
port 413 nsew signal input
flabel metal2 s 528990 -960 529102 480 0 FreeSans 448 90 0 0 la_oenb[113]
port 414 nsew signal input
flabel metal2 s 532486 -960 532598 480 0 FreeSans 448 90 0 0 la_oenb[114]
port 415 nsew signal input
flabel metal2 s 536074 -960 536186 480 0 FreeSans 448 90 0 0 la_oenb[115]
port 416 nsew signal input
flabel metal2 s 539570 -960 539682 480 0 FreeSans 448 90 0 0 la_oenb[116]
port 417 nsew signal input
flabel metal2 s 543158 -960 543270 480 0 FreeSans 448 90 0 0 la_oenb[117]
port 418 nsew signal input
flabel metal2 s 546654 -960 546766 480 0 FreeSans 448 90 0 0 la_oenb[118]
port 419 nsew signal input
flabel metal2 s 550242 -960 550354 480 0 FreeSans 448 90 0 0 la_oenb[119]
port 420 nsew signal input
flabel metal2 s 167154 -960 167266 480 0 FreeSans 448 90 0 0 la_oenb[11]
port 421 nsew signal input
flabel metal2 s 553738 -960 553850 480 0 FreeSans 448 90 0 0 la_oenb[120]
port 422 nsew signal input
flabel metal2 s 557326 -960 557438 480 0 FreeSans 448 90 0 0 la_oenb[121]
port 423 nsew signal input
flabel metal2 s 560822 -960 560934 480 0 FreeSans 448 90 0 0 la_oenb[122]
port 424 nsew signal input
flabel metal2 s 564410 -960 564522 480 0 FreeSans 448 90 0 0 la_oenb[123]
port 425 nsew signal input
flabel metal2 s 567998 -960 568110 480 0 FreeSans 448 90 0 0 la_oenb[124]
port 426 nsew signal input
flabel metal2 s 571494 -960 571606 480 0 FreeSans 448 90 0 0 la_oenb[125]
port 427 nsew signal input
flabel metal2 s 575082 -960 575194 480 0 FreeSans 448 90 0 0 la_oenb[126]
port 428 nsew signal input
flabel metal2 s 578578 -960 578690 480 0 FreeSans 448 90 0 0 la_oenb[127]
port 429 nsew signal input
flabel metal2 s 170742 -960 170854 480 0 FreeSans 448 90 0 0 la_oenb[12]
port 430 nsew signal input
flabel metal2 s 174238 -960 174350 480 0 FreeSans 448 90 0 0 la_oenb[13]
port 431 nsew signal input
flabel metal2 s 177826 -960 177938 480 0 FreeSans 448 90 0 0 la_oenb[14]
port 432 nsew signal input
flabel metal2 s 181414 -960 181526 480 0 FreeSans 448 90 0 0 la_oenb[15]
port 433 nsew signal input
flabel metal2 s 184910 -960 185022 480 0 FreeSans 448 90 0 0 la_oenb[16]
port 434 nsew signal input
flabel metal2 s 188498 -960 188610 480 0 FreeSans 448 90 0 0 la_oenb[17]
port 435 nsew signal input
flabel metal2 s 191994 -960 192106 480 0 FreeSans 448 90 0 0 la_oenb[18]
port 436 nsew signal input
flabel metal2 s 195582 -960 195694 480 0 FreeSans 448 90 0 0 la_oenb[19]
port 437 nsew signal input
flabel metal2 s 131734 -960 131846 480 0 FreeSans 448 90 0 0 la_oenb[1]
port 438 nsew signal input
flabel metal2 s 199078 -960 199190 480 0 FreeSans 448 90 0 0 la_oenb[20]
port 439 nsew signal input
flabel metal2 s 202666 -960 202778 480 0 FreeSans 448 90 0 0 la_oenb[21]
port 440 nsew signal input
flabel metal2 s 206162 -960 206274 480 0 FreeSans 448 90 0 0 la_oenb[22]
port 441 nsew signal input
flabel metal2 s 209750 -960 209862 480 0 FreeSans 448 90 0 0 la_oenb[23]
port 442 nsew signal input
flabel metal2 s 213338 -960 213450 480 0 FreeSans 448 90 0 0 la_oenb[24]
port 443 nsew signal input
flabel metal2 s 216834 -960 216946 480 0 FreeSans 448 90 0 0 la_oenb[25]
port 444 nsew signal input
flabel metal2 s 220422 -960 220534 480 0 FreeSans 448 90 0 0 la_oenb[26]
port 445 nsew signal input
flabel metal2 s 223918 -960 224030 480 0 FreeSans 448 90 0 0 la_oenb[27]
port 446 nsew signal input
flabel metal2 s 227506 -960 227618 480 0 FreeSans 448 90 0 0 la_oenb[28]
port 447 nsew signal input
flabel metal2 s 231002 -960 231114 480 0 FreeSans 448 90 0 0 la_oenb[29]
port 448 nsew signal input
flabel metal2 s 135230 -960 135342 480 0 FreeSans 448 90 0 0 la_oenb[2]
port 449 nsew signal input
flabel metal2 s 234590 -960 234702 480 0 FreeSans 448 90 0 0 la_oenb[30]
port 450 nsew signal input
flabel metal2 s 238086 -960 238198 480 0 FreeSans 448 90 0 0 la_oenb[31]
port 451 nsew signal input
flabel metal2 s 241674 -960 241786 480 0 FreeSans 448 90 0 0 la_oenb[32]
port 452 nsew signal input
flabel metal2 s 245170 -960 245282 480 0 FreeSans 448 90 0 0 la_oenb[33]
port 453 nsew signal input
flabel metal2 s 248758 -960 248870 480 0 FreeSans 448 90 0 0 la_oenb[34]
port 454 nsew signal input
flabel metal2 s 252346 -960 252458 480 0 FreeSans 448 90 0 0 la_oenb[35]
port 455 nsew signal input
flabel metal2 s 255842 -960 255954 480 0 FreeSans 448 90 0 0 la_oenb[36]
port 456 nsew signal input
flabel metal2 s 259430 -960 259542 480 0 FreeSans 448 90 0 0 la_oenb[37]
port 457 nsew signal input
flabel metal2 s 262926 -960 263038 480 0 FreeSans 448 90 0 0 la_oenb[38]
port 458 nsew signal input
flabel metal2 s 266514 -960 266626 480 0 FreeSans 448 90 0 0 la_oenb[39]
port 459 nsew signal input
flabel metal2 s 138818 -960 138930 480 0 FreeSans 448 90 0 0 la_oenb[3]
port 460 nsew signal input
flabel metal2 s 270010 -960 270122 480 0 FreeSans 448 90 0 0 la_oenb[40]
port 461 nsew signal input
flabel metal2 s 273598 -960 273710 480 0 FreeSans 448 90 0 0 la_oenb[41]
port 462 nsew signal input
flabel metal2 s 277094 -960 277206 480 0 FreeSans 448 90 0 0 la_oenb[42]
port 463 nsew signal input
flabel metal2 s 280682 -960 280794 480 0 FreeSans 448 90 0 0 la_oenb[43]
port 464 nsew signal input
flabel metal2 s 284270 -960 284382 480 0 FreeSans 448 90 0 0 la_oenb[44]
port 465 nsew signal input
flabel metal2 s 287766 -960 287878 480 0 FreeSans 448 90 0 0 la_oenb[45]
port 466 nsew signal input
flabel metal2 s 291354 -960 291466 480 0 FreeSans 448 90 0 0 la_oenb[46]
port 467 nsew signal input
flabel metal2 s 294850 -960 294962 480 0 FreeSans 448 90 0 0 la_oenb[47]
port 468 nsew signal input
flabel metal2 s 298438 -960 298550 480 0 FreeSans 448 90 0 0 la_oenb[48]
port 469 nsew signal input
flabel metal2 s 301934 -960 302046 480 0 FreeSans 448 90 0 0 la_oenb[49]
port 470 nsew signal input
flabel metal2 s 142406 -960 142518 480 0 FreeSans 448 90 0 0 la_oenb[4]
port 471 nsew signal input
flabel metal2 s 305522 -960 305634 480 0 FreeSans 448 90 0 0 la_oenb[50]
port 472 nsew signal input
flabel metal2 s 309018 -960 309130 480 0 FreeSans 448 90 0 0 la_oenb[51]
port 473 nsew signal input
flabel metal2 s 312606 -960 312718 480 0 FreeSans 448 90 0 0 la_oenb[52]
port 474 nsew signal input
flabel metal2 s 316194 -960 316306 480 0 FreeSans 448 90 0 0 la_oenb[53]
port 475 nsew signal input
flabel metal2 s 319690 -960 319802 480 0 FreeSans 448 90 0 0 la_oenb[54]
port 476 nsew signal input
flabel metal2 s 323278 -960 323390 480 0 FreeSans 448 90 0 0 la_oenb[55]
port 477 nsew signal input
flabel metal2 s 326774 -960 326886 480 0 FreeSans 448 90 0 0 la_oenb[56]
port 478 nsew signal input
flabel metal2 s 330362 -960 330474 480 0 FreeSans 448 90 0 0 la_oenb[57]
port 479 nsew signal input
flabel metal2 s 333858 -960 333970 480 0 FreeSans 448 90 0 0 la_oenb[58]
port 480 nsew signal input
flabel metal2 s 337446 -960 337558 480 0 FreeSans 448 90 0 0 la_oenb[59]
port 481 nsew signal input
flabel metal2 s 145902 -960 146014 480 0 FreeSans 448 90 0 0 la_oenb[5]
port 482 nsew signal input
flabel metal2 s 340942 -960 341054 480 0 FreeSans 448 90 0 0 la_oenb[60]
port 483 nsew signal input
flabel metal2 s 344530 -960 344642 480 0 FreeSans 448 90 0 0 la_oenb[61]
port 484 nsew signal input
flabel metal2 s 348026 -960 348138 480 0 FreeSans 448 90 0 0 la_oenb[62]
port 485 nsew signal input
flabel metal2 s 351614 -960 351726 480 0 FreeSans 448 90 0 0 la_oenb[63]
port 486 nsew signal input
flabel metal2 s 355202 -960 355314 480 0 FreeSans 448 90 0 0 la_oenb[64]
port 487 nsew signal input
flabel metal2 s 358698 -960 358810 480 0 FreeSans 448 90 0 0 la_oenb[65]
port 488 nsew signal input
flabel metal2 s 362286 -960 362398 480 0 FreeSans 448 90 0 0 la_oenb[66]
port 489 nsew signal input
flabel metal2 s 365782 -960 365894 480 0 FreeSans 448 90 0 0 la_oenb[67]
port 490 nsew signal input
flabel metal2 s 369370 -960 369482 480 0 FreeSans 448 90 0 0 la_oenb[68]
port 491 nsew signal input
flabel metal2 s 372866 -960 372978 480 0 FreeSans 448 90 0 0 la_oenb[69]
port 492 nsew signal input
flabel metal2 s 149490 -960 149602 480 0 FreeSans 448 90 0 0 la_oenb[6]
port 493 nsew signal input
flabel metal2 s 376454 -960 376566 480 0 FreeSans 448 90 0 0 la_oenb[70]
port 494 nsew signal input
flabel metal2 s 379950 -960 380062 480 0 FreeSans 448 90 0 0 la_oenb[71]
port 495 nsew signal input
flabel metal2 s 383538 -960 383650 480 0 FreeSans 448 90 0 0 la_oenb[72]
port 496 nsew signal input
flabel metal2 s 387126 -960 387238 480 0 FreeSans 448 90 0 0 la_oenb[73]
port 497 nsew signal input
flabel metal2 s 390622 -960 390734 480 0 FreeSans 448 90 0 0 la_oenb[74]
port 498 nsew signal input
flabel metal2 s 394210 -960 394322 480 0 FreeSans 448 90 0 0 la_oenb[75]
port 499 nsew signal input
flabel metal2 s 397706 -960 397818 480 0 FreeSans 448 90 0 0 la_oenb[76]
port 500 nsew signal input
flabel metal2 s 401294 -960 401406 480 0 FreeSans 448 90 0 0 la_oenb[77]
port 501 nsew signal input
flabel metal2 s 404790 -960 404902 480 0 FreeSans 448 90 0 0 la_oenb[78]
port 502 nsew signal input
flabel metal2 s 408378 -960 408490 480 0 FreeSans 448 90 0 0 la_oenb[79]
port 503 nsew signal input
flabel metal2 s 152986 -960 153098 480 0 FreeSans 448 90 0 0 la_oenb[7]
port 504 nsew signal input
flabel metal2 s 411874 -960 411986 480 0 FreeSans 448 90 0 0 la_oenb[80]
port 505 nsew signal input
flabel metal2 s 415462 -960 415574 480 0 FreeSans 448 90 0 0 la_oenb[81]
port 506 nsew signal input
flabel metal2 s 418958 -960 419070 480 0 FreeSans 448 90 0 0 la_oenb[82]
port 507 nsew signal input
flabel metal2 s 422546 -960 422658 480 0 FreeSans 448 90 0 0 la_oenb[83]
port 508 nsew signal input
flabel metal2 s 426134 -960 426246 480 0 FreeSans 448 90 0 0 la_oenb[84]
port 509 nsew signal input
flabel metal2 s 429630 -960 429742 480 0 FreeSans 448 90 0 0 la_oenb[85]
port 510 nsew signal input
flabel metal2 s 433218 -960 433330 480 0 FreeSans 448 90 0 0 la_oenb[86]
port 511 nsew signal input
flabel metal2 s 436714 -960 436826 480 0 FreeSans 448 90 0 0 la_oenb[87]
port 512 nsew signal input
flabel metal2 s 440302 -960 440414 480 0 FreeSans 448 90 0 0 la_oenb[88]
port 513 nsew signal input
flabel metal2 s 443798 -960 443910 480 0 FreeSans 448 90 0 0 la_oenb[89]
port 514 nsew signal input
flabel metal2 s 156574 -960 156686 480 0 FreeSans 448 90 0 0 la_oenb[8]
port 515 nsew signal input
flabel metal2 s 447386 -960 447498 480 0 FreeSans 448 90 0 0 la_oenb[90]
port 516 nsew signal input
flabel metal2 s 450882 -960 450994 480 0 FreeSans 448 90 0 0 la_oenb[91]
port 517 nsew signal input
flabel metal2 s 454470 -960 454582 480 0 FreeSans 448 90 0 0 la_oenb[92]
port 518 nsew signal input
flabel metal2 s 458058 -960 458170 480 0 FreeSans 448 90 0 0 la_oenb[93]
port 519 nsew signal input
flabel metal2 s 461554 -960 461666 480 0 FreeSans 448 90 0 0 la_oenb[94]
port 520 nsew signal input
flabel metal2 s 465142 -960 465254 480 0 FreeSans 448 90 0 0 la_oenb[95]
port 521 nsew signal input
flabel metal2 s 468638 -960 468750 480 0 FreeSans 448 90 0 0 la_oenb[96]
port 522 nsew signal input
flabel metal2 s 472226 -960 472338 480 0 FreeSans 448 90 0 0 la_oenb[97]
port 523 nsew signal input
flabel metal2 s 475722 -960 475834 480 0 FreeSans 448 90 0 0 la_oenb[98]
port 524 nsew signal input
flabel metal2 s 479310 -960 479422 480 0 FreeSans 448 90 0 0 la_oenb[99]
port 525 nsew signal input
flabel metal2 s 160070 -960 160182 480 0 FreeSans 448 90 0 0 la_oenb[9]
port 526 nsew signal input
flabel metal2 s 579774 -960 579886 480 0 FreeSans 448 90 0 0 user_clock2
port 527 nsew signal input
flabel metal2 s 580970 -960 581082 480 0 FreeSans 448 90 0 0 user_irq[0]
port 528 nsew signal tristate
flabel metal2 s 582166 -960 582278 480 0 FreeSans 448 90 0 0 user_irq[1]
port 529 nsew signal tristate
flabel metal2 s 583362 -960 583474 480 0 FreeSans 448 90 0 0 user_irq[2]
port 530 nsew signal tristate
flabel metal4 s -2006 -934 -1386 704870 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2006 -934 585930 -314 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2006 704250 585930 704870 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 585310 -934 585930 704870 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 1794 -7654 2414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 37794 -7654 38414 49367 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 37794 674393 38414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 73794 -7654 74414 49367 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 73794 674393 74414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 109794 -7654 110414 49367 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 109794 674393 110414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 145794 -7654 146414 49367 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 145794 674393 146414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 181794 -7654 182414 49367 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 181794 674393 182414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 217794 -7654 218414 49367 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 217794 674393 218414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 253794 -7654 254414 49367 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 253794 674393 254414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 289794 -7654 290414 49367 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 289794 674393 290414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 325794 -7654 326414 49367 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 325794 674393 326414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 361794 -7654 362414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 397794 -7654 398414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 433794 -7654 434414 127767 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 433794 157249 434414 422599 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 433794 442833 434414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 469794 -7654 470414 201919 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 469794 385580 470414 601103 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 469794 669073 470414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 505794 -7654 506414 82599 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 505794 139281 506414 201919 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 505794 259417 506414 601103 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 505794 669073 506414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 541794 -7654 542414 425068 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 541794 460836 542414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 577794 -7654 578414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 2866 592650 3486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 38866 592650 39486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 74866 592650 75486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 110866 592650 111486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 146866 592650 147486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 182866 592650 183486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 218866 592650 219486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 254866 592650 255486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 290866 592650 291486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 326866 592650 327486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 362866 592650 363486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 398866 592650 399486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 434866 592650 435486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 470866 592650 471486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 506866 592650 507486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 542866 592650 543486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 578866 592650 579486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 614866 592650 615486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 650866 592650 651486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 686866 592650 687486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s -3926 -2854 -3306 706790 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -3926 -2854 587850 -2234 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -3926 706170 587850 706790 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 587230 -2854 587850 706790 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 9234 -7654 9854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 45234 -7654 45854 49367 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 45234 674393 45854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 81234 -7654 81854 49367 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 81234 674393 81854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 117234 -7654 117854 49367 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 117234 674393 117854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 153234 -7654 153854 49367 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 153234 674393 153854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 189234 -7654 189854 49367 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 189234 674393 189854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 225234 -7654 225854 49367 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 225234 674393 225854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 261234 -7654 261854 49367 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 261234 674393 261854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 297234 -7654 297854 49367 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 297234 674393 297854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 333234 -7654 333854 49367 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 333234 674393 333854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 369234 -7654 369854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 405234 -7654 405854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 441234 -7654 441854 127767 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 441234 157249 441854 422599 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 441234 442833 441854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 477234 -7654 477854 201919 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 477234 259417 477854 322287 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 477234 385225 477854 601103 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 477234 669073 477854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 513234 -7654 513854 82599 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 513234 139281 513854 201919 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 513234 259417 513854 601103 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 513234 669073 513854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 549234 -7654 549854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 10306 592650 10926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 46306 592650 46926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 82306 592650 82926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 118306 592650 118926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 154306 592650 154926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 190306 592650 190926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 226306 592650 226926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 262306 592650 262926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 298306 592650 298926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 334306 592650 334926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 370306 592650 370926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 406306 592650 406926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 442306 592650 442926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 478306 592650 478926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 514306 592650 514926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 550306 592650 550926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 586306 592650 586926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 622306 592650 622926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 658306 592650 658926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 694306 592650 694926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s -5846 -4774 -5226 708710 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -5846 -4774 589770 -4154 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -5846 708090 589770 708710 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 589150 -4774 589770 708710 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 16674 -7654 17294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 52674 -7654 53294 49367 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 88674 -7654 89294 49367 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 124674 -7654 125294 49367 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 160674 -7654 161294 49367 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 196674 -7654 197294 49367 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 232674 -7654 233294 49367 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 268674 -7654 269294 49367 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 304674 -7654 305294 49367 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 340674 -7654 341294 49367 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 376674 -7654 377294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 412674 -7654 413294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 448674 -7654 449294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 484674 -7654 485294 201919 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 484674 259417 485294 322068 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 484674 385580 485294 500068 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 484674 517884 485294 601103 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 520674 -7654 521294 82599 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 520674 139281 521294 201919 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 520674 259417 521294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 556674 -7654 557294 360068 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 556674 377884 557294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 17746 592650 18366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 53746 592650 54366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 89746 592650 90366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 125746 592650 126366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 161746 592650 162366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 197746 592650 198366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 233746 592650 234366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 269746 592650 270366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 305746 592650 306366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 341746 592650 342366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 377746 592650 378366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 413746 592650 414366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 449746 592650 450366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 485746 592650 486366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 521746 592650 522366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 557746 592650 558366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 593746 592650 594366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 629746 592650 630366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 665746 592650 666366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s -7766 -6694 -7146 710630 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -7766 -6694 591690 -6074 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -7766 710010 591690 710630 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 591070 -6694 591690 710630 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 24114 -7654 24734 45068 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 60114 -7654 60734 49367 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 96114 -7654 96734 49367 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 132114 -7654 132734 49367 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 168114 -7654 168734 49367 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 204114 -7654 204734 49367 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 240114 -7654 240734 49367 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 276114 -7654 276734 49367 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 312114 -7654 312734 49367 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 348114 -7654 348734 49367 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 384114 -7654 384734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 420114 -7654 420734 127767 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 420114 157249 420734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 456114 -7654 456734 500068 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 456114 517884 456734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 492114 -7654 492734 82599 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 492114 259417 492734 322287 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 492114 385225 492734 601103 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 492114 669073 492734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 528114 -7654 528734 82599 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 528114 259417 528734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 564114 -7654 564734 360068 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 564114 377884 564734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 25186 592650 25806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 61186 592650 61806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 97186 592650 97806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 133186 592650 133806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 169186 592650 169806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 205186 592650 205806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 241186 592650 241806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 277186 592650 277806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 313186 592650 313806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 349186 592650 349806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 385186 592650 385806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 421186 592650 421806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 457186 592650 457806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 493186 592650 493806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 529186 592650 529806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 565186 592650 565806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 601186 592650 601806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 637186 592650 637806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 673186 592650 673806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s -6806 -5734 -6186 709670 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -6806 -5734 590730 -5114 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -6806 709050 590730 709670 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 590110 -5734 590730 709670 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 20394 -7654 21014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 56394 -7654 57014 49367 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 92394 -7654 93014 49367 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 128394 -7654 129014 49367 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 164394 -7654 165014 49367 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 200394 -7654 201014 49367 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 236394 -7654 237014 49367 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 272394 -7654 273014 49367 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 308394 -7654 309014 49367 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 344394 -7654 345014 49367 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 380394 -7654 381014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 416394 -7654 417014 127767 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 416394 157249 417014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 452394 -7654 453014 500068 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 452394 517884 453014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 488394 -7654 489014 82599 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 488394 139281 489014 201919 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 488394 259417 489014 322287 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 488394 453692 489014 500068 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 488394 517884 489014 601103 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 488394 669073 489014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 524394 -7654 525014 82599 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 524394 139281 525014 201919 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 524394 259417 525014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 560394 -7654 561014 30068 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 560394 51692 561014 360068 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 560394 377884 561014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 21466 592650 22086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 57466 592650 58086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 93466 592650 94086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 129466 592650 130086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 165466 592650 166086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 201466 592650 202086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 237466 592650 238086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 273466 592650 274086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 309466 592650 310086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 345466 592650 346086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 381466 592650 382086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 417466 592650 418086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 453466 592650 454086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 489466 592650 490086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 525466 592650 526086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 561466 592650 562086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 597466 592650 598086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 633466 592650 634086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 669466 592650 670086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s -8726 -7654 -8106 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 -7654 592650 -7034 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 710970 592650 711590 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 592030 -7654 592650 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 27834 -7654 28454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 63834 -7654 64454 49367 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 63834 674393 64454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 99834 -7654 100454 49367 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 99834 674393 100454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 135834 -7654 136454 49367 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 135834 674393 136454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 171834 -7654 172454 49367 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 171834 674393 172454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 207834 -7654 208454 49367 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 207834 674393 208454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 243834 -7654 244454 49367 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 243834 674393 244454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 279834 -7654 280454 49367 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 279834 674393 280454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 315834 -7654 316454 45068 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 351834 -7654 352454 49367 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 351834 674393 352454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 387834 -7654 388454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 423834 -7654 424454 127767 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 423834 157249 424454 420068 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 423834 444412 424454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 459834 -7654 460454 500068 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 459834 517884 460454 601103 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 459834 669073 460454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 495834 -7654 496454 82599 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 495834 259417 496454 601103 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 495834 669073 496454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 531834 -7654 532454 82599 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 531834 139281 532454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 567834 -7654 568454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 28906 592650 29526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 64906 592650 65526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 100906 592650 101526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 136906 592650 137526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 172906 592650 173526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 208906 592650 209526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 244906 592650 245526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 280906 592650 281526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 316906 592650 317526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 352906 592650 353526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 388906 592650 389526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 424906 592650 425526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 460906 592650 461526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 496906 592650 497526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 532906 592650 533526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 568906 592650 569526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 604906 592650 605526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 640906 592650 641526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 676906 592650 677526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s -2966 -1894 -2346 705830 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -2966 -1894 586890 -1274 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -2966 705210 586890 705830 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 586270 -1894 586890 705830 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 5514 -7654 6134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 41514 -7654 42134 49367 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 41514 674393 42134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 77514 -7654 78134 49367 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 77514 674393 78134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 113514 -7654 114134 49367 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 113514 674393 114134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 149514 -7654 150134 49367 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 149514 674393 150134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 185514 -7654 186134 49367 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 185514 674393 186134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 221514 -7654 222134 49367 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 221514 674393 222134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 257514 -7654 258134 49367 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 257514 674393 258134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 293514 -7654 294134 49367 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 293514 674393 294134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 329514 -7654 330134 49367 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 329514 674393 330134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 365514 -7654 366134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 401514 -7654 402134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 437514 -7654 438134 127767 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 437514 157249 438134 420068 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 437514 444412 438134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 473514 -7654 474134 201919 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 473514 453692 474134 601103 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 473514 669073 474134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 509514 -7654 510134 82599 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 509514 139281 510134 201919 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 509514 259417 510134 601103 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 509514 669073 510134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 545514 -7654 546134 30068 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 545514 51692 546134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 581514 -7654 582134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 6586 592650 7206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 42586 592650 43206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 78586 592650 79206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 114586 592650 115206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 150586 592650 151206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 186586 592650 187206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 222586 592650 223206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 258586 592650 259206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 294586 592650 295206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 330586 592650 331206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 366586 592650 367206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 402586 592650 403206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 438586 592650 439206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 474586 592650 475206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 510586 592650 511206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 546586 592650 547206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 582586 592650 583206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 618586 592650 619206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 654586 592650 655206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 690586 592650 691206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s -4886 -3814 -4266 707750 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -4886 -3814 588810 -3194 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -4886 707130 588810 707750 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 588190 -3814 588810 707750 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 12954 -7654 13574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 48954 -7654 49574 49367 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 48954 674393 49574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 84954 -7654 85574 49367 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 84954 674393 85574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 120954 -7654 121574 49367 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 120954 674393 121574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 156954 -7654 157574 49367 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 156954 674393 157574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 192954 -7654 193574 45068 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 192954 684676 193574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 228954 -7654 229574 49367 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 228954 674393 229574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 264954 -7654 265574 49367 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 264954 674393 265574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 300954 -7654 301574 45068 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 300954 684676 301574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 336954 -7654 337574 49367 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 336954 674393 337574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 372954 -7654 373574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 408954 -7654 409574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 444954 -7654 445574 120068 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 444954 159644 445574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 480954 -7654 481574 201919 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 480954 259417 481574 322287 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 480954 453692 481574 601103 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 480954 669073 481574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 516954 -7654 517574 82599 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 516954 139281 517574 201919 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 516954 259417 517574 601103 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 516954 669073 517574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 552954 -7654 553574 30068 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 552954 51692 553574 360068 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 552954 377884 553574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 14026 592650 14646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 50026 592650 50646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 86026 592650 86646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 122026 592650 122646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 158026 592650 158646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 194026 592650 194646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 230026 592650 230646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 266026 592650 266646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 302026 592650 302646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 338026 592650 338646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 374026 592650 374646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 410026 592650 410646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 446026 592650 446646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 482026 592650 482646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 518026 592650 518646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 554026 592650 554646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 590026 592650 590646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 626026 592650 626646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 662026 592650 662646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 698026 592650 698646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal2 s 542 -960 654 480 0 FreeSans 448 90 0 0 wb_clk_i
port 539 nsew signal input
flabel metal2 s 1646 -960 1758 480 0 FreeSans 448 90 0 0 wb_rst_i
port 540 nsew signal input
flabel metal2 s 2842 -960 2954 480 0 FreeSans 448 90 0 0 wbs_ack_o
port 541 nsew signal tristate
flabel metal2 s 7626 -960 7738 480 0 FreeSans 448 90 0 0 wbs_adr_i[0]
port 542 nsew signal input
flabel metal2 s 47830 -960 47942 480 0 FreeSans 448 90 0 0 wbs_adr_i[10]
port 543 nsew signal input
flabel metal2 s 51326 -960 51438 480 0 FreeSans 448 90 0 0 wbs_adr_i[11]
port 544 nsew signal input
flabel metal2 s 54914 -960 55026 480 0 FreeSans 448 90 0 0 wbs_adr_i[12]
port 545 nsew signal input
flabel metal2 s 58410 -960 58522 480 0 FreeSans 448 90 0 0 wbs_adr_i[13]
port 546 nsew signal input
flabel metal2 s 61998 -960 62110 480 0 FreeSans 448 90 0 0 wbs_adr_i[14]
port 547 nsew signal input
flabel metal2 s 65494 -960 65606 480 0 FreeSans 448 90 0 0 wbs_adr_i[15]
port 548 nsew signal input
flabel metal2 s 69082 -960 69194 480 0 FreeSans 448 90 0 0 wbs_adr_i[16]
port 549 nsew signal input
flabel metal2 s 72578 -960 72690 480 0 FreeSans 448 90 0 0 wbs_adr_i[17]
port 550 nsew signal input
flabel metal2 s 76166 -960 76278 480 0 FreeSans 448 90 0 0 wbs_adr_i[18]
port 551 nsew signal input
flabel metal2 s 79662 -960 79774 480 0 FreeSans 448 90 0 0 wbs_adr_i[19]
port 552 nsew signal input
flabel metal2 s 12318 -960 12430 480 0 FreeSans 448 90 0 0 wbs_adr_i[1]
port 553 nsew signal input
flabel metal2 s 83250 -960 83362 480 0 FreeSans 448 90 0 0 wbs_adr_i[20]
port 554 nsew signal input
flabel metal2 s 86838 -960 86950 480 0 FreeSans 448 90 0 0 wbs_adr_i[21]
port 555 nsew signal input
flabel metal2 s 90334 -960 90446 480 0 FreeSans 448 90 0 0 wbs_adr_i[22]
port 556 nsew signal input
flabel metal2 s 93922 -960 94034 480 0 FreeSans 448 90 0 0 wbs_adr_i[23]
port 557 nsew signal input
flabel metal2 s 97418 -960 97530 480 0 FreeSans 448 90 0 0 wbs_adr_i[24]
port 558 nsew signal input
flabel metal2 s 101006 -960 101118 480 0 FreeSans 448 90 0 0 wbs_adr_i[25]
port 559 nsew signal input
flabel metal2 s 104502 -960 104614 480 0 FreeSans 448 90 0 0 wbs_adr_i[26]
port 560 nsew signal input
flabel metal2 s 108090 -960 108202 480 0 FreeSans 448 90 0 0 wbs_adr_i[27]
port 561 nsew signal input
flabel metal2 s 111586 -960 111698 480 0 FreeSans 448 90 0 0 wbs_adr_i[28]
port 562 nsew signal input
flabel metal2 s 115174 -960 115286 480 0 FreeSans 448 90 0 0 wbs_adr_i[29]
port 563 nsew signal input
flabel metal2 s 17010 -960 17122 480 0 FreeSans 448 90 0 0 wbs_adr_i[2]
port 564 nsew signal input
flabel metal2 s 118762 -960 118874 480 0 FreeSans 448 90 0 0 wbs_adr_i[30]
port 565 nsew signal input
flabel metal2 s 122258 -960 122370 480 0 FreeSans 448 90 0 0 wbs_adr_i[31]
port 566 nsew signal input
flabel metal2 s 21794 -960 21906 480 0 FreeSans 448 90 0 0 wbs_adr_i[3]
port 567 nsew signal input
flabel metal2 s 26486 -960 26598 480 0 FreeSans 448 90 0 0 wbs_adr_i[4]
port 568 nsew signal input
flabel metal2 s 30074 -960 30186 480 0 FreeSans 448 90 0 0 wbs_adr_i[5]
port 569 nsew signal input
flabel metal2 s 33570 -960 33682 480 0 FreeSans 448 90 0 0 wbs_adr_i[6]
port 570 nsew signal input
flabel metal2 s 37158 -960 37270 480 0 FreeSans 448 90 0 0 wbs_adr_i[7]
port 571 nsew signal input
flabel metal2 s 40654 -960 40766 480 0 FreeSans 448 90 0 0 wbs_adr_i[8]
port 572 nsew signal input
flabel metal2 s 44242 -960 44354 480 0 FreeSans 448 90 0 0 wbs_adr_i[9]
port 573 nsew signal input
flabel metal2 s 4038 -960 4150 480 0 FreeSans 448 90 0 0 wbs_cyc_i
port 574 nsew signal input
flabel metal2 s 8730 -960 8842 480 0 FreeSans 448 90 0 0 wbs_dat_i[0]
port 575 nsew signal input
flabel metal2 s 48934 -960 49046 480 0 FreeSans 448 90 0 0 wbs_dat_i[10]
port 576 nsew signal input
flabel metal2 s 52522 -960 52634 480 0 FreeSans 448 90 0 0 wbs_dat_i[11]
port 577 nsew signal input
flabel metal2 s 56018 -960 56130 480 0 FreeSans 448 90 0 0 wbs_dat_i[12]
port 578 nsew signal input
flabel metal2 s 59606 -960 59718 480 0 FreeSans 448 90 0 0 wbs_dat_i[13]
port 579 nsew signal input
flabel metal2 s 63194 -960 63306 480 0 FreeSans 448 90 0 0 wbs_dat_i[14]
port 580 nsew signal input
flabel metal2 s 66690 -960 66802 480 0 FreeSans 448 90 0 0 wbs_dat_i[15]
port 581 nsew signal input
flabel metal2 s 70278 -960 70390 480 0 FreeSans 448 90 0 0 wbs_dat_i[16]
port 582 nsew signal input
flabel metal2 s 73774 -960 73886 480 0 FreeSans 448 90 0 0 wbs_dat_i[17]
port 583 nsew signal input
flabel metal2 s 77362 -960 77474 480 0 FreeSans 448 90 0 0 wbs_dat_i[18]
port 584 nsew signal input
flabel metal2 s 80858 -960 80970 480 0 FreeSans 448 90 0 0 wbs_dat_i[19]
port 585 nsew signal input
flabel metal2 s 13514 -960 13626 480 0 FreeSans 448 90 0 0 wbs_dat_i[1]
port 586 nsew signal input
flabel metal2 s 84446 -960 84558 480 0 FreeSans 448 90 0 0 wbs_dat_i[20]
port 587 nsew signal input
flabel metal2 s 87942 -960 88054 480 0 FreeSans 448 90 0 0 wbs_dat_i[21]
port 588 nsew signal input
flabel metal2 s 91530 -960 91642 480 0 FreeSans 448 90 0 0 wbs_dat_i[22]
port 589 nsew signal input
flabel metal2 s 95118 -960 95230 480 0 FreeSans 448 90 0 0 wbs_dat_i[23]
port 590 nsew signal input
flabel metal2 s 98614 -960 98726 480 0 FreeSans 448 90 0 0 wbs_dat_i[24]
port 591 nsew signal input
flabel metal2 s 102202 -960 102314 480 0 FreeSans 448 90 0 0 wbs_dat_i[25]
port 592 nsew signal input
flabel metal2 s 105698 -960 105810 480 0 FreeSans 448 90 0 0 wbs_dat_i[26]
port 593 nsew signal input
flabel metal2 s 109286 -960 109398 480 0 FreeSans 448 90 0 0 wbs_dat_i[27]
port 594 nsew signal input
flabel metal2 s 112782 -960 112894 480 0 FreeSans 448 90 0 0 wbs_dat_i[28]
port 595 nsew signal input
flabel metal2 s 116370 -960 116482 480 0 FreeSans 448 90 0 0 wbs_dat_i[29]
port 596 nsew signal input
flabel metal2 s 18206 -960 18318 480 0 FreeSans 448 90 0 0 wbs_dat_i[2]
port 597 nsew signal input
flabel metal2 s 119866 -960 119978 480 0 FreeSans 448 90 0 0 wbs_dat_i[30]
port 598 nsew signal input
flabel metal2 s 123454 -960 123566 480 0 FreeSans 448 90 0 0 wbs_dat_i[31]
port 599 nsew signal input
flabel metal2 s 22990 -960 23102 480 0 FreeSans 448 90 0 0 wbs_dat_i[3]
port 600 nsew signal input
flabel metal2 s 27682 -960 27794 480 0 FreeSans 448 90 0 0 wbs_dat_i[4]
port 601 nsew signal input
flabel metal2 s 31270 -960 31382 480 0 FreeSans 448 90 0 0 wbs_dat_i[5]
port 602 nsew signal input
flabel metal2 s 34766 -960 34878 480 0 FreeSans 448 90 0 0 wbs_dat_i[6]
port 603 nsew signal input
flabel metal2 s 38354 -960 38466 480 0 FreeSans 448 90 0 0 wbs_dat_i[7]
port 604 nsew signal input
flabel metal2 s 41850 -960 41962 480 0 FreeSans 448 90 0 0 wbs_dat_i[8]
port 605 nsew signal input
flabel metal2 s 45438 -960 45550 480 0 FreeSans 448 90 0 0 wbs_dat_i[9]
port 606 nsew signal input
flabel metal2 s 9926 -960 10038 480 0 FreeSans 448 90 0 0 wbs_dat_o[0]
port 607 nsew signal tristate
flabel metal2 s 50130 -960 50242 480 0 FreeSans 448 90 0 0 wbs_dat_o[10]
port 608 nsew signal tristate
flabel metal2 s 53718 -960 53830 480 0 FreeSans 448 90 0 0 wbs_dat_o[11]
port 609 nsew signal tristate
flabel metal2 s 57214 -960 57326 480 0 FreeSans 448 90 0 0 wbs_dat_o[12]
port 610 nsew signal tristate
flabel metal2 s 60802 -960 60914 480 0 FreeSans 448 90 0 0 wbs_dat_o[13]
port 611 nsew signal tristate
flabel metal2 s 64298 -960 64410 480 0 FreeSans 448 90 0 0 wbs_dat_o[14]
port 612 nsew signal tristate
flabel metal2 s 67886 -960 67998 480 0 FreeSans 448 90 0 0 wbs_dat_o[15]
port 613 nsew signal tristate
flabel metal2 s 71474 -960 71586 480 0 FreeSans 448 90 0 0 wbs_dat_o[16]
port 614 nsew signal tristate
flabel metal2 s 74970 -960 75082 480 0 FreeSans 448 90 0 0 wbs_dat_o[17]
port 615 nsew signal tristate
flabel metal2 s 78558 -960 78670 480 0 FreeSans 448 90 0 0 wbs_dat_o[18]
port 616 nsew signal tristate
flabel metal2 s 82054 -960 82166 480 0 FreeSans 448 90 0 0 wbs_dat_o[19]
port 617 nsew signal tristate
flabel metal2 s 14710 -960 14822 480 0 FreeSans 448 90 0 0 wbs_dat_o[1]
port 618 nsew signal tristate
flabel metal2 s 85642 -960 85754 480 0 FreeSans 448 90 0 0 wbs_dat_o[20]
port 619 nsew signal tristate
flabel metal2 s 89138 -960 89250 480 0 FreeSans 448 90 0 0 wbs_dat_o[21]
port 620 nsew signal tristate
flabel metal2 s 92726 -960 92838 480 0 FreeSans 448 90 0 0 wbs_dat_o[22]
port 621 nsew signal tristate
flabel metal2 s 96222 -960 96334 480 0 FreeSans 448 90 0 0 wbs_dat_o[23]
port 622 nsew signal tristate
flabel metal2 s 99810 -960 99922 480 0 FreeSans 448 90 0 0 wbs_dat_o[24]
port 623 nsew signal tristate
flabel metal2 s 103306 -960 103418 480 0 FreeSans 448 90 0 0 wbs_dat_o[25]
port 624 nsew signal tristate
flabel metal2 s 106894 -960 107006 480 0 FreeSans 448 90 0 0 wbs_dat_o[26]
port 625 nsew signal tristate
flabel metal2 s 110482 -960 110594 480 0 FreeSans 448 90 0 0 wbs_dat_o[27]
port 626 nsew signal tristate
flabel metal2 s 113978 -960 114090 480 0 FreeSans 448 90 0 0 wbs_dat_o[28]
port 627 nsew signal tristate
flabel metal2 s 117566 -960 117678 480 0 FreeSans 448 90 0 0 wbs_dat_o[29]
port 628 nsew signal tristate
flabel metal2 s 19402 -960 19514 480 0 FreeSans 448 90 0 0 wbs_dat_o[2]
port 629 nsew signal tristate
flabel metal2 s 121062 -960 121174 480 0 FreeSans 448 90 0 0 wbs_dat_o[30]
port 630 nsew signal tristate
flabel metal2 s 124650 -960 124762 480 0 FreeSans 448 90 0 0 wbs_dat_o[31]
port 631 nsew signal tristate
flabel metal2 s 24186 -960 24298 480 0 FreeSans 448 90 0 0 wbs_dat_o[3]
port 632 nsew signal tristate
flabel metal2 s 28878 -960 28990 480 0 FreeSans 448 90 0 0 wbs_dat_o[4]
port 633 nsew signal tristate
flabel metal2 s 32374 -960 32486 480 0 FreeSans 448 90 0 0 wbs_dat_o[5]
port 634 nsew signal tristate
flabel metal2 s 35962 -960 36074 480 0 FreeSans 448 90 0 0 wbs_dat_o[6]
port 635 nsew signal tristate
flabel metal2 s 39550 -960 39662 480 0 FreeSans 448 90 0 0 wbs_dat_o[7]
port 636 nsew signal tristate
flabel metal2 s 43046 -960 43158 480 0 FreeSans 448 90 0 0 wbs_dat_o[8]
port 637 nsew signal tristate
flabel metal2 s 46634 -960 46746 480 0 FreeSans 448 90 0 0 wbs_dat_o[9]
port 638 nsew signal tristate
flabel metal2 s 11122 -960 11234 480 0 FreeSans 448 90 0 0 wbs_sel_i[0]
port 639 nsew signal input
flabel metal2 s 15906 -960 16018 480 0 FreeSans 448 90 0 0 wbs_sel_i[1]
port 640 nsew signal input
flabel metal2 s 20598 -960 20710 480 0 FreeSans 448 90 0 0 wbs_sel_i[2]
port 641 nsew signal input
flabel metal2 s 25290 -960 25402 480 0 FreeSans 448 90 0 0 wbs_sel_i[3]
port 642 nsew signal input
flabel metal2 s 5234 -960 5346 480 0 FreeSans 448 90 0 0 wbs_stb_i
port 643 nsew signal input
flabel metal2 s 6430 -960 6542 480 0 FreeSans 448 90 0 0 wbs_we_i
port 644 nsew signal input
rlabel via4 331568 651336 331568 651336 0 vccd1
rlabel via4 333704 46776 333704 46776 0 vccd2
rlabel via4 521144 666216 521144 666216 0 vdda1
rlabel via4 528584 637656 528584 637656 0 vdda2
rlabel via4 20864 669936 20864 669936 0 vssa1
rlabel via4 352304 677376 352304 677376 0 vssa2
rlabel via4 346928 655056 346928 655056 0 vssd1
rlabel via4 481424 122496 481424 122496 0 vssd2
rlabel metal2 422510 446172 422510 446172 0 design_clk
rlabel metal2 411624 159868 411624 159868 0 dsi_all\[0\]
rlabel metal2 448362 161058 448362 161058 0 dsi_all\[10\]
rlabel metal2 447626 172142 447626 172142 0 dsi_all\[11\]
rlabel metal3 449106 332588 449106 332588 0 dsi_all\[12\]
rlabel metal2 447166 332945 447166 332945 0 dsi_all\[13\]
rlabel metal2 447258 333319 447258 333319 0 dsi_all\[14\]
rlabel metal2 447166 334305 447166 334305 0 dsi_all\[15\]
rlabel metal1 445464 334050 445464 334050 0 dsi_all\[16\]
rlabel metal1 445464 335682 445464 335682 0 dsi_all\[17\]
rlabel metal2 447442 336005 447442 336005 0 dsi_all\[18\]
rlabel metal2 447166 336821 447166 336821 0 dsi_all\[19\]
rlabel metal3 449934 503472 449934 503472 0 dsi_all\[1\]
rlabel metal3 448830 338028 448830 338028 0 dsi_all\[20\]
rlabel metal2 447166 338453 447166 338453 0 dsi_all\[21\]
rlabel metal2 447258 338759 447258 338759 0 dsi_all\[22\]
rlabel metal2 431250 322252 431250 322252 0 dsi_all\[23\]
rlabel metal2 371910 327726 371910 327726 0 dsi_all\[24\]
rlabel metal2 444222 338504 444222 338504 0 dsi_all\[25\]
rlabel metal2 447166 341513 447166 341513 0 dsi_all\[26\]
rlabel metal3 449842 342788 449842 342788 0 dsi_all\[27\]
rlabel metal3 450156 505531 450156 505531 0 dsi_all\[2\]
rlabel metal3 450087 326604 450087 326604 0 dsi_all\[3\]
rlabel metal2 425208 159868 425208 159868 0 dsi_all\[4\]
rlabel metal2 428184 159596 428184 159596 0 dsi_all\[5\]
rlabel metal2 431496 159324 431496 159324 0 dsi_all\[6\]
rlabel metal3 450156 329037 450156 329037 0 dsi_all\[7\]
rlabel metal3 448646 329868 448646 329868 0 dsi_all\[8\]
rlabel metal3 449060 330548 449060 330548 0 dsi_all\[9\]
rlabel metal2 488849 322116 488849 322116 0 dso_6502\[0\]
rlabel via2 452594 135133 452594 135133 0 dso_6502\[10\]
rlabel via2 452594 136493 452594 136493 0 dso_6502\[11\]
rlabel via2 452594 137853 452594 137853 0 dso_6502\[12\]
rlabel metal2 451582 139281 451582 139281 0 dso_6502\[13\]
rlabel metal2 452594 140607 452594 140607 0 dso_6502\[14\]
rlabel via2 452594 141933 452594 141933 0 dso_6502\[15\]
rlabel metal1 475410 271150 475410 271150 0 dso_6502\[16\]
rlabel via2 452594 144653 452594 144653 0 dso_6502\[17\]
rlabel metal2 452594 146081 452594 146081 0 dso_6502\[18\]
rlabel metal1 476008 275298 476008 275298 0 dso_6502\[19\]
rlabel metal2 451950 123063 451950 123063 0 dso_6502\[1\]
rlabel metal1 474674 311202 474674 311202 0 dso_6502\[20\]
rlabel metal1 474904 276658 474904 276658 0 dso_6502\[21\]
rlabel metal1 473432 309774 473432 309774 0 dso_6502\[22\]
rlabel metal3 451068 152796 451068 152796 0 dso_6502\[23\]
rlabel metal3 451114 154156 451114 154156 0 dso_6502\[24\]
rlabel metal2 452594 155601 452594 155601 0 dso_6502\[25\]
rlabel metal3 450884 156876 450884 156876 0 dso_6502\[26\]
rlabel metal2 489249 322116 489249 322116 0 dso_6502\[2\]
rlabel metal2 489525 322116 489525 322116 0 dso_6502\[3\]
rlabel metal2 489801 322116 489801 322116 0 dso_6502\[4\]
rlabel metal1 471132 272510 471132 272510 0 dso_6502\[5\]
rlabel metal1 471316 268430 471316 268430 0 dso_6502\[6\]
rlabel via2 452594 131053 452594 131053 0 dso_6502\[7\]
rlabel metal1 472052 307122 472052 307122 0 dso_6502\[8\]
rlabel via2 452594 133773 452594 133773 0 dso_6502\[9\]
rlabel metal2 503785 385900 503785 385900 0 dso_LCD\[0\]
rlabel metal2 504337 385900 504337 385900 0 dso_LCD\[1\]
rlabel metal2 505310 388576 505310 388576 0 dso_LCD\[2\]
rlabel metal2 505809 385900 505809 385900 0 dso_LCD\[3\]
rlabel metal2 506683 385900 506683 385900 0 dso_LCD\[4\]
rlabel metal2 507327 385900 507327 385900 0 dso_LCD\[5\]
rlabel metal2 508063 385900 508063 385900 0 dso_LCD\[6\]
rlabel metal2 508753 385900 508753 385900 0 dso_LCD\[7\]
rlabel via2 539603 82756 539603 82756 0 dso_as1802\[0\]
rlabel metal3 540630 102748 540630 102748 0 dso_as1802\[10\]
rlabel metal3 540078 104788 540078 104788 0 dso_as1802\[11\]
rlabel metal3 540676 106828 540676 106828 0 dso_as1802\[12\]
rlabel metal2 499889 322116 499889 322116 0 dso_as1802\[13\]
rlabel metal2 500158 301201 500158 301201 0 dso_as1802\[14\]
rlabel via2 539787 113220 539787 113220 0 dso_as1802\[15\]
rlabel metal3 540124 114988 540124 114988 0 dso_as1802\[16\]
rlabel metal3 540722 117028 540722 117028 0 dso_as1802\[17\]
rlabel via2 539925 119612 539925 119612 0 dso_as1802\[18\]
rlabel metal3 540538 121108 540538 121108 0 dso_as1802\[19\]
rlabel via2 539741 84932 539741 84932 0 dso_as1802\[1\]
rlabel metal1 540960 138550 540960 138550 0 dso_as1802\[20\]
rlabel metal2 502090 314291 502090 314291 0 dso_as1802\[21\]
rlabel metal2 502274 300077 502274 300077 0 dso_as1802\[22\]
rlabel metal2 502550 319474 502550 319474 0 dso_as1802\[23\]
rlabel metal2 502826 320698 502826 320698 0 dso_as1802\[24\]
rlabel metal3 541596 133348 541596 133348 0 dso_as1802\[25\]
rlabel via2 539373 135660 539373 135660 0 dso_as1802\[26\]
rlabel metal3 540492 86428 540492 86428 0 dso_as1802\[2\]
rlabel metal3 541343 88468 541343 88468 0 dso_as1802\[3\]
rlabel metal3 541642 90508 541642 90508 0 dso_as1802\[4\]
rlabel metal3 541228 92548 541228 92548 0 dso_as1802\[5\]
rlabel metal3 541412 94588 541412 94588 0 dso_as1802\[6\]
rlabel metal3 541366 96628 541366 96628 0 dso_as1802\[7\]
rlabel metal3 539948 98955 539948 98955 0 dso_as1802\[8\]
rlabel metal3 541458 100708 541458 100708 0 dso_as1802\[9\]
rlabel metal2 463121 385900 463121 385900 0 dso_as2650\[0\]
rlabel metal2 470665 385900 470665 385900 0 dso_as2650\[10\]
rlabel metal2 471217 385900 471217 385900 0 dso_as2650\[11\]
rlabel metal1 458850 604044 458850 604044 0 dso_as2650\[12\]
rlabel metal2 458988 603908 458988 603908 0 dso_as2650\[13\]
rlabel metal2 461610 493782 461610 493782 0 dso_as2650\[14\]
rlabel metal3 459609 637908 459609 637908 0 dso_as2650\[15\]
rlabel metal2 462990 494462 462990 494462 0 dso_as2650\[16\]
rlabel metal2 468510 494326 468510 494326 0 dso_as2650\[17\]
rlabel metal2 464370 494292 464370 494292 0 dso_as2650\[18\]
rlabel metal2 477105 385900 477105 385900 0 dso_as2650\[19\]
rlabel metal2 463903 385900 463903 385900 0 dso_as2650\[1\]
rlabel metal2 468602 492218 468602 492218 0 dso_as2650\[20\]
rlabel metal2 467130 491504 467130 491504 0 dso_as2650\[21\]
rlabel metal3 459617 655724 459617 655724 0 dso_as2650\[22\]
rlabel metal2 480286 387250 480286 387250 0 dso_as2650\[23\]
rlabel metal2 481022 387216 481022 387216 0 dso_as2650\[24\]
rlabel metal2 481758 387284 481758 387284 0 dso_as2650\[25\]
rlabel metal2 482494 387182 482494 387182 0 dso_as2650\[26\]
rlabel metal2 464593 385900 464593 385900 0 dso_as2650\[2\]
rlabel metal2 465375 385900 465375 385900 0 dso_as2650\[3\]
rlabel metal2 466111 385900 466111 385900 0 dso_as2650\[4\]
rlabel metal2 466801 385900 466801 385900 0 dso_as2650\[5\]
rlabel metal2 467583 385900 467583 385900 0 dso_as2650\[6\]
rlabel metal2 468273 385900 468273 385900 0 dso_as2650\[7\]
rlabel metal2 469246 492786 469246 492786 0 dso_as2650\[8\]
rlabel metal2 469745 385900 469745 385900 0 dso_as2650\[9\]
rlabel metal2 409906 367778 409906 367778 0 dso_as512512512\[0\]
rlabel metal2 447258 371909 447258 371909 0 dso_as512512512\[10\]
rlabel metal2 447166 372283 447166 372283 0 dso_as512512512\[11\]
rlabel metal2 447258 373303 447258 373303 0 dso_as512512512\[12\]
rlabel metal2 447166 373677 447166 373677 0 dso_as512512512\[13\]
rlabel metal2 407790 449854 407790 449854 0 dso_as512512512\[14\]
rlabel metal2 406410 455396 406410 455396 0 dso_as512512512\[15\]
rlabel metal2 447258 376023 447258 376023 0 dso_as512512512\[16\]
rlabel metal2 403650 467126 403650 467126 0 dso_as512512512\[17\]
rlabel metal2 447258 377451 447258 377451 0 dso_as512512512\[18\]
rlabel metal2 368046 478856 368046 478856 0 dso_as512512512\[19\]
rlabel metal1 445556 365602 445556 365602 0 dso_as512512512\[1\]
rlabel metal2 447350 378811 447350 378811 0 dso_as512512512\[20\]
rlabel metal2 370530 490552 370530 490552 0 dso_as512512512\[21\]
rlabel metal2 447442 380171 447442 380171 0 dso_as512512512\[22\]
rlabel metal2 371910 502282 371910 502282 0 dso_as512512512\[23\]
rlabel metal2 447258 380783 447258 380783 0 dso_as512512512\[24\]
rlabel metal2 447258 381871 447258 381871 0 dso_as512512512\[25\]
rlabel metal2 447166 382177 447166 382177 0 dso_as512512512\[26\]
rlabel metal2 447258 383231 447258 383231 0 dso_as512512512\[27\]
rlabel metal1 445510 366962 445510 366962 0 dso_as512512512\[2\]
rlabel metal2 447166 366809 447166 366809 0 dso_as512512512\[3\]
rlabel metal1 445464 368390 445464 368390 0 dso_as512512512\[4\]
rlabel metal2 447166 368203 447166 368203 0 dso_as512512512\[5\]
rlabel metal2 447258 369189 447258 369189 0 dso_as512512512\[6\]
rlabel metal2 447166 369563 447166 369563 0 dso_as512512512\[7\]
rlabel metal2 447258 370549 447258 370549 0 dso_as512512512\[8\]
rlabel metal2 447166 370923 447166 370923 0 dso_as512512512\[9\]
rlabel metal2 483421 385900 483421 385900 0 dso_as5401\[0\]
rlabel metal2 490590 387862 490590 387862 0 dso_as5401\[10\]
rlabel metal2 491471 385900 491471 385900 0 dso_as5401\[11\]
rlabel metal2 492253 385900 492253 385900 0 dso_as5401\[12\]
rlabel metal2 492989 385900 492989 385900 0 dso_as5401\[13\]
rlabel metal2 539067 425068 539067 425068 0 dso_as5401\[14\]
rlabel metal2 540355 425068 540355 425068 0 dso_as5401\[15\]
rlabel metal2 541834 422630 541834 422630 0 dso_as5401\[16\]
rlabel metal2 542931 425068 542931 425068 0 dso_as5401\[17\]
rlabel metal2 544219 425068 544219 425068 0 dso_as5401\[18\]
rlabel metal2 545698 424092 545698 424092 0 dso_as5401\[19\]
rlabel metal2 483966 387386 483966 387386 0 dso_as5401\[1\]
rlabel metal2 546795 425068 546795 425068 0 dso_as5401\[20\]
rlabel metal2 498877 385900 498877 385900 0 dso_as5401\[21\]
rlabel metal2 522330 406096 522330 406096 0 dso_as5401\[22\]
rlabel metal2 500349 385900 500349 385900 0 dso_as5401\[23\]
rlabel metal2 500894 387352 500894 387352 0 dso_as5401\[24\]
rlabel metal2 501821 385900 501821 385900 0 dso_as5401\[25\]
rlabel metal2 502366 387454 502366 387454 0 dso_as5401\[26\]
rlabel metal2 484702 387284 484702 387284 0 dso_as5401\[2\]
rlabel metal2 485438 387250 485438 387250 0 dso_as5401\[3\]
rlabel metal2 486319 385900 486319 385900 0 dso_as5401\[4\]
rlabel metal2 486910 389607 486910 389607 0 dso_as5401\[5\]
rlabel metal2 487837 385900 487837 385900 0 dso_as5401\[6\]
rlabel metal2 488382 387216 488382 387216 0 dso_as5401\[7\]
rlabel metal2 489309 385900 489309 385900 0 dso_as5401\[8\]
rlabel metal2 489854 387182 489854 387182 0 dso_as5401\[9\]
rlabel metal2 522330 369036 522330 369036 0 dso_counter\[0\]
rlabel metal2 565294 360009 565294 360009 0 dso_counter\[10\]
rlabel via1 566766 360077 566766 360077 0 dso_counter\[11\]
rlabel metal2 547262 369206 547262 369206 0 dso_counter\[1\]
rlabel metal3 511282 379780 511282 379780 0 dso_counter\[2\]
rlabel metal3 511650 380324 511650 380324 0 dso_counter\[3\]
rlabel metal3 511604 380868 511604 380868 0 dso_counter\[4\]
rlabel metal2 547170 370396 547170 370396 0 dso_counter\[5\]
rlabel metal2 544410 367268 544410 367268 0 dso_counter\[6\]
rlabel metal2 561154 359254 561154 359254 0 dso_counter\[7\]
rlabel metal2 562626 359322 562626 359322 0 dso_counter\[8\]
rlabel metal2 519754 370804 519754 370804 0 dso_counter\[9\]
rlabel metal2 456734 387522 456734 387522 0 dso_diceroll\[0\]
rlabel metal2 457661 385900 457661 385900 0 dso_diceroll\[1\]
rlabel metal2 458351 385900 458351 385900 0 dso_diceroll\[2\]
rlabel metal2 459133 385900 459133 385900 0 dso_diceroll\[3\]
rlabel metal1 481620 429182 481620 429182 0 dso_diceroll\[4\]
rlabel metal1 484334 429182 484334 429182 0 dso_diceroll\[5\]
rlabel metal2 461150 387352 461150 387352 0 dso_diceroll\[6\]
rlabel metal2 461886 386876 461886 386876 0 dso_diceroll\[7\]
rlabel metal3 449106 352308 449106 352308 0 dso_mc14500\[0\]
rlabel metal3 449014 352988 449014 352988 0 dso_mc14500\[1\]
rlabel metal3 448922 353668 448922 353668 0 dso_mc14500\[2\]
rlabel metal3 448968 354348 448968 354348 0 dso_mc14500\[3\]
rlabel metal2 485224 500140 485224 500140 0 dso_mc14500\[4\]
rlabel metal2 486420 500140 486420 500140 0 dso_mc14500\[5\]
rlabel metal2 487478 500140 487478 500140 0 dso_mc14500\[6\]
rlabel metal2 489102 500140 489102 500140 0 dso_mc14500\[7\]
rlabel metal3 449888 357748 449888 357748 0 dso_mc14500\[8\]
rlabel metal2 450701 500140 450701 500140 0 dso_multiplier\[0\]
rlabel metal2 451773 385900 451773 385900 0 dso_multiplier\[1\]
rlabel metal2 452463 385900 452463 385900 0 dso_multiplier\[2\]
rlabel metal2 453054 387522 453054 387522 0 dso_multiplier\[3\]
rlabel metal2 453889 385900 453889 385900 0 dso_multiplier\[4\]
rlabel metal2 454717 385900 454717 385900 0 dso_multiplier\[5\]
rlabel metal2 455262 389607 455262 389607 0 dso_multiplier\[6\]
rlabel metal2 461058 498552 461058 498552 0 dso_multiplier\[7\]
rlabel metal2 487469 322116 487469 322116 0 dso_posit\[0\]
rlabel metal1 508898 309842 508898 309842 0 dso_posit\[1\]
rlabel metal1 509864 287674 509864 287674 0 dso_posit\[2\]
rlabel metal2 488145 322116 488145 322116 0 dso_posit\[3\]
rlabel metal1 445556 358870 445556 358870 0 dso_tbb1143\[0\]
rlabel metal2 447166 359295 447166 359295 0 dso_tbb1143\[1\]
rlabel metal2 447166 360349 447166 360349 0 dso_tbb1143\[2\]
rlabel metal2 447258 360723 447258 360723 0 dso_tbb1143\[3\]
rlabel metal1 444774 361658 444774 361658 0 dso_tbb1143\[4\]
rlabel metal2 447166 362049 447166 362049 0 dso_tbb1143\[5\]
rlabel metal2 447166 363069 447166 363069 0 dso_tbb1143\[6\]
rlabel metal2 447258 363443 447258 363443 0 dso_tbb1143\[7\]
rlabel metal2 504489 322116 504489 322116 0 dso_tune
rlabel metal2 580198 6715 580198 6715 0 io_in[0]
rlabel metal2 580198 457453 580198 457453 0 io_in[10]
rlabel metal2 580198 510969 580198 510969 0 io_in[11]
rlabel metal2 580198 563703 580198 563703 0 io_in[12]
rlabel metal2 579646 617185 579646 617185 0 io_in[13]
rlabel metal3 581954 670684 581954 670684 0 io_in[14]
rlabel metal3 558923 699788 558923 699788 0 io_in[15]
rlabel metal3 446085 422348 446085 422348 0 io_in[16]
rlabel metal2 429870 702110 429870 702110 0 io_in[17]
rlabel metal2 365010 526704 365010 526704 0 io_in[18]
rlabel metal4 444268 510816 444268 510816 0 io_in[19]
rlabel metal2 566490 180404 566490 180404 0 io_in[1]
rlabel metal2 235198 702178 235198 702178 0 io_in[20]
rlabel metal2 446430 510952 446430 510952 0 io_in[21]
rlabel metal3 443877 421940 443877 421940 0 io_in[22]
rlabel metal2 40526 701974 40526 701974 0 io_in[23]
rlabel metal4 447764 502724 447764 502724 0 io_in[24]
rlabel metal3 1970 632060 1970 632060 0 io_in[25]
rlabel metal3 1786 579972 1786 579972 0 io_in[26]
rlabel metal3 2154 527884 2154 527884 0 io_in[27]
rlabel metal3 2016 475660 2016 475660 0 io_in[28]
rlabel metal3 1970 423572 1970 423572 0 io_in[29]
rlabel metal2 580198 86547 580198 86547 0 io_in[2]
rlabel metal3 2108 371348 2108 371348 0 io_in[30]
rlabel metal1 4554 253946 4554 253946 0 io_in[31]
rlabel metal3 1924 267172 1924 267172 0 io_in[32]
rlabel metal3 2108 214948 2108 214948 0 io_in[33]
rlabel metal3 1832 162860 1832 162860 0 io_in[34]
rlabel metal3 1855 110636 1855 110636 0 io_in[35]
rlabel metal3 1970 71604 1970 71604 0 io_in[36]
rlabel metal3 1602 32436 1602 32436 0 io_in[37]
rlabel metal2 580198 126463 580198 126463 0 io_in[3]
rlabel metal2 580198 166413 580198 166413 0 io_in[4]
rlabel metal2 579830 206329 579830 206329 0 io_in[5]
rlabel via2 580198 245565 580198 245565 0 io_in[6]
rlabel metal2 461610 307734 461610 307734 0 io_in[7]
rlabel metal3 582184 351900 582184 351900 0 io_in[8]
rlabel metal2 580198 404651 580198 404651 0 io_in[9]
rlabel via2 580198 33099 580198 33099 0 io_oeb[0]
rlabel metal2 580198 484517 580198 484517 0 io_oeb[10]
rlabel metal2 519570 428366 519570 428366 0 io_oeb[11]
rlabel metal2 580198 590835 580198 590835 0 io_oeb[12]
rlabel metal3 582046 644028 582046 644028 0 io_oeb[13]
rlabel metal3 581908 697204 581908 697204 0 io_oeb[14]
rlabel metal3 523457 502316 523457 502316 0 io_oeb[15]
rlabel metal2 462346 687065 462346 687065 0 io_oeb[16]
rlabel metal2 447718 329120 447718 329120 0 io_oeb[17]
rlabel metal2 332534 694460 332534 694460 0 io_oeb[18]
rlabel metal2 445142 510918 445142 510918 0 io_oeb[19]
rlabel metal2 544410 189652 544410 189652 0 io_oeb[1]
rlabel metal2 445326 502282 445326 502282 0 io_oeb[20]
rlabel metal2 137862 702042 137862 702042 0 io_oeb[21]
rlabel metal2 449374 502333 449374 502333 0 io_oeb[22]
rlabel metal2 445050 510782 445050 510782 0 io_oeb[23]
rlabel metal3 1740 658172 1740 658172 0 io_oeb[24]
rlabel metal3 1855 606084 1855 606084 0 io_oeb[25]
rlabel metal3 2200 553860 2200 553860 0 io_oeb[26]
rlabel metal3 2062 501772 2062 501772 0 io_oeb[27]
rlabel metal3 1878 449548 1878 449548 0 io_oeb[28]
rlabel metal1 366942 140794 366942 140794 0 io_oeb[29]
rlabel metal2 579830 112965 579830 112965 0 io_oeb[2]
rlabel metal1 4186 292570 4186 292570 0 io_oeb[30]
rlabel metal3 1970 293148 1970 293148 0 io_oeb[31]
rlabel metal3 2062 241060 2062 241060 0 io_oeb[32]
rlabel metal3 2200 188836 2200 188836 0 io_oeb[33]
rlabel metal3 3013 98668 3013 98668 0 io_oeb[34]
rlabel metal3 2039 84660 2039 84660 0 io_oeb[35]
rlabel metal3 1924 45492 1924 45492 0 io_oeb[36]
rlabel metal3 1878 6460 1878 6460 0 io_oeb[37]
rlabel metal2 580198 152915 580198 152915 0 io_oeb[3]
rlabel metal2 580198 192831 580198 192831 0 io_oeb[4]
rlabel metal2 580198 232781 580198 232781 0 io_oeb[5]
rlabel metal2 579922 272697 579922 272697 0 io_oeb[6]
rlabel metal2 500250 320824 500250 320824 0 io_oeb[7]
rlabel metal2 580198 378301 580198 378301 0 io_oeb[8]
rlabel metal3 582092 431596 582092 431596 0 io_oeb[9]
rlabel metal2 580014 20213 580014 20213 0 io_out[0]
rlabel metal3 582046 471444 582046 471444 0 io_out[10]
rlabel via2 580198 524467 580198 524467 0 io_out[11]
rlabel metal2 580014 577269 580014 577269 0 io_out[12]
rlabel metal3 582000 630836 582000 630836 0 io_out[13]
rlabel metal2 579646 683519 579646 683519 0 io_out[14]
rlabel metal2 543490 701957 543490 701957 0 io_out[15]
rlabel metal1 446108 422994 446108 422994 0 io_out[16]
rlabel metal2 449650 327964 449650 327964 0 io_out[17]
rlabel metal2 348818 695072 348818 695072 0 io_out[18]
rlabel metal2 446706 502758 446706 502758 0 io_out[19]
rlabel metal2 580198 60163 580198 60163 0 io_out[1]
rlabel metal2 219006 702144 219006 702144 0 io_out[20]
rlabel metal2 154146 702110 154146 702110 0 io_out[21]
rlabel metal2 89194 694392 89194 694392 0 io_out[22]
rlabel metal2 24334 695021 24334 695021 0 io_out[23]
rlabel metal3 2039 671228 2039 671228 0 io_out[24]
rlabel metal3 1947 619140 1947 619140 0 io_out[25]
rlabel metal3 1832 566916 1832 566916 0 io_out[26]
rlabel metal3 2108 514828 2108 514828 0 io_out[27]
rlabel metal3 1924 462604 1924 462604 0 io_out[28]
rlabel metal3 2154 410516 2154 410516 0 io_out[29]
rlabel metal2 580198 100079 580198 100079 0 io_out[2]
rlabel metal1 5336 59330 5336 59330 0 io_out[30]
rlabel metal3 2016 306204 2016 306204 0 io_out[31]
rlabel metal3 1878 254116 1878 254116 0 io_out[32]
rlabel metal3 2154 201892 2154 201892 0 io_out[33]
rlabel metal3 1786 149804 1786 149804 0 io_out[34]
rlabel metal3 1947 97580 1947 97580 0 io_out[35]
rlabel metal3 1924 58548 1924 58548 0 io_out[36]
rlabel metal3 1878 19380 1878 19380 0 io_out[37]
rlabel via2 580198 139349 580198 139349 0 io_out[3]
rlabel metal2 580198 179265 580198 179265 0 io_out[4]
rlabel metal3 581908 219028 581908 219028 0 io_out[5]
rlabel metal2 468786 292939 468786 292939 0 io_out[6]
rlabel metal2 580198 312647 580198 312647 0 io_out[7]
rlabel metal2 580198 364735 580198 364735 0 io_out[8]
rlabel metal1 580842 330514 580842 330514 0 io_out[9]
rlabel metal2 488421 322116 488421 322116 0 oeb_6502
rlabel metal3 539281 137972 539281 137972 0 oeb_as1802
rlabel metal2 462622 386910 462622 386910 0 oeb_as2650
rlabel via2 447166 383605 447166 383605 0 oeb_as512512512
rlabel metal2 503293 385900 503293 385900 0 oeb_as5401
rlabel metal3 449566 358428 449566 358428 0 oeb_mc14500
rlabel metal2 448346 159868 448346 159868 0 rst_6502
rlabel metal2 427478 446070 427478 446070 0 rst_LCD
rlabel metal3 449014 345508 449014 345508 0 rst_as1802
rlabel metal3 449129 346188 449129 346188 0 rst_as2650
rlabel metal2 447166 347633 447166 347633 0 rst_as512512512
rlabel metal3 449198 346868 449198 346868 0 rst_as5401
rlabel metal3 449796 348228 449796 348228 0 rst_counter
rlabel metal3 449152 348908 449152 348908 0 rst_diceroll
rlabel metal3 449980 349588 449980 349588 0 rst_mc14500
rlabel metal3 449934 350268 449934 350268 0 rst_posit
rlabel metal2 405957 334900 405957 334900 0 rst_tbb1143
rlabel metal3 448738 351628 448738 351628 0 rst_tune
rlabel metal2 598 1843 598 1843 0 wb_clk_i
rlabel metal2 1702 1911 1702 1911 0 wb_rst_i
rlabel metal2 2898 1979 2898 1979 0 wbs_ack_o
rlabel metal2 406686 175457 406686 175457 0 wbs_adr_i[0]
rlabel metal2 406778 175321 406778 175321 0 wbs_adr_i[10]
rlabel metal2 406502 175474 406502 175474 0 wbs_adr_i[11]
rlabel metal2 403834 175474 403834 175474 0 wbs_adr_i[12]
rlabel metal2 58466 22702 58466 22702 0 wbs_adr_i[13]
rlabel metal2 62054 22736 62054 22736 0 wbs_adr_i[14]
rlabel metal2 403742 175508 403742 175508 0 wbs_adr_i[15]
rlabel metal2 404018 174148 404018 174148 0 wbs_adr_i[16]
rlabel metal1 236900 42262 236900 42262 0 wbs_adr_i[17]
rlabel metal2 76222 21342 76222 21342 0 wbs_adr_i[18]
rlabel metal2 79718 21376 79718 21376 0 wbs_adr_i[19]
rlabel metal1 206816 42058 206816 42058 0 wbs_adr_i[1]
rlabel metal2 83306 21410 83306 21410 0 wbs_adr_i[20]
rlabel metal1 242650 42534 242650 42534 0 wbs_adr_i[21]
rlabel metal1 244260 42602 244260 42602 0 wbs_adr_i[22]
rlabel metal2 93978 21546 93978 21546 0 wbs_adr_i[23]
rlabel metal2 97474 21172 97474 21172 0 wbs_adr_i[24]
rlabel metal2 101062 21240 101062 21240 0 wbs_adr_i[25]
rlabel metal2 451122 178211 451122 178211 0 wbs_adr_i[26]
rlabel metal1 251988 44642 251988 44642 0 wbs_adr_i[27]
rlabel metal1 285936 42194 285936 42194 0 wbs_adr_i[28]
rlabel metal2 115230 19812 115230 19812 0 wbs_adr_i[29]
rlabel metal2 17066 1894 17066 1894 0 wbs_adr_i[2]
rlabel metal2 118818 20084 118818 20084 0 wbs_adr_i[30]
rlabel metal2 122314 19778 122314 19778 0 wbs_adr_i[31]
rlabel metal2 21850 1996 21850 1996 0 wbs_adr_i[3]
rlabel metal2 450938 178143 450938 178143 0 wbs_adr_i[4]
rlabel metal2 30130 1214 30130 1214 0 wbs_adr_i[5]
rlabel metal2 33626 2132 33626 2132 0 wbs_adr_i[6]
rlabel metal2 37214 2064 37214 2064 0 wbs_adr_i[7]
rlabel metal2 40710 19914 40710 19914 0 wbs_adr_i[8]
rlabel metal2 44298 19948 44298 19948 0 wbs_adr_i[9]
rlabel metal2 4094 19880 4094 19880 0 wbs_cyc_i
rlabel metal2 392610 152116 392610 152116 0 wbs_dat_i[0]
rlabel metal2 392886 170034 392886 170034 0 wbs_dat_i[10]
rlabel metal2 52578 1928 52578 1928 0 wbs_dat_i[11]
rlabel metal2 56074 20050 56074 20050 0 wbs_dat_i[12]
rlabel metal2 59662 20118 59662 20118 0 wbs_dat_i[13]
rlabel metal2 63250 18486 63250 18486 0 wbs_dat_i[14]
rlabel metal2 389942 168470 389942 168470 0 wbs_dat_i[15]
rlabel metal2 390126 167008 390126 167008 0 wbs_dat_i[16]
rlabel metal2 390034 167416 390034 167416 0 wbs_dat_i[17]
rlabel metal2 77418 18622 77418 18622 0 wbs_dat_i[18]
rlabel metal2 80914 21512 80914 21512 0 wbs_dat_i[19]
rlabel metal2 387090 150603 387090 150603 0 wbs_dat_i[1]
rlabel metal2 387550 171258 387550 171258 0 wbs_dat_i[20]
rlabel metal2 387274 167280 387274 167280 0 wbs_dat_i[21]
rlabel metal2 387182 167382 387182 167382 0 wbs_dat_i[22]
rlabel metal2 95174 18724 95174 18724 0 wbs_dat_i[23]
rlabel metal2 98670 18758 98670 18758 0 wbs_dat_i[24]
rlabel metal2 102258 20186 102258 20186 0 wbs_dat_i[25]
rlabel metal2 384514 167348 384514 167348 0 wbs_dat_i[26]
rlabel metal1 245548 36482 245548 36482 0 wbs_dat_i[27]
rlabel metal2 518926 333880 518926 333880 0 wbs_dat_i[28]
rlabel metal2 116426 17364 116426 17364 0 wbs_dat_i[29]
rlabel metal2 18262 17058 18262 17058 0 wbs_dat_i[2]
rlabel metal2 119922 17398 119922 17398 0 wbs_dat_i[30]
rlabel metal1 445694 386546 445694 386546 0 wbs_dat_i[31]
rlabel metal2 23046 17092 23046 17092 0 wbs_dat_i[3]
rlabel metal2 27738 2098 27738 2098 0 wbs_dat_i[4]
rlabel metal2 520858 314636 520858 314636 0 wbs_dat_i[5]
rlabel metal2 519754 316064 519754 316064 0 wbs_dat_i[6]
rlabel metal2 38410 22770 38410 22770 0 wbs_dat_i[7]
rlabel metal2 41906 17194 41906 17194 0 wbs_dat_i[8]
rlabel metal2 45494 17228 45494 17228 0 wbs_dat_i[9]
rlabel metal2 507518 308329 507518 308329 0 wbs_dat_o[0]
rlabel metal1 446292 294882 446292 294882 0 wbs_dat_o[10]
rlabel metal2 53774 2200 53774 2200 0 wbs_dat_o[11]
rlabel metal2 57270 17296 57270 17296 0 wbs_dat_o[12]
rlabel metal2 60858 17330 60858 17330 0 wbs_dat_o[13]
rlabel metal2 64354 15766 64354 15766 0 wbs_dat_o[14]
rlabel metal2 373382 161466 373382 161466 0 wbs_dat_o[15]
rlabel metal2 373566 166158 373566 166158 0 wbs_dat_o[16]
rlabel metal2 75026 15834 75026 15834 0 wbs_dat_o[17]
rlabel metal2 78614 15868 78614 15868 0 wbs_dat_o[18]
rlabel metal2 82110 2030 82110 2030 0 wbs_dat_o[19]
rlabel metal2 370714 161398 370714 161398 0 wbs_dat_o[1]
rlabel metal2 85698 2234 85698 2234 0 wbs_dat_o[20]
rlabel metal2 370530 161670 370530 161670 0 wbs_dat_o[21]
rlabel metal2 92782 1860 92782 1860 0 wbs_dat_o[22]
rlabel metal2 96278 15936 96278 15936 0 wbs_dat_o[23]
rlabel metal2 99866 15970 99866 15970 0 wbs_dat_o[24]
rlabel metal2 103362 1826 103362 1826 0 wbs_dat_o[25]
rlabel metal2 370990 166940 370990 166940 0 wbs_dat_o[26]
rlabel metal2 110538 1792 110538 1792 0 wbs_dat_o[27]
rlabel metal2 114034 16004 114034 16004 0 wbs_dat_o[28]
rlabel metal2 117622 16038 117622 16038 0 wbs_dat_o[29]
rlabel metal2 19458 15732 19458 15732 0 wbs_dat_o[2]
rlabel metal2 121118 15664 121118 15664 0 wbs_dat_o[30]
rlabel metal2 367862 208658 367862 208658 0 wbs_dat_o[31]
rlabel metal2 24242 1962 24242 1962 0 wbs_dat_o[3]
rlabel metal2 368230 162962 368230 162962 0 wbs_dat_o[4]
rlabel metal2 365194 158712 365194 158712 0 wbs_dat_o[5]
rlabel metal2 36018 14338 36018 14338 0 wbs_dat_o[6]
rlabel metal2 39606 2166 39606 2166 0 wbs_dat_o[7]
rlabel metal2 43102 14372 43102 14372 0 wbs_dat_o[8]
rlabel metal2 365286 158882 365286 158882 0 wbs_dat_o[9]
rlabel metal2 5290 1775 5290 1775 0 wbs_stb_i
rlabel metal2 6486 1758 6486 1758 0 wbs_we_i
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
