magic
tech sky130B
magscale 1 2
timestamp 1683540219
<< obsli1 >>
rect 1104 2159 68816 67473
<< obsm1 >>
rect 382 1844 68816 67504
<< metal2 >>
rect 3238 0 3294 800
rect 9586 0 9642 800
rect 15934 0 15990 800
rect 22282 0 22338 800
rect 28630 0 28686 800
rect 34978 0 35034 800
rect 41326 0 41382 800
rect 47674 0 47730 800
rect 54022 0 54078 800
rect 60370 0 60426 800
rect 66718 0 66774 800
<< obsm2 >>
rect 294 856 68060 67969
rect 294 800 3182 856
rect 3350 800 9530 856
rect 9698 800 15878 856
rect 16046 800 22226 856
rect 22394 800 28574 856
rect 28742 800 34922 856
rect 35090 800 41270 856
rect 41438 800 47618 856
rect 47786 800 53966 856
rect 54134 800 60314 856
rect 60482 800 66662 856
rect 66830 800 68060 856
<< metal3 >>
rect 0 67872 800 67992
rect 0 65424 800 65544
rect 0 62976 800 63096
rect 0 60528 800 60648
rect 0 58080 800 58200
rect 0 55632 800 55752
rect 0 53184 800 53304
rect 0 50736 800 50856
rect 0 48288 800 48408
rect 0 45840 800 45960
rect 0 43392 800 43512
rect 0 40944 800 41064
rect 0 38496 800 38616
rect 0 36048 800 36168
rect 0 33600 800 33720
rect 0 31152 800 31272
rect 0 28704 800 28824
rect 0 26256 800 26376
rect 0 23808 800 23928
rect 0 21360 800 21480
rect 0 18912 800 19032
rect 0 16464 800 16584
rect 0 14016 800 14136
rect 0 11568 800 11688
rect 0 9120 800 9240
rect 0 6672 800 6792
rect 0 4224 800 4344
rect 0 1776 800 1896
<< obsm3 >>
rect 880 67792 65966 67965
rect 289 65624 65966 67792
rect 880 65344 65966 65624
rect 289 63176 65966 65344
rect 880 62896 65966 63176
rect 289 60728 65966 62896
rect 880 60448 65966 60728
rect 289 58280 65966 60448
rect 880 58000 65966 58280
rect 289 55832 65966 58000
rect 880 55552 65966 55832
rect 289 53384 65966 55552
rect 880 53104 65966 53384
rect 289 50936 65966 53104
rect 880 50656 65966 50936
rect 289 48488 65966 50656
rect 880 48208 65966 48488
rect 289 46040 65966 48208
rect 880 45760 65966 46040
rect 289 43592 65966 45760
rect 880 43312 65966 43592
rect 289 41144 65966 43312
rect 880 40864 65966 41144
rect 289 38696 65966 40864
rect 880 38416 65966 38696
rect 289 36248 65966 38416
rect 880 35968 65966 36248
rect 289 33800 65966 35968
rect 880 33520 65966 33800
rect 289 31352 65966 33520
rect 880 31072 65966 31352
rect 289 28904 65966 31072
rect 880 28624 65966 28904
rect 289 26456 65966 28624
rect 880 26176 65966 26456
rect 289 24008 65966 26176
rect 880 23728 65966 24008
rect 289 21560 65966 23728
rect 880 21280 65966 21560
rect 289 19112 65966 21280
rect 880 18832 65966 19112
rect 289 16664 65966 18832
rect 880 16384 65966 16664
rect 289 14216 65966 16384
rect 880 13936 65966 14216
rect 289 11768 65966 13936
rect 880 11488 65966 11768
rect 289 9320 65966 11488
rect 880 9040 65966 9320
rect 289 6872 65966 9040
rect 880 6592 65966 6872
rect 289 4424 65966 6592
rect 880 4144 65966 4424
rect 289 1976 65966 4144
rect 880 1803 65966 1976
<< metal4 >>
rect 4208 2128 4528 67504
rect 19568 2128 19888 67504
rect 34928 2128 35248 67504
rect 50288 2128 50608 67504
rect 65648 2128 65968 67504
<< obsm4 >>
rect 795 2347 4128 66741
rect 4608 2347 19488 66741
rect 19968 2347 34848 66741
rect 35328 2347 50208 66741
rect 50688 2347 56245 66741
<< labels >>
rlabel metal2 s 60370 0 60426 800 6 clk
port 1 nsew signal input
rlabel metal2 s 3238 0 3294 800 6 io_in[0]
port 2 nsew signal input
rlabel metal2 s 9586 0 9642 800 6 io_in[1]
port 3 nsew signal input
rlabel metal2 s 15934 0 15990 800 6 io_in[2]
port 4 nsew signal input
rlabel metal2 s 22282 0 22338 800 6 io_in[3]
port 5 nsew signal input
rlabel metal2 s 28630 0 28686 800 6 io_in[4]
port 6 nsew signal input
rlabel metal2 s 34978 0 35034 800 6 io_in[5]
port 7 nsew signal input
rlabel metal2 s 41326 0 41382 800 6 io_in[6]
port 8 nsew signal input
rlabel metal2 s 47674 0 47730 800 6 io_in[7]
port 9 nsew signal input
rlabel metal2 s 54022 0 54078 800 6 io_in[8]
port 10 nsew signal input
rlabel metal3 s 0 67872 800 67992 6 io_oeb
port 11 nsew signal output
rlabel metal3 s 0 1776 800 1896 6 io_out[0]
port 12 nsew signal output
rlabel metal3 s 0 26256 800 26376 6 io_out[10]
port 13 nsew signal output
rlabel metal3 s 0 28704 800 28824 6 io_out[11]
port 14 nsew signal output
rlabel metal3 s 0 31152 800 31272 6 io_out[12]
port 15 nsew signal output
rlabel metal3 s 0 33600 800 33720 6 io_out[13]
port 16 nsew signal output
rlabel metal3 s 0 36048 800 36168 6 io_out[14]
port 17 nsew signal output
rlabel metal3 s 0 38496 800 38616 6 io_out[15]
port 18 nsew signal output
rlabel metal3 s 0 40944 800 41064 6 io_out[16]
port 19 nsew signal output
rlabel metal3 s 0 43392 800 43512 6 io_out[17]
port 20 nsew signal output
rlabel metal3 s 0 45840 800 45960 6 io_out[18]
port 21 nsew signal output
rlabel metal3 s 0 48288 800 48408 6 io_out[19]
port 22 nsew signal output
rlabel metal3 s 0 4224 800 4344 6 io_out[1]
port 23 nsew signal output
rlabel metal3 s 0 50736 800 50856 6 io_out[20]
port 24 nsew signal output
rlabel metal3 s 0 53184 800 53304 6 io_out[21]
port 25 nsew signal output
rlabel metal3 s 0 55632 800 55752 6 io_out[22]
port 26 nsew signal output
rlabel metal3 s 0 58080 800 58200 6 io_out[23]
port 27 nsew signal output
rlabel metal3 s 0 60528 800 60648 6 io_out[24]
port 28 nsew signal output
rlabel metal3 s 0 62976 800 63096 6 io_out[25]
port 29 nsew signal output
rlabel metal3 s 0 65424 800 65544 6 io_out[26]
port 30 nsew signal output
rlabel metal3 s 0 6672 800 6792 6 io_out[2]
port 31 nsew signal output
rlabel metal3 s 0 9120 800 9240 6 io_out[3]
port 32 nsew signal output
rlabel metal3 s 0 11568 800 11688 6 io_out[4]
port 33 nsew signal output
rlabel metal3 s 0 14016 800 14136 6 io_out[5]
port 34 nsew signal output
rlabel metal3 s 0 16464 800 16584 6 io_out[6]
port 35 nsew signal output
rlabel metal3 s 0 18912 800 19032 6 io_out[7]
port 36 nsew signal output
rlabel metal3 s 0 21360 800 21480 6 io_out[8]
port 37 nsew signal output
rlabel metal3 s 0 23808 800 23928 6 io_out[9]
port 38 nsew signal output
rlabel metal2 s 66718 0 66774 800 6 rst
port 39 nsew signal input
rlabel metal4 s 4208 2128 4528 67504 6 vccd1
port 40 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 67504 6 vccd1
port 40 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 67504 6 vccd1
port 40 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 67504 6 vssd1
port 41 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 67504 6 vssd1
port 41 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 70000 70000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 15943890
string GDS_FILE /media/lucah/e6042058-84c8-448b-be8a-b40bc065b34b/TMBoC/openlane/AS2650/runs/23_05_08_11_47/results/signoff/wrapped_as2650.magic.gds
string GDS_START 1385758
<< end >>

