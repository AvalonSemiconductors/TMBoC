magic
tech sky130B
magscale 1 2
timestamp 1681463552
<< metal1 >>
rect 397454 700816 397460 700868
rect 397512 700856 397518 700868
rect 444098 700856 444104 700868
rect 397512 700828 444104 700856
rect 397512 700816 397518 700828
rect 444098 700816 444104 700828
rect 444156 700816 444162 700868
rect 364978 700748 364984 700800
rect 365036 700788 365042 700800
rect 446490 700788 446496 700800
rect 365036 700760 446496 700788
rect 365036 700748 365042 700760
rect 446490 700748 446496 700760
rect 446548 700748 446554 700800
rect 332502 700680 332508 700732
rect 332560 700720 332566 700732
rect 445018 700720 445024 700732
rect 332560 700692 445024 700720
rect 332560 700680 332566 700692
rect 445018 700680 445024 700692
rect 445076 700680 445082 700732
rect 267642 700612 267648 700664
rect 267700 700652 267706 700664
rect 449250 700652 449256 700664
rect 267700 700624 449256 700652
rect 267700 700612 267706 700624
rect 449250 700612 449256 700624
rect 449308 700612 449314 700664
rect 235166 700544 235172 700596
rect 235224 700584 235230 700596
rect 449158 700584 449164 700596
rect 235224 700556 449164 700584
rect 235224 700544 235230 700556
rect 449158 700544 449164 700556
rect 449216 700544 449222 700596
rect 170306 700476 170312 700528
rect 170364 700516 170370 700528
rect 446398 700516 446404 700528
rect 170364 700488 446404 700516
rect 170364 700476 170370 700488
rect 446398 700476 446404 700488
rect 446456 700476 446462 700528
rect 154114 700408 154120 700460
rect 154172 700448 154178 700460
rect 445110 700448 445116 700460
rect 154172 700420 445116 700448
rect 154172 700408 154178 700420
rect 445110 700408 445116 700420
rect 445168 700408 445174 700460
rect 105446 700340 105452 700392
rect 105504 700380 105510 700392
rect 444190 700380 444196 700392
rect 105504 700352 444196 700380
rect 105504 700340 105510 700352
rect 444190 700340 444196 700352
rect 444248 700340 444254 700392
rect 445662 700340 445668 700392
rect 445720 700380 445726 700392
rect 478506 700380 478512 700392
rect 445720 700352 478512 700380
rect 445720 700340 445726 700352
rect 478506 700340 478512 700352
rect 478564 700340 478570 700392
rect 8110 700272 8116 700324
rect 8168 700312 8174 700324
rect 418798 700312 418804 700324
rect 8168 700284 418804 700312
rect 8168 700272 8174 700284
rect 418798 700272 418804 700284
rect 418856 700272 418862 700324
rect 447870 700272 447876 700324
rect 447928 700312 447934 700324
rect 494790 700312 494796 700324
rect 447928 700284 494796 700312
rect 447928 700272 447934 700284
rect 494790 700272 494796 700284
rect 494848 700272 494854 700324
rect 571978 696940 571984 696992
rect 572036 696980 572042 696992
rect 580166 696980 580172 696992
rect 572036 696952 580172 696980
rect 572036 696940 572042 696952
rect 580166 696940 580172 696952
rect 580224 696940 580230 696992
rect 218974 692044 218980 692096
rect 219032 692084 219038 692096
rect 446582 692084 446588 692096
rect 219032 692056 446588 692084
rect 219032 692044 219038 692056
rect 446582 692044 446588 692056
rect 446640 692044 446646 692096
rect 283834 687896 283840 687948
rect 283892 687936 283898 687948
rect 446674 687936 446680 687948
rect 283892 687908 446680 687936
rect 283892 687896 283898 687908
rect 446674 687896 446680 687908
rect 446732 687896 446738 687948
rect 348786 686468 348792 686520
rect 348844 686508 348850 686520
rect 445202 686508 445208 686520
rect 348844 686480 445208 686508
rect 348844 686468 348850 686480
rect 445202 686468 445208 686480
rect 445260 686468 445266 686520
rect 137830 685244 137836 685296
rect 137888 685284 137894 685296
rect 446766 685284 446772 685296
rect 137888 685256 446772 685284
rect 137888 685244 137894 685256
rect 446766 685244 446772 685256
rect 446824 685244 446830 685296
rect 89162 685176 89168 685228
rect 89220 685216 89226 685228
rect 416038 685216 416044 685228
rect 89220 685188 416044 685216
rect 89220 685176 89226 685188
rect 416038 685176 416044 685188
rect 416096 685176 416102 685228
rect 72970 685108 72976 685160
rect 73028 685148 73034 685160
rect 418890 685148 418896 685160
rect 73028 685120 418896 685148
rect 73028 685108 73034 685120
rect 418890 685108 418896 685120
rect 418948 685108 418954 685160
rect 3878 684496 3884 684548
rect 3936 684536 3942 684548
rect 445570 684536 445576 684548
rect 3936 684508 445576 684536
rect 3936 684496 3942 684508
rect 445570 684496 445576 684508
rect 445628 684496 445634 684548
rect 24118 683884 24124 683936
rect 24176 683924 24182 683936
rect 359458 683924 359464 683936
rect 24176 683896 359464 683924
rect 24176 683884 24182 683896
rect 359458 683884 359464 683896
rect 359516 683884 359522 683936
rect 19978 683816 19984 683868
rect 20036 683856 20042 683868
rect 418982 683856 418988 683868
rect 20036 683828 418988 683856
rect 20036 683816 20042 683828
rect 418982 683816 418988 683828
rect 419040 683816 419046 683868
rect 21358 683748 21364 683800
rect 21416 683788 21422 683800
rect 420638 683788 420644 683800
rect 21416 683760 420644 683788
rect 21416 683748 21422 683760
rect 420638 683748 420644 683760
rect 420696 683748 420702 683800
rect 4062 683680 4068 683732
rect 4120 683720 4126 683732
rect 420178 683720 420184 683732
rect 4120 683692 420184 683720
rect 4120 683680 4126 683692
rect 420178 683680 420184 683692
rect 420236 683680 420242 683732
rect 3510 683612 3516 683664
rect 3568 683652 3574 683664
rect 420362 683652 420368 683664
rect 3568 683624 420368 683652
rect 3568 683612 3574 683624
rect 420362 683612 420368 683624
rect 420420 683612 420426 683664
rect 3326 683544 3332 683596
rect 3384 683584 3390 683596
rect 420270 683584 420276 683596
rect 3384 683556 420276 683584
rect 3384 683544 3390 683556
rect 420270 683544 420276 683556
rect 420328 683544 420334 683596
rect 3694 683476 3700 683528
rect 3752 683516 3758 683528
rect 420730 683516 420736 683528
rect 3752 683488 420736 683516
rect 3752 683476 3758 683488
rect 420730 683476 420736 683488
rect 420788 683476 420794 683528
rect 3418 683408 3424 683460
rect 3476 683448 3482 683460
rect 420546 683448 420552 683460
rect 3476 683420 420552 683448
rect 3476 683408 3482 683420
rect 420546 683408 420552 683420
rect 420604 683408 420610 683460
rect 3602 683340 3608 683392
rect 3660 683380 3666 683392
rect 420822 683380 420828 683392
rect 3660 683352 420828 683380
rect 3660 683340 3666 683352
rect 420822 683340 420828 683352
rect 420880 683340 420886 683392
rect 3786 683272 3792 683324
rect 3844 683312 3850 683324
rect 445294 683312 445300 683324
rect 3844 683284 445300 683312
rect 3844 683272 3850 683284
rect 445294 683272 445300 683284
rect 445352 683272 445358 683324
rect 3970 683204 3976 683256
rect 4028 683244 4034 683256
rect 445478 683244 445484 683256
rect 4028 683216 445484 683244
rect 4028 683204 4034 683216
rect 445478 683204 445484 683216
rect 445536 683204 445542 683256
rect 3234 683136 3240 683188
rect 3292 683176 3298 683188
rect 445386 683176 445392 683188
rect 3292 683148 445392 683176
rect 3292 683136 3298 683148
rect 445386 683136 445392 683148
rect 445444 683136 445450 683188
rect 573358 683136 573364 683188
rect 573416 683176 573422 683188
rect 580166 683176 580172 683188
rect 573416 683148 580172 683176
rect 573416 683136 573422 683148
rect 580166 683136 580172 683148
rect 580224 683136 580230 683188
rect 19242 682728 19248 682780
rect 19300 682768 19306 682780
rect 24118 682768 24124 682780
rect 19300 682740 24124 682768
rect 19300 682728 19306 682740
rect 24118 682728 24124 682740
rect 24176 682728 24182 682780
rect 3234 682660 3240 682712
rect 3292 682700 3298 682712
rect 446950 682700 446956 682712
rect 3292 682672 446956 682700
rect 3292 682660 3298 682672
rect 446950 682660 446956 682672
rect 447008 682660 447014 682712
rect 17218 680348 17224 680400
rect 17276 680388 17282 680400
rect 19242 680388 19248 680400
rect 17276 680360 19248 680388
rect 17276 680348 17282 680360
rect 19242 680348 19248 680360
rect 19300 680348 19306 680400
rect 361758 678988 361764 679040
rect 361816 679028 361822 679040
rect 387058 679028 387064 679040
rect 361816 679000 387064 679028
rect 361816 678988 361822 679000
rect 387058 678988 387064 679000
rect 387116 678988 387122 679040
rect 570598 670692 570604 670744
rect 570656 670732 570662 670744
rect 580166 670732 580172 670744
rect 570656 670704 580172 670732
rect 570656 670692 570662 670704
rect 580166 670692 580172 670704
rect 580224 670692 580230 670744
rect 447778 669944 447784 669996
rect 447836 669984 447842 669996
rect 462314 669984 462320 669996
rect 447836 669956 462320 669984
rect 447836 669944 447842 669956
rect 462314 669944 462320 669956
rect 462372 669944 462378 669996
rect 361758 667904 361764 667956
rect 361816 667944 361822 667956
rect 382918 667944 382924 667956
rect 361816 667916 382924 667944
rect 361816 667904 361822 667916
rect 382918 667904 382924 667916
rect 382976 667904 382982 667956
rect 17218 661076 17224 661088
rect 16546 661048 17224 661076
rect 14182 660968 14188 661020
rect 14240 661008 14246 661020
rect 16546 661008 16574 661048
rect 17218 661036 17224 661048
rect 17276 661036 17282 661088
rect 14240 660980 16574 661008
rect 14240 660968 14246 660980
rect 3142 658180 3148 658232
rect 3200 658220 3206 658232
rect 19978 658220 19984 658232
rect 3200 658192 19984 658220
rect 3200 658180 3206 658192
rect 19978 658180 19984 658192
rect 20036 658180 20042 658232
rect 361758 656888 361764 656940
rect 361816 656928 361822 656940
rect 381538 656928 381544 656940
rect 361816 656900 381544 656928
rect 361816 656888 361822 656900
rect 381538 656888 381544 656900
rect 381596 656888 381602 656940
rect 11698 656616 11704 656668
rect 11756 656656 11762 656668
rect 14182 656656 14188 656668
rect 11756 656628 14188 656656
rect 11756 656616 11762 656628
rect 14182 656616 14188 656628
rect 14240 656616 14246 656668
rect 361758 645872 361764 645924
rect 361816 645912 361822 645924
rect 378778 645912 378784 645924
rect 361816 645884 378784 645912
rect 361816 645872 361822 645884
rect 378778 645872 378784 645884
rect 378836 645872 378842 645924
rect 10594 645804 10600 645856
rect 10652 645844 10658 645856
rect 11698 645844 11704 645856
rect 10652 645816 11704 645844
rect 10652 645804 10658 645816
rect 11698 645804 11704 645816
rect 11756 645804 11762 645856
rect 5534 643696 5540 643748
rect 5592 643736 5598 643748
rect 10594 643736 10600 643748
rect 5592 643708 10600 643736
rect 5592 643696 5598 643708
rect 10594 643696 10600 643708
rect 10652 643696 10658 643748
rect 4798 640296 4804 640348
rect 4856 640336 4862 640348
rect 5534 640336 5540 640348
rect 4856 640308 5540 640336
rect 4856 640296 4862 640308
rect 5534 640296 5540 640308
rect 5592 640296 5598 640348
rect 361574 634788 361580 634840
rect 361632 634828 361638 634840
rect 403618 634828 403624 634840
rect 361632 634800 403624 634828
rect 361632 634788 361638 634800
rect 403618 634788 403624 634800
rect 403676 634788 403682 634840
rect 3694 631320 3700 631372
rect 3752 631360 3758 631372
rect 20898 631360 20904 631372
rect 3752 631332 20904 631360
rect 3752 631320 3758 631332
rect 20898 631320 20904 631332
rect 20956 631320 20962 631372
rect 361574 623772 361580 623824
rect 361632 623812 361638 623824
rect 376018 623812 376024 623824
rect 361632 623784 376024 623812
rect 361632 623772 361638 623784
rect 376018 623772 376024 623784
rect 376076 623772 376082 623824
rect 569218 616836 569224 616888
rect 569276 616876 569282 616888
rect 580166 616876 580172 616888
rect 569276 616848 580172 616876
rect 569276 616836 569282 616848
rect 580166 616836 580172 616848
rect 580224 616836 580230 616888
rect 361574 612756 361580 612808
rect 361632 612796 361638 612808
rect 406378 612796 406384 612808
rect 361632 612768 406384 612796
rect 361632 612756 361638 612768
rect 406378 612756 406384 612768
rect 406436 612756 406442 612808
rect 361758 601672 361764 601724
rect 361816 601712 361822 601724
rect 374638 601712 374644 601724
rect 361816 601684 374644 601712
rect 361816 601672 361822 601684
rect 374638 601672 374644 601684
rect 374696 601672 374702 601724
rect 457622 600584 457628 600636
rect 457680 600624 457686 600636
rect 461578 600624 461584 600636
rect 457680 600596 461584 600624
rect 457680 600584 457686 600596
rect 461578 600584 461584 600596
rect 461636 600584 461642 600636
rect 457714 600244 457720 600296
rect 457772 600284 457778 600296
rect 461670 600284 461676 600296
rect 457772 600256 461676 600284
rect 457772 600244 457778 600256
rect 461670 600244 461676 600256
rect 461728 600244 461734 600296
rect 460014 599836 460020 599888
rect 460072 599876 460078 599888
rect 463694 599876 463700 599888
rect 460072 599848 463700 599876
rect 460072 599836 460078 599848
rect 463694 599836 463700 599848
rect 463752 599836 463758 599888
rect 458634 599700 458640 599752
rect 458692 599740 458698 599752
rect 465074 599740 465080 599752
rect 458692 599712 465080 599740
rect 458692 599700 458698 599712
rect 465074 599700 465080 599712
rect 465132 599700 465138 599752
rect 458818 599632 458824 599684
rect 458876 599672 458882 599684
rect 466454 599672 466460 599684
rect 458876 599644 466460 599672
rect 458876 599632 458882 599644
rect 466454 599632 466460 599644
rect 466512 599632 466518 599684
rect 457438 599564 457444 599616
rect 457496 599604 457502 599616
rect 469858 599604 469864 599616
rect 457496 599576 469864 599604
rect 457496 599564 457502 599576
rect 469858 599564 469864 599576
rect 469916 599564 469922 599616
rect 515398 599564 515404 599616
rect 515456 599604 515462 599616
rect 580258 599604 580264 599616
rect 515456 599576 580264 599604
rect 515456 599564 515462 599576
rect 580258 599564 580264 599576
rect 580316 599564 580322 599616
rect 458726 598340 458732 598392
rect 458784 598380 458790 598392
rect 465166 598380 465172 598392
rect 458784 598352 465172 598380
rect 458784 598340 458790 598352
rect 465166 598340 465172 598352
rect 465224 598340 465230 598392
rect 460106 598272 460112 598324
rect 460164 598312 460170 598324
rect 470594 598312 470600 598324
rect 460164 598284 470600 598312
rect 460164 598272 460170 598284
rect 470594 598272 470600 598284
rect 470652 598272 470658 598324
rect 457530 598204 457536 598256
rect 457588 598244 457594 598256
rect 468478 598244 468484 598256
rect 457588 598216 468484 598244
rect 457588 598204 457594 598216
rect 468478 598204 468484 598216
rect 468536 598204 468542 598256
rect 488626 598204 488632 598256
rect 488684 598244 488690 598256
rect 494054 598244 494060 598256
rect 488684 598216 494060 598244
rect 488684 598204 488690 598216
rect 494054 598204 494060 598216
rect 494112 598204 494118 598256
rect 459922 596980 459928 597032
rect 459980 597020 459986 597032
rect 463786 597020 463792 597032
rect 459980 596992 463792 597020
rect 459980 596980 459986 596992
rect 463786 596980 463792 596992
rect 463844 596980 463850 597032
rect 458910 596844 458916 596896
rect 458968 596884 458974 596896
rect 466546 596884 466552 596896
rect 458968 596856 466552 596884
rect 458968 596844 458974 596856
rect 466546 596844 466552 596856
rect 466604 596844 466610 596896
rect 450538 596776 450544 596828
rect 450596 596816 450602 596828
rect 494974 596816 494980 596828
rect 450596 596788 494980 596816
rect 450596 596776 450602 596788
rect 494974 596776 494980 596788
rect 495032 596776 495038 596828
rect 457346 596164 457352 596216
rect 457404 596204 457410 596216
rect 462958 596204 462964 596216
rect 457404 596176 462964 596204
rect 457404 596164 457410 596176
rect 462958 596164 462964 596176
rect 463016 596164 463022 596216
rect 457806 595416 457812 595468
rect 457864 595456 457870 595468
rect 468570 595456 468576 595468
rect 457864 595428 468576 595456
rect 457864 595416 457870 595428
rect 468570 595416 468576 595428
rect 468628 595416 468634 595468
rect 460198 594396 460204 594448
rect 460256 594436 460262 594448
rect 462314 594436 462320 594448
rect 460256 594408 462320 594436
rect 460256 594396 460262 594408
rect 462314 594396 462320 594408
rect 462372 594396 462378 594448
rect 457254 592628 457260 592680
rect 457312 592668 457318 592680
rect 465718 592668 465724 592680
rect 457312 592640 465724 592668
rect 457312 592628 457318 592640
rect 465718 592628 465724 592640
rect 465776 592628 465782 592680
rect 361758 590656 361764 590708
rect 361816 590696 361822 590708
rect 407758 590696 407764 590708
rect 361816 590668 407764 590696
rect 361816 590656 361822 590668
rect 407758 590656 407764 590668
rect 407816 590656 407822 590708
rect 519538 590656 519544 590708
rect 519596 590696 519602 590708
rect 580166 590696 580172 590708
rect 519596 590668 580172 590696
rect 519596 590656 519602 590668
rect 580166 590656 580172 590668
rect 580224 590656 580230 590708
rect 361758 579640 361764 579692
rect 361816 579680 361822 579692
rect 371878 579680 371884 579692
rect 361816 579652 371884 579680
rect 361816 579640 361822 579652
rect 371878 579640 371884 579652
rect 371936 579640 371942 579692
rect 574738 576852 574744 576904
rect 574796 576892 574802 576904
rect 580166 576892 580172 576904
rect 574796 576864 580172 576892
rect 574796 576852 574802 576864
rect 580166 576852 580172 576864
rect 580224 576852 580230 576904
rect 361574 568760 361580 568812
rect 361632 568800 361638 568812
rect 363598 568800 363604 568812
rect 361632 568772 363604 568800
rect 361632 568760 361638 568772
rect 363598 568760 363604 568772
rect 363656 568760 363662 568812
rect 359458 561620 359464 561672
rect 359516 561660 359522 561672
rect 362218 561660 362224 561672
rect 359516 561632 362224 561660
rect 359516 561620 359522 561632
rect 362218 561620 362224 561632
rect 362276 561620 362282 561672
rect 361666 557540 361672 557592
rect 361724 557580 361730 557592
rect 370498 557580 370504 557592
rect 361724 557552 370504 557580
rect 361724 557540 361730 557552
rect 370498 557540 370504 557552
rect 370556 557540 370562 557592
rect 362218 551284 362224 551336
rect 362276 551324 362282 551336
rect 369118 551324 369124 551336
rect 362276 551296 369124 551324
rect 362276 551284 362282 551296
rect 369118 551284 369124 551296
rect 369176 551284 369182 551336
rect 361758 546456 361764 546508
rect 361816 546496 361822 546508
rect 367738 546496 367744 546508
rect 361816 546468 367744 546496
rect 361816 546456 361822 546468
rect 367738 546456 367744 546468
rect 367796 546456 367802 546508
rect 459462 544348 459468 544400
rect 459520 544388 459526 544400
rect 470870 544388 470876 544400
rect 459520 544360 470876 544388
rect 459520 544348 459526 544360
rect 470870 544348 470876 544360
rect 470928 544348 470934 544400
rect 518158 536800 518164 536852
rect 518216 536840 518222 536852
rect 580166 536840 580172 536852
rect 518216 536812 580172 536840
rect 518216 536800 518222 536812
rect 580166 536800 580172 536812
rect 580224 536800 580230 536852
rect 361574 535440 361580 535492
rect 361632 535480 361638 535492
rect 363690 535480 363696 535492
rect 361632 535452 363696 535480
rect 361632 535440 361638 535452
rect 363690 535440 363696 535452
rect 363748 535440 363754 535492
rect 361574 524696 361580 524748
rect 361632 524736 361638 524748
rect 363782 524736 363788 524748
rect 361632 524708 363788 524736
rect 361632 524696 361638 524708
rect 363782 524696 363788 524708
rect 363840 524696 363846 524748
rect 369118 522248 369124 522300
rect 369176 522288 369182 522300
rect 378870 522288 378876 522300
rect 369176 522260 378876 522288
rect 369176 522248 369182 522260
rect 378870 522248 378876 522260
rect 378928 522248 378934 522300
rect 457898 520888 457904 520940
rect 457956 520928 457962 520940
rect 467926 520928 467932 520940
rect 457956 520900 467932 520928
rect 457956 520888 457962 520900
rect 467926 520888 467932 520900
rect 467984 520888 467990 520940
rect 482922 520888 482928 520940
rect 482980 520928 482986 520940
rect 520274 520928 520280 520940
rect 482980 520900 520280 520928
rect 482980 520888 482986 520900
rect 520274 520888 520280 520900
rect 520332 520888 520338 520940
rect 464338 520276 464344 520328
rect 464396 520316 464402 520328
rect 488626 520316 488632 520328
rect 464396 520288 488632 520316
rect 464396 520276 464402 520288
rect 488626 520276 488632 520288
rect 488684 520276 488690 520328
rect 458082 519528 458088 519580
rect 458140 519568 458146 519580
rect 465810 519568 465816 519580
rect 458140 519540 465816 519568
rect 458140 519528 458146 519540
rect 465810 519528 465816 519540
rect 465868 519528 465874 519580
rect 459830 518372 459836 518424
rect 459888 518412 459894 518424
rect 462406 518412 462412 518424
rect 459888 518384 462412 518412
rect 459888 518372 459894 518384
rect 462406 518372 462412 518384
rect 462464 518372 462470 518424
rect 457990 518236 457996 518288
rect 458048 518276 458054 518288
rect 469950 518276 469956 518288
rect 458048 518248 469956 518276
rect 458048 518236 458054 518248
rect 469950 518236 469956 518248
rect 470008 518236 470014 518288
rect 449802 518168 449808 518220
rect 449860 518208 449866 518220
rect 470042 518208 470048 518220
rect 449860 518180 470048 518208
rect 449860 518168 449866 518180
rect 470042 518168 470048 518180
rect 470100 518208 470106 518220
rect 494238 518208 494244 518220
rect 470100 518180 494244 518208
rect 470100 518168 470106 518180
rect 494238 518168 494244 518180
rect 494296 518168 494302 518220
rect 476022 517556 476028 517608
rect 476080 517596 476086 517608
rect 494146 517596 494152 517608
rect 476080 517568 494152 517596
rect 476080 517556 476086 517568
rect 494146 517556 494152 517568
rect 494204 517556 494210 517608
rect 450354 517488 450360 517540
rect 450412 517528 450418 517540
rect 494054 517528 494060 517540
rect 450412 517500 494060 517528
rect 450412 517488 450418 517500
rect 494054 517488 494060 517500
rect 494112 517488 494118 517540
rect 482278 517420 482284 517472
rect 482336 517420 482342 517472
rect 450630 516808 450636 516860
rect 450688 516848 450694 516860
rect 476022 516848 476028 516860
rect 450688 516820 476028 516848
rect 450688 516808 450694 516820
rect 476022 516808 476028 516820
rect 476080 516808 476086 516860
rect 449986 516740 449992 516792
rect 450044 516780 450050 516792
rect 482296 516780 482324 517420
rect 492122 516780 492128 516792
rect 450044 516752 492128 516780
rect 450044 516740 450050 516752
rect 492122 516740 492128 516752
rect 492180 516740 492186 516792
rect 3970 514768 3976 514820
rect 4028 514808 4034 514820
rect 4798 514808 4804 514820
rect 4028 514780 4804 514808
rect 4028 514768 4034 514780
rect 4798 514768 4804 514780
rect 4856 514768 4862 514820
rect 502242 514020 502248 514072
rect 502300 514060 502306 514072
rect 545114 514060 545120 514072
rect 502300 514032 545120 514060
rect 502300 514020 502306 514032
rect 545114 514020 545120 514032
rect 545172 514020 545178 514072
rect 361758 513340 361764 513392
rect 361816 513380 361822 513392
rect 410518 513380 410524 513392
rect 361816 513352 410524 513380
rect 361816 513340 361822 513352
rect 410518 513340 410524 513352
rect 410576 513340 410582 513392
rect 492122 512592 492128 512644
rect 492180 512632 492186 512644
rect 535454 512632 535460 512644
rect 492180 512604 535460 512632
rect 492180 512592 492186 512604
rect 535454 512592 535460 512604
rect 535512 512592 535518 512644
rect 494054 509872 494060 509924
rect 494112 509912 494118 509924
rect 538214 509912 538220 509924
rect 494112 509884 538220 509912
rect 494112 509872 494118 509884
rect 538214 509872 538220 509884
rect 538272 509872 538278 509924
rect 494146 508512 494152 508564
rect 494204 508552 494210 508564
rect 532694 508552 532700 508564
rect 494204 508524 532700 508552
rect 494204 508512 494210 508524
rect 532694 508512 532700 508524
rect 532752 508512 532758 508564
rect 378870 508444 378876 508496
rect 378928 508484 378934 508496
rect 381262 508484 381268 508496
rect 378928 508456 381268 508484
rect 378928 508444 378934 508456
rect 381262 508444 381268 508456
rect 381320 508444 381326 508496
rect 495066 505724 495072 505776
rect 495124 505764 495130 505776
rect 529934 505764 529940 505776
rect 495124 505736 529940 505764
rect 495124 505724 495130 505736
rect 529934 505724 529940 505736
rect 529992 505724 529998 505776
rect 361758 502324 361764 502376
rect 361816 502364 361822 502376
rect 411898 502364 411904 502376
rect 361816 502336 411904 502364
rect 361816 502324 361822 502336
rect 411898 502324 411904 502336
rect 411956 502324 411962 502376
rect 381262 501576 381268 501628
rect 381320 501616 381326 501628
rect 387334 501616 387340 501628
rect 381320 501588 387340 501616
rect 381320 501576 381326 501588
rect 387334 501576 387340 501588
rect 387392 501576 387398 501628
rect 387334 498108 387340 498160
rect 387392 498148 387398 498160
rect 393958 498148 393964 498160
rect 387392 498120 393964 498148
rect 387392 498108 387398 498120
rect 393958 498108 393964 498120
rect 394016 498108 394022 498160
rect 468662 497768 468668 497820
rect 468720 497808 468726 497820
rect 483842 497808 483848 497820
rect 468720 497780 483848 497808
rect 468720 497768 468726 497780
rect 483842 497768 483848 497780
rect 483900 497768 483906 497820
rect 464430 497700 464436 497752
rect 464488 497740 464494 497752
rect 485038 497740 485044 497752
rect 464488 497712 485044 497740
rect 464488 497700 464494 497712
rect 485038 497700 485044 497712
rect 485096 497700 485102 497752
rect 457622 497632 457628 497684
rect 457680 497672 457686 497684
rect 481634 497672 481640 497684
rect 457680 497644 481640 497672
rect 457680 497632 457686 497644
rect 481634 497632 481640 497644
rect 481692 497632 481698 497684
rect 457438 497564 457444 497616
rect 457496 497604 457502 497616
rect 482646 497604 482652 497616
rect 457496 497576 482652 497604
rect 457496 497564 457502 497576
rect 482646 497564 482652 497576
rect 482704 497564 482710 497616
rect 453298 497496 453304 497548
rect 453356 497536 453362 497548
rect 480254 497536 480260 497548
rect 453356 497508 480260 497536
rect 453356 497496 453362 497508
rect 480254 497496 480260 497508
rect 480312 497496 480318 497548
rect 458818 497428 458824 497480
rect 458876 497468 458882 497480
rect 486234 497468 486240 497480
rect 458876 497440 486240 497468
rect 458876 497428 458882 497440
rect 486234 497428 486240 497440
rect 486292 497428 486298 497480
rect 455322 497020 455328 497072
rect 455380 497060 455386 497072
rect 459554 497060 459560 497072
rect 455380 497032 459560 497060
rect 455380 497020 455386 497032
rect 459554 497020 459560 497032
rect 459612 497020 459618 497072
rect 456518 496952 456524 497004
rect 456576 496992 456582 497004
rect 461026 496992 461032 497004
rect 456576 496964 461032 496992
rect 456576 496952 456582 496964
rect 461026 496952 461032 496964
rect 461084 496952 461090 497004
rect 455138 496884 455144 496936
rect 455196 496924 455202 496936
rect 458082 496924 458088 496936
rect 455196 496896 458088 496924
rect 455196 496884 455202 496896
rect 458082 496884 458088 496896
rect 458140 496884 458146 496936
rect 452562 496816 452568 496868
rect 452620 496856 452626 496868
rect 453666 496856 453672 496868
rect 452620 496828 453672 496856
rect 452620 496816 452626 496828
rect 453666 496816 453672 496828
rect 453724 496816 453730 496868
rect 453942 496816 453948 496868
rect 454000 496856 454006 496868
rect 456610 496856 456616 496868
rect 454000 496828 456616 496856
rect 454000 496816 454006 496828
rect 456610 496816 456616 496828
rect 456668 496816 456674 496868
rect 361758 491308 361764 491360
rect 361816 491348 361822 491360
rect 414658 491348 414664 491360
rect 361816 491320 414664 491348
rect 361816 491308 361822 491320
rect 414658 491308 414664 491320
rect 414716 491308 414722 491360
rect 515490 484372 515496 484424
rect 515548 484412 515554 484424
rect 580166 484412 580172 484424
rect 515548 484384 580172 484412
rect 515548 484372 515554 484384
rect 580166 484372 580172 484384
rect 580224 484372 580230 484424
rect 361758 480224 361764 480276
rect 361816 480264 361822 480276
rect 419074 480264 419080 480276
rect 361816 480236 419080 480264
rect 361816 480224 361822 480236
rect 419074 480224 419080 480236
rect 419132 480224 419138 480276
rect 361758 469208 361764 469260
rect 361816 469248 361822 469260
rect 417418 469248 417424 469260
rect 361816 469220 417424 469248
rect 361816 469208 361822 469220
rect 417418 469208 417424 469220
rect 417476 469208 417482 469260
rect 393958 466284 393964 466336
rect 394016 466324 394022 466336
rect 398098 466324 398104 466336
rect 394016 466296 398104 466324
rect 394016 466284 394022 466296
rect 398098 466284 398104 466296
rect 398156 466284 398162 466336
rect 449802 464312 449808 464364
rect 449860 464352 449866 464364
rect 525794 464352 525800 464364
rect 449860 464324 525800 464352
rect 449860 464312 449866 464324
rect 525794 464312 525800 464324
rect 525852 464312 525858 464364
rect 494698 462408 494704 462460
rect 494756 462448 494762 462460
rect 527634 462448 527640 462460
rect 494756 462420 527640 462448
rect 494756 462408 494762 462420
rect 527634 462408 527640 462420
rect 527692 462408 527698 462460
rect 450538 462340 450544 462392
rect 450596 462380 450602 462392
rect 542354 462380 542360 462392
rect 450596 462352 542360 462380
rect 450596 462340 450602 462352
rect 542354 462340 542360 462352
rect 542412 462340 542418 462392
rect 449710 461048 449716 461100
rect 449768 461088 449774 461100
rect 524690 461088 524696 461100
rect 449768 461060 524696 461088
rect 449768 461048 449774 461060
rect 524690 461048 524696 461060
rect 524748 461048 524754 461100
rect 461854 460980 461860 461032
rect 461912 461020 461918 461032
rect 553854 461020 553860 461032
rect 461912 460992 553860 461020
rect 461912 460980 461918 460992
rect 553854 460980 553860 460992
rect 553912 460980 553918 461032
rect 458910 460912 458916 460964
rect 458968 460952 458974 460964
rect 550910 460952 550916 460964
rect 458968 460924 550916 460952
rect 458968 460912 458974 460924
rect 550910 460912 550916 460924
rect 550968 460912 550974 460964
rect 361758 458192 361764 458244
rect 361816 458232 361822 458244
rect 385770 458232 385776 458244
rect 361816 458204 385776 458232
rect 361816 458192 361822 458204
rect 385770 458192 385776 458204
rect 385828 458192 385834 458244
rect 576118 456764 576124 456816
rect 576176 456804 576182 456816
rect 580166 456804 580172 456816
rect 576176 456776 580172 456804
rect 576176 456764 576182 456776
rect 580166 456764 580172 456776
rect 580224 456764 580230 456816
rect 488258 456016 488264 456068
rect 488316 456056 488322 456068
rect 494698 456056 494704 456068
rect 488316 456028 494704 456056
rect 488316 456016 488322 456028
rect 494698 456016 494704 456028
rect 494756 456016 494762 456068
rect 460198 455472 460204 455524
rect 460256 455512 460262 455524
rect 488258 455512 488264 455524
rect 460256 455484 488264 455512
rect 460256 455472 460262 455484
rect 488258 455472 488264 455484
rect 488316 455472 488322 455524
rect 452010 455404 452016 455456
rect 452068 455444 452074 455456
rect 480990 455444 480996 455456
rect 452068 455416 480996 455444
rect 452068 455404 452074 455416
rect 480990 455404 480996 455416
rect 481048 455404 481054 455456
rect 449618 454724 449624 454776
rect 449676 454764 449682 454776
rect 487154 454764 487160 454776
rect 449676 454736 487160 454764
rect 449676 454724 449682 454736
rect 487154 454724 487160 454736
rect 487212 454724 487218 454776
rect 449526 454656 449532 454708
rect 449584 454696 449590 454708
rect 489914 454696 489920 454708
rect 449584 454668 489920 454696
rect 449584 454656 449590 454668
rect 489914 454656 489920 454668
rect 489972 454656 489978 454708
rect 461946 454044 461952 454096
rect 462004 454084 462010 454096
rect 473722 454084 473728 454096
rect 462004 454056 473728 454084
rect 462004 454044 462010 454056
rect 473722 454044 473728 454056
rect 473780 454044 473786 454096
rect 447318 447924 447324 447976
rect 447376 447964 447382 447976
rect 458910 447964 458916 447976
rect 447376 447936 458916 447964
rect 447376 447924 447382 447936
rect 458910 447924 458916 447936
rect 458968 447924 458974 447976
rect 447226 447856 447232 447908
rect 447284 447896 447290 447908
rect 448422 447896 448428 447908
rect 447284 447868 448428 447896
rect 447284 447856 447290 447868
rect 448422 447856 448428 447868
rect 448480 447896 448486 447908
rect 461946 447896 461952 447908
rect 448480 447868 461952 447896
rect 448480 447856 448486 447868
rect 461946 447856 461952 447868
rect 462004 447856 462010 447908
rect 447134 447788 447140 447840
rect 447192 447828 447198 447840
rect 448054 447828 448060 447840
rect 447192 447800 448060 447828
rect 447192 447788 447198 447800
rect 448054 447788 448060 447800
rect 448112 447828 448118 447840
rect 461854 447828 461860 447840
rect 448112 447800 461860 447828
rect 448112 447788 448118 447800
rect 461854 447788 461860 447800
rect 461912 447788 461918 447840
rect 422478 447312 422484 447364
rect 422536 447352 422542 447364
rect 447226 447352 447232 447364
rect 422536 447324 447232 447352
rect 422536 447312 422542 447324
rect 447226 447312 447232 447324
rect 447284 447312 447290 447364
rect 437382 447244 437388 447296
rect 437440 447284 437446 447296
rect 447134 447284 447140 447296
rect 437440 447256 447140 447284
rect 437440 447244 437446 447256
rect 447134 447244 447140 447256
rect 447192 447244 447198 447296
rect 432414 447176 432420 447228
rect 432472 447216 432478 447228
rect 447318 447216 447324 447228
rect 432472 447188 447324 447216
rect 432472 447176 432478 447188
rect 447318 447176 447324 447188
rect 447376 447216 447382 447228
rect 447962 447216 447968 447228
rect 447376 447188 447968 447216
rect 447376 447176 447382 447188
rect 447962 447176 447968 447188
rect 448020 447176 448026 447228
rect 427722 444388 427728 444440
rect 427780 444428 427786 444440
rect 446306 444428 446312 444440
rect 427780 444400 446312 444428
rect 427780 444388 427786 444400
rect 446306 444388 446312 444400
rect 446364 444388 446370 444440
rect 442626 444320 442632 444372
rect 442684 444360 442690 444372
rect 446214 444360 446220 444372
rect 442684 444332 446220 444360
rect 442684 444320 442690 444332
rect 446214 444320 446220 444332
rect 446272 444320 446278 444372
rect 361758 436092 361764 436144
rect 361816 436132 361822 436144
rect 419166 436132 419172 436144
rect 361816 436104 419172 436132
rect 361816 436092 361822 436104
rect 419166 436092 419172 436104
rect 419224 436092 419230 436144
rect 569310 430584 569316 430636
rect 569368 430624 569374 430636
rect 580166 430624 580172 430636
rect 569368 430596 580172 430624
rect 569368 430584 569374 430596
rect 580166 430584 580172 430596
rect 580224 430584 580230 430636
rect 458082 429904 458088 429956
rect 458140 429944 458146 429956
rect 474274 429944 474280 429956
rect 458140 429916 474280 429944
rect 458140 429904 458146 429916
rect 474274 429904 474280 429916
rect 474332 429904 474338 429956
rect 459462 429836 459468 429888
rect 459520 429876 459526 429888
rect 479610 429876 479616 429888
rect 459520 429848 479616 429876
rect 459520 429836 459526 429848
rect 479610 429836 479616 429848
rect 479668 429836 479674 429888
rect 475378 429156 475384 429208
rect 475436 429196 475442 429208
rect 476942 429196 476948 429208
rect 475436 429168 476948 429196
rect 475436 429156 475442 429168
rect 476942 429156 476948 429168
rect 477000 429156 477006 429208
rect 457530 427048 457536 427100
rect 457588 427088 457594 427100
rect 471606 427088 471612 427100
rect 457588 427060 471612 427088
rect 457588 427048 457594 427060
rect 471606 427048 471612 427060
rect 471664 427048 471670 427100
rect 503622 424328 503628 424380
rect 503680 424368 503686 424380
rect 557534 424368 557540 424380
rect 503680 424340 557540 424368
rect 503680 424328 503686 424340
rect 557534 424328 557540 424340
rect 557592 424328 557598 424380
rect 529198 423580 529204 423632
rect 529256 423620 529262 423632
rect 530210 423620 530216 423632
rect 529256 423592 530216 423620
rect 529256 423580 529262 423592
rect 530210 423580 530216 423592
rect 530268 423580 530274 423632
rect 530578 423580 530584 423632
rect 530636 423620 530642 423632
rect 532786 423620 532792 423632
rect 530636 423592 532792 423620
rect 530636 423580 530642 423592
rect 532786 423580 532792 423592
rect 532844 423580 532850 423632
rect 502978 423512 502984 423564
rect 503036 423552 503042 423564
rect 523770 423552 523776 423564
rect 503036 423524 523776 423552
rect 503036 423512 503042 423524
rect 523770 423512 523776 423524
rect 523828 423512 523834 423564
rect 522298 423444 522304 423496
rect 522356 423484 522362 423496
rect 549530 423484 549536 423496
rect 522356 423456 549536 423484
rect 522356 423444 522362 423456
rect 549530 423444 549536 423456
rect 549588 423444 549594 423496
rect 484302 423376 484308 423428
rect 484360 423416 484366 423428
rect 522482 423416 522488 423428
rect 484360 423388 522488 423416
rect 484360 423376 484366 423388
rect 522482 423376 522488 423388
rect 522540 423376 522546 423428
rect 523678 423376 523684 423428
rect 523736 423416 523742 423428
rect 552106 423416 552112 423428
rect 523736 423388 552112 423416
rect 523736 423376 523742 423388
rect 552106 423376 552112 423388
rect 552164 423376 552170 423428
rect 487062 423308 487068 423360
rect 487120 423348 487126 423360
rect 526346 423348 526352 423360
rect 487120 423320 526352 423348
rect 487120 423308 487126 423320
rect 526346 423308 526352 423320
rect 526404 423308 526410 423360
rect 526438 423308 526444 423360
rect 526496 423348 526502 423360
rect 554682 423348 554688 423360
rect 526496 423320 554688 423348
rect 526496 423308 526502 423320
rect 554682 423308 554688 423320
rect 554740 423308 554746 423360
rect 488258 423240 488264 423292
rect 488316 423280 488322 423292
rect 528922 423280 528928 423292
rect 488316 423252 528928 423280
rect 488316 423240 488322 423252
rect 528922 423240 528928 423252
rect 528980 423240 528986 423292
rect 489638 423172 489644 423224
rect 489696 423212 489702 423224
rect 531498 423212 531504 423224
rect 489696 423184 531504 423212
rect 489696 423172 489702 423184
rect 531498 423172 531504 423184
rect 531556 423172 531562 423224
rect 498102 423104 498108 423156
rect 498160 423144 498166 423156
rect 545666 423144 545672 423156
rect 498160 423116 545672 423144
rect 498160 423104 498166 423116
rect 545666 423104 545672 423116
rect 545724 423104 545730 423156
rect 499298 423036 499304 423088
rect 499356 423076 499362 423088
rect 548242 423076 548248 423088
rect 499356 423048 548248 423076
rect 499356 423036 499362 423048
rect 548242 423036 548248 423048
rect 548300 423036 548306 423088
rect 444282 422968 444288 423020
rect 444340 423008 444346 423020
rect 447870 423008 447876 423020
rect 444340 422980 447876 423008
rect 444340 422968 444346 422980
rect 447870 422968 447876 422980
rect 447928 422968 447934 423020
rect 500678 422968 500684 423020
rect 500736 423008 500742 423020
rect 550818 423008 550824 423020
rect 500736 422980 550824 423008
rect 500736 422968 500742 422980
rect 550818 422968 550824 422980
rect 550876 422968 550882 423020
rect 502242 422900 502248 422952
rect 502300 422940 502306 422952
rect 553394 422940 553400 422952
rect 502300 422912 553400 422940
rect 502300 422900 502306 422912
rect 553394 422900 553400 422912
rect 553452 422900 553458 422952
rect 484210 421540 484216 421592
rect 484268 421580 484274 421592
rect 521194 421580 521200 421592
rect 484268 421552 521200 421580
rect 484268 421540 484274 421552
rect 521194 421540 521200 421552
rect 521252 421540 521258 421592
rect 533430 421540 533436 421592
rect 533488 421580 533494 421592
rect 580350 421580 580356 421592
rect 533488 421552 580356 421580
rect 533488 421540 533494 421552
rect 580350 421540 580356 421552
rect 580408 421540 580414 421592
rect 495342 420180 495348 420232
rect 495400 420220 495406 420232
rect 541802 420220 541808 420232
rect 495400 420192 541808 420220
rect 495400 420180 495406 420192
rect 541802 420180 541808 420192
rect 541860 420180 541866 420232
rect 362310 418752 362316 418804
rect 362368 418792 362374 418804
rect 442258 418792 442264 418804
rect 362368 418764 442264 418792
rect 362368 418752 362374 418764
rect 442258 418752 442264 418764
rect 442316 418752 442322 418804
rect 425330 417732 425336 417784
rect 425388 417772 425394 417784
rect 507854 417772 507860 417784
rect 425388 417744 507860 417772
rect 425388 417732 425394 417744
rect 507854 417732 507860 417744
rect 507912 417732 507918 417784
rect 424686 417664 424692 417716
rect 424744 417704 424750 417716
rect 506474 417704 506480 417716
rect 424744 417676 506480 417704
rect 424744 417664 424750 417676
rect 506474 417664 506480 417676
rect 506532 417664 506538 417716
rect 422110 417596 422116 417648
rect 422168 417636 422174 417648
rect 503990 417636 503996 417648
rect 422168 417608 503996 417636
rect 422168 417596 422174 417608
rect 503990 417596 503996 417608
rect 504048 417596 504054 417648
rect 421466 417528 421472 417580
rect 421524 417568 421530 417580
rect 503714 417568 503720 417580
rect 421524 417540 503720 417568
rect 421524 417528 421530 417540
rect 503714 417528 503720 417540
rect 503772 417528 503778 417580
rect 424042 417460 424048 417512
rect 424100 417500 424106 417512
rect 506566 417500 506572 417512
rect 424100 417472 506572 417500
rect 424100 417460 424106 417472
rect 506566 417460 506572 417472
rect 506624 417460 506630 417512
rect 425974 417392 425980 417444
rect 426032 417432 426038 417444
rect 507946 417432 507952 417444
rect 426032 417404 507952 417432
rect 426032 417392 426038 417404
rect 507946 417392 507952 417404
rect 508004 417392 508010 417444
rect 398098 416100 398104 416152
rect 398156 416140 398162 416152
rect 409138 416140 409144 416152
rect 398156 416112 409144 416140
rect 398156 416100 398162 416112
rect 409138 416100 409144 416112
rect 409196 416100 409202 416152
rect 362218 416032 362224 416084
rect 362276 416072 362282 416084
rect 436738 416072 436744 416084
rect 362276 416044 436744 416072
rect 362276 416032 362282 416044
rect 436738 416032 436744 416044
rect 436796 416032 436802 416084
rect 486970 416032 486976 416084
rect 487028 416072 487034 416084
rect 527634 416072 527640 416084
rect 487028 416044 527640 416072
rect 487028 416032 487034 416044
rect 527634 416032 527640 416044
rect 527692 416032 527698 416084
rect 423122 415964 423128 416016
rect 423180 416004 423186 416016
rect 423582 416004 423588 416016
rect 423180 415976 423588 416004
rect 423180 415964 423186 415976
rect 423582 415964 423588 415976
rect 423640 415964 423646 416016
rect 361574 413992 361580 414044
rect 361632 414032 361638 414044
rect 443638 414032 443644 414044
rect 361632 414004 443644 414032
rect 361632 413992 361638 414004
rect 443638 413992 443644 414004
rect 443696 413992 443702 414044
rect 511258 404336 511264 404388
rect 511316 404376 511322 404388
rect 580166 404376 580172 404388
rect 511316 404348 580172 404376
rect 511316 404336 511322 404348
rect 580166 404336 580172 404348
rect 580224 404336 580230 404388
rect 361574 402976 361580 403028
rect 361632 403016 361638 403028
rect 439498 403016 439504 403028
rect 361632 402988 439504 403016
rect 361632 402976 361638 402988
rect 439498 402976 439504 402988
rect 439556 402976 439562 403028
rect 497918 400868 497924 400920
rect 497976 400908 497982 400920
rect 546494 400908 546500 400920
rect 497976 400880 546500 400908
rect 497976 400868 497982 400880
rect 546494 400868 546500 400880
rect 546552 400868 546558 400920
rect 496722 399440 496728 399492
rect 496780 399480 496786 399492
rect 543734 399480 543740 399492
rect 496780 399452 543740 399480
rect 496780 399440 496786 399452
rect 543734 399440 543740 399452
rect 543792 399440 543798 399492
rect 494606 398080 494612 398132
rect 494664 398120 494670 398132
rect 539594 398120 539600 398132
rect 494664 398092 539600 398120
rect 494664 398080 494670 398092
rect 539594 398080 539600 398092
rect 539652 398080 539658 398132
rect 493962 396720 493968 396772
rect 494020 396760 494026 396772
rect 538214 396760 538220 396772
rect 494020 396732 538220 396760
rect 494020 396720 494026 396732
rect 538214 396720 538220 396732
rect 538272 396720 538278 396772
rect 462222 395292 462228 395344
rect 462280 395332 462286 395344
rect 489914 395332 489920 395344
rect 462280 395304 489920 395332
rect 462280 395292 462286 395304
rect 489914 395292 489920 395304
rect 489972 395292 489978 395344
rect 493134 395292 493140 395344
rect 493192 395332 493198 395344
rect 536834 395332 536840 395344
rect 493192 395304 536840 395332
rect 493192 395292 493198 395304
rect 536834 395292 536840 395304
rect 536892 395292 536898 395344
rect 462590 393932 462596 393984
rect 462648 393972 462654 393984
rect 484394 393972 484400 393984
rect 462648 393944 484400 393972
rect 462648 393932 462654 393944
rect 484394 393932 484400 393944
rect 484452 393932 484458 393984
rect 491662 393932 491668 393984
rect 491720 393972 491726 393984
rect 534166 393972 534172 393984
rect 491720 393944 534172 393972
rect 491720 393932 491726 393944
rect 534166 393932 534172 393944
rect 534224 393932 534230 393984
rect 458174 392708 458180 392760
rect 458232 392748 458238 392760
rect 475378 392748 475384 392760
rect 458232 392720 475384 392748
rect 458232 392708 458238 392720
rect 475378 392708 475384 392720
rect 475436 392708 475442 392760
rect 448238 392640 448244 392692
rect 448296 392680 448302 392692
rect 464430 392680 464436 392692
rect 448296 392652 464436 392680
rect 448296 392640 448302 392652
rect 464430 392640 464436 392652
rect 464488 392640 464494 392692
rect 461118 392572 461124 392624
rect 461176 392612 461182 392624
rect 487154 392612 487160 392624
rect 461176 392584 487160 392612
rect 461176 392572 461182 392584
rect 487154 392572 487160 392584
rect 487212 392572 487218 392624
rect 490558 392572 490564 392624
rect 490616 392612 490622 392624
rect 534074 392612 534080 392624
rect 490616 392584 534080 392612
rect 490616 392572 490622 392584
rect 534074 392572 534080 392584
rect 534132 392572 534138 392624
rect 361574 391960 361580 392012
rect 361632 392000 361638 392012
rect 443730 392000 443736 392012
rect 361632 391972 443736 392000
rect 361632 391960 361638 391972
rect 443730 391960 443736 391972
rect 443788 391960 443794 392012
rect 495710 391280 495716 391332
rect 495768 391320 495774 391332
rect 542354 391320 542360 391332
rect 495768 391292 542360 391320
rect 495768 391280 495774 391292
rect 542354 391280 542360 391292
rect 542412 391280 542418 391332
rect 423490 391212 423496 391264
rect 423548 391252 423554 391264
rect 506014 391252 506020 391264
rect 423548 391224 506020 391252
rect 423548 391212 423554 391224
rect 506014 391212 506020 391224
rect 506072 391212 506078 391264
rect 462774 389852 462780 389904
rect 462832 389892 462838 389904
rect 481634 389892 481640 389904
rect 462832 389864 481640 389892
rect 462832 389852 462838 389864
rect 481634 389852 481640 389864
rect 481692 389852 481698 389904
rect 492030 389852 492036 389904
rect 492088 389892 492094 389904
rect 535454 389892 535460 389904
rect 492088 389864 535460 389892
rect 492088 389852 492094 389864
rect 535454 389852 535460 389864
rect 535512 389852 535518 389904
rect 423582 389784 423588 389836
rect 423640 389824 423646 389836
rect 505278 389824 505284 389836
rect 423640 389796 505284 389824
rect 423640 389784 423646 389796
rect 505278 389784 505284 389796
rect 505336 389784 505342 389836
rect 463694 389240 463700 389292
rect 463752 389280 463758 389292
rect 464430 389280 464436 389292
rect 463752 389252 464436 389280
rect 463752 389240 463758 389252
rect 464430 389240 464436 389252
rect 464488 389240 464494 389292
rect 466454 389240 466460 389292
rect 466512 389280 466518 389292
rect 467374 389280 467380 389292
rect 466512 389252 467380 389280
rect 466512 389240 466518 389252
rect 467374 389240 467380 389252
rect 467432 389240 467438 389292
rect 486418 389240 486424 389292
rect 486476 389280 486482 389292
rect 487062 389280 487068 389292
rect 486476 389252 487068 389280
rect 486476 389240 486482 389252
rect 487062 389240 487068 389252
rect 487120 389240 487126 389292
rect 497458 389240 497464 389292
rect 497516 389280 497522 389292
rect 498102 389280 498108 389292
rect 497516 389252 498108 389280
rect 497516 389240 497522 389252
rect 498102 389240 498108 389252
rect 498160 389240 498166 389292
rect 506474 389240 506480 389292
rect 506532 389280 506538 389292
rect 507118 389280 507124 389292
rect 506532 389252 507124 389280
rect 506532 389240 506538 389252
rect 507118 389240 507124 389252
rect 507176 389240 507182 389292
rect 453022 389104 453028 389156
rect 453080 389144 453086 389156
rect 454034 389144 454040 389156
rect 453080 389116 454040 389144
rect 453080 389104 453086 389116
rect 454034 389104 454040 389116
rect 454092 389104 454098 389156
rect 456702 389104 456708 389156
rect 456760 389144 456766 389156
rect 457530 389144 457536 389156
rect 456760 389116 457536 389144
rect 456760 389104 456766 389116
rect 457530 389104 457536 389116
rect 457588 389104 457594 389156
rect 460382 389104 460388 389156
rect 460440 389144 460446 389156
rect 462590 389144 462596 389156
rect 460440 389116 462596 389144
rect 460440 389104 460446 389116
rect 462590 389104 462596 389116
rect 462648 389104 462654 389156
rect 469950 388968 469956 389020
rect 470008 389008 470014 389020
rect 473630 389008 473636 389020
rect 470008 388980 473636 389008
rect 470008 388968 470014 388980
rect 473630 388968 473636 388980
rect 473688 388968 473694 389020
rect 465810 388900 465816 388952
rect 465868 388940 465874 388952
rect 469398 388940 469404 388952
rect 465868 388912 469404 388940
rect 465868 388900 465874 388912
rect 469398 388900 469404 388912
rect 469456 388900 469462 388952
rect 469858 388900 469864 388952
rect 469916 388940 469922 388952
rect 475838 388940 475844 388952
rect 469916 388912 475844 388940
rect 469916 388900 469922 388912
rect 475838 388900 475844 388912
rect 475896 388900 475902 388952
rect 502334 388900 502340 388952
rect 502392 388940 502398 388952
rect 502392 388912 509234 388940
rect 502392 388900 502398 388912
rect 468478 388832 468484 388884
rect 468536 388872 468542 388884
rect 476574 388872 476580 388884
rect 468536 388844 476580 388872
rect 468536 388832 468542 388844
rect 476574 388832 476580 388844
rect 476632 388832 476638 388884
rect 468570 388764 468576 388816
rect 468628 388804 468634 388816
rect 480254 388804 480260 388816
rect 468628 388776 480260 388804
rect 468628 388764 468634 388776
rect 480254 388764 480260 388776
rect 480312 388764 480318 388816
rect 484670 388764 484676 388816
rect 484728 388804 484734 388816
rect 502978 388804 502984 388816
rect 484728 388776 502984 388804
rect 484728 388764 484734 388776
rect 502978 388764 502984 388776
rect 503036 388764 503042 388816
rect 509206 388804 509234 388912
rect 526438 388804 526444 388816
rect 509206 388776 526444 388804
rect 526438 388764 526444 388776
rect 526496 388764 526502 388816
rect 467098 388696 467104 388748
rect 467156 388736 467162 388748
rect 467156 388708 469352 388736
rect 467156 388696 467162 388708
rect 465718 388628 465724 388680
rect 465776 388668 465782 388680
rect 469214 388668 469220 388680
rect 465776 388640 469220 388668
rect 465776 388628 465782 388640
rect 469214 388628 469220 388640
rect 469272 388628 469278 388680
rect 469324 388668 469352 388708
rect 469398 388696 469404 388748
rect 469456 388736 469462 388748
rect 480990 388736 480996 388748
rect 469456 388708 480996 388736
rect 469456 388696 469462 388708
rect 480990 388696 480996 388708
rect 481048 388696 481054 388748
rect 500862 388696 500868 388748
rect 500920 388736 500926 388748
rect 523678 388736 523684 388748
rect 500920 388708 523684 388736
rect 500920 388696 500926 388708
rect 523678 388696 523684 388708
rect 523736 388696 523742 388748
rect 481726 388668 481732 388680
rect 469324 388640 481732 388668
rect 481726 388628 481732 388640
rect 481784 388628 481790 388680
rect 499390 388628 499396 388680
rect 499448 388668 499454 388680
rect 522298 388668 522304 388680
rect 499448 388640 522304 388668
rect 499448 388628 499454 388640
rect 522298 388628 522304 388640
rect 522356 388628 522362 388680
rect 461670 388560 461676 388612
rect 461728 388600 461734 388612
rect 478782 388600 478788 388612
rect 461728 388572 478788 388600
rect 461728 388560 461734 388572
rect 478782 388560 478788 388572
rect 478840 388560 478846 388612
rect 485406 388560 485412 388612
rect 485464 388600 485470 388612
rect 524414 388600 524420 388612
rect 485464 388572 524420 388600
rect 485464 388560 485470 388572
rect 524414 388560 524420 388572
rect 524472 388560 524478 388612
rect 461578 388492 461584 388544
rect 461636 388532 461642 388544
rect 478046 388532 478052 388544
rect 461636 388504 478052 388532
rect 461636 388492 461642 388504
rect 478046 388492 478052 388504
rect 478104 388492 478110 388544
rect 489822 388492 489828 388544
rect 489880 388532 489886 388544
rect 530578 388532 530584 388544
rect 489880 388504 530584 388532
rect 489880 388492 489886 388504
rect 530578 388492 530584 388504
rect 530636 388492 530642 388544
rect 447410 388424 447416 388476
rect 447468 388464 447474 388476
rect 458818 388464 458824 388476
rect 447468 388436 458824 388464
rect 447468 388424 447474 388436
rect 458818 388424 458824 388436
rect 458876 388424 458882 388476
rect 461762 388424 461768 388476
rect 461820 388464 461826 388476
rect 482462 388464 482468 388476
rect 461820 388436 482468 388464
rect 461820 388424 461826 388436
rect 482462 388424 482468 388436
rect 482520 388424 482526 388476
rect 488350 388424 488356 388476
rect 488408 388464 488414 388476
rect 529198 388464 529204 388476
rect 488408 388436 529204 388464
rect 488408 388424 488414 388436
rect 529198 388424 529204 388436
rect 529256 388424 529262 388476
rect 462958 388356 462964 388408
rect 463016 388396 463022 388408
rect 469950 388396 469956 388408
rect 463016 388368 469956 388396
rect 463016 388356 463022 388368
rect 469950 388356 469956 388368
rect 470008 388356 470014 388408
rect 459646 388152 459652 388204
rect 459704 388192 459710 388204
rect 462774 388192 462780 388204
rect 459704 388164 462780 388192
rect 459704 388152 459710 388164
rect 462774 388152 462780 388164
rect 462832 388152 462838 388204
rect 450722 387336 450728 387388
rect 450780 387376 450786 387388
rect 460198 387376 460204 387388
rect 450780 387348 460204 387376
rect 450780 387336 450786 387348
rect 460198 387336 460204 387348
rect 460256 387336 460262 387388
rect 447594 387268 447600 387320
rect 447652 387308 447658 387320
rect 457438 387308 457444 387320
rect 447652 387280 457444 387308
rect 447652 387268 447658 387280
rect 457438 387268 457444 387280
rect 457496 387268 457502 387320
rect 447686 387200 447692 387252
rect 447744 387240 447750 387252
rect 468662 387240 468668 387252
rect 447744 387212 468668 387240
rect 447744 387200 447750 387212
rect 468662 387200 468668 387212
rect 468720 387200 468726 387252
rect 448974 387132 448980 387184
rect 449032 387172 449038 387184
rect 491294 387172 491300 387184
rect 449032 387144 491300 387172
rect 449032 387132 449038 387144
rect 491294 387132 491300 387144
rect 491352 387132 491358 387184
rect 441522 387064 441528 387116
rect 441580 387104 441586 387116
rect 447778 387104 447784 387116
rect 441580 387076 447784 387104
rect 441580 387064 441586 387076
rect 447778 387064 447784 387076
rect 447836 387064 447842 387116
rect 449434 387064 449440 387116
rect 449492 387104 449498 387116
rect 513374 387104 513380 387116
rect 449492 387076 513380 387104
rect 449492 387064 449498 387076
rect 513374 387064 513380 387076
rect 513432 387064 513438 387116
rect 448422 386588 448428 386640
rect 448480 386628 448486 386640
rect 553946 386628 553952 386640
rect 448480 386600 553952 386628
rect 448480 386588 448486 386600
rect 553946 386588 553952 386600
rect 554004 386588 554010 386640
rect 385678 386520 385684 386572
rect 385736 386560 385742 386572
rect 512086 386560 512092 386572
rect 385736 386532 512092 386560
rect 385736 386520 385742 386532
rect 512086 386520 512092 386532
rect 512144 386520 512150 386572
rect 380158 386452 380164 386504
rect 380216 386492 380222 386504
rect 512270 386492 512276 386504
rect 380216 386464 512276 386492
rect 380216 386452 380222 386464
rect 512270 386452 512276 386464
rect 512328 386452 512334 386504
rect 373258 386384 373264 386436
rect 373316 386424 373322 386436
rect 511994 386424 512000 386436
rect 373316 386396 512000 386424
rect 373316 386384 373322 386396
rect 511994 386384 512000 386396
rect 512052 386384 512058 386436
rect 448146 385976 448152 386028
rect 448204 386016 448210 386028
rect 453298 386016 453304 386028
rect 448204 385988 453304 386016
rect 448204 385976 448210 385988
rect 453298 385976 453304 385988
rect 453356 385976 453362 386028
rect 447870 385636 447876 385688
rect 447928 385676 447934 385688
rect 457346 385676 457352 385688
rect 447928 385648 457352 385676
rect 447928 385636 447934 385648
rect 457346 385636 457352 385648
rect 457404 385636 457410 385688
rect 448330 385500 448336 385552
rect 448388 385540 448394 385552
rect 452010 385540 452016 385552
rect 448388 385512 452016 385540
rect 448388 385500 448394 385512
rect 452010 385500 452016 385512
rect 452068 385500 452074 385552
rect 449342 385432 449348 385484
rect 449400 385472 449406 385484
rect 563422 385472 563428 385484
rect 449400 385444 563428 385472
rect 449400 385432 449406 385444
rect 563422 385432 563428 385444
rect 563480 385432 563486 385484
rect 377398 385364 377404 385416
rect 377456 385404 377462 385416
rect 512178 385404 512184 385416
rect 377456 385376 512184 385404
rect 377456 385364 377462 385376
rect 512178 385364 512184 385376
rect 512236 385364 512242 385416
rect 387058 384956 387064 385008
rect 387116 384996 387122 385008
rect 447134 384996 447140 385008
rect 387116 384968 447140 384996
rect 387116 384956 387122 384968
rect 447134 384956 447140 384968
rect 447192 384956 447198 385008
rect 513282 383732 513288 383784
rect 513340 383772 513346 383784
rect 534718 383772 534724 383784
rect 513340 383744 534724 383772
rect 513340 383732 513346 383744
rect 534718 383732 534724 383744
rect 534776 383732 534782 383784
rect 512454 383664 512460 383716
rect 512512 383704 512518 383716
rect 548518 383704 548524 383716
rect 512512 383676 548524 383704
rect 512512 383664 512518 383676
rect 548518 383664 548524 383676
rect 548576 383664 548582 383716
rect 381538 383596 381544 383648
rect 381596 383636 381602 383648
rect 447226 383636 447232 383648
rect 381596 383608 447232 383636
rect 381596 383596 381602 383608
rect 447226 383596 447232 383608
rect 447284 383596 447290 383648
rect 382918 383528 382924 383580
rect 382976 383568 382982 383580
rect 447134 383568 447140 383580
rect 382976 383540 447140 383568
rect 382976 383528 382982 383540
rect 447134 383528 447140 383540
rect 447192 383528 447198 383580
rect 512638 382984 512644 383036
rect 512696 383024 512702 383036
rect 519722 383024 519728 383036
rect 512696 382996 519728 383024
rect 512696 382984 512702 382996
rect 519722 382984 519728 382996
rect 519780 382984 519786 383036
rect 513006 382916 513012 382968
rect 513064 382956 513070 382968
rect 518250 382956 518256 382968
rect 513064 382928 518256 382956
rect 513064 382916 513070 382928
rect 518250 382916 518256 382928
rect 518308 382916 518314 382968
rect 512454 382440 512460 382492
rect 512512 382480 512518 382492
rect 515582 382480 515588 382492
rect 512512 382452 515588 382480
rect 512512 382440 512518 382452
rect 515582 382440 515588 382452
rect 515640 382440 515646 382492
rect 378778 382168 378784 382220
rect 378836 382208 378842 382220
rect 447134 382208 447140 382220
rect 378836 382180 447140 382208
rect 378836 382168 378842 382180
rect 447134 382168 447140 382180
rect 447192 382168 447198 382220
rect 403618 382100 403624 382152
rect 403676 382140 403682 382152
rect 447226 382140 447232 382152
rect 403676 382112 447232 382140
rect 403676 382100 403682 382112
rect 447226 382100 447232 382112
rect 447284 382100 447290 382152
rect 361574 380876 361580 380928
rect 361632 380916 361638 380928
rect 443822 380916 443828 380928
rect 361632 380888 443828 380916
rect 361632 380876 361638 380888
rect 443822 380876 443828 380888
rect 443880 380876 443886 380928
rect 513282 380876 513288 380928
rect 513340 380916 513346 380928
rect 547138 380916 547144 380928
rect 513340 380888 547144 380916
rect 513340 380876 513346 380888
rect 547138 380876 547144 380888
rect 547196 380876 547202 380928
rect 376018 380808 376024 380860
rect 376076 380848 376082 380860
rect 447134 380848 447140 380860
rect 376076 380820 447140 380848
rect 376076 380808 376082 380820
rect 447134 380808 447140 380820
rect 447192 380808 447198 380860
rect 406378 380740 406384 380792
rect 406436 380780 406442 380792
rect 447226 380780 447232 380792
rect 406436 380752 447232 380780
rect 406436 380740 406442 380752
rect 447226 380740 447232 380752
rect 447284 380740 447290 380792
rect 512546 379720 512552 379772
rect 512604 379760 512610 379772
rect 515674 379760 515680 379772
rect 512604 379732 515680 379760
rect 512604 379720 512610 379732
rect 515674 379720 515680 379732
rect 515732 379720 515738 379772
rect 513282 379516 513288 379568
rect 513340 379556 513346 379568
rect 549898 379556 549904 379568
rect 513340 379528 549904 379556
rect 513340 379516 513346 379528
rect 549898 379516 549904 379528
rect 549956 379516 549962 379568
rect 374638 379448 374644 379500
rect 374696 379488 374702 379500
rect 447134 379488 447140 379500
rect 374696 379460 447140 379488
rect 374696 379448 374702 379460
rect 447134 379448 447140 379460
rect 447192 379448 447198 379500
rect 407758 379380 407764 379432
rect 407816 379420 407822 379432
rect 447226 379420 447232 379432
rect 407816 379392 447232 379420
rect 407816 379380 407822 379392
rect 447226 379380 447232 379392
rect 447284 379380 447290 379432
rect 512454 378224 512460 378276
rect 512512 378264 512518 378276
rect 522298 378264 522304 378276
rect 512512 378236 522304 378264
rect 512512 378224 512518 378236
rect 522298 378224 522304 378236
rect 522356 378224 522362 378276
rect 512914 378156 512920 378208
rect 512972 378196 512978 378208
rect 547230 378196 547236 378208
rect 512972 378168 547236 378196
rect 512972 378156 512978 378168
rect 547230 378156 547236 378168
rect 547288 378156 547294 378208
rect 363598 378088 363604 378140
rect 363656 378128 363662 378140
rect 447226 378128 447232 378140
rect 363656 378100 447232 378128
rect 363656 378088 363662 378100
rect 447226 378088 447232 378100
rect 447284 378088 447290 378140
rect 371878 378020 371884 378072
rect 371936 378060 371942 378072
rect 447134 378060 447140 378072
rect 371936 378032 447140 378060
rect 371936 378020 371942 378032
rect 447134 378020 447140 378032
rect 447192 378020 447198 378072
rect 513190 377408 513196 377460
rect 513248 377448 513254 377460
rect 548610 377448 548616 377460
rect 513248 377420 548616 377448
rect 513248 377408 513254 377420
rect 548610 377408 548616 377420
rect 548668 377408 548674 377460
rect 512638 376728 512644 376780
rect 512696 376768 512702 376780
rect 516410 376768 516416 376780
rect 512696 376740 516416 376768
rect 512696 376728 512702 376740
rect 516410 376728 516416 376740
rect 516468 376728 516474 376780
rect 367738 376660 367744 376712
rect 367796 376700 367802 376712
rect 447226 376700 447232 376712
rect 367796 376672 447232 376700
rect 367796 376660 367802 376672
rect 447226 376660 447232 376672
rect 447284 376660 447290 376712
rect 370498 376592 370504 376644
rect 370556 376632 370562 376644
rect 447134 376632 447140 376644
rect 370556 376604 447140 376632
rect 370556 376592 370562 376604
rect 447134 376592 447140 376604
rect 447192 376592 447198 376644
rect 513098 375980 513104 376032
rect 513156 376020 513162 376032
rect 544378 376020 544384 376032
rect 513156 375992 544384 376020
rect 513156 375980 513162 375992
rect 544378 375980 544384 375992
rect 544436 375980 544442 376032
rect 512822 375436 512828 375488
rect 512880 375476 512886 375488
rect 516226 375476 516232 375488
rect 512880 375448 516232 375476
rect 512880 375436 512886 375448
rect 516226 375436 516232 375448
rect 516284 375436 516290 375488
rect 512638 375368 512644 375420
rect 512696 375408 512702 375420
rect 520274 375408 520280 375420
rect 512696 375380 520280 375408
rect 512696 375368 512702 375380
rect 520274 375368 520280 375380
rect 520332 375368 520338 375420
rect 363690 375300 363696 375352
rect 363748 375340 363754 375352
rect 447134 375340 447140 375352
rect 363748 375312 447140 375340
rect 363748 375300 363754 375312
rect 447134 375300 447140 375312
rect 447192 375300 447198 375352
rect 363782 375232 363788 375284
rect 363840 375272 363846 375284
rect 447226 375272 447232 375284
rect 363840 375244 447232 375272
rect 363840 375232 363846 375244
rect 447226 375232 447232 375244
rect 447284 375232 447290 375284
rect 513282 374008 513288 374060
rect 513340 374048 513346 374060
rect 520366 374048 520372 374060
rect 513340 374020 520372 374048
rect 513340 374008 513346 374020
rect 520366 374008 520372 374020
rect 520424 374008 520430 374060
rect 410518 373940 410524 373992
rect 410576 373980 410582 373992
rect 447134 373980 447140 373992
rect 410576 373952 447140 373980
rect 410576 373940 410582 373952
rect 447134 373940 447140 373952
rect 447192 373940 447198 373992
rect 411898 373872 411904 373924
rect 411956 373912 411962 373924
rect 447226 373912 447232 373924
rect 411956 373884 447232 373912
rect 411956 373872 411962 373884
rect 447226 373872 447232 373884
rect 447284 373872 447290 373924
rect 512638 373736 512644 373788
rect 512696 373776 512702 373788
rect 516318 373776 516324 373788
rect 512696 373748 516324 373776
rect 512696 373736 512702 373748
rect 516318 373736 516324 373748
rect 516376 373736 516382 373788
rect 512454 372716 512460 372768
rect 512512 372756 512518 372768
rect 523034 372756 523040 372768
rect 512512 372728 523040 372756
rect 512512 372716 512518 372728
rect 523034 372716 523040 372728
rect 523092 372716 523098 372768
rect 512086 372648 512092 372700
rect 512144 372688 512150 372700
rect 514754 372688 514760 372700
rect 512144 372660 514760 372688
rect 512144 372648 512150 372660
rect 514754 372648 514760 372660
rect 514812 372648 514818 372700
rect 414658 372512 414664 372564
rect 414716 372552 414722 372564
rect 447134 372552 447140 372564
rect 414716 372524 447140 372552
rect 414716 372512 414722 372524
rect 447134 372512 447140 372524
rect 447192 372512 447198 372564
rect 419074 372444 419080 372496
rect 419132 372484 419138 372496
rect 447226 372484 447232 372496
rect 419132 372456 447232 372484
rect 419132 372444 419138 372456
rect 447226 372444 447232 372456
rect 447284 372444 447290 372496
rect 512822 371220 512828 371272
rect 512880 371260 512886 371272
rect 517514 371260 517520 371272
rect 512880 371232 517520 371260
rect 512880 371220 512886 371232
rect 517514 371220 517520 371232
rect 517572 371220 517578 371272
rect 385770 371152 385776 371204
rect 385828 371192 385834 371204
rect 447226 371192 447232 371204
rect 385828 371164 447232 371192
rect 385828 371152 385834 371164
rect 447226 371152 447232 371164
rect 447284 371152 447290 371204
rect 417418 371084 417424 371136
rect 417476 371124 417482 371136
rect 447134 371124 447140 371136
rect 417476 371096 447140 371124
rect 417476 371084 417482 371096
rect 447134 371084 447140 371096
rect 447192 371084 447198 371136
rect 512638 369928 512644 369980
rect 512696 369968 512702 369980
rect 516962 369968 516968 369980
rect 512696 369940 516968 369968
rect 512696 369928 512702 369940
rect 516962 369928 516968 369940
rect 517020 369928 517026 369980
rect 361574 369860 361580 369912
rect 361632 369900 361638 369912
rect 409874 369900 409880 369912
rect 361632 369872 409880 369900
rect 361632 369860 361638 369872
rect 409874 369860 409880 369872
rect 409932 369860 409938 369912
rect 513282 369860 513288 369912
rect 513340 369900 513346 369912
rect 521654 369900 521660 369912
rect 513340 369872 521660 369900
rect 513340 369860 513346 369872
rect 521654 369860 521660 369872
rect 521712 369860 521718 369912
rect 419166 369792 419172 369844
rect 419224 369832 419230 369844
rect 447226 369832 447232 369844
rect 419224 369804 447232 369832
rect 419224 369792 419230 369804
rect 447226 369792 447232 369804
rect 447284 369792 447290 369844
rect 436738 369724 436744 369776
rect 436796 369764 436802 369776
rect 447134 369764 447140 369776
rect 436796 369736 447140 369764
rect 436796 369724 436802 369736
rect 447134 369724 447140 369736
rect 447192 369724 447198 369776
rect 513282 368568 513288 368620
rect 513340 368608 513346 368620
rect 520458 368608 520464 368620
rect 513340 368580 520464 368608
rect 513340 368568 513346 368580
rect 520458 368568 520464 368580
rect 520516 368568 520522 368620
rect 512822 368500 512828 368552
rect 512880 368540 512886 368552
rect 516502 368540 516508 368552
rect 512880 368512 516508 368540
rect 512880 368500 512886 368512
rect 516502 368500 516508 368512
rect 516560 368500 516566 368552
rect 443638 368432 443644 368484
rect 443696 368472 443702 368484
rect 447134 368472 447140 368484
rect 443696 368444 447140 368472
rect 443696 368432 443702 368444
rect 447134 368432 447140 368444
rect 447192 368432 447198 368484
rect 442258 368364 442264 368416
rect 442316 368404 442322 368416
rect 447226 368404 447232 368416
rect 442316 368376 447232 368404
rect 442316 368364 442322 368376
rect 447226 368364 447232 368376
rect 447284 368364 447290 368416
rect 511994 367344 512000 367396
rect 512052 367384 512058 367396
rect 514110 367384 514116 367396
rect 512052 367356 514116 367384
rect 512052 367344 512058 367356
rect 514110 367344 514116 367356
rect 514168 367344 514174 367396
rect 513282 367208 513288 367260
rect 513340 367248 513346 367260
rect 517882 367248 517888 367260
rect 513340 367220 517888 367248
rect 513340 367208 513346 367220
rect 517882 367208 517888 367220
rect 517940 367208 517946 367260
rect 439498 367004 439504 367056
rect 439556 367044 439562 367056
rect 447134 367044 447140 367056
rect 439556 367016 447140 367044
rect 439556 367004 439562 367016
rect 447134 367004 447140 367016
rect 447192 367004 447198 367056
rect 443730 366936 443736 366988
rect 443788 366976 443794 366988
rect 447226 366976 447232 366988
rect 443788 366948 447232 366976
rect 443788 366936 443794 366948
rect 447226 366936 447232 366948
rect 447284 366936 447290 366988
rect 511994 366120 512000 366172
rect 512052 366160 512058 366172
rect 514202 366160 514208 366172
rect 512052 366132 514208 366160
rect 512052 366120 512058 366132
rect 514202 366120 514208 366132
rect 514260 366120 514266 366172
rect 513282 365712 513288 365764
rect 513340 365752 513346 365764
rect 523126 365752 523132 365764
rect 513340 365724 523132 365752
rect 513340 365712 513346 365724
rect 523126 365712 523132 365724
rect 523184 365712 523190 365764
rect 409874 365644 409880 365696
rect 409932 365684 409938 365696
rect 447134 365684 447140 365696
rect 409932 365656 447140 365684
rect 409932 365644 409938 365656
rect 447134 365644 447140 365656
rect 447192 365644 447198 365696
rect 443822 365576 443828 365628
rect 443880 365616 443886 365628
rect 447226 365616 447232 365628
rect 443880 365588 447232 365616
rect 443880 365576 443886 365588
rect 447226 365576 447232 365588
rect 447284 365576 447290 365628
rect 513282 364488 513288 364540
rect 513340 364528 513346 364540
rect 520550 364528 520556 364540
rect 513340 364500 520556 364528
rect 513340 364488 513346 364500
rect 520550 364488 520556 364500
rect 520608 364488 520614 364540
rect 512638 364352 512644 364404
rect 512696 364392 512702 364404
rect 521746 364392 521752 364404
rect 512696 364364 521752 364392
rect 512696 364352 512702 364364
rect 521746 364352 521752 364364
rect 521804 364352 521810 364404
rect 569402 364352 569408 364404
rect 569460 364392 569466 364404
rect 580166 364392 580172 364404
rect 569460 364364 580172 364392
rect 569460 364352 569466 364364
rect 580166 364352 580172 364364
rect 580224 364352 580230 364404
rect 409138 363604 409144 363656
rect 409196 363644 409202 363656
rect 416130 363644 416136 363656
rect 409196 363616 416136 363644
rect 409196 363604 409202 363616
rect 416130 363604 416136 363616
rect 416188 363604 416194 363656
rect 512178 363264 512184 363316
rect 512236 363304 512242 363316
rect 514846 363304 514852 363316
rect 512236 363276 514852 363304
rect 512236 363264 512242 363276
rect 514846 363264 514852 363276
rect 514904 363264 514910 363316
rect 432690 362992 432696 363044
rect 432748 363032 432754 363044
rect 447134 363032 447140 363044
rect 432748 363004 447140 363032
rect 432748 362992 432754 363004
rect 447134 362992 447140 363004
rect 447192 362992 447198 363044
rect 432782 362924 432788 362976
rect 432840 362964 432846 362976
rect 447226 362964 447232 362976
rect 432840 362936 447232 362964
rect 432840 362924 432846 362936
rect 447226 362924 447232 362936
rect 447284 362924 447290 362976
rect 513282 362924 513288 362976
rect 513340 362964 513346 362976
rect 523218 362964 523224 362976
rect 513340 362936 523224 362964
rect 513340 362924 513346 362936
rect 523218 362924 523224 362936
rect 523276 362924 523282 362976
rect 512178 362312 512184 362364
rect 512236 362352 512242 362364
rect 513650 362352 513656 362364
rect 512236 362324 513656 362352
rect 512236 362312 512242 362324
rect 513650 362312 513656 362324
rect 513708 362312 513714 362364
rect 443914 361632 443920 361684
rect 443972 361672 443978 361684
rect 447226 361672 447232 361684
rect 443972 361644 447232 361672
rect 443972 361632 443978 361644
rect 447226 361632 447232 361644
rect 447284 361632 447290 361684
rect 513006 361632 513012 361684
rect 513064 361672 513070 361684
rect 517606 361672 517612 361684
rect 513064 361644 517612 361672
rect 513064 361632 513070 361644
rect 517606 361632 517612 361644
rect 517664 361632 517670 361684
rect 432598 361564 432604 361616
rect 432656 361604 432662 361616
rect 447134 361604 447140 361616
rect 432656 361576 447140 361604
rect 432656 361564 432662 361576
rect 447134 361564 447140 361576
rect 447192 361564 447198 361616
rect 442258 360272 442264 360324
rect 442316 360312 442322 360324
rect 447226 360312 447232 360324
rect 442316 360284 447232 360312
rect 442316 360272 442322 360284
rect 447226 360272 447232 360284
rect 447284 360272 447290 360324
rect 513006 360272 513012 360324
rect 513064 360312 513070 360324
rect 517698 360312 517704 360324
rect 513064 360284 517704 360312
rect 513064 360272 513070 360284
rect 517698 360272 517704 360284
rect 517756 360272 517762 360324
rect 436922 360204 436928 360256
rect 436980 360244 436986 360256
rect 447134 360244 447140 360256
rect 436980 360216 447140 360244
rect 436980 360204 436986 360216
rect 447134 360204 447140 360216
rect 447192 360204 447198 360256
rect 513282 360204 513288 360256
rect 513340 360244 513346 360256
rect 518894 360244 518900 360256
rect 513340 360216 518900 360244
rect 513340 360204 513346 360216
rect 518894 360204 518900 360216
rect 518952 360204 518958 360256
rect 547230 360136 547236 360188
rect 547288 360176 547294 360188
rect 552014 360176 552020 360188
rect 547288 360148 552020 360176
rect 547288 360136 547294 360148
rect 552014 360136 552020 360148
rect 552072 360136 552078 360188
rect 534718 360068 534724 360120
rect 534776 360108 534782 360120
rect 566734 360108 566740 360120
rect 534776 360080 566740 360108
rect 534776 360068 534782 360080
rect 566734 360068 566740 360080
rect 566792 360068 566798 360120
rect 549898 360000 549904 360052
rect 549956 360040 549962 360052
rect 554958 360040 554964 360052
rect 549956 360012 554964 360040
rect 549956 360000 549962 360012
rect 554958 360000 554964 360012
rect 555016 360000 555022 360052
rect 548518 359932 548524 359984
rect 548576 359972 548582 359984
rect 565262 359972 565268 359984
rect 548576 359944 565268 359972
rect 548576 359932 548582 359944
rect 565262 359932 565268 359944
rect 565320 359932 565326 359984
rect 547138 359864 547144 359916
rect 547196 359904 547202 359916
rect 558178 359904 558184 359916
rect 547196 359876 558184 359904
rect 547196 359864 547202 359876
rect 558178 359864 558184 359876
rect 558236 359864 558242 359916
rect 515674 359796 515680 359848
rect 515732 359836 515738 359848
rect 553762 359836 553768 359848
rect 515732 359808 553768 359836
rect 515732 359796 515738 359808
rect 553762 359796 553768 359808
rect 553820 359796 553826 359848
rect 522298 359728 522304 359780
rect 522356 359768 522362 359780
rect 550818 359768 550824 359780
rect 522356 359740 550824 359768
rect 522356 359728 522362 359740
rect 550818 359728 550824 359740
rect 550876 359728 550882 359780
rect 443822 358844 443828 358896
rect 443880 358884 443886 358896
rect 447226 358884 447232 358896
rect 443880 358856 447232 358884
rect 443880 358844 443886 358856
rect 447226 358844 447232 358856
rect 447284 358844 447290 358896
rect 435358 358776 435364 358828
rect 435416 358816 435422 358828
rect 447134 358816 447140 358828
rect 435416 358788 447140 358816
rect 435416 358776 435422 358788
rect 447134 358776 447140 358788
rect 447192 358776 447198 358828
rect 548610 358708 548616 358760
rect 548668 358748 548674 358760
rect 556706 358748 556712 358760
rect 548668 358720 556712 358748
rect 548668 358708 548674 358720
rect 556706 358708 556712 358720
rect 556764 358708 556770 358760
rect 518250 358640 518256 358692
rect 518308 358680 518314 358692
rect 562594 358680 562600 358692
rect 518308 358652 562600 358680
rect 518308 358640 518314 358652
rect 562594 358640 562600 358652
rect 562652 358640 562658 358692
rect 519722 358572 519728 358624
rect 519780 358612 519786 358624
rect 564066 358612 564072 358624
rect 519780 358584 564072 358612
rect 519780 358572 519786 358584
rect 564066 358572 564072 358584
rect 564124 358572 564130 358624
rect 544378 358504 544384 358556
rect 544436 358544 544442 358556
rect 559650 358544 559656 358556
rect 544436 358516 559656 358544
rect 544436 358504 544442 358516
rect 559650 358504 559656 358516
rect 559708 358504 559714 358556
rect 515582 358436 515588 358488
rect 515640 358476 515646 358488
rect 561122 358476 561128 358488
rect 515640 358448 561128 358476
rect 515640 358436 515646 358448
rect 561122 358436 561128 358448
rect 561180 358436 561186 358488
rect 512178 357688 512184 357740
rect 512236 357728 512242 357740
rect 514018 357728 514024 357740
rect 512236 357700 514024 357728
rect 512236 357688 512242 357700
rect 514018 357688 514024 357700
rect 514076 357688 514082 357740
rect 512178 357552 512184 357604
rect 512236 357592 512242 357604
rect 512362 357592 512368 357604
rect 512236 357564 512368 357592
rect 512236 357552 512242 357564
rect 512362 357552 512368 357564
rect 512420 357552 512426 357604
rect 513282 356056 513288 356108
rect 513340 356096 513346 356108
rect 521838 356096 521844 356108
rect 513340 356068 521844 356096
rect 513340 356056 513346 356068
rect 521838 356056 521844 356068
rect 521896 356056 521902 356108
rect 513282 354696 513288 354748
rect 513340 354736 513346 354748
rect 517974 354736 517980 354748
rect 513340 354708 517980 354736
rect 513340 354696 513346 354708
rect 517974 354696 517980 354708
rect 518032 354696 518038 354748
rect 512454 353608 512460 353660
rect 512512 353648 512518 353660
rect 513742 353648 513748 353660
rect 512512 353620 513748 353648
rect 512512 353608 512518 353620
rect 513742 353608 513748 353620
rect 513800 353608 513806 353660
rect 513190 353472 513196 353524
rect 513248 353512 513254 353524
rect 517790 353512 517796 353524
rect 513248 353484 517796 353512
rect 513248 353472 513254 353484
rect 517790 353472 517796 353484
rect 517848 353472 517854 353524
rect 446214 352656 446220 352708
rect 446272 352696 446278 352708
rect 447778 352696 447784 352708
rect 446272 352668 447784 352696
rect 446272 352656 446278 352668
rect 447778 352656 447784 352668
rect 447836 352656 447842 352708
rect 512454 352520 512460 352572
rect 512512 352560 512518 352572
rect 515030 352560 515036 352572
rect 512512 352532 515036 352560
rect 512512 352520 512518 352532
rect 515030 352520 515036 352532
rect 515088 352520 515094 352572
rect 511350 352044 511356 352096
rect 511408 352084 511414 352096
rect 580166 352084 580172 352096
rect 511408 352056 580172 352084
rect 511408 352044 511414 352056
rect 580166 352044 580172 352056
rect 580224 352044 580230 352096
rect 513282 351976 513288 352028
rect 513340 352016 513346 352028
rect 523310 352016 523316 352028
rect 513340 351988 523316 352016
rect 513340 351976 513346 351988
rect 523310 351976 523316 351988
rect 523368 351976 523374 352028
rect 395982 351908 395988 351960
rect 396040 351948 396046 351960
rect 447134 351948 447140 351960
rect 396040 351920 447140 351948
rect 396040 351908 396046 351920
rect 447134 351908 447140 351920
rect 447192 351908 447198 351960
rect 513282 350888 513288 350940
rect 513340 350928 513346 350940
rect 518986 350928 518992 350940
rect 513340 350900 518992 350928
rect 513340 350888 513346 350900
rect 518986 350888 518992 350900
rect 519044 350888 519050 350940
rect 512454 350752 512460 350804
rect 512512 350792 512518 350804
rect 515122 350792 515128 350804
rect 512512 350764 515128 350792
rect 512512 350752 512518 350764
rect 515122 350752 515128 350764
rect 515180 350752 515186 350804
rect 407022 350548 407028 350600
rect 407080 350588 407086 350600
rect 447134 350588 447140 350600
rect 407080 350560 447140 350588
rect 407080 350548 407086 350560
rect 447134 350548 447140 350560
rect 447192 350548 447198 350600
rect 509786 349800 509792 349852
rect 509844 349840 509850 349852
rect 510062 349840 510068 349852
rect 509844 349812 510068 349840
rect 509844 349800 509850 349812
rect 510062 349800 510068 349812
rect 510120 349800 510126 349852
rect 513282 349664 513288 349716
rect 513340 349704 513346 349716
rect 519170 349704 519176 349716
rect 513340 349676 519176 349704
rect 513340 349664 513346 349676
rect 519170 349664 519176 349676
rect 519228 349664 519234 349716
rect 512454 349528 512460 349580
rect 512512 349568 512518 349580
rect 514938 349568 514944 349580
rect 512512 349540 514944 349568
rect 512512 349528 512518 349540
rect 514938 349528 514944 349540
rect 514996 349528 515002 349580
rect 512454 349120 512460 349172
rect 512512 349160 512518 349172
rect 513834 349160 513840 349172
rect 512512 349132 513840 349160
rect 512512 349120 512518 349132
rect 513834 349120 513840 349132
rect 513892 349120 513898 349172
rect 513006 347896 513012 347948
rect 513064 347936 513070 347948
rect 516686 347936 516692 347948
rect 513064 347908 516692 347936
rect 513064 347896 513070 347908
rect 516686 347896 516692 347908
rect 516744 347896 516750 347948
rect 361758 347760 361764 347812
rect 361816 347800 361822 347812
rect 402238 347800 402244 347812
rect 361816 347772 402244 347800
rect 361816 347760 361822 347772
rect 402238 347760 402244 347772
rect 402296 347760 402302 347812
rect 362218 347692 362224 347744
rect 362276 347732 362282 347744
rect 447134 347732 447140 347744
rect 362276 347704 447140 347732
rect 362276 347692 362282 347704
rect 447134 347692 447140 347704
rect 447192 347692 447198 347744
rect 512454 347624 512460 347676
rect 512512 347664 512518 347676
rect 513926 347664 513932 347676
rect 512512 347636 513932 347664
rect 512512 347624 512518 347636
rect 513926 347624 513932 347636
rect 513984 347624 513990 347676
rect 513282 346536 513288 346588
rect 513340 346576 513346 346588
rect 518066 346576 518072 346588
rect 513340 346548 518072 346576
rect 513340 346536 513346 346548
rect 518066 346536 518072 346548
rect 518124 346536 518130 346588
rect 416130 346400 416136 346452
rect 416188 346440 416194 346452
rect 423674 346440 423680 346452
rect 416188 346412 423680 346440
rect 416188 346400 416194 346412
rect 423674 346400 423680 346412
rect 423732 346400 423738 346452
rect 512822 346400 512828 346452
rect 512880 346440 512886 346452
rect 516594 346440 516600 346452
rect 512880 346412 516600 346440
rect 512880 346400 512886 346412
rect 516594 346400 516600 346412
rect 516652 346400 516658 346452
rect 512454 345584 512460 345636
rect 512512 345624 512518 345636
rect 515214 345624 515220 345636
rect 512512 345596 515220 345624
rect 512512 345584 512518 345596
rect 515214 345584 515220 345596
rect 515272 345584 515278 345636
rect 446306 344700 446312 344752
rect 446364 344740 446370 344752
rect 448330 344740 448336 344752
rect 446364 344712 448336 344740
rect 446364 344700 446370 344712
rect 448330 344700 448336 344712
rect 448388 344700 448394 344752
rect 513282 344360 513288 344412
rect 513340 344400 513346 344412
rect 519078 344400 519084 344412
rect 513340 344372 519084 344400
rect 513340 344360 513346 344372
rect 519078 344360 519084 344372
rect 519136 344360 519142 344412
rect 513006 343680 513012 343732
rect 513064 343720 513070 343732
rect 518250 343720 518256 343732
rect 513064 343692 518256 343720
rect 513064 343680 513070 343692
rect 518250 343680 518256 343692
rect 518308 343680 518314 343732
rect 513006 343136 513012 343188
rect 513064 343176 513070 343188
rect 518342 343176 518348 343188
rect 513064 343148 518348 343176
rect 513064 343136 513070 343148
rect 518342 343136 518348 343148
rect 518400 343136 518406 343188
rect 423674 341572 423680 341624
rect 423732 341612 423738 341624
rect 429838 341612 429844 341624
rect 423732 341584 429844 341612
rect 423732 341572 423738 341584
rect 429838 341572 429844 341584
rect 429896 341572 429902 341624
rect 513282 341232 513288 341284
rect 513340 341272 513346 341284
rect 520642 341272 520648 341284
rect 513340 341244 520648 341272
rect 513340 341232 513346 341244
rect 520642 341232 520648 341244
rect 520700 341232 520706 341284
rect 513282 341096 513288 341148
rect 513340 341136 513346 341148
rect 519354 341136 519360 341148
rect 513340 341108 519360 341136
rect 513340 341096 513346 341108
rect 519354 341096 519360 341108
rect 519412 341096 519418 341148
rect 438854 340960 438860 341012
rect 438912 341000 438918 341012
rect 447134 341000 447140 341012
rect 438912 340972 447140 341000
rect 438912 340960 438918 340972
rect 447134 340960 447140 340972
rect 447192 340960 447198 341012
rect 361758 340892 361764 340944
rect 361816 340932 361822 340944
rect 447226 340932 447232 340944
rect 361816 340904 447232 340932
rect 361816 340892 361822 340904
rect 447226 340892 447232 340904
rect 447284 340892 447290 340944
rect 513098 339600 513104 339652
rect 513156 339640 513162 339652
rect 516778 339640 516784 339652
rect 513156 339612 516784 339640
rect 513156 339600 513162 339612
rect 516778 339600 516784 339612
rect 516836 339600 516842 339652
rect 435450 339532 435456 339584
rect 435508 339572 435514 339584
rect 447134 339572 447140 339584
rect 435508 339544 447140 339572
rect 435508 339532 435514 339544
rect 447134 339532 447140 339544
rect 447192 339532 447198 339584
rect 513282 339532 513288 339584
rect 513340 339572 513346 339584
rect 519722 339572 519728 339584
rect 513340 339544 519728 339572
rect 513340 339532 513346 339544
rect 519722 339532 519728 339544
rect 519780 339532 519786 339584
rect 374638 339464 374644 339516
rect 374696 339504 374702 339516
rect 447226 339504 447232 339516
rect 374696 339476 447232 339504
rect 374696 339464 374702 339476
rect 447226 339464 447232 339476
rect 447284 339464 447290 339516
rect 513006 338648 513012 338700
rect 513064 338688 513070 338700
rect 519262 338688 519268 338700
rect 513064 338660 519268 338688
rect 513064 338648 513070 338660
rect 519262 338648 519268 338660
rect 519320 338648 519326 338700
rect 439682 338172 439688 338224
rect 439740 338212 439746 338224
rect 447134 338212 447140 338224
rect 439740 338184 447140 338212
rect 439740 338172 439746 338184
rect 447134 338172 447140 338184
rect 447192 338172 447198 338224
rect 436830 338104 436836 338156
rect 436888 338144 436894 338156
rect 447226 338144 447232 338156
rect 436888 338116 447232 338144
rect 436888 338104 436894 338116
rect 447226 338104 447232 338116
rect 447284 338104 447290 338156
rect 450078 337424 450084 337476
rect 450136 337464 450142 337476
rect 450354 337464 450360 337476
rect 450136 337436 450360 337464
rect 450136 337424 450142 337436
rect 450354 337424 450360 337436
rect 450412 337424 450418 337476
rect 402238 337356 402244 337408
rect 402296 337396 402302 337408
rect 447318 337396 447324 337408
rect 402296 337368 447324 337396
rect 402296 337356 402302 337368
rect 447318 337356 447324 337368
rect 447376 337396 447382 337408
rect 448422 337396 448428 337408
rect 447376 337368 448428 337396
rect 447376 337356 447382 337368
rect 448422 337356 448428 337368
rect 448480 337356 448486 337408
rect 513282 337152 513288 337204
rect 513340 337192 513346 337204
rect 520734 337192 520740 337204
rect 513340 337164 520740 337192
rect 513340 337152 513346 337164
rect 520734 337152 520740 337164
rect 520792 337152 520798 337204
rect 512730 337016 512736 337068
rect 512788 337056 512794 337068
rect 515306 337056 515312 337068
rect 512788 337028 515312 337056
rect 512788 337016 512794 337028
rect 515306 337016 515312 337028
rect 515364 337016 515370 337068
rect 512822 336948 512828 337000
rect 512880 336988 512886 337000
rect 516134 336988 516140 337000
rect 512880 336960 516140 336988
rect 512880 336948 512886 336960
rect 516134 336948 516140 336960
rect 516192 336948 516198 337000
rect 416774 336880 416780 336932
rect 416832 336920 416838 336932
rect 450354 336920 450360 336932
rect 416832 336892 450360 336920
rect 416832 336880 416838 336892
rect 450354 336880 450360 336892
rect 450412 336880 450418 336932
rect 413094 336812 413100 336864
rect 413152 336852 413158 336864
rect 450170 336852 450176 336864
rect 413152 336824 450176 336852
rect 413152 336812 413158 336824
rect 450170 336812 450176 336824
rect 450228 336812 450234 336864
rect 409414 336744 409420 336796
rect 409472 336784 409478 336796
rect 450722 336784 450728 336796
rect 409472 336756 450728 336784
rect 409472 336744 409478 336756
rect 450722 336744 450728 336756
rect 450780 336744 450786 336796
rect 438118 336472 438124 336524
rect 438176 336512 438182 336524
rect 447134 336512 447140 336524
rect 438176 336484 447140 336512
rect 438176 336472 438182 336484
rect 447134 336472 447140 336484
rect 447192 336472 447198 336524
rect 418982 336404 418988 336456
rect 419040 336444 419046 336456
rect 442350 336444 442356 336456
rect 419040 336416 442356 336444
rect 419040 336404 419046 336416
rect 442350 336404 442356 336416
rect 442408 336404 442414 336456
rect 418890 336336 418896 336388
rect 418948 336376 418954 336388
rect 442442 336376 442448 336388
rect 418948 336348 442448 336376
rect 418948 336336 418954 336348
rect 442442 336336 442448 336348
rect 442500 336336 442506 336388
rect 418798 336268 418804 336320
rect 418856 336308 418862 336320
rect 442718 336308 442724 336320
rect 418856 336280 442724 336308
rect 418856 336268 418862 336280
rect 442718 336268 442724 336280
rect 442776 336268 442782 336320
rect 416038 336200 416044 336252
rect 416096 336240 416102 336252
rect 439958 336240 439964 336252
rect 416096 336212 439964 336240
rect 416096 336200 416102 336212
rect 439958 336200 439964 336212
rect 440016 336200 440022 336252
rect 413646 336132 413652 336184
rect 413704 336172 413710 336184
rect 449434 336172 449440 336184
rect 413704 336144 449440 336172
rect 413704 336132 413710 336144
rect 449434 336132 449440 336144
rect 449492 336132 449498 336184
rect 399478 336064 399484 336116
rect 399536 336104 399542 336116
rect 447226 336104 447232 336116
rect 399536 336076 447232 336104
rect 399536 336064 399542 336076
rect 447226 336064 447232 336076
rect 447284 336064 447290 336116
rect 362218 335996 362224 336048
rect 362276 336036 362282 336048
rect 438854 336036 438860 336048
rect 362276 336008 438860 336036
rect 362276 335996 362282 336008
rect 438854 335996 438860 336008
rect 438912 335996 438918 336048
rect 512730 335928 512736 335980
rect 512788 335968 512794 335980
rect 515582 335968 515588 335980
rect 512788 335940 515588 335968
rect 512788 335928 512794 335940
rect 515582 335928 515588 335940
rect 515640 335928 515646 335980
rect 443730 335656 443736 335708
rect 443788 335696 443794 335708
rect 447134 335696 447140 335708
rect 443788 335668 447140 335696
rect 443788 335656 443794 335668
rect 447134 335656 447140 335668
rect 447192 335656 447198 335708
rect 439590 335316 439596 335368
rect 439648 335356 439654 335368
rect 447134 335356 447140 335368
rect 439648 335328 447140 335356
rect 439648 335316 439654 335328
rect 447134 335316 447140 335328
rect 447192 335316 447198 335368
rect 420546 335044 420552 335096
rect 420604 335084 420610 335096
rect 439774 335084 439780 335096
rect 420604 335056 439780 335084
rect 420604 335044 420610 335056
rect 439774 335044 439780 335056
rect 439832 335044 439838 335096
rect 420178 334976 420184 335028
rect 420236 335016 420242 335028
rect 439866 335016 439872 335028
rect 420236 334988 439872 335016
rect 420236 334976 420242 334988
rect 439866 334976 439872 334988
rect 439924 334976 439930 335028
rect 420822 334908 420828 334960
rect 420880 334948 420886 334960
rect 442534 334948 442540 334960
rect 420880 334920 442540 334948
rect 420880 334908 420886 334920
rect 442534 334908 442540 334920
rect 442592 334908 442598 334960
rect 420638 334840 420644 334892
rect 420696 334880 420702 334892
rect 442626 334880 442632 334892
rect 420696 334852 442632 334880
rect 420696 334840 420702 334852
rect 442626 334840 442632 334852
rect 442684 334840 442690 334892
rect 420270 334772 420276 334824
rect 420328 334812 420334 334824
rect 442810 334812 442816 334824
rect 420328 334784 442816 334812
rect 420328 334772 420334 334784
rect 442810 334772 442816 334784
rect 442868 334772 442874 334824
rect 420730 334704 420736 334756
rect 420788 334744 420794 334756
rect 444006 334744 444012 334756
rect 420788 334716 444012 334744
rect 420788 334704 420794 334716
rect 444006 334704 444012 334716
rect 444064 334704 444070 334756
rect 513006 334704 513012 334756
rect 513064 334744 513070 334756
rect 519446 334744 519452 334756
rect 513064 334716 519452 334744
rect 513064 334704 513070 334716
rect 519446 334704 519452 334716
rect 519504 334704 519510 334756
rect 420270 334636 420276 334688
rect 420328 334676 420334 334688
rect 444926 334676 444932 334688
rect 420328 334648 444932 334676
rect 420328 334636 420334 334648
rect 444926 334636 444932 334648
rect 444984 334636 444990 334688
rect 420086 334568 420092 334620
rect 420144 334608 420150 334620
rect 444834 334608 444840 334620
rect 420144 334580 444840 334608
rect 420144 334568 420150 334580
rect 444834 334568 444840 334580
rect 444892 334568 444898 334620
rect 513282 334568 513288 334620
rect 513340 334608 513346 334620
rect 520918 334608 520924 334620
rect 513340 334580 520924 334608
rect 513340 334568 513346 334580
rect 520918 334568 520924 334580
rect 520976 334568 520982 334620
rect 443638 334024 443644 334076
rect 443696 334064 443702 334076
rect 447226 334064 447232 334076
rect 443696 334036 447232 334064
rect 443696 334024 443702 334036
rect 447226 334024 447232 334036
rect 447284 334024 447290 334076
rect 364058 333956 364064 334008
rect 364116 333996 364122 334008
rect 447134 333996 447140 334008
rect 364116 333968 447140 333996
rect 364116 333956 364122 333968
rect 447134 333956 447140 333968
rect 447192 333956 447198 334008
rect 436738 332664 436744 332716
rect 436796 332704 436802 332716
rect 447226 332704 447232 332716
rect 436796 332676 447232 332704
rect 436796 332664 436802 332676
rect 447226 332664 447232 332676
rect 447284 332664 447290 332716
rect 431218 332596 431224 332648
rect 431276 332636 431282 332648
rect 447134 332636 447140 332648
rect 431276 332608 447140 332636
rect 431276 332596 431282 332608
rect 447134 332596 447140 332608
rect 447192 332596 447198 332648
rect 432782 331848 432788 331900
rect 432840 331888 432846 331900
rect 443914 331888 443920 331900
rect 432840 331860 443920 331888
rect 432840 331848 432846 331860
rect 443914 331848 443920 331860
rect 443972 331848 443978 331900
rect 512822 331576 512828 331628
rect 512880 331616 512886 331628
rect 520826 331616 520832 331628
rect 512880 331588 520832 331616
rect 512880 331576 512886 331588
rect 520826 331576 520832 331588
rect 520884 331576 520890 331628
rect 450078 330488 450084 330540
rect 450136 330528 450142 330540
rect 450722 330528 450728 330540
rect 450136 330500 450728 330528
rect 450136 330488 450142 330500
rect 450722 330488 450728 330500
rect 450780 330488 450786 330540
rect 442902 330080 442908 330132
rect 442960 330120 442966 330132
rect 447134 330120 447140 330132
rect 442960 330092 447140 330120
rect 442960 330080 442966 330092
rect 447134 330080 447140 330092
rect 447192 330080 447198 330132
rect 512822 329128 512828 329180
rect 512880 329168 512886 329180
rect 516870 329168 516876 329180
rect 512880 329140 516876 329168
rect 512880 329128 512886 329140
rect 516870 329128 516876 329140
rect 516928 329128 516934 329180
rect 439498 329060 439504 329112
rect 439556 329100 439562 329112
rect 447134 329100 447140 329112
rect 439556 329072 447140 329100
rect 439556 329060 439562 329072
rect 447134 329060 447140 329072
rect 447192 329060 447198 329112
rect 436002 328448 436008 328500
rect 436060 328488 436066 328500
rect 449894 328488 449900 328500
rect 436060 328460 449900 328488
rect 436060 328448 436066 328460
rect 449894 328448 449900 328460
rect 449952 328448 449958 328500
rect 431862 327088 431868 327140
rect 431920 327128 431926 327140
rect 449894 327128 449900 327140
rect 431920 327100 449900 327128
rect 431920 327088 431926 327100
rect 449894 327088 449900 327100
rect 449952 327088 449958 327140
rect 509786 326408 509792 326460
rect 509844 326448 509850 326460
rect 510062 326448 510068 326460
rect 509844 326420 510068 326448
rect 509844 326408 509850 326420
rect 510062 326408 510068 326420
rect 510120 326408 510126 326460
rect 432690 324912 432696 324964
rect 432748 324952 432754 324964
rect 442258 324952 442264 324964
rect 432748 324924 442264 324952
rect 432748 324912 432754 324924
rect 442258 324912 442264 324924
rect 442316 324912 442322 324964
rect 511902 324912 511908 324964
rect 511960 324952 511966 324964
rect 580626 324952 580632 324964
rect 511960 324924 580632 324952
rect 511960 324912 511966 324924
rect 580626 324912 580632 324924
rect 580684 324912 580690 324964
rect 510430 323552 510436 323604
rect 510488 323592 510494 323604
rect 580350 323592 580356 323604
rect 510488 323564 580356 323592
rect 510488 323552 510494 323564
rect 580350 323552 580356 323564
rect 580408 323552 580414 323604
rect 432598 322940 432604 322992
rect 432656 322980 432662 322992
rect 436922 322980 436928 322992
rect 432656 322952 436928 322980
rect 432656 322940 432662 322952
rect 436922 322940 436928 322952
rect 436980 322940 436986 322992
rect 429838 322192 429844 322244
rect 429896 322232 429902 322244
rect 448514 322232 448520 322244
rect 429896 322204 448520 322232
rect 429896 322192 429902 322204
rect 448514 322192 448520 322204
rect 448572 322192 448578 322244
rect 510522 322192 510528 322244
rect 510580 322232 510586 322244
rect 580442 322232 580448 322244
rect 510580 322204 580448 322232
rect 510580 322192 510586 322204
rect 580442 322192 580448 322204
rect 580500 322192 580506 322244
rect 471790 321960 471796 321972
rect 451246 321932 471796 321960
rect 442810 321852 442816 321904
rect 442868 321892 442874 321904
rect 451246 321892 451274 321932
rect 471790 321920 471796 321932
rect 471848 321920 471854 321972
rect 574738 321960 574744 321972
rect 471992 321932 574744 321960
rect 442868 321864 451274 321892
rect 442868 321852 442874 321864
rect 454540 321852 454546 321904
rect 454598 321892 454604 321904
rect 454954 321892 454960 321904
rect 454598 321864 454960 321892
rect 454598 321852 454604 321864
rect 454954 321852 454960 321864
rect 455012 321852 455018 321904
rect 468294 321852 468300 321904
rect 468352 321892 468358 321904
rect 471992 321892 472020 321932
rect 574738 321920 574744 321932
rect 574796 321920 574802 321972
rect 468352 321864 472020 321892
rect 468352 321852 468358 321864
rect 477494 321852 477500 321904
rect 477552 321892 477558 321904
rect 580166 321892 580172 321904
rect 477552 321864 580172 321892
rect 477552 321852 477558 321864
rect 580166 321852 580172 321864
rect 580224 321852 580230 321904
rect 449250 321784 449256 321836
rect 449308 321824 449314 321836
rect 480714 321824 480720 321836
rect 449308 321796 480720 321824
rect 449308 321784 449314 321796
rect 480714 321784 480720 321796
rect 480772 321784 480778 321836
rect 507210 321784 507216 321836
rect 507268 321824 507274 321836
rect 511166 321824 511172 321836
rect 507268 321796 511172 321824
rect 507268 321784 507274 321796
rect 511166 321784 511172 321796
rect 511224 321784 511230 321836
rect 445570 321716 445576 321768
rect 445628 321756 445634 321768
rect 472434 321756 472440 321768
rect 445628 321728 472440 321756
rect 445628 321716 445634 321728
rect 472434 321716 472440 321728
rect 472492 321716 472498 321768
rect 507394 321716 507400 321768
rect 507452 321756 507458 321768
rect 513466 321756 513472 321768
rect 507452 321728 513472 321756
rect 507452 321716 507458 321728
rect 513466 321716 513472 321728
rect 513524 321716 513530 321768
rect 457806 321580 457812 321632
rect 457864 321620 457870 321632
rect 457864 321592 463694 321620
rect 457864 321580 457870 321592
rect 458358 321512 458364 321564
rect 458416 321552 458422 321564
rect 463666 321552 463694 321592
rect 580258 321552 580264 321564
rect 458416 321524 461440 321552
rect 463666 321524 580264 321552
rect 458416 321512 458422 321524
rect 446490 321444 446496 321496
rect 446548 321484 446554 321496
rect 459462 321484 459468 321496
rect 446548 321456 459468 321484
rect 446548 321444 446554 321456
rect 459462 321444 459468 321456
rect 459520 321444 459526 321496
rect 461412 321484 461440 321524
rect 580258 321512 580264 321524
rect 580316 321512 580322 321564
rect 570598 321484 570604 321496
rect 461412 321456 570604 321484
rect 570598 321444 570604 321456
rect 570656 321444 570662 321496
rect 449158 321376 449164 321428
rect 449216 321416 449222 321428
rect 449216 321388 455644 321416
rect 449216 321376 449222 321388
rect 446398 321308 446404 321360
rect 446456 321348 446462 321360
rect 455616 321348 455644 321388
rect 468846 321376 468852 321428
rect 468904 321416 468910 321428
rect 573358 321416 573364 321428
rect 468904 321388 573364 321416
rect 468904 321376 468910 321388
rect 573358 321376 573364 321388
rect 573416 321376 573422 321428
rect 460014 321348 460020 321360
rect 446456 321320 451274 321348
rect 455616 321320 460020 321348
rect 446456 321308 446462 321320
rect 451246 321280 451274 321320
rect 460014 321308 460020 321320
rect 460072 321308 460078 321360
rect 467190 321308 467196 321360
rect 467248 321348 467254 321360
rect 569402 321348 569408 321360
rect 467248 321320 569408 321348
rect 467248 321308 467254 321320
rect 569402 321308 569408 321320
rect 569460 321308 569466 321360
rect 460290 321280 460296 321292
rect 451246 321252 460296 321280
rect 460290 321240 460296 321252
rect 460348 321240 460354 321292
rect 477954 321240 477960 321292
rect 478012 321280 478018 321292
rect 569310 321280 569316 321292
rect 478012 321252 569316 321280
rect 478012 321240 478018 321252
rect 569310 321240 569316 321252
rect 569368 321240 569374 321292
rect 456702 321172 456708 321224
rect 456760 321212 456766 321224
rect 511350 321212 511356 321224
rect 456760 321184 511356 321212
rect 456760 321172 456766 321184
rect 511350 321172 511356 321184
rect 511408 321172 511414 321224
rect 456978 321104 456984 321156
rect 457036 321144 457042 321156
rect 511258 321144 511264 321156
rect 457036 321116 511264 321144
rect 457036 321104 457042 321116
rect 511258 321104 511264 321116
rect 511316 321104 511322 321156
rect 444098 321036 444104 321088
rect 444156 321076 444162 321088
rect 480162 321076 480168 321088
rect 444156 321048 480168 321076
rect 444156 321036 444162 321048
rect 480162 321036 480168 321048
rect 480220 321036 480226 321088
rect 445018 320968 445024 321020
rect 445076 321008 445082 321020
rect 480438 321008 480444 321020
rect 445076 320980 480444 321008
rect 445076 320968 445082 320980
rect 480438 320968 480444 320980
rect 480496 320968 480502 321020
rect 446950 320900 446956 320952
rect 447008 320940 447014 320952
rect 461670 320940 461676 320952
rect 447008 320912 461676 320940
rect 447008 320900 447014 320912
rect 461670 320900 461676 320912
rect 461728 320900 461734 320952
rect 477678 320900 477684 320952
rect 477736 320940 477742 320952
rect 580718 320940 580724 320952
rect 477736 320912 580724 320940
rect 477736 320900 477742 320912
rect 580718 320900 580724 320912
rect 580776 320900 580782 320952
rect 457530 320832 457536 320884
rect 457588 320872 457594 320884
rect 580534 320872 580540 320884
rect 457588 320844 580540 320872
rect 457588 320832 457594 320844
rect 580534 320832 580540 320844
rect 580592 320832 580598 320884
rect 445478 320764 445484 320816
rect 445536 320804 445542 320816
rect 461946 320804 461952 320816
rect 445536 320776 461952 320804
rect 445536 320764 445542 320776
rect 461946 320764 461952 320776
rect 462004 320764 462010 320816
rect 445386 320696 445392 320748
rect 445444 320736 445450 320748
rect 461118 320736 461124 320748
rect 445444 320708 461124 320736
rect 445444 320696 445450 320708
rect 461118 320696 461124 320708
rect 461176 320696 461182 320748
rect 444006 320628 444012 320680
rect 444064 320668 444070 320680
rect 461394 320668 461400 320680
rect 444064 320640 461400 320668
rect 444064 320628 444070 320640
rect 461394 320628 461400 320640
rect 461452 320628 461458 320680
rect 445110 320560 445116 320612
rect 445168 320600 445174 320612
rect 470778 320600 470784 320612
rect 445168 320572 470784 320600
rect 445168 320560 445174 320572
rect 470778 320560 470784 320572
rect 470836 320560 470842 320612
rect 441522 320492 441528 320544
rect 441580 320532 441586 320544
rect 479886 320532 479892 320544
rect 441580 320504 479892 320532
rect 441580 320492 441586 320504
rect 479886 320492 479892 320504
rect 479944 320492 479950 320544
rect 507670 320288 507676 320340
rect 507728 320328 507734 320340
rect 514018 320328 514024 320340
rect 507728 320300 514024 320328
rect 507728 320288 507734 320300
rect 514018 320288 514024 320300
rect 514076 320288 514082 320340
rect 507762 320220 507768 320272
rect 507820 320260 507826 320272
rect 511074 320260 511080 320272
rect 507820 320232 511080 320260
rect 507820 320220 507826 320232
rect 511074 320220 511080 320232
rect 511132 320220 511138 320272
rect 507486 320152 507492 320204
rect 507544 320192 507550 320204
rect 510246 320192 510252 320204
rect 507544 320164 510252 320192
rect 507544 320152 507550 320164
rect 510246 320152 510252 320164
rect 510304 320152 510310 320204
rect 479334 320084 479340 320136
rect 479392 320124 479398 320136
rect 571978 320124 571984 320136
rect 479392 320096 571984 320124
rect 479392 320084 479398 320096
rect 571978 320084 571984 320096
rect 572036 320084 572042 320136
rect 442626 320016 442632 320068
rect 442684 320056 442690 320068
rect 462498 320056 462504 320068
rect 442684 320028 462504 320056
rect 442684 320016 442690 320028
rect 462498 320016 462504 320028
rect 462556 320016 462562 320068
rect 468570 320016 468576 320068
rect 468628 320056 468634 320068
rect 533430 320056 533436 320068
rect 468628 320028 533436 320056
rect 468628 320016 468634 320028
rect 533430 320016 533436 320028
rect 533488 320016 533494 320068
rect 442534 319948 442540 320000
rect 442592 319988 442598 320000
rect 462222 319988 462228 320000
rect 442592 319960 462228 319988
rect 442592 319948 442598 319960
rect 462222 319948 462228 319960
rect 462280 319948 462286 320000
rect 467742 319948 467748 320000
rect 467800 319988 467806 320000
rect 511902 319988 511908 320000
rect 467800 319960 511908 319988
rect 467800 319948 467806 319960
rect 511902 319948 511908 319960
rect 511960 319948 511966 320000
rect 444282 319880 444288 319932
rect 444340 319920 444346 319932
rect 458910 319920 458916 319932
rect 444340 319892 458916 319920
rect 444340 319880 444346 319892
rect 458910 319880 458916 319892
rect 458968 319880 458974 319932
rect 467466 319880 467472 319932
rect 467524 319920 467530 319932
rect 510430 319920 510436 319932
rect 467524 319892 510436 319920
rect 467524 319880 467530 319892
rect 510430 319880 510436 319892
rect 510488 319880 510494 319932
rect 468018 319812 468024 319864
rect 468076 319852 468082 319864
rect 510522 319852 510528 319864
rect 468076 319824 510528 319852
rect 468076 319812 468082 319824
rect 510522 319812 510528 319824
rect 510580 319812 510586 319864
rect 446674 319744 446680 319796
rect 446732 319784 446738 319796
rect 470226 319784 470232 319796
rect 446732 319756 470232 319784
rect 446732 319744 446738 319756
rect 470226 319744 470232 319756
rect 470284 319744 470290 319796
rect 478782 319744 478788 319796
rect 478840 319784 478846 319796
rect 519538 319784 519544 319796
rect 478840 319756 519544 319784
rect 478840 319744 478846 319756
rect 519538 319744 519544 319756
rect 519596 319744 519602 319796
rect 446582 319676 446588 319728
rect 446640 319716 446646 319728
rect 470502 319716 470508 319728
rect 446640 319688 470508 319716
rect 446640 319676 446646 319688
rect 470502 319676 470508 319688
rect 470560 319676 470566 319728
rect 479610 319676 479616 319728
rect 479668 319716 479674 319728
rect 519630 319716 519636 319728
rect 479668 319688 519636 319716
rect 479668 319676 479674 319688
rect 519630 319676 519636 319688
rect 519688 319676 519694 319728
rect 448514 319608 448520 319660
rect 448572 319648 448578 319660
rect 472986 319648 472992 319660
rect 448572 319620 472992 319648
rect 448572 319608 448578 319620
rect 472986 319608 472992 319620
rect 473044 319608 473050 319660
rect 478506 319608 478512 319660
rect 478564 319648 478570 319660
rect 518158 319648 518164 319660
rect 478564 319620 518164 319648
rect 478564 319608 478570 319620
rect 518158 319608 518164 319620
rect 518216 319608 518222 319660
rect 445202 319540 445208 319592
rect 445260 319580 445266 319592
rect 469950 319580 469956 319592
rect 445260 319552 469956 319580
rect 445260 319540 445266 319552
rect 469950 319540 469956 319552
rect 470008 319540 470014 319592
rect 478230 319540 478236 319592
rect 478288 319580 478294 319592
rect 515490 319580 515496 319592
rect 478288 319552 515496 319580
rect 478288 319540 478294 319552
rect 515490 319540 515496 319552
rect 515548 319540 515554 319592
rect 446858 319472 446864 319524
rect 446916 319512 446922 319524
rect 471606 319512 471612 319524
rect 446916 319484 471612 319512
rect 446916 319472 446922 319484
rect 471606 319472 471612 319484
rect 471664 319472 471670 319524
rect 479058 319472 479064 319524
rect 479116 319512 479122 319524
rect 515398 319512 515404 319524
rect 479116 319484 515404 319512
rect 479116 319472 479122 319484
rect 515398 319472 515404 319484
rect 515456 319472 515462 319524
rect 449434 319404 449440 319456
rect 449492 319444 449498 319456
rect 469674 319444 469680 319456
rect 449492 319416 469680 319444
rect 449492 319404 449498 319416
rect 469674 319404 469680 319416
rect 469732 319404 469738 319456
rect 479518 319404 479524 319456
rect 479576 319444 479582 319456
rect 483474 319444 483480 319456
rect 479576 319416 483480 319444
rect 479576 319404 479582 319416
rect 483474 319404 483480 319416
rect 483532 319404 483538 319456
rect 502518 319404 502524 319456
rect 502576 319444 502582 319456
rect 543734 319444 543740 319456
rect 502576 319416 543740 319444
rect 502576 319404 502582 319416
rect 543734 319404 543740 319416
rect 543792 319404 543798 319456
rect 497274 319336 497280 319388
rect 497332 319376 497338 319388
rect 533338 319376 533344 319388
rect 497332 319348 533344 319376
rect 497332 319336 497338 319348
rect 533338 319336 533344 319348
rect 533396 319336 533402 319388
rect 445294 319268 445300 319320
rect 445352 319308 445358 319320
rect 482922 319308 482928 319320
rect 445352 319280 482928 319308
rect 445352 319268 445358 319280
rect 482922 319268 482928 319280
rect 482980 319268 482986 319320
rect 439866 319200 439872 319252
rect 439924 319240 439930 319252
rect 482646 319240 482652 319252
rect 439924 319212 482652 319240
rect 439924 319200 439930 319212
rect 482646 319200 482652 319212
rect 482704 319200 482710 319252
rect 446766 319132 446772 319184
rect 446824 319172 446830 319184
rect 481266 319172 481272 319184
rect 446824 319144 481272 319172
rect 446824 319132 446830 319144
rect 481266 319132 481272 319144
rect 481324 319132 481330 319184
rect 480898 319064 480904 319116
rect 480956 319104 480962 319116
rect 483750 319104 483756 319116
rect 480956 319076 483756 319104
rect 480956 319064 480962 319076
rect 483750 319064 483756 319076
rect 483808 319064 483814 319116
rect 485866 319064 485872 319116
rect 485924 319104 485930 319116
rect 487062 319104 487068 319116
rect 485924 319076 487068 319104
rect 485924 319064 485930 319076
rect 487062 319064 487068 319076
rect 487120 319064 487126 319116
rect 502702 319064 502708 319116
rect 502760 319104 502766 319116
rect 503622 319104 503628 319116
rect 502760 319076 503628 319104
rect 502760 319064 502766 319076
rect 503622 319064 503628 319076
rect 503680 319064 503686 319116
rect 447594 318724 447600 318776
rect 447652 318764 447658 318776
rect 449158 318764 449164 318776
rect 447652 318736 449164 318764
rect 447652 318724 447658 318736
rect 449158 318724 449164 318736
rect 449216 318724 449222 318776
rect 457254 318724 457260 318776
rect 457312 318764 457318 318776
rect 576118 318764 576124 318776
rect 457312 318736 576124 318764
rect 457312 318724 457318 318736
rect 576118 318724 576124 318736
rect 576176 318724 576182 318776
rect 458082 318656 458088 318708
rect 458140 318696 458146 318708
rect 569218 318696 569224 318708
rect 458140 318668 569224 318696
rect 458140 318656 458146 318668
rect 569218 318656 569224 318668
rect 569276 318656 569282 318708
rect 439774 318588 439780 318640
rect 439832 318628 439838 318640
rect 483198 318628 483204 318640
rect 439832 318600 483204 318628
rect 439832 318588 439838 318600
rect 483198 318588 483204 318600
rect 483256 318588 483262 318640
rect 432046 318520 432052 318572
rect 432104 318560 432110 318572
rect 435358 318560 435364 318572
rect 432104 318532 435364 318560
rect 432104 318520 432110 318532
rect 435358 318520 435364 318532
rect 435416 318520 435422 318572
rect 442350 318520 442356 318572
rect 442408 318560 442414 318572
rect 482094 318560 482100 318572
rect 442408 318532 482100 318560
rect 442408 318520 442414 318532
rect 482094 318520 482100 318532
rect 482152 318520 482158 318572
rect 444926 318452 444932 318504
rect 444984 318492 444990 318504
rect 472710 318492 472716 318504
rect 444984 318464 472716 318492
rect 444984 318452 444990 318464
rect 472710 318452 472716 318464
rect 472768 318452 472774 318504
rect 445662 318384 445668 318436
rect 445720 318424 445726 318436
rect 469398 318424 469404 318436
rect 445720 318396 469404 318424
rect 445720 318384 445726 318396
rect 469398 318384 469404 318396
rect 469456 318384 469462 318436
rect 458910 318248 458916 318300
rect 458968 318288 458974 318300
rect 490098 318288 490104 318300
rect 458968 318260 490104 318288
rect 458968 318248 458974 318260
rect 490098 318248 490104 318260
rect 490156 318248 490162 318300
rect 496446 318248 496452 318300
rect 496504 318288 496510 318300
rect 539594 318288 539600 318300
rect 496504 318260 539600 318288
rect 496504 318248 496510 318260
rect 539594 318248 539600 318260
rect 539652 318248 539658 318300
rect 459094 318180 459100 318232
rect 459152 318220 459158 318232
rect 492582 318220 492588 318232
rect 459152 318192 492588 318220
rect 459152 318180 459158 318192
rect 492582 318180 492588 318192
rect 492640 318180 492646 318232
rect 494790 318180 494796 318232
rect 494848 318220 494854 318232
rect 540974 318220 540980 318232
rect 494848 318192 540980 318220
rect 494848 318180 494854 318192
rect 540974 318180 540980 318192
rect 541032 318180 541038 318232
rect 460750 318112 460756 318164
rect 460808 318152 460814 318164
rect 513374 318152 513380 318164
rect 460808 318124 513380 318152
rect 460808 318112 460814 318124
rect 513374 318112 513380 318124
rect 513432 318112 513438 318164
rect 450630 318044 450636 318096
rect 450688 318084 450694 318096
rect 457714 318084 457720 318096
rect 450688 318056 457720 318084
rect 450688 318044 450694 318056
rect 457714 318044 457720 318056
rect 457772 318044 457778 318096
rect 460658 318044 460664 318096
rect 460716 318084 460722 318096
rect 516134 318084 516140 318096
rect 460716 318056 516140 318084
rect 460716 318044 460722 318056
rect 516134 318044 516140 318056
rect 516192 318044 516198 318096
rect 497734 317704 497740 317756
rect 497792 317744 497798 317756
rect 498102 317744 498108 317756
rect 497792 317716 498108 317744
rect 497792 317704 497798 317716
rect 498102 317704 498108 317716
rect 498160 317704 498166 317756
rect 498654 317024 498660 317076
rect 498712 317064 498718 317076
rect 541066 317064 541072 317076
rect 498712 317036 541072 317064
rect 498712 317024 498718 317036
rect 541066 317024 541072 317036
rect 541124 317024 541130 317076
rect 459002 316956 459008 317008
rect 459060 316996 459066 317008
rect 491478 316996 491484 317008
rect 459060 316968 491484 316996
rect 459060 316956 459066 316968
rect 491478 316956 491484 316968
rect 491536 316956 491542 317008
rect 499758 316956 499764 317008
rect 499816 316996 499822 317008
rect 543090 316996 543096 317008
rect 499816 316968 543096 316996
rect 499816 316956 499822 316968
rect 543090 316956 543096 316968
rect 543148 316956 543154 317008
rect 485958 316888 485964 316940
rect 486016 316928 486022 316940
rect 529934 316928 529940 316940
rect 486016 316900 529940 316928
rect 486016 316888 486022 316900
rect 529934 316888 529940 316900
rect 529992 316888 529998 316940
rect 453298 316820 453304 316872
rect 453356 316860 453362 316872
rect 488994 316860 489000 316872
rect 453356 316832 489000 316860
rect 453356 316820 453362 316832
rect 488994 316820 489000 316832
rect 489052 316820 489058 316872
rect 495618 316820 495624 316872
rect 495676 316860 495682 316872
rect 543182 316860 543188 316872
rect 495676 316832 543188 316860
rect 495676 316820 495682 316832
rect 543182 316820 543188 316832
rect 543240 316820 543246 316872
rect 454678 316752 454684 316804
rect 454736 316792 454742 316804
rect 503346 316792 503352 316804
rect 454736 316764 503352 316792
rect 454736 316752 454742 316764
rect 503346 316752 503352 316764
rect 503404 316752 503410 316804
rect 450538 316684 450544 316736
rect 450596 316724 450602 316736
rect 504174 316724 504180 316736
rect 450596 316696 504180 316724
rect 450596 316684 450602 316696
rect 504174 316684 504180 316696
rect 504232 316684 504238 316736
rect 456426 316004 456432 316056
rect 456484 316044 456490 316056
rect 461578 316044 461584 316056
rect 456484 316016 461584 316044
rect 456484 316004 456490 316016
rect 461578 316004 461584 316016
rect 461636 316004 461642 316056
rect 499022 316004 499028 316056
rect 499080 316044 499086 316056
rect 499206 316044 499212 316056
rect 499080 316016 499212 316044
rect 499080 316004 499086 316016
rect 499206 316004 499212 316016
rect 499264 316004 499270 316056
rect 361758 315936 361764 315988
rect 361816 315976 361822 315988
rect 374638 315976 374644 315988
rect 361816 315948 374644 315976
rect 361816 315936 361822 315948
rect 374638 315936 374644 315948
rect 374696 315936 374702 315988
rect 457438 315392 457444 315444
rect 457496 315432 457502 315444
rect 491754 315432 491760 315444
rect 457496 315404 491760 315432
rect 457496 315392 457502 315404
rect 491754 315392 491760 315404
rect 491812 315392 491818 315444
rect 453390 315324 453396 315376
rect 453448 315364 453454 315376
rect 489546 315364 489552 315376
rect 453448 315336 489552 315364
rect 453448 315324 453454 315336
rect 489546 315324 489552 315336
rect 489604 315324 489610 315376
rect 499114 315324 499120 315376
rect 499172 315364 499178 315376
rect 539870 315364 539876 315376
rect 499172 315336 539876 315364
rect 499172 315324 499178 315336
rect 539870 315324 539876 315336
rect 539928 315324 539934 315376
rect 450630 315256 450636 315308
rect 450688 315296 450694 315308
rect 502702 315296 502708 315308
rect 450688 315268 502708 315296
rect 450688 315256 450694 315268
rect 502702 315256 502708 315268
rect 502760 315256 502766 315308
rect 509786 314168 509792 314220
rect 509844 314208 509850 314220
rect 510062 314208 510068 314220
rect 509844 314180 510068 314208
rect 509844 314168 509850 314180
rect 510062 314168 510068 314180
rect 510120 314168 510126 314220
rect 448514 314100 448520 314152
rect 448572 314140 448578 314152
rect 462774 314140 462780 314152
rect 448572 314112 462780 314140
rect 448572 314100 448578 314112
rect 462774 314100 462780 314112
rect 462832 314100 462838 314152
rect 452010 314032 452016 314084
rect 452068 314072 452074 314084
rect 492858 314072 492864 314084
rect 452068 314044 492864 314072
rect 452068 314032 452074 314044
rect 492858 314032 492864 314044
rect 492916 314032 492922 314084
rect 500310 314032 500316 314084
rect 500368 314072 500374 314084
rect 542722 314072 542728 314084
rect 500368 314044 542728 314072
rect 500368 314032 500374 314044
rect 542722 314032 542728 314044
rect 542780 314032 542786 314084
rect 450722 313964 450728 314016
rect 450780 314004 450786 314016
rect 503898 314004 503904 314016
rect 450780 313976 503904 314004
rect 450780 313964 450786 313976
rect 503898 313964 503904 313976
rect 503956 313964 503962 314016
rect 432690 313896 432696 313948
rect 432748 313936 432754 313948
rect 443822 313936 443828 313948
rect 432748 313908 443828 313936
rect 432748 313896 432754 313908
rect 443822 313896 443828 313908
rect 443880 313896 443886 313948
rect 455230 313896 455236 313948
rect 455288 313936 455294 313948
rect 463050 313936 463056 313948
rect 455288 313908 463056 313936
rect 455288 313896 455294 313908
rect 463050 313896 463056 313908
rect 463108 313896 463114 313948
rect 533430 313936 533436 313948
rect 470566 313908 533436 313936
rect 455598 313828 455604 313880
rect 455656 313868 455662 313880
rect 470566 313868 470594 313908
rect 533430 313896 533436 313908
rect 533488 313896 533494 313948
rect 455656 313840 470594 313868
rect 455656 313828 455662 313840
rect 466914 313216 466920 313268
rect 466972 313256 466978 313268
rect 580166 313256 580172 313268
rect 466972 313228 580172 313256
rect 466972 313216 466978 313228
rect 580166 313216 580172 313228
rect 580224 313216 580230 313268
rect 500034 312604 500040 312656
rect 500092 312644 500098 312656
rect 542630 312644 542636 312656
rect 500092 312616 542636 312644
rect 500092 312604 500098 312616
rect 542630 312604 542636 312616
rect 542688 312604 542694 312656
rect 496354 312536 496360 312588
rect 496412 312576 496418 312588
rect 539686 312576 539692 312588
rect 496412 312548 539692 312576
rect 496412 312536 496418 312548
rect 539686 312536 539692 312548
rect 539744 312536 539750 312588
rect 472618 311312 472624 311364
rect 472676 311352 472682 311364
rect 480898 311352 480904 311364
rect 472676 311324 480904 311352
rect 472676 311312 472682 311324
rect 480898 311312 480904 311324
rect 480956 311312 480962 311364
rect 452194 311244 452200 311296
rect 452252 311284 452258 311296
rect 494238 311284 494244 311296
rect 452252 311256 494244 311284
rect 452252 311244 452258 311256
rect 494238 311244 494244 311256
rect 494296 311244 494302 311296
rect 501966 311244 501972 311296
rect 502024 311284 502030 311296
rect 538858 311284 538864 311296
rect 502024 311256 538864 311284
rect 502024 311244 502030 311256
rect 538858 311244 538864 311256
rect 538916 311244 538922 311296
rect 450814 311176 450820 311228
rect 450872 311216 450878 311228
rect 504450 311216 504456 311228
rect 450872 311188 504456 311216
rect 450872 311176 450878 311188
rect 504450 311176 504456 311188
rect 504508 311176 504514 311228
rect 440878 311108 440884 311160
rect 440936 311148 440942 311160
rect 448514 311148 448520 311160
rect 440936 311120 448520 311148
rect 440936 311108 440942 311120
rect 448514 311108 448520 311120
rect 448572 311108 448578 311160
rect 475746 311108 475752 311160
rect 475804 311148 475810 311160
rect 544378 311148 544384 311160
rect 475804 311120 544384 311148
rect 475804 311108 475810 311120
rect 544378 311108 544384 311120
rect 544436 311108 544442 311160
rect 458818 309816 458824 309868
rect 458876 309856 458882 309868
rect 488442 309856 488448 309868
rect 458876 309828 488448 309856
rect 458876 309816 458882 309828
rect 488442 309816 488448 309828
rect 488500 309816 488506 309868
rect 495894 309816 495900 309868
rect 495952 309856 495958 309868
rect 542446 309856 542452 309868
rect 495952 309828 542452 309856
rect 495952 309816 495958 309828
rect 542446 309816 542452 309828
rect 542504 309816 542510 309868
rect 476298 309748 476304 309800
rect 476356 309788 476362 309800
rect 537478 309788 537484 309800
rect 476356 309760 537484 309788
rect 476356 309748 476362 309760
rect 537478 309748 537484 309760
rect 537536 309748 537542 309800
rect 451918 308456 451924 308508
rect 451976 308496 451982 308508
rect 488718 308496 488724 308508
rect 451976 308468 488724 308496
rect 451976 308456 451982 308468
rect 488718 308456 488724 308468
rect 488776 308456 488782 308508
rect 496998 308456 497004 308508
rect 497056 308496 497062 308508
rect 539778 308496 539784 308508
rect 497056 308468 539784 308496
rect 497056 308456 497062 308468
rect 539778 308456 539784 308468
rect 539836 308456 539842 308508
rect 465258 308388 465264 308440
rect 465316 308428 465322 308440
rect 548518 308428 548524 308440
rect 465316 308400 548524 308428
rect 465316 308388 465322 308400
rect 548518 308388 548524 308400
rect 548576 308388 548582 308440
rect 3510 307708 3516 307760
rect 3568 307748 3574 307760
rect 4798 307748 4804 307760
rect 3568 307720 4804 307748
rect 3568 307708 3574 307720
rect 4798 307708 4804 307720
rect 4856 307708 4862 307760
rect 455874 307096 455880 307148
rect 455932 307136 455938 307148
rect 576118 307136 576124 307148
rect 455932 307108 576124 307136
rect 455932 307096 455938 307108
rect 576118 307096 576124 307108
rect 576176 307096 576182 307148
rect 383010 307028 383016 307080
rect 383068 307068 383074 307080
rect 520918 307068 520924 307080
rect 383068 307040 520924 307068
rect 383068 307028 383074 307040
rect 520918 307028 520924 307040
rect 520976 307028 520982 307080
rect 383102 306280 383108 306332
rect 383160 306320 383166 306332
rect 464706 306320 464712 306332
rect 383160 306292 464712 306320
rect 383160 306280 383166 306292
rect 464706 306280 464712 306292
rect 464764 306280 464770 306332
rect 381998 306212 382004 306264
rect 382056 306252 382062 306264
rect 463878 306252 463884 306264
rect 382056 306224 463884 306252
rect 382056 306212 382062 306224
rect 463878 306212 463884 306224
rect 463936 306212 463942 306264
rect 378870 306144 378876 306196
rect 378928 306184 378934 306196
rect 463602 306184 463608 306196
rect 378928 306156 463608 306184
rect 378928 306144 378934 306156
rect 463602 306144 463608 306156
rect 463660 306144 463666 306196
rect 384482 306076 384488 306128
rect 384540 306116 384546 306128
rect 474642 306116 474648 306128
rect 384540 306088 474648 306116
rect 384540 306076 384546 306088
rect 474642 306076 474648 306088
rect 474700 306076 474706 306128
rect 381906 306008 381912 306060
rect 381964 306048 381970 306060
rect 474366 306048 474372 306060
rect 381964 306020 474372 306048
rect 381964 306008 381970 306020
rect 474366 306008 474372 306020
rect 474424 306008 474430 306060
rect 382090 305940 382096 305992
rect 382148 305980 382154 305992
rect 474918 305980 474924 305992
rect 382148 305952 474924 305980
rect 382148 305940 382154 305952
rect 474918 305940 474924 305952
rect 474976 305940 474982 305992
rect 378962 305872 378968 305924
rect 379020 305912 379026 305924
rect 474090 305912 474096 305924
rect 379020 305884 474096 305912
rect 379020 305872 379026 305884
rect 474090 305872 474096 305884
rect 474148 305872 474154 305924
rect 475470 305872 475476 305924
rect 475528 305912 475534 305924
rect 562318 305912 562324 305924
rect 475528 305884 562324 305912
rect 475528 305872 475534 305884
rect 562318 305872 562324 305884
rect 562376 305872 562382 305924
rect 384758 305804 384764 305856
rect 384816 305844 384822 305856
rect 484854 305844 484860 305856
rect 384816 305816 484860 305844
rect 384816 305804 384822 305816
rect 484854 305804 484860 305816
rect 484912 305804 484918 305856
rect 384574 305736 384580 305788
rect 384632 305776 384638 305788
rect 485130 305776 485136 305788
rect 384632 305748 485136 305776
rect 384632 305736 384638 305748
rect 485130 305736 485136 305748
rect 485188 305736 485194 305788
rect 381814 305668 381820 305720
rect 381872 305708 381878 305720
rect 484578 305708 484584 305720
rect 381872 305680 484584 305708
rect 381872 305668 381878 305680
rect 484578 305668 484584 305680
rect 484636 305668 484642 305720
rect 362310 305600 362316 305652
rect 362368 305640 362374 305652
rect 516410 305640 516416 305652
rect 362368 305612 516416 305640
rect 362368 305600 362374 305612
rect 516410 305600 516416 305612
rect 516468 305600 516474 305652
rect 384390 305532 384396 305584
rect 384448 305572 384454 305584
rect 464430 305572 464436 305584
rect 384448 305544 464436 305572
rect 384448 305532 384454 305544
rect 464430 305532 464436 305544
rect 464488 305532 464494 305584
rect 384298 305464 384304 305516
rect 384356 305504 384362 305516
rect 464154 305504 464160 305516
rect 384356 305476 464160 305504
rect 384356 305464 384362 305476
rect 464154 305464 464160 305476
rect 464212 305464 464218 305516
rect 457530 305396 457536 305448
rect 457588 305436 457594 305448
rect 490650 305436 490656 305448
rect 457588 305408 490656 305436
rect 457588 305396 457594 305408
rect 490650 305396 490656 305408
rect 490708 305396 490714 305448
rect 361758 304920 361764 304972
rect 361816 304960 361822 304972
rect 435450 304960 435456 304972
rect 361816 304932 435456 304960
rect 361816 304920 361822 304932
rect 435450 304920 435456 304932
rect 435508 304920 435514 304972
rect 486234 304444 486240 304496
rect 486292 304484 486298 304496
rect 530026 304484 530032 304496
rect 486292 304456 530032 304484
rect 486292 304444 486298 304456
rect 530026 304444 530032 304456
rect 530084 304444 530090 304496
rect 385770 304376 385776 304428
rect 385828 304416 385834 304428
rect 520826 304416 520832 304428
rect 385828 304388 520832 304416
rect 385828 304376 385834 304388
rect 520826 304376 520832 304388
rect 520884 304376 520890 304428
rect 363598 304308 363604 304360
rect 363656 304348 363662 304360
rect 512730 304348 512736 304360
rect 363656 304320 512736 304348
rect 363656 304308 363662 304320
rect 512730 304308 512736 304320
rect 512788 304308 512794 304360
rect 360930 304240 360936 304292
rect 360988 304280 360994 304292
rect 512638 304280 512644 304292
rect 360988 304252 512644 304280
rect 360988 304240 360994 304252
rect 512638 304240 512644 304252
rect 512696 304240 512702 304292
rect 475378 303628 475384 303680
rect 475436 303668 475442 303680
rect 479518 303668 479524 303680
rect 475436 303640 479524 303668
rect 475436 303628 475442 303640
rect 479518 303628 479524 303640
rect 479576 303628 479582 303680
rect 378594 303560 378600 303612
rect 378652 303600 378658 303612
rect 484302 303600 484308 303612
rect 378652 303572 484308 303600
rect 378652 303560 378658 303572
rect 484302 303560 484308 303572
rect 484360 303560 484366 303612
rect 376662 303492 376668 303544
rect 376720 303532 376726 303544
rect 484026 303532 484032 303544
rect 376720 303504 484032 303532
rect 376720 303492 376726 303504
rect 484026 303492 484032 303504
rect 484084 303492 484090 303544
rect 379330 303424 379336 303476
rect 379388 303464 379394 303476
rect 510982 303464 510988 303476
rect 379388 303436 510988 303464
rect 379388 303424 379394 303436
rect 510982 303424 510988 303436
rect 511040 303424 511046 303476
rect 378686 303356 378692 303408
rect 378744 303396 378750 303408
rect 510890 303396 510896 303408
rect 378744 303368 510896 303396
rect 378744 303356 378750 303368
rect 510890 303356 510896 303368
rect 510948 303356 510954 303408
rect 379238 303288 379244 303340
rect 379296 303328 379302 303340
rect 513926 303328 513932 303340
rect 379296 303300 513932 303328
rect 379296 303288 379302 303300
rect 513926 303288 513932 303300
rect 513984 303288 513990 303340
rect 379422 303220 379428 303272
rect 379480 303260 379486 303272
rect 515214 303260 515220 303272
rect 379480 303232 515220 303260
rect 379480 303220 379486 303232
rect 515214 303220 515220 303232
rect 515272 303220 515278 303272
rect 376570 303152 376576 303204
rect 376628 303192 376634 303204
rect 513742 303192 513748 303204
rect 376628 303164 513748 303192
rect 376628 303152 376634 303164
rect 513742 303152 513748 303164
rect 513800 303152 513806 303204
rect 376386 303084 376392 303136
rect 376444 303124 376450 303136
rect 513834 303124 513840 303136
rect 376444 303096 513840 303124
rect 376444 303084 376450 303096
rect 513834 303084 513840 303096
rect 513892 303084 513898 303136
rect 376478 303016 376484 303068
rect 376536 303056 376542 303068
rect 515030 303056 515036 303068
rect 376536 303028 515036 303056
rect 376536 303016 376542 303028
rect 515030 303016 515036 303028
rect 515088 303016 515094 303068
rect 376294 302948 376300 303000
rect 376352 302988 376358 303000
rect 515122 302988 515128 303000
rect 376352 302960 515128 302988
rect 376352 302948 376358 302960
rect 515122 302948 515128 302960
rect 515180 302948 515186 303000
rect 364978 302880 364984 302932
rect 365036 302920 365042 302932
rect 512454 302920 512460 302932
rect 365036 302892 512460 302920
rect 365036 302880 365042 302892
rect 512454 302880 512460 302892
rect 512512 302880 512518 302932
rect 373626 302812 373632 302864
rect 373684 302852 373690 302864
rect 473538 302852 473544 302864
rect 373684 302824 473544 302852
rect 373684 302812 373690 302824
rect 473538 302812 473544 302824
rect 473596 302812 473602 302864
rect 476574 302812 476580 302864
rect 476632 302852 476638 302864
rect 547138 302852 547144 302864
rect 476632 302824 547144 302852
rect 476632 302812 476638 302824
rect 547138 302812 547144 302824
rect 547196 302812 547202 302864
rect 376018 302744 376024 302796
rect 376076 302784 376082 302796
rect 473814 302784 473820 302796
rect 376076 302756 473820 302784
rect 376076 302744 376082 302756
rect 473814 302744 473820 302756
rect 473872 302744 473878 302796
rect 375926 302676 375932 302728
rect 375984 302716 375990 302728
rect 463326 302716 463332 302728
rect 375984 302688 463332 302716
rect 375984 302676 375990 302688
rect 463326 302676 463332 302688
rect 463384 302676 463390 302728
rect 465534 301656 465540 301708
rect 465592 301696 465598 301708
rect 559558 301696 559564 301708
rect 465592 301668 559564 301696
rect 465592 301656 465598 301668
rect 559558 301656 559564 301668
rect 559616 301656 559622 301708
rect 408402 301588 408408 301640
rect 408460 301628 408466 301640
rect 503070 301628 503076 301640
rect 408460 301600 503076 301628
rect 408460 301588 408466 301600
rect 503070 301588 503076 301600
rect 503128 301588 503134 301640
rect 370498 301520 370504 301572
rect 370556 301560 370562 301572
rect 512270 301560 512276 301572
rect 370556 301532 512276 301560
rect 370556 301520 370562 301532
rect 512270 301520 512276 301532
rect 512328 301520 512334 301572
rect 367738 301452 367744 301504
rect 367796 301492 367802 301504
rect 512362 301492 512368 301504
rect 367796 301464 512368 301492
rect 367796 301452 367802 301464
rect 512362 301452 512368 301464
rect 512420 301452 512426 301504
rect 471238 301044 471244 301096
rect 471296 301084 471302 301096
rect 473262 301084 473268 301096
rect 471296 301056 473268 301084
rect 471296 301044 471302 301056
rect 473262 301044 473268 301056
rect 473320 301044 473326 301096
rect 373718 300772 373724 300824
rect 373776 300812 373782 300824
rect 510798 300812 510804 300824
rect 373776 300784 510804 300812
rect 373776 300772 373782 300784
rect 510798 300772 510804 300784
rect 510856 300772 510862 300824
rect 370774 300704 370780 300756
rect 370832 300744 370838 300756
rect 509878 300744 509884 300756
rect 370832 300716 509884 300744
rect 370832 300704 370838 300716
rect 509878 300704 509884 300716
rect 509936 300704 509942 300756
rect 370682 300636 370688 300688
rect 370740 300676 370746 300688
rect 510614 300676 510620 300688
rect 370740 300648 510620 300676
rect 370740 300636 370746 300648
rect 510614 300636 510620 300648
rect 510672 300636 510678 300688
rect 367922 300568 367928 300620
rect 367980 300608 367986 300620
rect 509694 300608 509700 300620
rect 367980 300580 509700 300608
rect 367980 300568 367986 300580
rect 509694 300568 509700 300580
rect 509752 300568 509758 300620
rect 370866 300500 370872 300552
rect 370924 300540 370930 300552
rect 513650 300540 513656 300552
rect 370924 300512 513656 300540
rect 370924 300500 370930 300512
rect 513650 300500 513656 300512
rect 513708 300500 513714 300552
rect 370958 300432 370964 300484
rect 371016 300472 371022 300484
rect 514846 300472 514852 300484
rect 371016 300444 514852 300472
rect 371016 300432 371022 300444
rect 514846 300432 514852 300444
rect 514904 300432 514910 300484
rect 368106 300364 368112 300416
rect 368164 300404 368170 300416
rect 513558 300404 513564 300416
rect 368164 300376 513564 300404
rect 368164 300364 368170 300376
rect 513558 300364 513564 300376
rect 513616 300364 513622 300416
rect 368014 300296 368020 300348
rect 368072 300336 368078 300348
rect 516502 300336 516508 300348
rect 368072 300308 516508 300336
rect 368072 300296 368078 300308
rect 516502 300296 516508 300308
rect 516560 300296 516566 300348
rect 361022 300228 361028 300280
rect 361080 300268 361086 300280
rect 511994 300268 512000 300280
rect 361080 300240 512000 300268
rect 361080 300228 361086 300240
rect 511994 300228 512000 300240
rect 512052 300228 512058 300280
rect 365346 300160 365352 300212
rect 365404 300200 365410 300212
rect 516318 300200 516324 300212
rect 365404 300172 516324 300200
rect 365404 300160 365410 300172
rect 516318 300160 516324 300172
rect 516376 300160 516382 300212
rect 365254 300092 365260 300144
rect 365312 300132 365318 300144
rect 517514 300132 517520 300144
rect 365312 300104 517520 300132
rect 365312 300092 365318 300104
rect 517514 300092 517520 300104
rect 517572 300092 517578 300144
rect 373442 300024 373448 300076
rect 373500 300064 373506 300076
rect 509970 300064 509976 300076
rect 373500 300036 509976 300064
rect 373500 300024 373506 300036
rect 509970 300024 509976 300036
rect 510028 300024 510034 300076
rect 373534 299956 373540 300008
rect 373592 299996 373598 300008
rect 510338 299996 510344 300008
rect 373592 299968 510344 299996
rect 373592 299956 373598 299968
rect 510338 299956 510344 299968
rect 510396 299956 510402 300008
rect 466086 299888 466092 299940
rect 466144 299928 466150 299940
rect 551278 299928 551284 299940
rect 466144 299900 551284 299928
rect 466144 299888 466150 299900
rect 551278 299888 551284 299900
rect 551336 299888 551342 299940
rect 461578 299412 461584 299464
rect 461636 299452 461642 299464
rect 580166 299452 580172 299464
rect 461636 299424 580172 299452
rect 461636 299412 461642 299424
rect 580166 299412 580172 299424
rect 580224 299412 580230 299464
rect 403618 298800 403624 298852
rect 403676 298840 403682 298852
rect 502794 298840 502800 298852
rect 403676 298812 502800 298840
rect 403676 298800 403682 298812
rect 502794 298800 502800 298812
rect 502852 298800 502858 298852
rect 381630 298732 381636 298784
rect 381688 298772 381694 298784
rect 485682 298772 485688 298784
rect 381688 298744 485688 298772
rect 381688 298732 381694 298744
rect 485682 298732 485688 298744
rect 485740 298732 485746 298784
rect 454954 298052 454960 298104
rect 455012 298092 455018 298104
rect 566458 298092 566464 298104
rect 455012 298064 566464 298092
rect 455012 298052 455018 298064
rect 566458 298052 566464 298064
rect 566516 298052 566522 298104
rect 382918 297984 382924 298036
rect 382976 298024 382982 298036
rect 519354 298024 519360 298036
rect 382976 297996 519360 298024
rect 382976 297984 382982 297996
rect 519354 297984 519360 297996
rect 519412 297984 519418 298036
rect 370590 297916 370596 297968
rect 370648 297956 370654 297968
rect 518066 297956 518072 297968
rect 370648 297928 518072 297956
rect 370648 297916 370654 297928
rect 518066 297916 518072 297928
rect 518124 297916 518130 297968
rect 369210 297848 369216 297900
rect 369268 297888 369274 297900
rect 518250 297888 518256 297900
rect 369268 297860 518256 297888
rect 369268 297848 369274 297860
rect 518250 297848 518256 297860
rect 518308 297848 518314 297900
rect 361114 297780 361120 297832
rect 361172 297820 361178 297832
rect 512178 297820 512184 297832
rect 361172 297792 512184 297820
rect 361172 297780 361178 297792
rect 512178 297780 512184 297792
rect 512236 297780 512242 297832
rect 363966 297712 363972 297764
rect 364024 297752 364030 297764
rect 515306 297752 515312 297764
rect 364024 297724 515312 297752
rect 364024 297712 364030 297724
rect 515306 297712 515312 297724
rect 515364 297712 515370 297764
rect 366542 297644 366548 297696
rect 366600 297684 366606 297696
rect 518342 297684 518348 297696
rect 366600 297656 518348 297684
rect 366600 297644 366606 297656
rect 518342 297644 518348 297656
rect 518400 297644 518406 297696
rect 365070 297576 365076 297628
rect 365128 297616 365134 297628
rect 516870 297616 516876 297628
rect 365128 297588 516876 297616
rect 365128 297576 365134 297588
rect 516870 297576 516876 297588
rect 516928 297576 516934 297628
rect 362402 297508 362408 297560
rect 362460 297548 362466 297560
rect 515582 297548 515588 297560
rect 362460 297520 515588 297548
rect 362460 297508 362466 297520
rect 515582 297508 515588 297520
rect 515640 297508 515646 297560
rect 366450 297440 366456 297492
rect 366508 297480 366514 297492
rect 519722 297480 519728 297492
rect 366508 297452 519728 297480
rect 366508 297440 366514 297452
rect 519722 297440 519728 297452
rect 519780 297440 519786 297492
rect 362494 297372 362500 297424
rect 362552 297412 362558 297424
rect 516226 297412 516232 297424
rect 362552 297384 516232 297412
rect 362552 297372 362558 297384
rect 516226 297372 516232 297384
rect 516284 297372 516290 297424
rect 454770 295944 454776 295996
rect 454828 295984 454834 295996
rect 573358 295984 573364 295996
rect 454828 295956 573364 295984
rect 454828 295944 454834 295956
rect 573358 295944 573364 295956
rect 573416 295944 573422 295996
rect 435358 295332 435364 295384
rect 435416 295372 435422 295384
rect 440878 295372 440884 295384
rect 435416 295344 440884 295372
rect 435416 295332 435422 295344
rect 440878 295332 440884 295344
rect 440936 295332 440942 295384
rect 469858 295332 469864 295384
rect 469916 295372 469922 295384
rect 471238 295372 471244 295384
rect 469916 295344 471244 295372
rect 469916 295332 469922 295344
rect 471238 295332 471244 295344
rect 471296 295332 471302 295384
rect 374638 295264 374644 295316
rect 374696 295304 374702 295316
rect 507578 295304 507584 295316
rect 374696 295276 507584 295304
rect 374696 295264 374702 295276
rect 507578 295264 507584 295276
rect 507636 295264 507642 295316
rect 379146 295196 379152 295248
rect 379204 295236 379210 295248
rect 514202 295236 514208 295248
rect 379204 295208 514208 295236
rect 379204 295196 379210 295208
rect 514202 295196 514208 295208
rect 514260 295196 514266 295248
rect 372062 295128 372068 295180
rect 372120 295168 372126 295180
rect 509786 295168 509792 295180
rect 372120 295140 509792 295168
rect 372120 295128 372126 295140
rect 509786 295128 509792 295140
rect 509844 295128 509850 295180
rect 371970 295060 371976 295112
rect 372028 295100 372034 295112
rect 510706 295100 510712 295112
rect 372028 295072 510712 295100
rect 372028 295060 372034 295072
rect 510706 295060 510712 295072
rect 510764 295060 510770 295112
rect 375098 294992 375104 295044
rect 375156 295032 375162 295044
rect 517606 295032 517612 295044
rect 375156 295004 517612 295032
rect 375156 294992 375162 295004
rect 517606 294992 517612 295004
rect 517664 294992 517670 295044
rect 375006 294924 375012 294976
rect 375064 294964 375070 294976
rect 517698 294964 517704 294976
rect 375064 294936 517704 294964
rect 375064 294924 375070 294936
rect 517698 294924 517704 294936
rect 517756 294924 517762 294976
rect 377582 294856 377588 294908
rect 377640 294896 377646 294908
rect 520550 294896 520556 294908
rect 377640 294868 520556 294896
rect 377640 294856 377646 294868
rect 520550 294856 520556 294868
rect 520608 294856 520614 294908
rect 373350 294788 373356 294840
rect 373408 294828 373414 294840
rect 517974 294828 517980 294840
rect 373408 294800 517980 294828
rect 373408 294788 373414 294800
rect 517974 294788 517980 294800
rect 518032 294788 518038 294840
rect 372338 294720 372344 294772
rect 372396 294760 372402 294772
rect 519170 294760 519176 294772
rect 372396 294732 519176 294760
rect 372396 294720 372402 294732
rect 519170 294720 519176 294732
rect 519228 294720 519234 294772
rect 371878 294652 371884 294704
rect 371936 294692 371942 294704
rect 518986 294692 518992 294704
rect 371936 294664 518992 294692
rect 371936 294652 371942 294664
rect 518986 294652 518992 294664
rect 519044 294652 519050 294704
rect 369394 294584 369400 294636
rect 369452 294624 369458 294636
rect 516686 294624 516692 294636
rect 369452 294596 516692 294624
rect 369452 294584 369458 294596
rect 516686 294584 516692 294596
rect 516744 294584 516750 294636
rect 374914 294516 374920 294568
rect 374972 294556 374978 294568
rect 507670 294556 507676 294568
rect 374972 294528 507676 294556
rect 374972 294516 374978 294528
rect 507670 294516 507676 294528
rect 507728 294516 507734 294568
rect 376202 294448 376208 294500
rect 376260 294488 376266 294500
rect 507762 294488 507768 294500
rect 376260 294460 507768 294488
rect 376260 294448 376266 294460
rect 507762 294448 507768 294460
rect 507820 294448 507826 294500
rect 455046 294380 455052 294432
rect 455104 294420 455110 294432
rect 570598 294420 570604 294432
rect 455104 294392 570604 294420
rect 455104 294380 455110 294392
rect 570598 294380 570604 294392
rect 570656 294380 570662 294432
rect 361758 293904 361764 293956
rect 361816 293944 361822 293956
rect 436830 293944 436836 293956
rect 361816 293916 436836 293944
rect 361816 293904 361822 293916
rect 436830 293904 436836 293916
rect 436888 293904 436894 293956
rect 476850 293224 476856 293276
rect 476908 293264 476914 293276
rect 558178 293264 558184 293276
rect 476908 293236 558184 293264
rect 476908 293224 476914 293236
rect 558178 293224 558184 293236
rect 558236 293224 558242 293276
rect 3418 292544 3424 292596
rect 3476 292584 3482 292596
rect 4890 292584 4896 292596
rect 3476 292556 4896 292584
rect 3476 292544 3482 292556
rect 4890 292544 4896 292556
rect 4948 292544 4954 292596
rect 383470 292476 383476 292528
rect 383528 292516 383534 292528
rect 507486 292516 507492 292528
rect 383528 292488 507492 292516
rect 383528 292476 383534 292488
rect 507486 292476 507492 292488
rect 507544 292476 507550 292528
rect 386046 292408 386052 292460
rect 386104 292448 386110 292460
rect 520274 292448 520280 292460
rect 386104 292420 520280 292448
rect 386104 292408 386110 292420
rect 520274 292408 520280 292420
rect 520332 292408 520338 292460
rect 380434 292340 380440 292392
rect 380492 292380 380498 292392
rect 514754 292380 514760 292392
rect 380492 292352 514760 292380
rect 380492 292340 380498 292352
rect 514754 292340 514760 292352
rect 514812 292340 514818 292392
rect 381354 292272 381360 292324
rect 381412 292312 381418 292324
rect 516962 292312 516968 292324
rect 381412 292284 516968 292312
rect 381412 292272 381418 292284
rect 516962 292272 516968 292284
rect 517020 292272 517026 292324
rect 377766 292204 377772 292256
rect 377824 292244 377830 292256
rect 514110 292244 514116 292256
rect 377824 292216 514116 292244
rect 377824 292204 377830 292216
rect 514110 292204 514116 292216
rect 514168 292204 514174 292256
rect 383378 292136 383384 292188
rect 383436 292176 383442 292188
rect 520366 292176 520372 292188
rect 383436 292148 520372 292176
rect 383436 292136 383442 292148
rect 520366 292136 520372 292148
rect 520424 292136 520430 292188
rect 380526 292068 380532 292120
rect 380584 292108 380590 292120
rect 520458 292108 520464 292120
rect 380584 292080 520464 292108
rect 380584 292068 380590 292080
rect 520458 292068 520464 292080
rect 520516 292068 520522 292120
rect 369118 292000 369124 292052
rect 369176 292040 369182 292052
rect 516778 292040 516784 292052
rect 369176 292012 516784 292040
rect 369176 292000 369182 292012
rect 516778 292000 516784 292012
rect 516836 292000 516842 292052
rect 366358 291932 366364 291984
rect 366416 291972 366422 291984
rect 519262 291972 519268 291984
rect 366416 291944 519268 291972
rect 366416 291932 366422 291944
rect 519262 291932 519268 291944
rect 519320 291932 519326 291984
rect 363874 291864 363880 291916
rect 363932 291904 363938 291916
rect 520734 291904 520740 291916
rect 363932 291876 520740 291904
rect 363932 291864 363938 291876
rect 520734 291864 520740 291876
rect 520792 291864 520798 291916
rect 361206 291796 361212 291848
rect 361264 291836 361270 291848
rect 519446 291836 519452 291848
rect 361264 291808 519452 291836
rect 361264 291796 361270 291808
rect 519446 291796 519452 291808
rect 519504 291796 519510 291848
rect 385862 291728 385868 291780
rect 385920 291768 385926 291780
rect 507394 291768 507400 291780
rect 385920 291740 507400 291768
rect 385920 291728 385926 291740
rect 507394 291728 507400 291740
rect 507452 291728 507458 291780
rect 456150 291660 456156 291712
rect 456208 291700 456214 291712
rect 572070 291700 572076 291712
rect 456208 291672 572076 291700
rect 456208 291660 456214 291672
rect 572070 291660 572076 291672
rect 572128 291660 572134 291712
rect 454954 290504 454960 290556
rect 455012 290544 455018 290556
rect 485866 290544 485872 290556
rect 455012 290516 485872 290544
rect 455012 290504 455018 290516
rect 485866 290504 485872 290516
rect 485924 290504 485930 290556
rect 476022 290436 476028 290488
rect 476080 290476 476086 290488
rect 569218 290476 569224 290488
rect 476080 290448 569224 290476
rect 476080 290436 476086 290448
rect 569218 290436 569224 290448
rect 569276 290436 569282 290488
rect 374822 289756 374828 289808
rect 374880 289796 374886 289808
rect 507118 289796 507124 289808
rect 374880 289768 507124 289796
rect 374880 289756 374886 289768
rect 507118 289756 507124 289768
rect 507176 289756 507182 289808
rect 383194 289688 383200 289740
rect 383252 289728 383258 289740
rect 517790 289728 517796 289740
rect 383252 289700 517796 289728
rect 383252 289688 383258 289700
rect 517790 289688 517796 289700
rect 517848 289688 517854 289740
rect 385954 289620 385960 289672
rect 386012 289660 386018 289672
rect 521838 289660 521844 289672
rect 386012 289632 521844 289660
rect 386012 289620 386018 289632
rect 521838 289620 521844 289632
rect 521896 289620 521902 289672
rect 380342 289552 380348 289604
rect 380400 289592 380406 289604
rect 516594 289592 516600 289604
rect 380400 289564 516600 289592
rect 380400 289552 380406 289564
rect 516594 289552 516600 289564
rect 516652 289552 516658 289604
rect 382182 289484 382188 289536
rect 382240 289524 382246 289536
rect 518894 289524 518900 289536
rect 382240 289496 518900 289524
rect 382240 289484 382246 289496
rect 518894 289484 518900 289496
rect 518952 289484 518958 289536
rect 377490 289416 377496 289468
rect 377548 289456 377554 289468
rect 514938 289456 514944 289468
rect 377548 289428 514944 289456
rect 377548 289416 377554 289428
rect 514938 289416 514944 289428
rect 514996 289416 515002 289468
rect 377674 289348 377680 289400
rect 377732 289388 377738 289400
rect 519078 289388 519084 289400
rect 377732 289360 519084 289388
rect 377732 289348 377738 289360
rect 519078 289348 519084 289360
rect 519136 289348 519142 289400
rect 380250 289280 380256 289332
rect 380308 289320 380314 289332
rect 523310 289320 523316 289332
rect 380308 289292 523316 289320
rect 380308 289280 380314 289292
rect 523310 289280 523316 289292
rect 523368 289280 523374 289332
rect 379054 289212 379060 289264
rect 379112 289252 379118 289264
rect 523218 289252 523224 289264
rect 379112 289224 523224 289252
rect 379112 289212 379118 289224
rect 523218 289212 523224 289224
rect 523276 289212 523282 289264
rect 376110 289144 376116 289196
rect 376168 289184 376174 289196
rect 521746 289184 521752 289196
rect 376168 289156 521752 289184
rect 376168 289144 376174 289156
rect 521746 289144 521752 289156
rect 521804 289144 521810 289196
rect 372246 289076 372252 289128
rect 372304 289116 372310 289128
rect 520642 289116 520648 289128
rect 372304 289088 520648 289116
rect 372304 289076 372310 289088
rect 520642 289076 520648 289088
rect 520700 289076 520706 289128
rect 383286 289008 383292 289060
rect 383344 289048 383350 289060
rect 507210 289048 507216 289060
rect 383344 289020 507216 289048
rect 383344 289008 383350 289020
rect 507210 289008 507216 289020
rect 507268 289008 507274 289060
rect 384666 288940 384672 288992
rect 384724 288980 384730 288992
rect 507302 288980 507308 288992
rect 384724 288952 507308 288980
rect 384724 288940 384730 288952
rect 507302 288940 507308 288952
rect 507360 288940 507366 288992
rect 450354 288872 450360 288924
rect 450412 288912 450418 288924
rect 455138 288912 455144 288924
rect 450412 288884 455144 288912
rect 450412 288872 450418 288884
rect 455138 288872 455144 288884
rect 455196 288872 455202 288924
rect 455322 288872 455328 288924
rect 455380 288912 455386 288924
rect 574738 288912 574744 288924
rect 455380 288884 574744 288912
rect 455380 288872 455386 288884
rect 574738 288872 574744 288884
rect 574796 288872 574802 288924
rect 502242 287716 502248 287768
rect 502300 287756 502306 287768
rect 538950 287756 538956 287768
rect 502300 287728 538956 287756
rect 502300 287716 502306 287728
rect 538950 287716 538956 287728
rect 539008 287716 539014 287768
rect 451182 287648 451188 287700
rect 451240 287688 451246 287700
rect 505002 287688 505008 287700
rect 451240 287660 505008 287688
rect 451240 287648 451246 287660
rect 505002 287648 505008 287660
rect 505060 287648 505066 287700
rect 452102 286628 452108 286680
rect 452160 286668 452166 286680
rect 487890 286668 487896 286680
rect 452160 286640 487896 286668
rect 452160 286628 452166 286640
rect 487890 286628 487896 286640
rect 487948 286628 487954 286680
rect 378778 286560 378784 286612
rect 378836 286600 378842 286612
rect 475194 286600 475200 286612
rect 378836 286572 475200 286600
rect 378836 286560 378842 286572
rect 475194 286560 475200 286572
rect 475252 286560 475258 286612
rect 486510 286560 486516 286612
rect 486568 286600 486574 286612
rect 531314 286600 531320 286612
rect 486568 286572 531320 286600
rect 486568 286560 486574 286572
rect 531314 286560 531320 286572
rect 531372 286560 531378 286612
rect 464982 286492 464988 286544
rect 465040 286532 465046 286544
rect 571978 286532 571984 286544
rect 465040 286504 571984 286532
rect 465040 286492 465046 286504
rect 571978 286492 571984 286504
rect 572036 286492 572042 286544
rect 372154 286424 372160 286476
rect 372212 286464 372218 286476
rect 523034 286464 523040 286476
rect 372212 286436 523040 286464
rect 372212 286424 372218 286436
rect 523034 286424 523040 286436
rect 523092 286424 523098 286476
rect 369302 286356 369308 286408
rect 369360 286396 369366 286408
rect 521654 286396 521660 286408
rect 369360 286368 521660 286396
rect 369360 286356 369366 286368
rect 521654 286356 521660 286368
rect 521712 286356 521718 286408
rect 366634 286288 366640 286340
rect 366692 286328 366698 286340
rect 523126 286328 523132 286340
rect 366692 286300 523132 286328
rect 366692 286288 366698 286300
rect 523126 286288 523132 286300
rect 523184 286288 523190 286340
rect 455046 284996 455052 285048
rect 455104 285036 455110 285048
rect 494514 285036 494520 285048
rect 455104 285008 494520 285036
rect 455104 284996 455110 285008
rect 494514 284996 494520 285008
rect 494572 284996 494578 285048
rect 449802 284928 449808 284980
rect 449860 284968 449866 284980
rect 536834 284968 536840 284980
rect 449860 284940 536840 284968
rect 449860 284928 449866 284940
rect 536834 284928 536840 284940
rect 536892 284928 536898 284980
rect 453574 283636 453580 283688
rect 453632 283676 453638 283688
rect 493962 283676 493968 283688
rect 453632 283648 493968 283676
rect 453632 283636 453638 283648
rect 493962 283636 493968 283648
rect 494020 283636 494026 283688
rect 501414 283636 501420 283688
rect 501472 283676 501478 283688
rect 540238 283676 540244 283688
rect 501472 283648 540244 283676
rect 501472 283636 501478 283648
rect 540238 283636 540244 283648
rect 540296 283636 540302 283688
rect 477218 283568 477224 283620
rect 477276 283608 477282 283620
rect 580258 283608 580264 283620
rect 477276 283580 580264 283608
rect 477276 283568 477282 283580
rect 580258 283568 580264 283580
rect 580316 283568 580322 283620
rect 361758 282820 361764 282872
rect 361816 282860 361822 282872
rect 439682 282860 439688 282872
rect 361816 282832 439688 282860
rect 361816 282820 361822 282832
rect 439682 282820 439688 282832
rect 439740 282820 439746 282872
rect 459278 282140 459284 282192
rect 459336 282180 459342 282192
rect 492306 282180 492312 282192
rect 459336 282152 492312 282180
rect 459336 282140 459342 282152
rect 492306 282140 492312 282152
rect 492364 282140 492370 282192
rect 432598 282072 432604 282124
rect 432656 282112 432662 282124
rect 435358 282112 435364 282124
rect 432656 282084 435364 282112
rect 432656 282072 432662 282084
rect 435358 282072 435364 282084
rect 435416 282072 435422 282124
rect 452378 280848 452384 280900
rect 452436 280888 452442 280900
rect 493134 280888 493140 280900
rect 452436 280860 493140 280888
rect 452436 280848 452442 280860
rect 493134 280848 493140 280860
rect 493192 280848 493198 280900
rect 500862 280848 500868 280900
rect 500920 280888 500926 280900
rect 540146 280888 540152 280900
rect 500920 280860 540152 280888
rect 500920 280848 500926 280860
rect 540146 280848 540152 280860
rect 540204 280848 540210 280900
rect 458082 280780 458088 280832
rect 458140 280820 458146 280832
rect 505278 280820 505284 280832
rect 458140 280792 505284 280820
rect 458140 280780 458146 280792
rect 505278 280780 505284 280792
rect 505336 280780 505342 280832
rect 453666 279420 453672 279472
rect 453724 279460 453730 279472
rect 493686 279460 493692 279472
rect 453724 279432 493692 279460
rect 453724 279420 453730 279432
rect 493686 279420 493692 279432
rect 493744 279420 493750 279472
rect 471974 279012 471980 279064
rect 472032 279052 472038 279064
rect 475378 279052 475384 279064
rect 472032 279024 475384 279052
rect 472032 279012 472038 279024
rect 475378 279012 475384 279024
rect 475436 279012 475442 279064
rect 457622 277992 457628 278044
rect 457680 278032 457686 278044
rect 493410 278032 493416 278044
rect 457680 278004 493416 278032
rect 457680 277992 457686 278004
rect 493410 277992 493416 278004
rect 493468 277992 493474 278044
rect 499206 277992 499212 278044
rect 499264 278032 499270 278044
rect 541434 278032 541440 278044
rect 499264 278004 541440 278032
rect 499264 277992 499270 278004
rect 541434 277992 541440 278004
rect 541492 277992 541498 278044
rect 467098 277380 467104 277432
rect 467156 277420 467162 277432
rect 472618 277420 472624 277432
rect 467156 277392 472624 277420
rect 467156 277380 467162 277392
rect 472618 277380 472624 277392
rect 472676 277380 472682 277432
rect 466454 276836 466460 276888
rect 466512 276876 466518 276888
rect 471974 276876 471980 276888
rect 466512 276848 471980 276876
rect 466512 276836 466518 276848
rect 471974 276836 471980 276848
rect 472032 276836 472038 276888
rect 456426 276700 456432 276752
rect 456484 276740 456490 276752
rect 492030 276740 492036 276752
rect 456484 276712 492036 276740
rect 456484 276700 456490 276712
rect 492030 276700 492036 276712
rect 492088 276700 492094 276752
rect 375834 276632 375840 276684
rect 375892 276672 375898 276684
rect 485406 276672 485412 276684
rect 375892 276644 485412 276672
rect 375892 276632 375898 276644
rect 485406 276632 485412 276644
rect 485464 276632 485470 276684
rect 497734 276632 497740 276684
rect 497792 276672 497798 276684
rect 541342 276672 541348 276684
rect 497792 276644 541348 276672
rect 497792 276632 497798 276644
rect 541342 276632 541348 276644
rect 541400 276632 541406 276684
rect 453482 275340 453488 275392
rect 453540 275380 453546 275392
rect 488166 275380 488172 275392
rect 453540 275352 488172 275380
rect 453540 275340 453546 275352
rect 488166 275340 488172 275352
rect 488224 275340 488230 275392
rect 500494 275340 500500 275392
rect 500552 275380 500558 275392
rect 540330 275380 540336 275392
rect 500552 275352 540336 275380
rect 500552 275340 500558 275352
rect 540330 275340 540336 275352
rect 540388 275340 540394 275392
rect 454862 275272 454868 275324
rect 454920 275312 454926 275324
rect 491202 275312 491208 275324
rect 454920 275284 491208 275312
rect 454920 275272 454926 275284
rect 491202 275272 491208 275284
rect 491260 275272 491266 275324
rect 497826 275272 497832 275324
rect 497884 275312 497890 275324
rect 541250 275312 541256 275324
rect 497884 275284 541256 275312
rect 497884 275272 497890 275284
rect 541250 275272 541256 275284
rect 541308 275272 541314 275324
rect 429194 274592 429200 274644
rect 429252 274632 429258 274644
rect 432598 274632 432604 274644
rect 429252 274604 432604 274632
rect 429252 274592 429258 274604
rect 432598 274592 432604 274604
rect 432656 274592 432662 274644
rect 459186 273980 459192 274032
rect 459244 274020 459250 274032
rect 487338 274020 487344 274032
rect 459244 273992 487344 274020
rect 459244 273980 459250 273992
rect 487338 273980 487344 273992
rect 487396 273980 487402 274032
rect 498930 273980 498936 274032
rect 498988 274020 498994 274032
rect 540054 274020 540060 274032
rect 498988 273992 540060 274020
rect 498988 273980 498994 273992
rect 540054 273980 540060 273992
rect 540112 273980 540118 274032
rect 456334 273912 456340 273964
rect 456392 273952 456398 273964
rect 490926 273952 490932 273964
rect 456392 273924 490932 273952
rect 456392 273912 456398 273924
rect 490926 273912 490932 273924
rect 490984 273912 490990 273964
rect 497550 273912 497556 273964
rect 497608 273952 497614 273964
rect 541158 273952 541164 273964
rect 497608 273924 541164 273952
rect 497608 273912 497614 273924
rect 541158 273912 541164 273924
rect 541216 273912 541222 273964
rect 462222 273232 462228 273284
rect 462280 273272 462286 273284
rect 466454 273272 466460 273284
rect 462280 273244 466460 273272
rect 462280 273232 462286 273244
rect 466454 273232 466460 273244
rect 466512 273232 466518 273284
rect 454770 272552 454776 272604
rect 454828 272592 454834 272604
rect 487614 272592 487620 272604
rect 454828 272564 487620 272592
rect 454828 272552 454834 272564
rect 487614 272552 487620 272564
rect 487672 272552 487678 272604
rect 498378 272552 498384 272604
rect 498436 272592 498442 272604
rect 539962 272592 539968 272604
rect 498436 272564 539968 272592
rect 498436 272552 498442 272564
rect 539962 272552 539968 272564
rect 540020 272552 540026 272604
rect 456242 272484 456248 272536
rect 456300 272524 456306 272536
rect 490374 272524 490380 272536
rect 456300 272496 490380 272524
rect 456300 272484 456306 272496
rect 490374 272484 490380 272496
rect 490432 272484 490438 272536
rect 496170 272484 496176 272536
rect 496228 272524 496234 272536
rect 542998 272524 543004 272536
rect 496228 272496 543004 272524
rect 496228 272484 496234 272496
rect 542998 272484 543004 272496
rect 543056 272484 543062 272536
rect 361758 271804 361764 271856
rect 361816 271844 361822 271856
rect 438118 271844 438124 271856
rect 361816 271816 438124 271844
rect 361816 271804 361822 271816
rect 438118 271804 438124 271816
rect 438176 271804 438182 271856
rect 452286 271192 452292 271244
rect 452344 271232 452350 271244
rect 489822 271232 489828 271244
rect 452344 271204 489828 271232
rect 452344 271192 452350 271204
rect 489822 271192 489828 271204
rect 489880 271192 489886 271244
rect 495066 271192 495072 271244
rect 495124 271232 495130 271244
rect 542814 271232 542820 271244
rect 495124 271204 542820 271232
rect 495124 271192 495130 271204
rect 542814 271192 542820 271204
rect 542872 271192 542878 271244
rect 466638 271124 466644 271176
rect 466696 271164 466702 271176
rect 580350 271164 580356 271176
rect 466696 271136 580356 271164
rect 466696 271124 466702 271136
rect 580350 271124 580356 271136
rect 580408 271124 580414 271176
rect 456518 270920 456524 270972
rect 456576 270960 456582 270972
rect 462222 270960 462228 270972
rect 456576 270932 462228 270960
rect 456576 270920 456582 270932
rect 462222 270920 462228 270932
rect 462280 270920 462286 270972
rect 465810 269832 465816 269884
rect 465868 269872 465874 269884
rect 555418 269872 555424 269884
rect 465868 269844 555424 269872
rect 465868 269832 465874 269844
rect 555418 269832 555424 269844
rect 555476 269832 555482 269884
rect 450446 269764 450452 269816
rect 450504 269804 450510 269816
rect 457806 269804 457812 269816
rect 450504 269776 457812 269804
rect 450504 269764 450510 269776
rect 457806 269764 457812 269776
rect 457864 269764 457870 269816
rect 466362 269764 466368 269816
rect 466420 269804 466426 269816
rect 580258 269804 580264 269816
rect 466420 269776 580264 269804
rect 466420 269764 466426 269776
rect 580258 269764 580264 269776
rect 580316 269764 580322 269816
rect 427078 269016 427084 269068
rect 427136 269056 427142 269068
rect 429194 269056 429200 269068
rect 427136 269028 429200 269056
rect 427136 269016 427142 269028
rect 429194 269016 429200 269028
rect 429252 269016 429258 269068
rect 449894 268540 449900 268592
rect 449952 268580 449958 268592
rect 469858 268580 469864 268592
rect 449952 268552 469864 268580
rect 449952 268540 449958 268552
rect 469858 268540 469864 268552
rect 469916 268540 469922 268592
rect 442258 268472 442264 268524
rect 442316 268512 442322 268524
rect 467098 268512 467104 268524
rect 442316 268484 467104 268512
rect 442316 268472 442322 268484
rect 467098 268472 467104 268484
rect 467156 268472 467162 268524
rect 486878 268472 486884 268524
rect 486936 268512 486942 268524
rect 531222 268512 531228 268524
rect 486936 268484 531228 268512
rect 486936 268472 486942 268484
rect 531222 268472 531228 268484
rect 531280 268472 531286 268524
rect 456150 268404 456156 268456
rect 456208 268444 456214 268456
rect 489270 268444 489276 268456
rect 456208 268416 489276 268444
rect 456208 268404 456214 268416
rect 489270 268404 489276 268416
rect 489328 268404 489334 268456
rect 495342 268404 495348 268456
rect 495400 268444 495406 268456
rect 542906 268444 542912 268456
rect 495400 268416 542912 268444
rect 495400 268404 495406 268416
rect 542906 268404 542912 268416
rect 542964 268404 542970 268456
rect 450906 268336 450912 268388
rect 450964 268376 450970 268388
rect 504726 268376 504732 268388
rect 450964 268348 504732 268376
rect 450964 268336 450970 268348
rect 504726 268336 504732 268348
rect 504784 268336 504790 268388
rect 443178 266976 443184 267028
rect 443236 267016 443242 267028
rect 456518 267016 456524 267028
rect 443236 266988 456524 267016
rect 443236 266976 443242 266988
rect 456518 266976 456524 266988
rect 456576 266976 456582 267028
rect 449158 263508 449164 263560
rect 449216 263548 449222 263560
rect 456794 263548 456800 263560
rect 449216 263520 456800 263548
rect 449216 263508 449222 263520
rect 456794 263508 456800 263520
rect 456852 263508 456858 263560
rect 438118 261808 438124 261860
rect 438176 261848 438182 261860
rect 443178 261848 443184 261860
rect 438176 261820 443184 261848
rect 438176 261808 438182 261820
rect 443178 261808 443184 261820
rect 443236 261808 443242 261860
rect 361758 260788 361764 260840
rect 361816 260828 361822 260840
rect 399478 260828 399484 260840
rect 361816 260800 399484 260828
rect 361816 260788 361822 260800
rect 399478 260788 399484 260800
rect 399536 260788 399542 260840
rect 447778 260788 447784 260840
rect 447836 260828 447842 260840
rect 449802 260828 449808 260840
rect 447836 260800 449808 260828
rect 447836 260788 447842 260800
rect 449802 260788 449808 260800
rect 449860 260788 449866 260840
rect 431310 258680 431316 258732
rect 431368 258720 431374 258732
rect 455230 258720 455236 258732
rect 431368 258692 455236 258720
rect 431368 258680 431374 258692
rect 455230 258680 455236 258692
rect 455288 258680 455294 258732
rect 3970 253920 3976 253972
rect 4028 253960 4034 253972
rect 5074 253960 5080 253972
rect 4028 253932 5080 253960
rect 4028 253920 4034 253932
rect 5074 253920 5080 253932
rect 5132 253920 5138 253972
rect 421558 250452 421564 250504
rect 421616 250492 421622 250504
rect 427078 250492 427084 250504
rect 421616 250464 427084 250492
rect 421616 250452 421622 250464
rect 427078 250452 427084 250464
rect 427136 250452 427142 250504
rect 361758 249704 361764 249756
rect 361816 249744 361822 249756
rect 443730 249744 443736 249756
rect 361816 249716 443736 249744
rect 361816 249704 361822 249716
rect 443730 249704 443736 249716
rect 443788 249704 443794 249756
rect 447134 249704 447140 249756
rect 447192 249744 447198 249756
rect 456794 249744 456800 249756
rect 447192 249716 456800 249744
rect 447192 249704 447198 249716
rect 456794 249704 456800 249716
rect 456852 249704 456858 249756
rect 446398 248888 446404 248940
rect 446456 248928 446462 248940
rect 447134 248928 447140 248940
rect 446456 248900 447140 248928
rect 446456 248888 446462 248900
rect 447134 248888 447140 248900
rect 447192 248888 447198 248940
rect 443730 245624 443736 245676
rect 443788 245664 443794 245676
rect 447778 245664 447784 245676
rect 443788 245636 447784 245664
rect 443788 245624 443794 245636
rect 447778 245624 447784 245636
rect 447836 245624 447842 245676
rect 572070 245556 572076 245608
rect 572128 245596 572134 245608
rect 580166 245596 580172 245608
rect 572128 245568 580172 245596
rect 572128 245556 572134 245568
rect 580166 245556 580172 245568
rect 580224 245556 580230 245608
rect 425698 244264 425704 244316
rect 425756 244304 425762 244316
rect 431310 244304 431316 244316
rect 425756 244276 431316 244304
rect 425756 244264 425762 244276
rect 431310 244264 431316 244276
rect 431368 244264 431374 244316
rect 3786 243924 3792 243976
rect 3844 243964 3850 243976
rect 4982 243964 4988 243976
rect 3844 243936 4988 243964
rect 3844 243924 3850 243936
rect 4982 243924 4988 243936
rect 5040 243924 5046 243976
rect 418522 238960 418528 239012
rect 418580 239000 418586 239012
rect 421558 239000 421564 239012
rect 418580 238972 421564 239000
rect 418580 238960 418586 238972
rect 421558 238960 421564 238972
rect 421616 238960 421622 239012
rect 361758 238688 361764 238740
rect 361816 238728 361822 238740
rect 439590 238728 439596 238740
rect 361816 238700 439596 238728
rect 361816 238688 361822 238700
rect 439590 238688 439596 238700
rect 439648 238688 439654 238740
rect 406378 236648 406384 236700
rect 406436 236688 406442 236700
rect 418522 236688 418528 236700
rect 406436 236660 418528 236688
rect 406436 236648 406442 236660
rect 418522 236648 418528 236660
rect 418580 236648 418586 236700
rect 558178 233180 558184 233232
rect 558236 233220 558242 233232
rect 580166 233220 580172 233232
rect 558236 233192 580172 233220
rect 558236 233180 558242 233192
rect 580166 233180 580172 233192
rect 580224 233180 580230 233232
rect 422938 232908 422944 232960
rect 422996 232948 423002 232960
rect 425698 232948 425704 232960
rect 422996 232920 425704 232948
rect 422996 232908 423002 232920
rect 425698 232908 425704 232920
rect 425756 232908 425762 232960
rect 361758 227672 361764 227724
rect 361816 227712 361822 227724
rect 443638 227712 443644 227724
rect 361816 227684 443644 227712
rect 361816 227672 361822 227684
rect 443638 227672 443644 227684
rect 443696 227672 443702 227724
rect 439590 224068 439596 224120
rect 439648 224108 439654 224120
rect 443730 224108 443736 224120
rect 439648 224080 443736 224108
rect 439648 224068 439654 224080
rect 443730 224068 443736 224080
rect 443788 224068 443794 224120
rect 3878 222096 3884 222148
rect 3936 222136 3942 222148
rect 5166 222136 5172 222148
rect 3936 222108 5172 222136
rect 3936 222096 3942 222108
rect 5166 222096 5172 222108
rect 5224 222096 5230 222148
rect 455138 222096 455144 222148
rect 455196 222136 455202 222148
rect 457806 222136 457812 222148
rect 455196 222108 457812 222136
rect 455196 222096 455202 222108
rect 457806 222096 457812 222108
rect 457864 222096 457870 222148
rect 439682 218016 439688 218068
rect 439740 218056 439746 218068
rect 442258 218056 442264 218068
rect 439740 218028 442264 218056
rect 439740 218016 439746 218028
rect 442258 218016 442264 218028
rect 442316 218016 442322 218068
rect 361666 216316 361672 216368
rect 361724 216356 361730 216368
rect 364058 216356 364064 216368
rect 361724 216328 364064 216356
rect 361724 216316 361730 216328
rect 364058 216316 364064 216328
rect 364116 216316 364122 216368
rect 432598 213868 432604 213920
rect 432656 213908 432662 213920
rect 438118 213908 438124 213920
rect 432656 213880 438124 213908
rect 432656 213868 432662 213880
rect 438118 213868 438124 213880
rect 438176 213868 438182 213920
rect 423030 209040 423036 209092
rect 423088 209080 423094 209092
rect 432598 209080 432604 209092
rect 423088 209052 432604 209080
rect 423088 209040 423094 209052
rect 432598 209040 432604 209052
rect 432656 209040 432662 209092
rect 457714 207884 457720 207936
rect 457772 207924 457778 207936
rect 459554 207924 459560 207936
rect 457772 207896 459560 207924
rect 457772 207884 457778 207896
rect 459554 207884 459560 207896
rect 459612 207884 459618 207936
rect 576118 206932 576124 206984
rect 576176 206972 576182 206984
rect 579798 206972 579804 206984
rect 576176 206944 579804 206972
rect 576176 206932 576182 206944
rect 579798 206932 579804 206944
rect 579856 206932 579862 206984
rect 361758 205572 361764 205624
rect 361816 205612 361822 205624
rect 436738 205612 436744 205624
rect 361816 205584 436744 205612
rect 361816 205572 361822 205584
rect 436738 205572 436744 205584
rect 436796 205572 436802 205624
rect 460566 201084 460572 201136
rect 460624 201124 460630 201136
rect 462406 201124 462412 201136
rect 460624 201096 462412 201124
rect 460624 201084 460630 201096
rect 462406 201084 462412 201096
rect 462464 201084 462470 201136
rect 460750 200676 460756 200728
rect 460808 200716 460814 200728
rect 462314 200716 462320 200728
rect 460808 200688 462320 200716
rect 460808 200676 460814 200688
rect 462314 200676 462320 200688
rect 462372 200676 462378 200728
rect 459462 200132 459468 200184
rect 459520 200172 459526 200184
rect 460934 200172 460940 200184
rect 459520 200144 460940 200172
rect 459520 200132 459526 200144
rect 460934 200132 460940 200144
rect 460992 200132 460998 200184
rect 448238 199384 448244 199436
rect 448296 199424 448302 199436
rect 461578 199424 461584 199436
rect 448296 199396 461584 199424
rect 448296 199384 448302 199396
rect 461578 199384 461584 199396
rect 461636 199384 461642 199436
rect 404078 197344 404084 197396
rect 404136 197384 404142 197396
rect 406378 197384 406384 197396
rect 404136 197356 406384 197384
rect 404136 197344 404142 197356
rect 406378 197344 406384 197356
rect 406436 197344 406442 197396
rect 438026 197344 438032 197396
rect 438084 197384 438090 197396
rect 439590 197384 439596 197396
rect 438084 197356 439596 197384
rect 438084 197344 438090 197356
rect 439590 197344 439596 197356
rect 439648 197344 439654 197396
rect 429194 195236 429200 195288
rect 429252 195276 429258 195288
rect 439682 195276 439688 195288
rect 429252 195248 439688 195276
rect 429252 195236 429258 195248
rect 439682 195236 439688 195248
rect 439740 195236 439746 195288
rect 361758 194488 361764 194540
rect 361816 194528 361822 194540
rect 431218 194528 431224 194540
rect 361816 194500 431224 194528
rect 361816 194488 361822 194500
rect 431218 194488 431224 194500
rect 431276 194488 431282 194540
rect 417418 194284 417424 194336
rect 417476 194324 417482 194336
rect 422938 194324 422944 194336
rect 417476 194296 422944 194324
rect 417476 194284 417482 194296
rect 422938 194284 422944 194296
rect 422996 194284 423002 194336
rect 547138 193128 547144 193180
rect 547196 193168 547202 193180
rect 580166 193168 580172 193180
rect 547196 193140 580172 193168
rect 547196 193128 547202 193140
rect 580166 193128 580172 193140
rect 580224 193128 580230 193180
rect 418062 192448 418068 192500
rect 418120 192488 418126 192500
rect 429194 192488 429200 192500
rect 418120 192460 429200 192488
rect 418120 192448 418126 192460
rect 429194 192448 429200 192460
rect 429252 192448 429258 192500
rect 419534 191836 419540 191888
rect 419592 191876 419598 191888
rect 423030 191876 423036 191888
rect 419592 191848 423036 191876
rect 419592 191836 419598 191848
rect 423030 191836 423036 191848
rect 423088 191836 423094 191888
rect 436370 191496 436376 191548
rect 436428 191536 436434 191548
rect 438026 191536 438032 191548
rect 436428 191508 438032 191536
rect 436428 191496 436434 191508
rect 438026 191496 438032 191508
rect 438084 191496 438090 191548
rect 394694 191088 394700 191140
rect 394752 191128 394758 191140
rect 404078 191128 404084 191140
rect 394752 191100 404084 191128
rect 394752 191088 394758 191100
rect 404078 191088 404084 191100
rect 404136 191088 404142 191140
rect 395338 189728 395344 189780
rect 395396 189768 395402 189780
rect 418062 189768 418068 189780
rect 395396 189740 418068 189768
rect 395396 189728 395402 189740
rect 418062 189728 418068 189740
rect 418120 189728 418126 189780
rect 433058 187688 433064 187740
rect 433116 187728 433122 187740
rect 436370 187728 436376 187740
rect 433116 187700 436376 187728
rect 433116 187688 433122 187700
rect 436370 187688 436376 187700
rect 436428 187688 436434 187740
rect 414658 186328 414664 186380
rect 414716 186368 414722 186380
rect 417418 186368 417424 186380
rect 414716 186340 417424 186368
rect 414716 186328 414722 186340
rect 417418 186328 417424 186340
rect 417476 186328 417482 186380
rect 391198 185376 391204 185428
rect 391256 185416 391262 185428
rect 394694 185416 394700 185428
rect 391256 185388 394700 185416
rect 391256 185376 391262 185388
rect 394694 185376 394700 185388
rect 394752 185376 394758 185428
rect 413922 183608 413928 183660
rect 413980 183648 413986 183660
rect 419534 183648 419540 183660
rect 413980 183620 419540 183648
rect 413980 183608 413986 183620
rect 419534 183608 419540 183620
rect 419592 183608 419598 183660
rect 361758 183472 361764 183524
rect 361816 183512 361822 183524
rect 447594 183512 447600 183524
rect 361816 183484 447600 183512
rect 361816 183472 361822 183484
rect 447594 183472 447600 183484
rect 447652 183512 447658 183524
rect 448146 183512 448152 183524
rect 447652 183484 448152 183512
rect 447652 183472 447658 183484
rect 448146 183472 448152 183484
rect 448204 183472 448210 183524
rect 447594 182792 447600 182844
rect 447652 182832 447658 182844
rect 528554 182832 528560 182844
rect 447652 182804 528560 182832
rect 447652 182792 447658 182804
rect 528554 182792 528560 182804
rect 528612 182792 528618 182844
rect 430574 182180 430580 182232
rect 430632 182220 430638 182232
rect 433058 182220 433064 182232
rect 430632 182192 433064 182220
rect 430632 182180 430638 182192
rect 433058 182180 433064 182192
rect 433116 182180 433122 182232
rect 400582 181432 400588 181484
rect 400640 181472 400646 181484
rect 413922 181472 413928 181484
rect 400640 181444 413928 181472
rect 400640 181432 400646 181444
rect 413922 181432 413928 181444
rect 413980 181432 413986 181484
rect 551278 179324 551284 179376
rect 551336 179364 551342 179376
rect 580166 179364 580172 179376
rect 551336 179336 580172 179364
rect 551336 179324 551342 179336
rect 580166 179324 580172 179336
rect 580224 179324 580230 179376
rect 398098 176672 398104 176724
rect 398156 176712 398162 176724
rect 400582 176712 400588 176724
rect 398156 176684 400588 176712
rect 398156 176672 398162 176684
rect 400582 176672 400588 176684
rect 400640 176672 400646 176724
rect 430574 176712 430580 176724
rect 426452 176684 430580 176712
rect 422938 176604 422944 176656
rect 422996 176644 423002 176656
rect 426452 176644 426480 176684
rect 430574 176672 430580 176684
rect 430632 176672 430638 176724
rect 422996 176616 426480 176644
rect 422996 176604 423002 176616
rect 361758 172456 361764 172508
rect 361816 172496 361822 172508
rect 447134 172496 447140 172508
rect 361816 172468 447140 172496
rect 361816 172456 361822 172468
rect 447134 172456 447140 172468
rect 447192 172456 447198 172508
rect 447134 171776 447140 171828
rect 447192 171816 447198 171828
rect 448330 171816 448336 171828
rect 447192 171788 448336 171816
rect 447192 171776 447198 171788
rect 448330 171776 448336 171788
rect 448388 171816 448394 171828
rect 524414 171816 524420 171828
rect 448388 171788 524420 171816
rect 448388 171776 448394 171788
rect 524414 171776 524420 171788
rect 524472 171776 524478 171828
rect 391290 171096 391296 171148
rect 391348 171136 391354 171148
rect 395338 171136 395344 171148
rect 391348 171108 395344 171136
rect 391348 171096 391354 171108
rect 395338 171096 395344 171108
rect 395396 171096 395402 171148
rect 420178 169736 420184 169788
rect 420236 169776 420242 169788
rect 422938 169776 422944 169788
rect 420236 169748 422944 169776
rect 420236 169736 420242 169748
rect 422938 169736 422944 169748
rect 422996 169736 423002 169788
rect 533430 166948 533436 167000
rect 533488 166988 533494 167000
rect 580166 166988 580172 167000
rect 533488 166960 580172 166988
rect 533488 166948 533494 166960
rect 580166 166948 580172 166960
rect 580224 166948 580230 167000
rect 388530 166268 388536 166320
rect 388588 166308 388594 166320
rect 391198 166308 391204 166320
rect 388588 166280 391204 166308
rect 388588 166268 388594 166280
rect 391198 166268 391204 166280
rect 391256 166268 391262 166320
rect 388438 164840 388444 164892
rect 388496 164880 388502 164892
rect 398098 164880 398104 164892
rect 388496 164852 398104 164880
rect 388496 164840 388502 164852
rect 398098 164840 398104 164852
rect 398156 164840 398162 164892
rect 448422 164160 448428 164212
rect 448480 164200 448486 164212
rect 449342 164200 449348 164212
rect 448480 164172 449348 164200
rect 448480 164160 448486 164172
rect 449342 164160 449348 164172
rect 449400 164160 449406 164212
rect 438578 163616 438584 163668
rect 438636 163656 438642 163668
rect 439498 163656 439504 163668
rect 438636 163628 439504 163656
rect 438636 163616 438642 163628
rect 439498 163616 439504 163628
rect 439556 163616 439562 163668
rect 445202 163616 445208 163668
rect 445260 163656 445266 163668
rect 446398 163656 446404 163668
rect 445260 163628 446404 163656
rect 445260 163616 445266 163628
rect 446398 163616 446404 163628
rect 446456 163616 446462 163668
rect 407022 162868 407028 162920
rect 407080 162908 407086 162920
rect 414658 162908 414664 162920
rect 407080 162880 414664 162908
rect 407080 162868 407086 162880
rect 414658 162868 414664 162880
rect 414716 162868 414722 162920
rect 456794 162256 456800 162308
rect 456852 162296 456858 162308
rect 457806 162296 457812 162308
rect 456852 162268 457812 162296
rect 456852 162256 456858 162268
rect 457806 162256 457812 162268
rect 457864 162296 457870 162308
rect 485774 162296 485780 162308
rect 457864 162268 485780 162296
rect 457864 162256 457870 162268
rect 485774 162256 485780 162268
rect 485832 162256 485838 162308
rect 418706 162188 418712 162240
rect 418764 162228 418770 162240
rect 457990 162228 457996 162240
rect 418764 162200 457996 162228
rect 418764 162188 418770 162200
rect 457990 162188 457996 162200
rect 458048 162228 458054 162240
rect 458048 162200 460934 162228
rect 458048 162188 458054 162200
rect 415118 162120 415124 162172
rect 415176 162160 415182 162172
rect 456794 162160 456800 162172
rect 415176 162132 456800 162160
rect 415176 162120 415182 162132
rect 456794 162120 456800 162132
rect 456852 162120 456858 162172
rect 460906 162160 460934 162200
rect 489914 162160 489920 162172
rect 460906 162132 489920 162160
rect 489914 162120 489920 162132
rect 489972 162120 489978 162172
rect 375190 161508 375196 161560
rect 375248 161548 375254 161560
rect 418706 161548 418712 161560
rect 375248 161520 418712 161548
rect 375248 161508 375254 161520
rect 418706 161508 418712 161520
rect 418764 161508 418770 161560
rect 445202 161508 445208 161560
rect 445260 161548 445266 161560
rect 450998 161548 451004 161560
rect 445260 161520 451004 161548
rect 445260 161508 445266 161520
rect 450998 161508 451004 161520
rect 451056 161508 451062 161560
rect 412082 161440 412088 161492
rect 412140 161480 412146 161492
rect 459554 161480 459560 161492
rect 412140 161452 459560 161480
rect 412140 161440 412146 161452
rect 459554 161440 459560 161452
rect 459612 161480 459618 161492
rect 460198 161480 460204 161492
rect 459612 161452 460204 161480
rect 459612 161440 459618 161452
rect 460198 161440 460204 161452
rect 460256 161440 460262 161492
rect 361758 161372 361764 161424
rect 361816 161412 361822 161424
rect 448330 161412 448336 161424
rect 361816 161384 448336 161412
rect 361816 161372 361822 161384
rect 448330 161372 448336 161384
rect 448388 161372 448394 161424
rect 359458 160692 359464 160744
rect 359516 160732 359522 160744
rect 388530 160732 388536 160744
rect 359516 160704 388536 160732
rect 359516 160692 359522 160704
rect 388530 160692 388536 160704
rect 388588 160692 388594 160744
rect 448330 160692 448336 160744
rect 448388 160732 448394 160744
rect 521654 160732 521660 160744
rect 448388 160704 521660 160732
rect 448388 160692 448394 160704
rect 521654 160692 521660 160704
rect 521712 160692 521718 160744
rect 425330 160488 425336 160540
rect 425388 160528 425394 160540
rect 425882 160528 425888 160540
rect 425388 160500 425888 160528
rect 425388 160488 425394 160500
rect 425882 160488 425888 160500
rect 425940 160528 425946 160540
rect 496814 160528 496820 160540
rect 425940 160500 496820 160528
rect 425940 160488 425946 160500
rect 496814 160488 496820 160500
rect 496872 160488 496878 160540
rect 428642 160420 428648 160472
rect 428700 160460 428706 160472
rect 500954 160460 500960 160472
rect 428700 160432 500960 160460
rect 428700 160420 428706 160432
rect 500954 160420 500960 160432
rect 501012 160420 501018 160472
rect 421834 160352 421840 160404
rect 421892 160392 421898 160404
rect 494054 160392 494060 160404
rect 421892 160364 494060 160392
rect 421892 160352 421898 160364
rect 494054 160352 494060 160364
rect 494112 160352 494118 160404
rect 435266 160284 435272 160336
rect 435324 160324 435330 160336
rect 436002 160324 436008 160336
rect 435324 160296 436008 160324
rect 435324 160284 435330 160296
rect 436002 160284 436008 160296
rect 436060 160324 436066 160336
rect 509234 160324 509240 160336
rect 436060 160296 509240 160324
rect 436060 160284 436066 160296
rect 509234 160284 509240 160296
rect 509292 160284 509298 160336
rect 431770 160216 431776 160268
rect 431828 160256 431834 160268
rect 505094 160256 505100 160268
rect 431828 160228 505100 160256
rect 431828 160216 431834 160228
rect 505094 160216 505100 160228
rect 505152 160216 505158 160268
rect 386138 160148 386144 160200
rect 386196 160188 386202 160200
rect 415118 160188 415124 160200
rect 386196 160160 415124 160188
rect 386196 160148 386202 160160
rect 415118 160148 415124 160160
rect 415176 160148 415182 160200
rect 438578 160148 438584 160200
rect 438636 160188 438642 160200
rect 513374 160188 513380 160200
rect 438636 160160 513380 160188
rect 438636 160148 438642 160160
rect 513374 160148 513380 160160
rect 513432 160148 513438 160200
rect 387794 160080 387800 160132
rect 387852 160120 387858 160132
rect 391290 160120 391296 160132
rect 387852 160092 391296 160120
rect 387852 160080 387858 160092
rect 391290 160080 391296 160092
rect 391348 160080 391354 160132
rect 409506 160080 409512 160132
rect 409564 160120 409570 160132
rect 441568 160120 441574 160132
rect 409564 160092 441574 160120
rect 409564 160080 409570 160092
rect 441568 160080 441574 160092
rect 441626 160120 441632 160132
rect 442902 160120 442908 160132
rect 441626 160092 442908 160120
rect 441626 160080 441632 160092
rect 442902 160080 442908 160092
rect 442960 160120 442966 160132
rect 517514 160120 517520 160132
rect 442960 160092 517520 160120
rect 442960 160080 442966 160092
rect 517514 160080 517520 160092
rect 517572 160080 517578 160132
rect 409874 159740 409880 159792
rect 409932 159780 409938 159792
rect 420178 159780 420184 159792
rect 409932 159752 420184 159780
rect 409932 159740 409938 159752
rect 420178 159740 420184 159752
rect 420236 159740 420242 159792
rect 409138 159672 409144 159724
rect 409196 159712 409202 159724
rect 427998 159712 428004 159724
rect 409196 159684 428004 159712
rect 409196 159672 409202 159684
rect 427998 159672 428004 159684
rect 428056 159672 428062 159724
rect 409230 159604 409236 159656
rect 409288 159644 409294 159656
rect 431310 159644 431316 159656
rect 409288 159616 431316 159644
rect 409288 159604 409294 159616
rect 431310 159604 431316 159616
rect 431368 159604 431374 159656
rect 409322 159536 409328 159588
rect 409380 159576 409386 159588
rect 434806 159576 434812 159588
rect 409380 159548 434812 159576
rect 409380 159536 409386 159548
rect 434806 159536 434812 159548
rect 434864 159536 434870 159588
rect 409414 159468 409420 159520
rect 409472 159508 409478 159520
rect 437934 159508 437940 159520
rect 409472 159480 437940 159508
rect 409472 159468 409478 159480
rect 437934 159468 437940 159480
rect 437992 159468 437998 159520
rect 384206 159400 384212 159452
rect 384264 159440 384270 159452
rect 421374 159440 421380 159452
rect 384264 159412 421380 159440
rect 384264 159400 384270 159412
rect 421374 159400 421380 159412
rect 421432 159400 421438 159452
rect 386230 159332 386236 159384
rect 386288 159372 386294 159384
rect 425146 159372 425152 159384
rect 386288 159344 425152 159372
rect 386288 159332 386294 159344
rect 425146 159332 425152 159344
rect 425204 159332 425210 159384
rect 451734 158652 451740 158704
rect 451792 158692 451798 158704
rect 454954 158692 454960 158704
rect 451792 158664 454960 158692
rect 451792 158652 451798 158664
rect 454954 158652 454960 158664
rect 455012 158652 455018 158704
rect 361574 157972 361580 158024
rect 361632 158012 361638 158024
rect 387794 158012 387800 158024
rect 361632 157984 387800 158012
rect 361632 157972 361638 157984
rect 387794 157972 387800 157984
rect 387852 157972 387858 158024
rect 398834 157972 398840 158024
rect 398892 158012 398898 158024
rect 409874 158012 409880 158024
rect 398892 157984 409880 158012
rect 398892 157972 398898 157984
rect 409874 157972 409880 157984
rect 409932 157972 409938 158024
rect 451734 157292 451740 157344
rect 451792 157332 451798 157344
rect 455046 157332 455052 157344
rect 451792 157304 455052 157332
rect 451792 157292 451798 157304
rect 455046 157292 455052 157304
rect 455104 157292 455110 157344
rect 402238 155184 402244 155236
rect 402296 155224 402302 155236
rect 407022 155224 407028 155236
rect 402296 155196 407028 155224
rect 402296 155184 402302 155196
rect 407022 155184 407028 155196
rect 407080 155184 407086 155236
rect 452470 154436 452476 154488
rect 452528 154476 452534 154488
rect 453574 154476 453580 154488
rect 452528 154448 453580 154476
rect 452528 154436 452534 154448
rect 453574 154436 453580 154448
rect 453632 154436 453638 154488
rect 389266 153824 389272 153876
rect 389324 153864 389330 153876
rect 398742 153864 398748 153876
rect 389324 153836 398748 153864
rect 389324 153824 389330 153836
rect 398742 153824 398748 153836
rect 398800 153824 398806 153876
rect 537478 153144 537484 153196
rect 537536 153184 537542 153196
rect 580166 153184 580172 153196
rect 537536 153156 580172 153184
rect 537536 153144 537542 153156
rect 580166 153144 580172 153156
rect 580224 153144 580230 153196
rect 452470 152940 452476 152992
rect 452528 152980 452534 152992
rect 453666 152980 453672 152992
rect 452528 152952 453672 152980
rect 452528 152940 452534 152952
rect 453666 152940 453672 152952
rect 453724 152940 453730 152992
rect 452562 151444 452568 151496
rect 452620 151484 452626 151496
rect 457622 151484 457628 151496
rect 452620 151456 457628 151484
rect 452620 151444 452626 151456
rect 457622 151444 457628 151456
rect 457680 151444 457686 151496
rect 386506 150560 386512 150612
rect 386564 150600 386570 150612
rect 389266 150600 389272 150612
rect 386564 150572 389272 150600
rect 386564 150560 386570 150572
rect 389266 150560 389272 150572
rect 389324 150560 389330 150612
rect 361758 150356 361764 150408
rect 361816 150396 361822 150408
rect 409506 150396 409512 150408
rect 361816 150368 409512 150396
rect 361816 150356 361822 150368
rect 409506 150356 409512 150368
rect 409564 150356 409570 150408
rect 371234 149744 371240 149796
rect 371292 149784 371298 149796
rect 386506 149784 386512 149796
rect 371292 149756 386512 149784
rect 371292 149744 371298 149756
rect 386506 149744 386512 149756
rect 386564 149744 386570 149796
rect 368290 149676 368296 149728
rect 368348 149716 368354 149728
rect 388438 149716 388444 149728
rect 368348 149688 388444 149716
rect 368348 149676 368354 149688
rect 388438 149676 388444 149688
rect 388496 149676 388502 149728
rect 365714 147636 365720 147688
rect 365772 147676 365778 147688
rect 371234 147676 371240 147688
rect 365772 147648 371240 147676
rect 365772 147636 365778 147648
rect 371234 147636 371240 147648
rect 371292 147636 371298 147688
rect 452562 147364 452568 147416
rect 452620 147404 452626 147416
rect 459094 147404 459100 147416
rect 452620 147376 459100 147404
rect 452620 147364 452626 147376
rect 459094 147364 459100 147376
rect 459152 147364 459158 147416
rect 393958 146956 393964 147008
rect 394016 146996 394022 147008
rect 402238 146996 402244 147008
rect 394016 146968 402244 146996
rect 394016 146956 394022 146968
rect 402238 146956 402244 146968
rect 402296 146956 402302 147008
rect 451826 146208 451832 146260
rect 451884 146248 451890 146260
rect 459278 146248 459284 146260
rect 451884 146220 459284 146248
rect 451884 146208 451890 146220
rect 459278 146208 459284 146220
rect 459336 146208 459342 146260
rect 364334 144848 364340 144900
rect 364392 144888 364398 144900
rect 368290 144888 368296 144900
rect 364392 144860 368296 144888
rect 364392 144848 364398 144860
rect 368290 144848 368296 144860
rect 368348 144848 368354 144900
rect 451550 144780 451556 144832
rect 451608 144820 451614 144832
rect 456426 144820 456432 144832
rect 451608 144792 456432 144820
rect 451608 144780 451614 144792
rect 456426 144780 456432 144792
rect 456484 144780 456490 144832
rect 362954 143556 362960 143608
rect 363012 143596 363018 143608
rect 365622 143596 365628 143608
rect 363012 143568 365628 143596
rect 363012 143556 363018 143568
rect 365622 143556 365628 143568
rect 365680 143556 365686 143608
rect 460198 143488 460204 143540
rect 460256 143528 460262 143540
rect 460842 143528 460848 143540
rect 460256 143500 460848 143528
rect 460256 143488 460262 143500
rect 460842 143488 460848 143500
rect 460900 143488 460906 143540
rect 452562 143420 452568 143472
rect 452620 143460 452626 143472
rect 457438 143460 457444 143472
rect 452620 143432 457444 143460
rect 452620 143420 452626 143432
rect 457438 143420 457444 143432
rect 457496 143420 457502 143472
rect 460842 142196 460848 142248
rect 460900 142236 460906 142248
rect 481910 142236 481916 142248
rect 460900 142208 481916 142236
rect 460900 142196 460906 142208
rect 481910 142196 481916 142208
rect 481968 142196 481974 142248
rect 450998 142128 451004 142180
rect 451056 142168 451062 142180
rect 533982 142168 533988 142180
rect 451056 142140 533988 142168
rect 451056 142128 451062 142140
rect 533982 142128 533988 142140
rect 534040 142168 534046 142180
rect 540422 142168 540428 142180
rect 534040 142140 540428 142168
rect 534040 142128 534046 142140
rect 540422 142128 540428 142140
rect 540480 142128 540486 142180
rect 452562 141924 452568 141976
rect 452620 141964 452626 141976
rect 459002 141964 459008 141976
rect 452620 141936 459008 141964
rect 452620 141924 452626 141936
rect 459002 141924 459008 141936
rect 459060 141924 459066 141976
rect 452562 140700 452568 140752
rect 452620 140740 452626 140752
rect 454862 140740 454868 140752
rect 452620 140712 454868 140740
rect 452620 140700 452626 140712
rect 454862 140700 454868 140712
rect 454920 140700 454926 140752
rect 359642 140020 359648 140072
rect 359700 140060 359706 140072
rect 393958 140060 393964 140072
rect 359700 140032 393964 140060
rect 359700 140020 359706 140032
rect 393958 140020 393964 140032
rect 394016 140020 394022 140072
rect 533338 140020 533344 140072
rect 533396 140060 533402 140072
rect 542538 140060 542544 140072
rect 533396 140032 542544 140060
rect 533396 140020 533402 140032
rect 542538 140020 542544 140032
rect 542596 140020 542602 140072
rect 359550 139544 359556 139596
rect 359608 139584 359614 139596
rect 364334 139584 364340 139596
rect 359608 139556 364340 139584
rect 359608 139544 359614 139556
rect 364334 139544 364340 139556
rect 364392 139544 364398 139596
rect 361758 139340 361764 139392
rect 361816 139380 361822 139392
rect 409414 139380 409420 139392
rect 361816 139352 409420 139380
rect 361816 139340 361822 139352
rect 409414 139340 409420 139352
rect 409472 139340 409478 139392
rect 555418 139340 555424 139392
rect 555476 139380 555482 139392
rect 580166 139380 580172 139392
rect 555476 139352 580172 139380
rect 555476 139340 555482 139352
rect 580166 139340 580172 139352
rect 580224 139340 580230 139392
rect 451550 139204 451556 139256
rect 451608 139244 451614 139256
rect 456334 139244 456340 139256
rect 451608 139216 456340 139244
rect 451608 139204 451614 139216
rect 456334 139204 456340 139216
rect 456392 139204 456398 139256
rect 452562 137844 452568 137896
rect 452620 137884 452626 137896
rect 457530 137884 457536 137896
rect 452620 137856 457536 137884
rect 452620 137844 452626 137856
rect 457530 137844 457536 137856
rect 457588 137844 457594 137896
rect 538950 136552 538956 136604
rect 539008 136592 539014 136604
rect 539502 136592 539508 136604
rect 539008 136564 539508 136592
rect 539008 136552 539014 136564
rect 539502 136552 539508 136564
rect 539560 136552 539566 136604
rect 451550 136484 451556 136536
rect 451608 136524 451614 136536
rect 456242 136524 456248 136536
rect 451608 136496 456248 136524
rect 451608 136484 451614 136496
rect 456242 136484 456248 136496
rect 456300 136484 456306 136536
rect 452010 135124 452016 135176
rect 452068 135164 452074 135176
rect 458910 135164 458916 135176
rect 452068 135136 458916 135164
rect 452068 135124 452074 135136
rect 458910 135124 458916 135136
rect 458968 135124 458974 135176
rect 452286 132404 452292 132456
rect 452344 132444 452350 132456
rect 453390 132444 453396 132456
rect 452344 132416 453396 132444
rect 452344 132404 452350 132416
rect 453390 132404 453396 132416
rect 453448 132404 453454 132456
rect 361390 131112 361396 131164
rect 361448 131152 361454 131164
rect 362586 131152 362592 131164
rect 361448 131124 362592 131152
rect 361448 131112 361454 131124
rect 362586 131112 362592 131124
rect 362644 131112 362650 131164
rect 452562 131044 452568 131096
rect 452620 131084 452626 131096
rect 456150 131084 456156 131096
rect 452620 131056 456156 131084
rect 452620 131044 452626 131056
rect 456150 131044 456156 131056
rect 456208 131044 456214 131096
rect 452102 129684 452108 129736
rect 452160 129724 452166 129736
rect 453298 129724 453304 129736
rect 452160 129696 453304 129724
rect 452160 129684 452166 129696
rect 453298 129684 453304 129696
rect 453356 129684 453362 129736
rect 361758 128256 361764 128308
rect 361816 128296 361822 128308
rect 409322 128296 409328 128308
rect 361816 128268 409328 128296
rect 361816 128256 361822 128268
rect 409322 128256 409328 128268
rect 409380 128256 409386 128308
rect 452562 126896 452568 126948
rect 452620 126936 452626 126948
rect 458818 126936 458824 126948
rect 452620 126908 458824 126936
rect 452620 126896 452626 126908
rect 458818 126896 458824 126908
rect 458876 126896 458882 126948
rect 574738 126896 574744 126948
rect 574796 126936 574802 126948
rect 580166 126936 580172 126948
rect 574796 126908 580172 126936
rect 574796 126896 574802 126908
rect 580166 126896 580172 126908
rect 580224 126896 580230 126948
rect 451734 126760 451740 126812
rect 451792 126800 451798 126812
rect 453482 126800 453488 126812
rect 451792 126772 453488 126800
rect 451792 126760 451798 126772
rect 453482 126760 453488 126772
rect 453540 126760 453546 126812
rect 451734 123088 451740 123140
rect 451792 123128 451798 123140
rect 454770 123128 454776 123140
rect 451792 123100 454776 123128
rect 451792 123088 451798 123100
rect 454770 123088 454776 123100
rect 454828 123088 454834 123140
rect 451918 122000 451924 122052
rect 451976 122040 451982 122052
rect 459186 122040 459192 122052
rect 451976 122012 459192 122040
rect 451976 122000 451982 122012
rect 459186 122000 459192 122012
rect 459244 122000 459250 122052
rect 384942 119348 384948 119400
rect 385000 119388 385006 119400
rect 456058 119388 456064 119400
rect 385000 119360 456064 119388
rect 385000 119348 385006 119360
rect 456058 119348 456064 119360
rect 456116 119348 456122 119400
rect 361758 117240 361764 117292
rect 361816 117280 361822 117292
rect 409230 117280 409236 117292
rect 361816 117252 409236 117280
rect 361816 117240 361822 117252
rect 409230 117240 409236 117252
rect 409288 117240 409294 117292
rect 569218 113092 569224 113144
rect 569276 113132 569282 113144
rect 579798 113132 579804 113144
rect 569276 113104 579804 113132
rect 569276 113092 569282 113104
rect 579798 113092 579804 113104
rect 579856 113092 579862 113144
rect 402146 107584 402152 107636
rect 402204 107624 402210 107636
rect 403618 107624 403624 107636
rect 402204 107596 403624 107624
rect 402204 107584 402210 107596
rect 403618 107584 403624 107596
rect 403676 107584 403682 107636
rect 439130 107244 439136 107296
rect 439188 107284 439194 107296
rect 450814 107284 450820 107296
rect 439188 107256 450820 107284
rect 439188 107244 439194 107256
rect 450814 107244 450820 107256
rect 450872 107244 450878 107296
rect 432966 107176 432972 107228
rect 433024 107216 433030 107228
rect 450538 107216 450544 107228
rect 433024 107188 450544 107216
rect 433024 107176 433030 107188
rect 450538 107176 450544 107188
rect 450596 107176 450602 107228
rect 426802 107108 426808 107160
rect 426860 107148 426866 107160
rect 450722 107148 450728 107160
rect 426860 107120 450728 107148
rect 426860 107108 426866 107120
rect 450722 107108 450728 107120
rect 450780 107108 450786 107160
rect 420638 107040 420644 107092
rect 420696 107080 420702 107092
rect 450630 107080 450636 107092
rect 420696 107052 450636 107080
rect 420696 107040 420702 107052
rect 450630 107040 450636 107052
rect 450688 107040 450694 107092
rect 414474 106972 414480 107024
rect 414532 107012 414538 107024
rect 454678 107012 454684 107024
rect 414532 106984 454684 107012
rect 414532 106972 414538 106984
rect 454678 106972 454684 106984
rect 454736 106972 454742 107024
rect 389818 106904 389824 106956
rect 389876 106944 389882 106956
rect 450998 106944 451004 106956
rect 389876 106916 451004 106944
rect 389876 106904 389882 106916
rect 450998 106904 451004 106916
rect 451056 106904 451062 106956
rect 445294 106496 445300 106548
rect 445352 106536 445358 106548
rect 450906 106536 450912 106548
rect 445352 106508 450912 106536
rect 445352 106496 445358 106508
rect 450906 106496 450912 106508
rect 450964 106496 450970 106548
rect 361758 106224 361764 106276
rect 361816 106264 361822 106276
rect 409138 106264 409144 106276
rect 361816 106236 409144 106264
rect 361816 106224 361822 106236
rect 409138 106224 409144 106236
rect 409196 106224 409202 106276
rect 559558 100648 559564 100700
rect 559616 100688 559622 100700
rect 580166 100688 580172 100700
rect 559616 100660 580172 100688
rect 559616 100648 559622 100660
rect 580166 100648 580172 100660
rect 580224 100648 580230 100700
rect 3602 98608 3608 98660
rect 3660 98648 3666 98660
rect 20898 98648 20904 98660
rect 3660 98620 20904 98648
rect 3660 98608 3666 98620
rect 20898 98608 20904 98620
rect 20956 98608 20962 98660
rect 361758 95140 361764 95192
rect 361816 95180 361822 95192
rect 386230 95180 386236 95192
rect 361816 95152 386236 95180
rect 361816 95140 361822 95152
rect 386230 95140 386236 95152
rect 386288 95140 386294 95192
rect 570598 86912 570604 86964
rect 570656 86952 570662 86964
rect 580166 86952 580172 86964
rect 570656 86924 580172 86952
rect 570656 86912 570662 86924
rect 580166 86912 580172 86924
rect 580224 86912 580230 86964
rect 3694 86232 3700 86284
rect 3752 86272 3758 86284
rect 20898 86272 20904 86284
rect 3752 86244 20904 86272
rect 3752 86232 3758 86244
rect 20898 86232 20904 86244
rect 20956 86232 20962 86284
rect 361758 84124 361764 84176
rect 361816 84164 361822 84176
rect 384206 84164 384212 84176
rect 361816 84136 384212 84164
rect 361816 84124 361822 84136
rect 384206 84124 384212 84136
rect 384264 84124 384270 84176
rect 361758 73108 361764 73160
rect 361816 73148 361822 73160
rect 375190 73148 375196 73160
rect 361816 73120 375196 73148
rect 361816 73108 361822 73120
rect 375190 73108 375196 73120
rect 375248 73108 375254 73160
rect 544378 73108 544384 73160
rect 544436 73148 544442 73160
rect 580166 73148 580172 73160
rect 544436 73120 580172 73148
rect 544436 73108 544442 73120
rect 580166 73108 580172 73120
rect 580224 73108 580230 73160
rect 5074 71680 5080 71732
rect 5132 71720 5138 71732
rect 5534 71720 5540 71732
rect 5132 71692 5540 71720
rect 5132 71680 5138 71692
rect 5534 71680 5540 71692
rect 5592 71680 5598 71732
rect 3602 70388 3608 70440
rect 3660 70428 3666 70440
rect 19978 70428 19984 70440
rect 3660 70400 19984 70428
rect 3660 70388 3666 70400
rect 19978 70388 19984 70400
rect 20036 70388 20042 70440
rect 5534 70320 5540 70372
rect 5592 70360 5598 70372
rect 7558 70360 7564 70372
rect 5592 70332 7564 70360
rect 5592 70320 5598 70332
rect 7558 70320 7564 70332
rect 7616 70320 7622 70372
rect 361758 62024 361764 62076
rect 361816 62064 361822 62076
rect 386138 62064 386144 62076
rect 361816 62036 386144 62064
rect 361816 62024 361822 62036
rect 386138 62024 386144 62036
rect 386196 62024 386202 62076
rect 7558 60732 7564 60784
rect 7616 60772 7622 60784
rect 7616 60744 8340 60772
rect 7616 60732 7622 60744
rect 8312 60704 8340 60744
rect 10042 60704 10048 60716
rect 8312 60676 10048 60704
rect 10042 60664 10048 60676
rect 10100 60664 10106 60716
rect 548518 60664 548524 60716
rect 548576 60704 548582 60716
rect 580166 60704 580172 60716
rect 548576 60676 580172 60704
rect 548576 60664 548582 60676
rect 580166 60664 580172 60676
rect 580224 60664 580230 60716
rect 4798 59304 4804 59356
rect 4856 59344 4862 59356
rect 5810 59344 5816 59356
rect 4856 59316 5816 59344
rect 4856 59304 4862 59316
rect 5810 59304 5816 59316
rect 5868 59304 5874 59356
rect 3602 57944 3608 57996
rect 3660 57984 3666 57996
rect 20070 57984 20076 57996
rect 3660 57956 20076 57984
rect 3660 57944 3666 57956
rect 20070 57944 20076 57956
rect 20128 57944 20134 57996
rect 5810 57196 5816 57248
rect 5868 57236 5874 57248
rect 9766 57236 9772 57248
rect 5868 57208 9772 57236
rect 5868 57196 5874 57208
rect 9766 57196 9772 57208
rect 9824 57196 9830 57248
rect 4890 56516 4896 56568
rect 4948 56556 4954 56568
rect 7282 56556 7288 56568
rect 4948 56528 7288 56556
rect 4948 56516 4954 56528
rect 7282 56516 7288 56528
rect 7340 56516 7346 56568
rect 10042 56516 10048 56568
rect 10100 56556 10106 56568
rect 12342 56556 12348 56568
rect 10100 56528 12348 56556
rect 10100 56516 10106 56528
rect 12342 56516 12348 56528
rect 12400 56516 12406 56568
rect 9766 56108 9772 56160
rect 9824 56148 9830 56160
rect 12802 56148 12808 56160
rect 9824 56120 12808 56148
rect 9824 56108 9830 56120
rect 12802 56108 12808 56120
rect 12860 56108 12866 56160
rect 5534 54476 5540 54528
rect 5592 54516 5598 54528
rect 12250 54516 12256 54528
rect 5592 54488 12256 54516
rect 5592 54476 5598 54488
rect 12250 54476 12256 54488
rect 12308 54476 12314 54528
rect 7282 54068 7288 54120
rect 7340 54108 7346 54120
rect 11974 54108 11980 54120
rect 7340 54080 11980 54108
rect 7340 54068 7346 54080
rect 11974 54068 11980 54080
rect 12032 54068 12038 54120
rect 12342 53388 12348 53440
rect 12400 53428 12406 53440
rect 15194 53428 15200 53440
rect 12400 53400 15200 53428
rect 12400 53388 12406 53400
rect 15194 53388 15200 53400
rect 15252 53388 15258 53440
rect 11974 52436 11980 52488
rect 12032 52476 12038 52488
rect 12032 52448 13860 52476
rect 12032 52436 12038 52448
rect 13832 52408 13860 52448
rect 19242 52408 19248 52420
rect 13832 52380 19248 52408
rect 19242 52368 19248 52380
rect 19300 52368 19306 52420
rect 361758 51076 361764 51128
rect 361816 51116 361822 51128
rect 386138 51116 386144 51128
rect 361816 51088 386144 51116
rect 361816 51076 361822 51088
rect 386138 51076 386144 51088
rect 386196 51076 386202 51128
rect 540606 51076 540612 51128
rect 540664 51116 540670 51128
rect 543734 51116 543740 51128
rect 540664 51088 543740 51116
rect 540664 51076 540670 51088
rect 543734 51076 543740 51088
rect 543792 51076 543798 51128
rect 4982 50328 4988 50380
rect 5040 50368 5046 50380
rect 11698 50368 11704 50380
rect 5040 50340 11704 50368
rect 5040 50328 5046 50340
rect 11698 50328 11704 50340
rect 11756 50328 11762 50380
rect 12802 50328 12808 50380
rect 12860 50368 12866 50380
rect 20622 50368 20628 50380
rect 12860 50340 20628 50368
rect 12860 50328 12866 50340
rect 20622 50328 20628 50340
rect 20680 50328 20686 50380
rect 15194 49716 15200 49768
rect 15252 49756 15258 49768
rect 15252 49728 16574 49756
rect 15252 49716 15258 49728
rect 16546 49688 16574 49728
rect 18966 49688 18972 49700
rect 16546 49660 18972 49688
rect 18966 49648 18972 49660
rect 19024 49648 19030 49700
rect 18966 47812 18972 47864
rect 19024 47852 19030 47864
rect 20898 47852 20904 47864
rect 19024 47824 20904 47852
rect 19024 47812 19030 47824
rect 20898 47812 20904 47824
rect 20956 47812 20962 47864
rect 3050 46996 3056 47048
rect 3108 47036 3114 47048
rect 384758 47036 384764 47048
rect 3108 47008 384764 47036
rect 3108 46996 3114 47008
rect 384758 46996 384764 47008
rect 384816 46996 384822 47048
rect 3694 46860 3700 46912
rect 3752 46900 3758 46912
rect 384574 46900 384580 46912
rect 3752 46872 384580 46900
rect 3752 46860 3758 46872
rect 384574 46860 384580 46872
rect 384632 46860 384638 46912
rect 573358 46860 573364 46912
rect 573416 46900 573422 46912
rect 580166 46900 580172 46912
rect 573416 46872 580172 46900
rect 573416 46860 573422 46872
rect 580166 46860 580172 46872
rect 580224 46860 580230 46912
rect 3234 46792 3240 46844
rect 3292 46832 3298 46844
rect 381906 46832 381912 46844
rect 3292 46804 381912 46832
rect 3292 46792 3298 46804
rect 381906 46792 381912 46804
rect 381964 46792 381970 46844
rect 3326 46724 3332 46776
rect 3384 46764 3390 46776
rect 381998 46764 382004 46776
rect 3384 46736 382004 46764
rect 3384 46724 3390 46736
rect 381998 46724 382004 46736
rect 382056 46724 382062 46776
rect 3970 46656 3976 46708
rect 4028 46696 4034 46708
rect 378962 46696 378968 46708
rect 4028 46668 378968 46696
rect 4028 46656 4034 46668
rect 378962 46656 378968 46668
rect 379020 46656 379026 46708
rect 3878 46588 3884 46640
rect 3936 46628 3942 46640
rect 378870 46628 378876 46640
rect 3936 46600 378876 46628
rect 3936 46588 3942 46600
rect 378870 46588 378876 46600
rect 378928 46588 378934 46640
rect 3786 46520 3792 46572
rect 3844 46560 3850 46572
rect 378594 46560 378600 46572
rect 3844 46532 378600 46560
rect 3844 46520 3850 46532
rect 378594 46520 378600 46532
rect 378652 46520 378658 46572
rect 3418 46452 3424 46504
rect 3476 46492 3482 46504
rect 375926 46492 375932 46504
rect 3476 46464 375932 46492
rect 3476 46452 3482 46464
rect 375926 46452 375932 46464
rect 375984 46452 375990 46504
rect 19978 46384 19984 46436
rect 20036 46424 20042 46436
rect 384390 46424 384396 46436
rect 20036 46396 384396 46424
rect 20036 46384 20042 46396
rect 384390 46384 384396 46396
rect 384448 46384 384454 46436
rect 20070 46316 20076 46368
rect 20128 46356 20134 46368
rect 382090 46356 382096 46368
rect 20128 46328 382096 46356
rect 20128 46316 20134 46328
rect 382090 46316 382096 46328
rect 382148 46316 382154 46368
rect 21450 46248 21456 46300
rect 21508 46288 21514 46300
rect 376662 46288 376668 46300
rect 21508 46260 376668 46288
rect 21508 46248 21514 46260
rect 376662 46248 376668 46260
rect 376720 46248 376726 46300
rect 21358 46180 21364 46232
rect 21416 46220 21422 46232
rect 373626 46220 373632 46232
rect 21416 46192 373632 46220
rect 21416 46180 21422 46192
rect 373626 46180 373632 46192
rect 373684 46180 373690 46232
rect 12434 46112 12440 46164
rect 12492 46152 12498 46164
rect 359458 46152 359464 46164
rect 12492 46124 359464 46152
rect 12492 46112 12498 46124
rect 359458 46112 359464 46124
rect 359516 46112 359522 46164
rect 20898 46044 20904 46096
rect 20956 46084 20962 46096
rect 359642 46084 359648 46096
rect 20956 46056 359648 46084
rect 20956 46044 20962 46056
rect 359642 46044 359648 46056
rect 359700 46044 359706 46096
rect 4062 45500 4068 45552
rect 4120 45540 4126 45552
rect 381814 45540 381820 45552
rect 4120 45512 381820 45540
rect 4120 45500 4126 45512
rect 381814 45500 381820 45512
rect 381872 45500 381878 45552
rect 3510 45432 3516 45484
rect 3568 45472 3574 45484
rect 376018 45472 376024 45484
rect 3568 45444 376024 45472
rect 3568 45432 3574 45444
rect 376018 45432 376024 45444
rect 376076 45432 376082 45484
rect 3418 45364 3424 45416
rect 3476 45404 3482 45416
rect 375834 45404 375840 45416
rect 3476 45376 375840 45404
rect 3476 45364 3482 45376
rect 375834 45364 375840 45376
rect 375892 45364 375898 45416
rect 20898 45296 20904 45348
rect 20956 45336 20962 45348
rect 361390 45336 361396 45348
rect 20956 45308 361396 45336
rect 20956 45296 20962 45308
rect 361390 45296 361396 45308
rect 361448 45296 361454 45348
rect 65518 45228 65524 45280
rect 65576 45268 65582 45280
rect 376294 45268 376300 45280
rect 65576 45240 376300 45268
rect 65576 45228 65582 45240
rect 376294 45228 376300 45240
rect 376352 45228 376358 45280
rect 62022 45160 62028 45212
rect 62080 45200 62086 45212
rect 376386 45200 376392 45212
rect 62080 45172 376392 45200
rect 62080 45160 62086 45172
rect 376386 45160 376392 45172
rect 376444 45160 376450 45212
rect 58434 45092 58440 45144
rect 58492 45132 58498 45144
rect 379238 45132 379244 45144
rect 58492 45104 379244 45132
rect 58492 45092 58498 45104
rect 379238 45092 379244 45104
rect 379296 45092 379302 45144
rect 54938 45024 54944 45076
rect 54996 45064 55002 45076
rect 379422 45064 379428 45076
rect 54996 45036 379428 45064
rect 54996 45024 55002 45036
rect 379422 45024 379428 45036
rect 379480 45024 379486 45076
rect 51350 44956 51356 45008
rect 51408 44996 51414 45008
rect 378686 44996 378692 45008
rect 51408 44968 378692 44996
rect 51408 44956 51414 44968
rect 378686 44956 378692 44968
rect 378744 44956 378750 45008
rect 47854 44888 47860 44940
rect 47912 44928 47918 44940
rect 379330 44928 379336 44940
rect 47912 44900 379336 44928
rect 47912 44888 47918 44900
rect 379330 44888 379336 44900
rect 379388 44888 379394 44940
rect 7650 44820 7656 44872
rect 7708 44860 7714 44872
rect 381446 44860 381452 44872
rect 7708 44832 381452 44860
rect 7708 44820 7714 44832
rect 381446 44820 381452 44832
rect 381504 44820 381510 44872
rect 69106 44752 69112 44804
rect 69164 44792 69170 44804
rect 376478 44792 376484 44804
rect 69164 44764 376484 44792
rect 69164 44752 69170 44764
rect 376478 44752 376484 44764
rect 376536 44752 376542 44804
rect 72602 44684 72608 44736
rect 72660 44724 72666 44736
rect 376570 44724 376576 44736
rect 72660 44696 376576 44724
rect 72660 44684 72666 44696
rect 376570 44684 376576 44696
rect 376628 44684 376634 44736
rect 76190 44616 76196 44668
rect 76248 44656 76254 44668
rect 373718 44656 373724 44668
rect 76248 44628 373724 44656
rect 76248 44616 76254 44628
rect 373718 44616 373724 44628
rect 373776 44616 373782 44668
rect 111610 42712 111616 42764
rect 111668 42752 111674 42764
rect 365254 42752 365260 42764
rect 111668 42724 365260 42752
rect 111668 42712 111674 42724
rect 365254 42712 365260 42724
rect 365312 42712 365318 42764
rect 108114 42644 108120 42696
rect 108172 42684 108178 42696
rect 367922 42684 367928 42696
rect 108172 42656 367928 42684
rect 108172 42644 108178 42656
rect 367922 42644 367928 42656
rect 367980 42644 367986 42696
rect 104526 42576 104532 42628
rect 104584 42616 104590 42628
rect 368014 42616 368020 42628
rect 104584 42588 368020 42616
rect 104584 42576 104590 42588
rect 368014 42576 368020 42588
rect 368072 42576 368078 42628
rect 101030 42508 101036 42560
rect 101088 42548 101094 42560
rect 367830 42548 367836 42560
rect 101088 42520 367836 42548
rect 101088 42508 101094 42520
rect 367830 42508 367836 42520
rect 367888 42508 367894 42560
rect 97442 42440 97448 42492
rect 97500 42480 97506 42492
rect 368106 42480 368112 42492
rect 97500 42452 368112 42480
rect 97500 42440 97506 42452
rect 368106 42440 368112 42452
rect 368164 42440 368170 42492
rect 93946 42372 93952 42424
rect 94004 42412 94010 42424
rect 370958 42412 370964 42424
rect 94004 42384 370964 42412
rect 94004 42372 94010 42384
rect 370958 42372 370964 42384
rect 371016 42372 371022 42424
rect 90358 42304 90364 42356
rect 90416 42344 90422 42356
rect 370866 42344 370872 42356
rect 90416 42316 370872 42344
rect 90416 42304 90422 42316
rect 370866 42304 370872 42316
rect 370924 42304 370930 42356
rect 86862 42236 86868 42288
rect 86920 42276 86926 42288
rect 370774 42276 370780 42288
rect 86920 42248 370780 42276
rect 86920 42236 86926 42248
rect 370774 42236 370780 42248
rect 370832 42236 370838 42288
rect 83274 42168 83280 42220
rect 83332 42208 83338 42220
rect 370682 42208 370688 42220
rect 83332 42180 370688 42208
rect 83332 42168 83338 42180
rect 370682 42168 370688 42180
rect 370740 42168 370746 42220
rect 79686 42100 79692 42152
rect 79744 42140 79750 42152
rect 373442 42140 373448 42152
rect 79744 42112 373448 42140
rect 79744 42100 79750 42112
rect 373442 42100 373448 42112
rect 373500 42100 373506 42152
rect 12342 42032 12348 42084
rect 12400 42072 12406 42084
rect 373534 42072 373540 42084
rect 12400 42044 373540 42072
rect 12400 42032 12406 42044
rect 373534 42032 373540 42044
rect 373592 42032 373598 42084
rect 115198 41964 115204 42016
rect 115256 42004 115262 42016
rect 365346 42004 365352 42016
rect 115256 41976 365352 42004
rect 115256 41964 115262 41976
rect 365346 41964 365352 41976
rect 365404 41964 365410 42016
rect 461578 41352 461584 41404
rect 461636 41392 461642 41404
rect 536834 41392 536840 41404
rect 461636 41364 536840 41392
rect 461636 41352 461642 41364
rect 536834 41352 536840 41364
rect 536892 41352 536898 41404
rect 118786 39992 118792 40044
rect 118844 40032 118850 40044
rect 362494 40032 362500 40044
rect 118844 40004 362500 40032
rect 118844 39992 118850 40004
rect 362494 39992 362500 40004
rect 362552 39992 362558 40044
rect 63218 39924 63224 39976
rect 63276 39964 63282 39976
rect 372338 39964 372344 39976
rect 63276 39936 372344 39964
rect 63276 39924 63282 39936
rect 372338 39924 372344 39936
rect 372396 39924 372402 39976
rect 59630 39856 59636 39908
rect 59688 39896 59694 39908
rect 369394 39896 369400 39908
rect 59688 39868 369400 39896
rect 59688 39856 59694 39868
rect 369394 39856 369400 39868
rect 369452 39856 369458 39908
rect 56042 39788 56048 39840
rect 56100 39828 56106 39840
rect 370590 39828 370596 39840
rect 56100 39800 370596 39828
rect 56100 39788 56106 39800
rect 370590 39788 370596 39800
rect 370648 39788 370654 39840
rect 52546 39720 52552 39772
rect 52604 39760 52610 39772
rect 369210 39760 369216 39772
rect 52604 39732 369216 39760
rect 52604 39720 52610 39732
rect 369210 39720 369216 39732
rect 369268 39720 369274 39772
rect 48958 39652 48964 39704
rect 49016 39692 49022 39704
rect 366542 39692 366548 39704
rect 49016 39664 366548 39692
rect 49016 39652 49022 39664
rect 366542 39652 366548 39664
rect 366600 39652 366606 39704
rect 40678 39584 40684 39636
rect 40736 39624 40742 39636
rect 366450 39624 366456 39636
rect 40736 39596 366456 39624
rect 40736 39584 40742 39596
rect 366450 39584 366456 39596
rect 366508 39584 366514 39636
rect 37182 39516 37188 39568
rect 37240 39556 37246 39568
rect 363966 39556 363972 39568
rect 37240 39528 363972 39556
rect 37240 39516 37246 39528
rect 363966 39516 363972 39528
rect 364024 39516 364030 39568
rect 33594 39448 33600 39500
rect 33652 39488 33658 39500
rect 362402 39488 362408 39500
rect 33652 39460 362408 39488
rect 33652 39448 33658 39460
rect 362402 39448 362408 39460
rect 362460 39448 362466 39500
rect 26510 39380 26516 39432
rect 26568 39420 26574 39432
rect 365162 39420 365168 39432
rect 26568 39392 365168 39420
rect 26568 39380 26574 39392
rect 365162 39380 365168 39392
rect 365220 39380 365226 39432
rect 4062 39312 4068 39364
rect 4120 39352 4126 39364
rect 368198 39352 368204 39364
rect 4120 39324 368204 39352
rect 4120 39312 4126 39324
rect 368198 39312 368204 39324
rect 368256 39312 368262 39364
rect 122282 39244 122288 39296
rect 122340 39284 122346 39296
rect 362310 39284 362316 39296
rect 122340 39256 362316 39284
rect 122340 39244 122346 39256
rect 362310 39244 362316 39256
rect 362368 39244 362374 39296
rect 102226 37204 102232 37256
rect 102284 37244 102290 37256
rect 377766 37244 377772 37256
rect 102284 37216 377772 37244
rect 102284 37204 102290 37216
rect 377766 37204 377772 37216
rect 377824 37204 377830 37256
rect 98638 37136 98644 37188
rect 98696 37176 98702 37188
rect 379146 37176 379152 37188
rect 98696 37148 379152 37176
rect 98696 37136 98702 37148
rect 379146 37136 379152 37148
rect 379204 37136 379210 37188
rect 95142 37068 95148 37120
rect 95200 37108 95206 37120
rect 377582 37108 377588 37120
rect 95200 37080 377588 37108
rect 95200 37068 95206 37080
rect 377582 37068 377588 37080
rect 377640 37068 377646 37120
rect 91554 37000 91560 37052
rect 91612 37040 91618 37052
rect 375098 37040 375104 37052
rect 91612 37012 375104 37040
rect 91612 37000 91618 37012
rect 375098 37000 375104 37012
rect 375156 37000 375162 37052
rect 87966 36932 87972 36984
rect 88024 36972 88030 36984
rect 375006 36972 375012 36984
rect 88024 36944 375012 36972
rect 88024 36932 88030 36944
rect 375006 36932 375012 36944
rect 375064 36932 375070 36984
rect 84470 36864 84476 36916
rect 84528 36904 84534 36916
rect 376202 36904 376208 36916
rect 84528 36876 376208 36904
rect 84528 36864 84534 36876
rect 376202 36864 376208 36876
rect 376260 36864 376266 36916
rect 80882 36796 80888 36848
rect 80940 36836 80946 36848
rect 374914 36836 374920 36848
rect 80940 36808 374920 36836
rect 80940 36796 80946 36808
rect 374914 36796 374920 36808
rect 374972 36796 374978 36848
rect 77386 36728 77392 36780
rect 77444 36768 77450 36780
rect 372062 36768 372068 36780
rect 77444 36740 372068 36768
rect 77444 36728 77450 36740
rect 372062 36728 372068 36740
rect 372120 36728 372126 36780
rect 73798 36660 73804 36712
rect 73856 36700 73862 36712
rect 373350 36700 373356 36712
rect 73856 36672 373356 36700
rect 73856 36660 73862 36672
rect 373350 36660 373356 36672
rect 373408 36660 373414 36712
rect 70302 36592 70308 36644
rect 70360 36632 70366 36644
rect 371970 36632 371976 36644
rect 70360 36604 371976 36632
rect 70360 36592 70366 36604
rect 371970 36592 371976 36604
rect 372028 36592 372034 36644
rect 66714 36524 66720 36576
rect 66772 36564 66778 36576
rect 371878 36564 371884 36576
rect 66772 36536 371884 36564
rect 66772 36524 66778 36536
rect 371878 36524 371884 36536
rect 371936 36524 371942 36576
rect 105722 36456 105728 36508
rect 105780 36496 105786 36508
rect 380526 36496 380532 36508
rect 105780 36468 380532 36496
rect 105780 36456 105786 36468
rect 380526 36456 380532 36468
rect 380584 36456 380590 36508
rect 119890 34416 119896 34468
rect 119948 34456 119954 34468
rect 386046 34456 386052 34468
rect 119948 34428 386052 34456
rect 119948 34416 119954 34428
rect 386046 34416 386052 34428
rect 386104 34416 386110 34468
rect 116394 34348 116400 34400
rect 116452 34388 116458 34400
rect 383378 34388 383384 34400
rect 116452 34360 383384 34388
rect 116452 34348 116458 34360
rect 383378 34348 383384 34360
rect 383436 34348 383442 34400
rect 112806 34280 112812 34332
rect 112864 34320 112870 34332
rect 380434 34320 380440 34332
rect 112864 34292 380440 34320
rect 112864 34280 112870 34292
rect 380434 34280 380440 34292
rect 380492 34280 380498 34332
rect 109310 34212 109316 34264
rect 109368 34252 109374 34264
rect 381354 34252 381360 34264
rect 109368 34224 381360 34252
rect 109368 34212 109374 34224
rect 381354 34212 381360 34224
rect 381412 34212 381418 34264
rect 45462 34144 45468 34196
rect 45520 34184 45526 34196
rect 372246 34184 372252 34196
rect 45520 34156 372252 34184
rect 45520 34144 45526 34156
rect 372246 34144 372252 34156
rect 372304 34144 372310 34196
rect 41874 34076 41880 34128
rect 41932 34116 41938 34128
rect 369118 34116 369124 34128
rect 41932 34088 369124 34116
rect 41932 34076 41938 34088
rect 369118 34076 369124 34088
rect 369176 34076 369182 34128
rect 50154 34008 50160 34060
rect 50212 34048 50218 34060
rect 377674 34048 377680 34060
rect 50212 34020 377680 34048
rect 50212 34008 50218 34020
rect 377674 34008 377680 34020
rect 377732 34008 377738 34060
rect 34790 33940 34796 33992
rect 34848 33980 34854 33992
rect 363874 33980 363880 33992
rect 34848 33952 363880 33980
rect 34848 33940 34854 33952
rect 363874 33940 363880 33952
rect 363932 33940 363938 33992
rect 31294 33872 31300 33924
rect 31352 33912 31358 33924
rect 361206 33912 361212 33924
rect 31352 33884 361212 33912
rect 31352 33872 31358 33884
rect 361206 33872 361212 33884
rect 361264 33872 361270 33924
rect 23014 33804 23020 33856
rect 23072 33844 23078 33856
rect 384850 33844 384856 33856
rect 23072 33816 384856 33844
rect 23072 33804 23078 33816
rect 384850 33804 384856 33816
rect 384908 33804 384914 33856
rect 18230 33736 18236 33788
rect 18288 33776 18294 33788
rect 383470 33776 383476 33788
rect 18288 33748 383476 33776
rect 18288 33736 18294 33748
rect 383470 33736 383476 33748
rect 383528 33736 383534 33788
rect 123478 33668 123484 33720
rect 123536 33708 123542 33720
rect 385678 33708 385684 33720
rect 123536 33680 385684 33708
rect 123536 33668 123542 33680
rect 385678 33668 385684 33680
rect 385736 33668 385742 33720
rect 2866 33056 2872 33108
rect 2924 33096 2930 33108
rect 383102 33096 383108 33108
rect 2924 33068 383108 33096
rect 2924 33056 2930 33068
rect 383102 33056 383108 33068
rect 383160 33056 383166 33108
rect 562318 33056 562324 33108
rect 562376 33096 562382 33108
rect 580166 33096 580172 33108
rect 562376 33068 580172 33096
rect 562376 33056 562382 33068
rect 580166 33056 580172 33068
rect 580224 33056 580230 33108
rect 99834 31696 99840 31748
rect 99892 31736 99898 31748
rect 366634 31736 366640 31748
rect 99892 31708 366640 31736
rect 99892 31696 99898 31708
rect 366634 31696 366640 31708
rect 366692 31696 366698 31748
rect 386138 31696 386144 31748
rect 386196 31736 386202 31748
rect 460198 31736 460204 31748
rect 386196 31708 460204 31736
rect 386196 31696 386202 31708
rect 460198 31696 460204 31708
rect 460256 31696 460262 31748
rect 96246 31628 96252 31680
rect 96304 31668 96310 31680
rect 376110 31668 376116 31680
rect 96304 31640 376116 31668
rect 96304 31628 96310 31640
rect 376110 31628 376116 31640
rect 376168 31628 376174 31680
rect 92750 31560 92756 31612
rect 92808 31600 92814 31612
rect 379054 31600 379060 31612
rect 92808 31572 379060 31600
rect 92808 31560 92814 31572
rect 379054 31560 379060 31572
rect 379112 31560 379118 31612
rect 85666 31492 85672 31544
rect 85724 31532 85730 31544
rect 382182 31532 382188 31544
rect 85724 31504 382188 31532
rect 85724 31492 85730 31504
rect 382182 31492 382188 31504
rect 382240 31492 382246 31544
rect 78582 31424 78588 31476
rect 78640 31464 78646 31476
rect 385954 31464 385960 31476
rect 78640 31436 385960 31464
rect 78640 31424 78646 31436
rect 385954 31424 385960 31436
rect 386012 31424 386018 31476
rect 71498 31356 71504 31408
rect 71556 31396 71562 31408
rect 383194 31396 383200 31408
rect 71556 31368 383200 31396
rect 71556 31356 71562 31368
rect 383194 31356 383200 31368
rect 383252 31356 383258 31408
rect 67910 31288 67916 31340
rect 67968 31328 67974 31340
rect 380250 31328 380256 31340
rect 67968 31300 380256 31328
rect 67968 31288 67974 31300
rect 380250 31288 380256 31300
rect 380308 31288 380314 31340
rect 64322 31220 64328 31272
rect 64380 31260 64386 31272
rect 377490 31260 377496 31272
rect 64380 31232 377496 31260
rect 64380 31220 64386 31232
rect 377490 31220 377496 31232
rect 377548 31220 377554 31272
rect 60826 31152 60832 31204
rect 60884 31192 60890 31204
rect 383286 31192 383292 31204
rect 60884 31164 383292 31192
rect 60884 31152 60890 31164
rect 383286 31152 383292 31164
rect 383344 31152 383350 31204
rect 57238 31084 57244 31136
rect 57296 31124 57302 31136
rect 380342 31124 380348 31136
rect 57296 31096 380348 31124
rect 57296 31084 57302 31096
rect 380342 31084 380348 31096
rect 380400 31084 380406 31136
rect 14734 31016 14740 31068
rect 14792 31056 14798 31068
rect 384666 31056 384672 31068
rect 14792 31028 384672 31056
rect 14792 31016 14798 31028
rect 384666 31016 384672 31028
rect 384724 31016 384730 31068
rect 106918 30948 106924 31000
rect 106976 30988 106982 31000
rect 369302 30988 369308 31000
rect 106976 30960 369308 30988
rect 106976 30948 106982 30960
rect 369302 30948 369308 30960
rect 369360 30948 369366 31000
rect 124674 28908 124680 28960
rect 124732 28948 124738 28960
rect 380158 28948 380164 28960
rect 124732 28920 380164 28948
rect 124732 28908 124738 28920
rect 380158 28908 380164 28920
rect 380216 28908 380222 28960
rect 117590 28840 117596 28892
rect 117648 28880 117654 28892
rect 373258 28880 373264 28892
rect 117648 28852 373264 28880
rect 117648 28840 117654 28852
rect 373258 28840 373264 28852
rect 373316 28840 373322 28892
rect 121086 28772 121092 28824
rect 121144 28812 121150 28824
rect 377398 28812 377404 28824
rect 121144 28784 377404 28812
rect 121144 28772 121150 28784
rect 377398 28772 377404 28784
rect 377456 28772 377462 28824
rect 114002 28704 114008 28756
rect 114060 28744 114066 28756
rect 372154 28744 372160 28756
rect 114060 28716 372160 28744
rect 114060 28704 114066 28716
rect 372154 28704 372160 28716
rect 372212 28704 372218 28756
rect 109678 28636 109684 28688
rect 109736 28676 109742 28688
rect 384942 28676 384948 28688
rect 109736 28648 384948 28676
rect 109736 28636 109742 28648
rect 384942 28636 384948 28648
rect 385000 28636 385006 28688
rect 28902 28568 28908 28620
rect 28960 28608 28966 28620
rect 383010 28608 383016 28620
rect 28960 28580 383016 28608
rect 28960 28568 28966 28580
rect 383010 28568 383016 28580
rect 383068 28568 383074 28620
rect 19426 28500 19432 28552
rect 19484 28540 19490 28552
rect 374730 28540 374736 28552
rect 19484 28512 374736 28540
rect 19484 28500 19490 28512
rect 374730 28500 374736 28512
rect 374788 28500 374794 28552
rect 43070 28432 43076 28484
rect 43128 28472 43134 28484
rect 462314 28472 462320 28484
rect 43128 28444 462320 28472
rect 43128 28432 43134 28444
rect 462314 28432 462320 28444
rect 462372 28432 462378 28484
rect 35986 28364 35992 28416
rect 36044 28404 36050 28416
rect 461026 28404 461032 28416
rect 36044 28376 461032 28404
rect 36044 28364 36050 28376
rect 461026 28364 461032 28376
rect 461084 28364 461090 28416
rect 32398 28296 32404 28348
rect 32456 28336 32462 28348
rect 462406 28336 462412 28348
rect 32456 28308 462412 28336
rect 32456 28296 32462 28308
rect 462406 28296 462412 28308
rect 462464 28296 462470 28348
rect 5258 28228 5264 28280
rect 5316 28268 5322 28280
rect 460934 28268 460940 28280
rect 5316 28240 460940 28268
rect 5316 28228 5322 28240
rect 460934 28228 460940 28240
rect 460992 28228 460998 28280
rect 3418 20612 3424 20664
rect 3476 20652 3482 20664
rect 378778 20652 378784 20664
rect 3476 20624 378784 20652
rect 3476 20612 3482 20624
rect 378778 20612 378784 20624
rect 378836 20612 378842 20664
rect 571978 20612 571984 20664
rect 572036 20652 572042 20664
rect 579982 20652 579988 20664
rect 572036 20624 579988 20652
rect 572036 20612 572042 20624
rect 579982 20612 579988 20624
rect 580040 20612 580046 20664
rect 3418 6808 3424 6860
rect 3476 6848 3482 6860
rect 381630 6848 381636 6860
rect 3476 6820 381636 6848
rect 3476 6808 3482 6820
rect 381630 6808 381636 6820
rect 381688 6808 381694 6860
rect 566458 6808 566464 6860
rect 566516 6848 566522 6860
rect 580166 6848 580172 6860
rect 566516 6820 580172 6848
rect 566516 6808 566522 6820
rect 580166 6808 580172 6820
rect 580224 6808 580230 6860
rect 82078 4088 82084 4140
rect 82136 4128 82142 4140
rect 370498 4128 370504 4140
rect 82136 4100 370504 4128
rect 82136 4088 82142 4100
rect 370498 4088 370504 4100
rect 370556 4088 370562 4140
rect 74994 4020 75000 4072
rect 75052 4060 75058 4072
rect 367738 4060 367744 4072
rect 75052 4032 367744 4060
rect 75052 4020 75058 4032
rect 367738 4020 367744 4032
rect 367796 4020 367802 4072
rect 53742 3952 53748 4004
rect 53800 3992 53806 4004
rect 364978 3992 364984 4004
rect 53800 3964 364984 3992
rect 53800 3952 53806 3964
rect 364978 3952 364984 3964
rect 365036 3952 365042 4004
rect 46658 3884 46664 3936
rect 46716 3924 46722 3936
rect 363690 3924 363696 3936
rect 46716 3896 363696 3924
rect 46716 3884 46722 3896
rect 363690 3884 363696 3896
rect 363748 3884 363754 3936
rect 39574 3816 39580 3868
rect 39632 3856 39638 3868
rect 360930 3856 360936 3868
rect 39632 3828 360936 3856
rect 39632 3816 39638 3828
rect 360930 3816 360936 3828
rect 360988 3816 360994 3868
rect 38378 3748 38384 3800
rect 38436 3788 38442 3800
rect 366358 3788 366364 3800
rect 38436 3760 366364 3788
rect 38436 3748 38442 3760
rect 366358 3748 366364 3760
rect 366416 3748 366422 3800
rect 30098 3680 30104 3732
rect 30156 3720 30162 3732
rect 363598 3720 363604 3732
rect 30156 3692 363604 3720
rect 30156 3680 30162 3692
rect 363598 3680 363604 3692
rect 363656 3680 363662 3732
rect 44266 3612 44272 3664
rect 44324 3652 44330 3664
rect 382918 3652 382924 3664
rect 44324 3624 382924 3652
rect 44324 3612 44330 3624
rect 382918 3612 382924 3624
rect 382976 3612 382982 3664
rect 21818 3544 21824 3596
rect 21876 3584 21882 3596
rect 363782 3584 363788 3596
rect 21876 3556 363788 3584
rect 21876 3544 21882 3556
rect 363782 3544 363788 3556
rect 363840 3544 363846 3596
rect 27706 3476 27712 3528
rect 27764 3516 27770 3528
rect 385862 3516 385868 3528
rect 27764 3488 385868 3516
rect 27764 3476 27770 3488
rect 385862 3476 385868 3488
rect 385920 3476 385926 3528
rect 24210 3408 24216 3460
rect 24268 3448 24274 3460
rect 385770 3448 385776 3460
rect 24268 3420 385776 3448
rect 24268 3408 24274 3420
rect 385770 3408 385776 3420
rect 385828 3408 385834 3460
rect 89162 3340 89168 3392
rect 89220 3380 89226 3392
rect 361114 3380 361120 3392
rect 89220 3352 361120 3380
rect 89220 3340 89226 3352
rect 361114 3340 361120 3352
rect 361172 3340 361178 3392
rect 103330 3272 103336 3324
rect 103388 3312 103394 3324
rect 361022 3312 361028 3324
rect 103388 3284 361028 3312
rect 103388 3272 103394 3284
rect 361022 3272 361028 3284
rect 361080 3272 361086 3324
rect 6454 3204 6460 3256
rect 6512 3244 6518 3256
rect 109678 3244 109684 3256
rect 6512 3216 109684 3244
rect 6512 3204 6518 3216
rect 109678 3204 109684 3216
rect 109736 3204 109742 3256
rect 110506 3204 110512 3256
rect 110564 3244 110570 3256
rect 360838 3244 360844 3256
rect 110564 3216 360844 3244
rect 110564 3204 110570 3216
rect 360838 3204 360844 3216
rect 360896 3204 360902 3256
<< via1 >>
rect 397460 700816 397512 700868
rect 444104 700816 444156 700868
rect 364984 700748 365036 700800
rect 446496 700748 446548 700800
rect 332508 700680 332560 700732
rect 445024 700680 445076 700732
rect 267648 700612 267700 700664
rect 449256 700612 449308 700664
rect 235172 700544 235224 700596
rect 449164 700544 449216 700596
rect 170312 700476 170364 700528
rect 446404 700476 446456 700528
rect 154120 700408 154172 700460
rect 445116 700408 445168 700460
rect 105452 700340 105504 700392
rect 444196 700340 444248 700392
rect 445668 700340 445720 700392
rect 478512 700340 478564 700392
rect 8116 700272 8168 700324
rect 418804 700272 418856 700324
rect 447876 700272 447928 700324
rect 494796 700272 494848 700324
rect 571984 696940 572036 696992
rect 580172 696940 580224 696992
rect 218980 692044 219032 692096
rect 446588 692044 446640 692096
rect 283840 687896 283892 687948
rect 446680 687896 446732 687948
rect 348792 686468 348844 686520
rect 445208 686468 445260 686520
rect 137836 685244 137888 685296
rect 446772 685244 446824 685296
rect 89168 685176 89220 685228
rect 416044 685176 416096 685228
rect 72976 685108 73028 685160
rect 418896 685108 418948 685160
rect 3884 684496 3936 684548
rect 445576 684496 445628 684548
rect 24124 683884 24176 683936
rect 359464 683884 359516 683936
rect 19984 683816 20036 683868
rect 418988 683816 419040 683868
rect 21364 683748 21416 683800
rect 420644 683748 420696 683800
rect 4068 683680 4120 683732
rect 420184 683680 420236 683732
rect 3516 683612 3568 683664
rect 420368 683612 420420 683664
rect 3332 683544 3384 683596
rect 420276 683544 420328 683596
rect 3700 683476 3752 683528
rect 420736 683476 420788 683528
rect 3424 683408 3476 683460
rect 420552 683408 420604 683460
rect 3608 683340 3660 683392
rect 420828 683340 420880 683392
rect 3792 683272 3844 683324
rect 445300 683272 445352 683324
rect 3976 683204 4028 683256
rect 445484 683204 445536 683256
rect 3240 683136 3292 683188
rect 445392 683136 445444 683188
rect 573364 683136 573416 683188
rect 580172 683136 580224 683188
rect 19248 682728 19300 682780
rect 24124 682728 24176 682780
rect 3240 682660 3292 682712
rect 446956 682660 447008 682712
rect 17224 680348 17276 680400
rect 19248 680348 19300 680400
rect 361764 678988 361816 679040
rect 387064 678988 387116 679040
rect 570604 670692 570656 670744
rect 580172 670692 580224 670744
rect 447784 669944 447836 669996
rect 462320 669944 462372 669996
rect 361764 667904 361816 667956
rect 382924 667904 382976 667956
rect 14188 660968 14240 661020
rect 17224 661036 17276 661088
rect 3148 658180 3200 658232
rect 19984 658180 20036 658232
rect 361764 656888 361816 656940
rect 381544 656888 381596 656940
rect 11704 656616 11756 656668
rect 14188 656616 14240 656668
rect 361764 645872 361816 645924
rect 378784 645872 378836 645924
rect 10600 645804 10652 645856
rect 11704 645804 11756 645856
rect 5540 643696 5592 643748
rect 10600 643696 10652 643748
rect 4804 640296 4856 640348
rect 5540 640296 5592 640348
rect 361580 634788 361632 634840
rect 403624 634788 403676 634840
rect 3700 631320 3752 631372
rect 20904 631320 20956 631372
rect 361580 623772 361632 623824
rect 376024 623772 376076 623824
rect 569224 616836 569276 616888
rect 580172 616836 580224 616888
rect 361580 612756 361632 612808
rect 406384 612756 406436 612808
rect 361764 601672 361816 601724
rect 374644 601672 374696 601724
rect 457628 600584 457680 600636
rect 461584 600584 461636 600636
rect 457720 600244 457772 600296
rect 461676 600244 461728 600296
rect 460020 599836 460072 599888
rect 463700 599836 463752 599888
rect 458640 599700 458692 599752
rect 465080 599700 465132 599752
rect 458824 599632 458876 599684
rect 466460 599632 466512 599684
rect 457444 599564 457496 599616
rect 469864 599564 469916 599616
rect 515404 599564 515456 599616
rect 580264 599564 580316 599616
rect 458732 598340 458784 598392
rect 465172 598340 465224 598392
rect 460112 598272 460164 598324
rect 470600 598272 470652 598324
rect 457536 598204 457588 598256
rect 468484 598204 468536 598256
rect 488632 598204 488684 598256
rect 494060 598204 494112 598256
rect 459928 596980 459980 597032
rect 463792 596980 463844 597032
rect 458916 596844 458968 596896
rect 466552 596844 466604 596896
rect 450544 596776 450596 596828
rect 494980 596776 495032 596828
rect 457352 596164 457404 596216
rect 462964 596164 463016 596216
rect 457812 595416 457864 595468
rect 468576 595416 468628 595468
rect 460204 594396 460256 594448
rect 462320 594396 462372 594448
rect 457260 592628 457312 592680
rect 465724 592628 465776 592680
rect 361764 590656 361816 590708
rect 407764 590656 407816 590708
rect 519544 590656 519596 590708
rect 580172 590656 580224 590708
rect 361764 579640 361816 579692
rect 371884 579640 371936 579692
rect 574744 576852 574796 576904
rect 580172 576852 580224 576904
rect 361580 568760 361632 568812
rect 363604 568760 363656 568812
rect 359464 561620 359516 561672
rect 362224 561620 362276 561672
rect 361672 557540 361724 557592
rect 370504 557540 370556 557592
rect 362224 551284 362276 551336
rect 369124 551284 369176 551336
rect 361764 546456 361816 546508
rect 367744 546456 367796 546508
rect 459468 544348 459520 544400
rect 470876 544348 470928 544400
rect 518164 536800 518216 536852
rect 580172 536800 580224 536852
rect 361580 535440 361632 535492
rect 363696 535440 363748 535492
rect 361580 524696 361632 524748
rect 363788 524696 363840 524748
rect 369124 522248 369176 522300
rect 378876 522248 378928 522300
rect 457904 520888 457956 520940
rect 467932 520888 467984 520940
rect 482928 520888 482980 520940
rect 520280 520888 520332 520940
rect 464344 520276 464396 520328
rect 488632 520276 488684 520328
rect 458088 519528 458140 519580
rect 465816 519528 465868 519580
rect 459836 518372 459888 518424
rect 462412 518372 462464 518424
rect 457996 518236 458048 518288
rect 469956 518236 470008 518288
rect 449808 518168 449860 518220
rect 470048 518168 470100 518220
rect 494244 518168 494296 518220
rect 476028 517556 476080 517608
rect 494152 517556 494204 517608
rect 450360 517488 450412 517540
rect 494060 517488 494112 517540
rect 482284 517420 482336 517472
rect 450636 516808 450688 516860
rect 476028 516808 476080 516860
rect 449992 516740 450044 516792
rect 492128 516740 492180 516792
rect 3976 514768 4028 514820
rect 4804 514768 4856 514820
rect 502248 514020 502300 514072
rect 545120 514020 545172 514072
rect 361764 513340 361816 513392
rect 410524 513340 410576 513392
rect 492128 512592 492180 512644
rect 535460 512592 535512 512644
rect 494060 509872 494112 509924
rect 538220 509872 538272 509924
rect 494152 508512 494204 508564
rect 532700 508512 532752 508564
rect 378876 508444 378928 508496
rect 381268 508444 381320 508496
rect 495072 505724 495124 505776
rect 529940 505724 529992 505776
rect 361764 502324 361816 502376
rect 411904 502324 411956 502376
rect 381268 501576 381320 501628
rect 387340 501576 387392 501628
rect 387340 498108 387392 498160
rect 393964 498108 394016 498160
rect 468668 497768 468720 497820
rect 483848 497768 483900 497820
rect 464436 497700 464488 497752
rect 485044 497700 485096 497752
rect 457628 497632 457680 497684
rect 481640 497632 481692 497684
rect 457444 497564 457496 497616
rect 482652 497564 482704 497616
rect 453304 497496 453356 497548
rect 480260 497496 480312 497548
rect 458824 497428 458876 497480
rect 486240 497428 486292 497480
rect 455328 497020 455380 497072
rect 459560 497020 459612 497072
rect 456524 496952 456576 497004
rect 461032 496952 461084 497004
rect 455144 496884 455196 496936
rect 458088 496884 458140 496936
rect 452568 496816 452620 496868
rect 453672 496816 453724 496868
rect 453948 496816 454000 496868
rect 456616 496816 456668 496868
rect 361764 491308 361816 491360
rect 414664 491308 414716 491360
rect 515496 484372 515548 484424
rect 580172 484372 580224 484424
rect 361764 480224 361816 480276
rect 419080 480224 419132 480276
rect 361764 469208 361816 469260
rect 417424 469208 417476 469260
rect 393964 466284 394016 466336
rect 398104 466284 398156 466336
rect 449808 464312 449860 464364
rect 525800 464312 525852 464364
rect 494704 462408 494756 462460
rect 527640 462408 527692 462460
rect 450544 462340 450596 462392
rect 542360 462340 542412 462392
rect 449716 461048 449768 461100
rect 524696 461048 524748 461100
rect 461860 460980 461912 461032
rect 553860 460980 553912 461032
rect 458916 460912 458968 460964
rect 550916 460912 550968 460964
rect 361764 458192 361816 458244
rect 385776 458192 385828 458244
rect 576124 456764 576176 456816
rect 580172 456764 580224 456816
rect 488264 456016 488316 456068
rect 494704 456016 494756 456068
rect 460204 455472 460256 455524
rect 488264 455472 488316 455524
rect 452016 455404 452068 455456
rect 480996 455404 481048 455456
rect 449624 454724 449676 454776
rect 487160 454724 487212 454776
rect 449532 454656 449584 454708
rect 489920 454656 489972 454708
rect 461952 454044 462004 454096
rect 473728 454044 473780 454096
rect 447324 447924 447376 447976
rect 458916 447924 458968 447976
rect 447232 447856 447284 447908
rect 448428 447856 448480 447908
rect 461952 447856 462004 447908
rect 447140 447788 447192 447840
rect 448060 447788 448112 447840
rect 461860 447788 461912 447840
rect 422484 447312 422536 447364
rect 447232 447312 447284 447364
rect 437388 447244 437440 447296
rect 447140 447244 447192 447296
rect 432420 447176 432472 447228
rect 447324 447176 447376 447228
rect 447968 447176 448020 447228
rect 427728 444388 427780 444440
rect 446312 444388 446364 444440
rect 442632 444320 442684 444372
rect 446220 444320 446272 444372
rect 361764 436092 361816 436144
rect 419172 436092 419224 436144
rect 569316 430584 569368 430636
rect 580172 430584 580224 430636
rect 458088 429904 458140 429956
rect 474280 429904 474332 429956
rect 459468 429836 459520 429888
rect 479616 429836 479668 429888
rect 475384 429156 475436 429208
rect 476948 429156 477000 429208
rect 457536 427048 457588 427100
rect 471612 427048 471664 427100
rect 503628 424328 503680 424380
rect 557540 424328 557592 424380
rect 529204 423580 529256 423632
rect 530216 423580 530268 423632
rect 530584 423580 530636 423632
rect 532792 423580 532844 423632
rect 502984 423512 503036 423564
rect 523776 423512 523828 423564
rect 522304 423444 522356 423496
rect 549536 423444 549588 423496
rect 484308 423376 484360 423428
rect 522488 423376 522540 423428
rect 523684 423376 523736 423428
rect 552112 423376 552164 423428
rect 487068 423308 487120 423360
rect 526352 423308 526404 423360
rect 526444 423308 526496 423360
rect 554688 423308 554740 423360
rect 488264 423240 488316 423292
rect 528928 423240 528980 423292
rect 489644 423172 489696 423224
rect 531504 423172 531556 423224
rect 498108 423104 498160 423156
rect 545672 423104 545724 423156
rect 499304 423036 499356 423088
rect 548248 423036 548300 423088
rect 444288 422968 444340 423020
rect 447876 422968 447928 423020
rect 500684 422968 500736 423020
rect 550824 422968 550876 423020
rect 502248 422900 502300 422952
rect 553400 422900 553452 422952
rect 484216 421540 484268 421592
rect 521200 421540 521252 421592
rect 533436 421540 533488 421592
rect 580356 421540 580408 421592
rect 495348 420180 495400 420232
rect 541808 420180 541860 420232
rect 362316 418752 362368 418804
rect 442264 418752 442316 418804
rect 425336 417732 425388 417784
rect 507860 417732 507912 417784
rect 424692 417664 424744 417716
rect 506480 417664 506532 417716
rect 422116 417596 422168 417648
rect 503996 417596 504048 417648
rect 421472 417528 421524 417580
rect 503720 417528 503772 417580
rect 424048 417460 424100 417512
rect 506572 417460 506624 417512
rect 425980 417392 426032 417444
rect 507952 417392 508004 417444
rect 398104 416100 398156 416152
rect 409144 416100 409196 416152
rect 362224 416032 362276 416084
rect 436744 416032 436796 416084
rect 486976 416032 487028 416084
rect 527640 416032 527692 416084
rect 423128 415964 423180 416016
rect 423588 415964 423640 416016
rect 361580 413992 361632 414044
rect 443644 413992 443696 414044
rect 511264 404336 511316 404388
rect 580172 404336 580224 404388
rect 361580 402976 361632 403028
rect 439504 402976 439556 403028
rect 497924 400868 497976 400920
rect 546500 400868 546552 400920
rect 496728 399440 496780 399492
rect 543740 399440 543792 399492
rect 494612 398080 494664 398132
rect 539600 398080 539652 398132
rect 493968 396720 494020 396772
rect 538220 396720 538272 396772
rect 462228 395292 462280 395344
rect 489920 395292 489972 395344
rect 493140 395292 493192 395344
rect 536840 395292 536892 395344
rect 462596 393932 462648 393984
rect 484400 393932 484452 393984
rect 491668 393932 491720 393984
rect 534172 393932 534224 393984
rect 458180 392708 458232 392760
rect 475384 392708 475436 392760
rect 448244 392640 448296 392692
rect 464436 392640 464488 392692
rect 461124 392572 461176 392624
rect 487160 392572 487212 392624
rect 490564 392572 490616 392624
rect 534080 392572 534132 392624
rect 361580 391960 361632 392012
rect 443736 391960 443788 392012
rect 495716 391280 495768 391332
rect 542360 391280 542412 391332
rect 423496 391212 423548 391264
rect 506020 391212 506072 391264
rect 462780 389852 462832 389904
rect 481640 389852 481692 389904
rect 492036 389852 492088 389904
rect 535460 389852 535512 389904
rect 423588 389784 423640 389836
rect 505284 389784 505336 389836
rect 463700 389240 463752 389292
rect 464436 389240 464488 389292
rect 466460 389240 466512 389292
rect 467380 389240 467432 389292
rect 486424 389240 486476 389292
rect 487068 389240 487120 389292
rect 497464 389240 497516 389292
rect 498108 389240 498160 389292
rect 506480 389240 506532 389292
rect 507124 389240 507176 389292
rect 453028 389104 453080 389156
rect 454040 389104 454092 389156
rect 456708 389104 456760 389156
rect 457536 389104 457588 389156
rect 460388 389104 460440 389156
rect 462596 389104 462648 389156
rect 469956 388968 470008 389020
rect 473636 388968 473688 389020
rect 465816 388900 465868 388952
rect 469404 388900 469456 388952
rect 469864 388900 469916 388952
rect 475844 388900 475896 388952
rect 502340 388900 502392 388952
rect 468484 388832 468536 388884
rect 476580 388832 476632 388884
rect 468576 388764 468628 388816
rect 480260 388764 480312 388816
rect 484676 388764 484728 388816
rect 502984 388764 503036 388816
rect 526444 388764 526496 388816
rect 467104 388696 467156 388748
rect 465724 388628 465776 388680
rect 469220 388628 469272 388680
rect 469404 388696 469456 388748
rect 480996 388696 481048 388748
rect 500868 388696 500920 388748
rect 523684 388696 523736 388748
rect 481732 388628 481784 388680
rect 499396 388628 499448 388680
rect 522304 388628 522356 388680
rect 461676 388560 461728 388612
rect 478788 388560 478840 388612
rect 485412 388560 485464 388612
rect 524420 388560 524472 388612
rect 461584 388492 461636 388544
rect 478052 388492 478104 388544
rect 489828 388492 489880 388544
rect 530584 388492 530636 388544
rect 447416 388424 447468 388476
rect 458824 388424 458876 388476
rect 461768 388424 461820 388476
rect 482468 388424 482520 388476
rect 488356 388424 488408 388476
rect 529204 388424 529256 388476
rect 462964 388356 463016 388408
rect 469956 388356 470008 388408
rect 459652 388152 459704 388204
rect 462780 388152 462832 388204
rect 450728 387336 450780 387388
rect 460204 387336 460256 387388
rect 447600 387268 447652 387320
rect 457444 387268 457496 387320
rect 447692 387200 447744 387252
rect 468668 387200 468720 387252
rect 448980 387132 449032 387184
rect 491300 387132 491352 387184
rect 441528 387064 441580 387116
rect 447784 387064 447836 387116
rect 449440 387064 449492 387116
rect 513380 387064 513432 387116
rect 448428 386588 448480 386640
rect 553952 386588 554004 386640
rect 385684 386520 385736 386572
rect 512092 386520 512144 386572
rect 380164 386452 380216 386504
rect 512276 386452 512328 386504
rect 373264 386384 373316 386436
rect 512000 386384 512052 386436
rect 448152 385976 448204 386028
rect 453304 385976 453356 386028
rect 447876 385636 447928 385688
rect 457352 385636 457404 385688
rect 448336 385500 448388 385552
rect 452016 385500 452068 385552
rect 449348 385432 449400 385484
rect 563428 385432 563480 385484
rect 377404 385364 377456 385416
rect 512184 385364 512236 385416
rect 387064 384956 387116 385008
rect 447140 384956 447192 385008
rect 513288 383732 513340 383784
rect 534724 383732 534776 383784
rect 512460 383664 512512 383716
rect 548524 383664 548576 383716
rect 381544 383596 381596 383648
rect 447232 383596 447284 383648
rect 382924 383528 382976 383580
rect 447140 383528 447192 383580
rect 512644 382984 512696 383036
rect 519728 382984 519780 383036
rect 513012 382916 513064 382968
rect 518256 382916 518308 382968
rect 512460 382440 512512 382492
rect 515588 382440 515640 382492
rect 378784 382168 378836 382220
rect 447140 382168 447192 382220
rect 403624 382100 403676 382152
rect 447232 382100 447284 382152
rect 361580 380876 361632 380928
rect 443828 380876 443880 380928
rect 513288 380876 513340 380928
rect 547144 380876 547196 380928
rect 376024 380808 376076 380860
rect 447140 380808 447192 380860
rect 406384 380740 406436 380792
rect 447232 380740 447284 380792
rect 512552 379720 512604 379772
rect 515680 379720 515732 379772
rect 513288 379516 513340 379568
rect 549904 379516 549956 379568
rect 374644 379448 374696 379500
rect 447140 379448 447192 379500
rect 407764 379380 407816 379432
rect 447232 379380 447284 379432
rect 512460 378224 512512 378276
rect 522304 378224 522356 378276
rect 512920 378156 512972 378208
rect 547236 378156 547288 378208
rect 363604 378088 363656 378140
rect 447232 378088 447284 378140
rect 371884 378020 371936 378072
rect 447140 378020 447192 378072
rect 513196 377408 513248 377460
rect 548616 377408 548668 377460
rect 512644 376728 512696 376780
rect 516416 376728 516468 376780
rect 367744 376660 367796 376712
rect 447232 376660 447284 376712
rect 370504 376592 370556 376644
rect 447140 376592 447192 376644
rect 513104 375980 513156 376032
rect 544384 375980 544436 376032
rect 512828 375436 512880 375488
rect 516232 375436 516284 375488
rect 512644 375368 512696 375420
rect 520280 375368 520332 375420
rect 363696 375300 363748 375352
rect 447140 375300 447192 375352
rect 363788 375232 363840 375284
rect 447232 375232 447284 375284
rect 513288 374008 513340 374060
rect 520372 374008 520424 374060
rect 410524 373940 410576 373992
rect 447140 373940 447192 373992
rect 411904 373872 411956 373924
rect 447232 373872 447284 373924
rect 512644 373736 512696 373788
rect 516324 373736 516376 373788
rect 512460 372716 512512 372768
rect 523040 372716 523092 372768
rect 512092 372648 512144 372700
rect 514760 372648 514812 372700
rect 414664 372512 414716 372564
rect 447140 372512 447192 372564
rect 419080 372444 419132 372496
rect 447232 372444 447284 372496
rect 512828 371220 512880 371272
rect 517520 371220 517572 371272
rect 385776 371152 385828 371204
rect 447232 371152 447284 371204
rect 417424 371084 417476 371136
rect 447140 371084 447192 371136
rect 512644 369928 512696 369980
rect 516968 369928 517020 369980
rect 361580 369860 361632 369912
rect 409880 369860 409932 369912
rect 513288 369860 513340 369912
rect 521660 369860 521712 369912
rect 419172 369792 419224 369844
rect 447232 369792 447284 369844
rect 436744 369724 436796 369776
rect 447140 369724 447192 369776
rect 513288 368568 513340 368620
rect 520464 368568 520516 368620
rect 512828 368500 512880 368552
rect 516508 368500 516560 368552
rect 443644 368432 443696 368484
rect 447140 368432 447192 368484
rect 442264 368364 442316 368416
rect 447232 368364 447284 368416
rect 512000 367344 512052 367396
rect 514116 367344 514168 367396
rect 513288 367208 513340 367260
rect 517888 367208 517940 367260
rect 439504 367004 439556 367056
rect 447140 367004 447192 367056
rect 443736 366936 443788 366988
rect 447232 366936 447284 366988
rect 512000 366120 512052 366172
rect 514208 366120 514260 366172
rect 513288 365712 513340 365764
rect 523132 365712 523184 365764
rect 409880 365644 409932 365696
rect 447140 365644 447192 365696
rect 443828 365576 443880 365628
rect 447232 365576 447284 365628
rect 513288 364488 513340 364540
rect 520556 364488 520608 364540
rect 512644 364352 512696 364404
rect 521752 364352 521804 364404
rect 569408 364352 569460 364404
rect 580172 364352 580224 364404
rect 409144 363604 409196 363656
rect 416136 363604 416188 363656
rect 512184 363264 512236 363316
rect 514852 363264 514904 363316
rect 432696 362992 432748 363044
rect 447140 362992 447192 363044
rect 432788 362924 432840 362976
rect 447232 362924 447284 362976
rect 513288 362924 513340 362976
rect 523224 362924 523276 362976
rect 512184 362312 512236 362364
rect 513656 362312 513708 362364
rect 443920 361632 443972 361684
rect 447232 361632 447284 361684
rect 513012 361632 513064 361684
rect 517612 361632 517664 361684
rect 432604 361564 432656 361616
rect 447140 361564 447192 361616
rect 442264 360272 442316 360324
rect 447232 360272 447284 360324
rect 513012 360272 513064 360324
rect 517704 360272 517756 360324
rect 436928 360204 436980 360256
rect 447140 360204 447192 360256
rect 513288 360204 513340 360256
rect 518900 360204 518952 360256
rect 547236 360136 547288 360188
rect 552020 360136 552072 360188
rect 534724 360068 534776 360120
rect 566740 360068 566792 360120
rect 549904 360000 549956 360052
rect 554964 360000 555016 360052
rect 548524 359932 548576 359984
rect 565268 359932 565320 359984
rect 547144 359864 547196 359916
rect 558184 359864 558236 359916
rect 515680 359796 515732 359848
rect 553768 359796 553820 359848
rect 522304 359728 522356 359780
rect 550824 359728 550876 359780
rect 443828 358844 443880 358896
rect 447232 358844 447284 358896
rect 435364 358776 435416 358828
rect 447140 358776 447192 358828
rect 548616 358708 548668 358760
rect 556712 358708 556764 358760
rect 518256 358640 518308 358692
rect 562600 358640 562652 358692
rect 519728 358572 519780 358624
rect 564072 358572 564124 358624
rect 544384 358504 544436 358556
rect 559656 358504 559708 358556
rect 515588 358436 515640 358488
rect 561128 358436 561180 358488
rect 512184 357688 512236 357740
rect 514024 357688 514076 357740
rect 512184 357552 512236 357604
rect 512368 357552 512420 357604
rect 513288 356056 513340 356108
rect 521844 356056 521896 356108
rect 513288 354696 513340 354748
rect 517980 354696 518032 354748
rect 512460 353608 512512 353660
rect 513748 353608 513800 353660
rect 513196 353472 513248 353524
rect 517796 353472 517848 353524
rect 446220 352656 446272 352708
rect 447784 352656 447836 352708
rect 512460 352520 512512 352572
rect 515036 352520 515088 352572
rect 511356 352044 511408 352096
rect 580172 352044 580224 352096
rect 513288 351976 513340 352028
rect 523316 351976 523368 352028
rect 395988 351908 396040 351960
rect 447140 351908 447192 351960
rect 513288 350888 513340 350940
rect 518992 350888 519044 350940
rect 512460 350752 512512 350804
rect 515128 350752 515180 350804
rect 407028 350548 407080 350600
rect 447140 350548 447192 350600
rect 509792 349800 509844 349852
rect 510068 349800 510120 349852
rect 513288 349664 513340 349716
rect 519176 349664 519228 349716
rect 512460 349528 512512 349580
rect 514944 349528 514996 349580
rect 512460 349120 512512 349172
rect 513840 349120 513892 349172
rect 513012 347896 513064 347948
rect 516692 347896 516744 347948
rect 361764 347760 361816 347812
rect 402244 347760 402296 347812
rect 362224 347692 362276 347744
rect 447140 347692 447192 347744
rect 512460 347624 512512 347676
rect 513932 347624 513984 347676
rect 513288 346536 513340 346588
rect 518072 346536 518124 346588
rect 416136 346400 416188 346452
rect 423680 346400 423732 346452
rect 512828 346400 512880 346452
rect 516600 346400 516652 346452
rect 512460 345584 512512 345636
rect 515220 345584 515272 345636
rect 446312 344700 446364 344752
rect 448336 344700 448388 344752
rect 513288 344360 513340 344412
rect 519084 344360 519136 344412
rect 513012 343680 513064 343732
rect 518256 343680 518308 343732
rect 513012 343136 513064 343188
rect 518348 343136 518400 343188
rect 423680 341572 423732 341624
rect 429844 341572 429896 341624
rect 513288 341232 513340 341284
rect 520648 341232 520700 341284
rect 513288 341096 513340 341148
rect 519360 341096 519412 341148
rect 438860 340960 438912 341012
rect 447140 340960 447192 341012
rect 361764 340892 361816 340944
rect 447232 340892 447284 340944
rect 513104 339600 513156 339652
rect 516784 339600 516836 339652
rect 435456 339532 435508 339584
rect 447140 339532 447192 339584
rect 513288 339532 513340 339584
rect 519728 339532 519780 339584
rect 374644 339464 374696 339516
rect 447232 339464 447284 339516
rect 513012 338648 513064 338700
rect 519268 338648 519320 338700
rect 439688 338172 439740 338224
rect 447140 338172 447192 338224
rect 436836 338104 436888 338156
rect 447232 338104 447284 338156
rect 450084 337424 450136 337476
rect 450360 337424 450412 337476
rect 402244 337356 402296 337408
rect 447324 337356 447376 337408
rect 448428 337356 448480 337408
rect 513288 337152 513340 337204
rect 520740 337152 520792 337204
rect 512736 337016 512788 337068
rect 515312 337016 515364 337068
rect 512828 336948 512880 337000
rect 516140 336948 516192 337000
rect 416780 336880 416832 336932
rect 450360 336880 450412 336932
rect 413100 336812 413152 336864
rect 450176 336812 450228 336864
rect 409420 336744 409472 336796
rect 450728 336744 450780 336796
rect 438124 336472 438176 336524
rect 447140 336472 447192 336524
rect 418988 336404 419040 336456
rect 442356 336404 442408 336456
rect 418896 336336 418948 336388
rect 442448 336336 442500 336388
rect 418804 336268 418856 336320
rect 442724 336268 442776 336320
rect 416044 336200 416096 336252
rect 439964 336200 440016 336252
rect 413652 336132 413704 336184
rect 449440 336132 449492 336184
rect 399484 336064 399536 336116
rect 447232 336064 447284 336116
rect 362224 335996 362276 336048
rect 438860 335996 438912 336048
rect 512736 335928 512788 335980
rect 515588 335928 515640 335980
rect 443736 335656 443788 335708
rect 447140 335656 447192 335708
rect 439596 335316 439648 335368
rect 447140 335316 447192 335368
rect 420552 335044 420604 335096
rect 439780 335044 439832 335096
rect 420184 334976 420236 335028
rect 439872 334976 439924 335028
rect 420828 334908 420880 334960
rect 442540 334908 442592 334960
rect 420644 334840 420696 334892
rect 442632 334840 442684 334892
rect 420276 334772 420328 334824
rect 442816 334772 442868 334824
rect 420736 334704 420788 334756
rect 444012 334704 444064 334756
rect 513012 334704 513064 334756
rect 519452 334704 519504 334756
rect 420276 334636 420328 334688
rect 444932 334636 444984 334688
rect 420092 334568 420144 334620
rect 444840 334568 444892 334620
rect 513288 334568 513340 334620
rect 520924 334568 520976 334620
rect 443644 334024 443696 334076
rect 447232 334024 447284 334076
rect 364064 333956 364116 334008
rect 447140 333956 447192 334008
rect 436744 332664 436796 332716
rect 447232 332664 447284 332716
rect 431224 332596 431276 332648
rect 447140 332596 447192 332648
rect 432788 331848 432840 331900
rect 443920 331848 443972 331900
rect 512828 331576 512880 331628
rect 520832 331576 520884 331628
rect 450084 330488 450136 330540
rect 450728 330488 450780 330540
rect 442908 330080 442960 330132
rect 447140 330080 447192 330132
rect 512828 329128 512880 329180
rect 516876 329128 516928 329180
rect 439504 329060 439556 329112
rect 447140 329060 447192 329112
rect 436008 328448 436060 328500
rect 449900 328448 449952 328500
rect 431868 327088 431920 327140
rect 449900 327088 449952 327140
rect 509792 326408 509844 326460
rect 510068 326408 510120 326460
rect 432696 324912 432748 324964
rect 442264 324912 442316 324964
rect 511908 324912 511960 324964
rect 580632 324912 580684 324964
rect 510436 323552 510488 323604
rect 580356 323552 580408 323604
rect 432604 322940 432656 322992
rect 436928 322940 436980 322992
rect 429844 322192 429896 322244
rect 448520 322192 448572 322244
rect 510528 322192 510580 322244
rect 580448 322192 580500 322244
rect 442816 321852 442868 321904
rect 471796 321920 471848 321972
rect 454546 321852 454598 321904
rect 454960 321852 455012 321904
rect 468300 321852 468352 321904
rect 574744 321920 574796 321972
rect 477500 321852 477552 321904
rect 580172 321852 580224 321904
rect 449256 321784 449308 321836
rect 480720 321784 480772 321836
rect 507216 321784 507268 321836
rect 511172 321784 511224 321836
rect 445576 321716 445628 321768
rect 472440 321716 472492 321768
rect 507400 321716 507452 321768
rect 513472 321716 513524 321768
rect 457812 321580 457864 321632
rect 458364 321512 458416 321564
rect 446496 321444 446548 321496
rect 459468 321444 459520 321496
rect 580264 321512 580316 321564
rect 570604 321444 570656 321496
rect 449164 321376 449216 321428
rect 446404 321308 446456 321360
rect 468852 321376 468904 321428
rect 573364 321376 573416 321428
rect 460020 321308 460072 321360
rect 467196 321308 467248 321360
rect 569408 321308 569460 321360
rect 460296 321240 460348 321292
rect 477960 321240 478012 321292
rect 569316 321240 569368 321292
rect 456708 321172 456760 321224
rect 511356 321172 511408 321224
rect 456984 321104 457036 321156
rect 511264 321104 511316 321156
rect 444104 321036 444156 321088
rect 480168 321036 480220 321088
rect 445024 320968 445076 321020
rect 480444 320968 480496 321020
rect 446956 320900 447008 320952
rect 461676 320900 461728 320952
rect 477684 320900 477736 320952
rect 580724 320900 580776 320952
rect 457536 320832 457588 320884
rect 580540 320832 580592 320884
rect 445484 320764 445536 320816
rect 461952 320764 462004 320816
rect 445392 320696 445444 320748
rect 461124 320696 461176 320748
rect 444012 320628 444064 320680
rect 461400 320628 461452 320680
rect 445116 320560 445168 320612
rect 470784 320560 470836 320612
rect 441528 320492 441580 320544
rect 479892 320492 479944 320544
rect 507676 320288 507728 320340
rect 514024 320288 514076 320340
rect 507768 320220 507820 320272
rect 511080 320220 511132 320272
rect 507492 320152 507544 320204
rect 510252 320152 510304 320204
rect 479340 320084 479392 320136
rect 571984 320084 572036 320136
rect 442632 320016 442684 320068
rect 462504 320016 462556 320068
rect 468576 320016 468628 320068
rect 533436 320016 533488 320068
rect 442540 319948 442592 320000
rect 462228 319948 462280 320000
rect 467748 319948 467800 320000
rect 511908 319948 511960 320000
rect 444288 319880 444340 319932
rect 458916 319880 458968 319932
rect 467472 319880 467524 319932
rect 510436 319880 510488 319932
rect 468024 319812 468076 319864
rect 510528 319812 510580 319864
rect 446680 319744 446732 319796
rect 470232 319744 470284 319796
rect 478788 319744 478840 319796
rect 519544 319744 519596 319796
rect 446588 319676 446640 319728
rect 470508 319676 470560 319728
rect 479616 319676 479668 319728
rect 519636 319676 519688 319728
rect 448520 319608 448572 319660
rect 472992 319608 473044 319660
rect 478512 319608 478564 319660
rect 518164 319608 518216 319660
rect 445208 319540 445260 319592
rect 469956 319540 470008 319592
rect 478236 319540 478288 319592
rect 515496 319540 515548 319592
rect 446864 319472 446916 319524
rect 471612 319472 471664 319524
rect 479064 319472 479116 319524
rect 515404 319472 515456 319524
rect 449440 319404 449492 319456
rect 469680 319404 469732 319456
rect 479524 319404 479576 319456
rect 483480 319404 483532 319456
rect 502524 319404 502576 319456
rect 543740 319404 543792 319456
rect 497280 319336 497332 319388
rect 533344 319336 533396 319388
rect 445300 319268 445352 319320
rect 482928 319268 482980 319320
rect 439872 319200 439924 319252
rect 482652 319200 482704 319252
rect 446772 319132 446824 319184
rect 481272 319132 481324 319184
rect 480904 319064 480956 319116
rect 483756 319064 483808 319116
rect 485872 319064 485924 319116
rect 487068 319064 487120 319116
rect 502708 319064 502760 319116
rect 503628 319064 503680 319116
rect 447600 318724 447652 318776
rect 449164 318724 449216 318776
rect 457260 318724 457312 318776
rect 576124 318724 576176 318776
rect 458088 318656 458140 318708
rect 569224 318656 569276 318708
rect 439780 318588 439832 318640
rect 483204 318588 483256 318640
rect 432052 318520 432104 318572
rect 435364 318520 435416 318572
rect 442356 318520 442408 318572
rect 482100 318520 482152 318572
rect 444932 318452 444984 318504
rect 472716 318452 472768 318504
rect 445668 318384 445720 318436
rect 469404 318384 469456 318436
rect 458916 318248 458968 318300
rect 490104 318248 490156 318300
rect 496452 318248 496504 318300
rect 539600 318248 539652 318300
rect 459100 318180 459152 318232
rect 492588 318180 492640 318232
rect 494796 318180 494848 318232
rect 540980 318180 541032 318232
rect 460756 318112 460808 318164
rect 513380 318112 513432 318164
rect 450636 318044 450688 318096
rect 457720 318044 457772 318096
rect 460664 318044 460716 318096
rect 516140 318044 516192 318096
rect 497740 317704 497792 317756
rect 498108 317704 498160 317756
rect 498660 317024 498712 317076
rect 541072 317024 541124 317076
rect 459008 316956 459060 317008
rect 491484 316956 491536 317008
rect 499764 316956 499816 317008
rect 543096 316956 543148 317008
rect 485964 316888 486016 316940
rect 529940 316888 529992 316940
rect 453304 316820 453356 316872
rect 489000 316820 489052 316872
rect 495624 316820 495676 316872
rect 543188 316820 543240 316872
rect 454684 316752 454736 316804
rect 503352 316752 503404 316804
rect 450544 316684 450596 316736
rect 504180 316684 504232 316736
rect 456432 316004 456484 316056
rect 461584 316004 461636 316056
rect 499028 316004 499080 316056
rect 499212 316004 499264 316056
rect 361764 315936 361816 315988
rect 374644 315936 374696 315988
rect 457444 315392 457496 315444
rect 491760 315392 491812 315444
rect 453396 315324 453448 315376
rect 489552 315324 489604 315376
rect 499120 315324 499172 315376
rect 539876 315324 539928 315376
rect 450636 315256 450688 315308
rect 502708 315256 502760 315308
rect 509792 314168 509844 314220
rect 510068 314168 510120 314220
rect 448520 314100 448572 314152
rect 462780 314100 462832 314152
rect 452016 314032 452068 314084
rect 492864 314032 492916 314084
rect 500316 314032 500368 314084
rect 542728 314032 542780 314084
rect 450728 313964 450780 314016
rect 503904 313964 503956 314016
rect 432696 313896 432748 313948
rect 443828 313896 443880 313948
rect 455236 313896 455288 313948
rect 463056 313896 463108 313948
rect 455604 313828 455656 313880
rect 533436 313896 533488 313948
rect 466920 313216 466972 313268
rect 580172 313216 580224 313268
rect 500040 312604 500092 312656
rect 542636 312604 542688 312656
rect 496360 312536 496412 312588
rect 539692 312536 539744 312588
rect 472624 311312 472676 311364
rect 480904 311312 480956 311364
rect 452200 311244 452252 311296
rect 494244 311244 494296 311296
rect 501972 311244 502024 311296
rect 538864 311244 538916 311296
rect 450820 311176 450872 311228
rect 504456 311176 504508 311228
rect 440884 311108 440936 311160
rect 448520 311108 448572 311160
rect 475752 311108 475804 311160
rect 544384 311108 544436 311160
rect 458824 309816 458876 309868
rect 488448 309816 488500 309868
rect 495900 309816 495952 309868
rect 542452 309816 542504 309868
rect 476304 309748 476356 309800
rect 537484 309748 537536 309800
rect 451924 308456 451976 308508
rect 488724 308456 488776 308508
rect 497004 308456 497056 308508
rect 539784 308456 539836 308508
rect 465264 308388 465316 308440
rect 548524 308388 548576 308440
rect 3516 307708 3568 307760
rect 4804 307708 4856 307760
rect 455880 307096 455932 307148
rect 576124 307096 576176 307148
rect 383016 307028 383068 307080
rect 520924 307028 520976 307080
rect 383108 306280 383160 306332
rect 464712 306280 464764 306332
rect 382004 306212 382056 306264
rect 463884 306212 463936 306264
rect 378876 306144 378928 306196
rect 463608 306144 463660 306196
rect 384488 306076 384540 306128
rect 474648 306076 474700 306128
rect 381912 306008 381964 306060
rect 474372 306008 474424 306060
rect 382096 305940 382148 305992
rect 474924 305940 474976 305992
rect 378968 305872 379020 305924
rect 474096 305872 474148 305924
rect 475476 305872 475528 305924
rect 562324 305872 562376 305924
rect 384764 305804 384816 305856
rect 484860 305804 484912 305856
rect 384580 305736 384632 305788
rect 485136 305736 485188 305788
rect 381820 305668 381872 305720
rect 484584 305668 484636 305720
rect 362316 305600 362368 305652
rect 516416 305600 516468 305652
rect 384396 305532 384448 305584
rect 464436 305532 464488 305584
rect 384304 305464 384356 305516
rect 464160 305464 464212 305516
rect 457536 305396 457588 305448
rect 490656 305396 490708 305448
rect 361764 304920 361816 304972
rect 435456 304920 435508 304972
rect 486240 304444 486292 304496
rect 530032 304444 530084 304496
rect 385776 304376 385828 304428
rect 520832 304376 520884 304428
rect 363604 304308 363656 304360
rect 512736 304308 512788 304360
rect 360936 304240 360988 304292
rect 512644 304240 512696 304292
rect 475384 303628 475436 303680
rect 479524 303628 479576 303680
rect 378600 303560 378652 303612
rect 484308 303560 484360 303612
rect 376668 303492 376720 303544
rect 484032 303492 484084 303544
rect 379336 303424 379388 303476
rect 510988 303424 511040 303476
rect 378692 303356 378744 303408
rect 510896 303356 510948 303408
rect 379244 303288 379296 303340
rect 513932 303288 513984 303340
rect 379428 303220 379480 303272
rect 515220 303220 515272 303272
rect 376576 303152 376628 303204
rect 513748 303152 513800 303204
rect 376392 303084 376444 303136
rect 513840 303084 513892 303136
rect 376484 303016 376536 303068
rect 515036 303016 515088 303068
rect 376300 302948 376352 303000
rect 515128 302948 515180 303000
rect 364984 302880 365036 302932
rect 512460 302880 512512 302932
rect 373632 302812 373684 302864
rect 473544 302812 473596 302864
rect 476580 302812 476632 302864
rect 547144 302812 547196 302864
rect 376024 302744 376076 302796
rect 473820 302744 473872 302796
rect 375932 302676 375984 302728
rect 463332 302676 463384 302728
rect 465540 301656 465592 301708
rect 559564 301656 559616 301708
rect 408408 301588 408460 301640
rect 503076 301588 503128 301640
rect 370504 301520 370556 301572
rect 512276 301520 512328 301572
rect 367744 301452 367796 301504
rect 512368 301452 512420 301504
rect 471244 301044 471296 301096
rect 473268 301044 473320 301096
rect 373724 300772 373776 300824
rect 510804 300772 510856 300824
rect 370780 300704 370832 300756
rect 509884 300704 509936 300756
rect 370688 300636 370740 300688
rect 510620 300636 510672 300688
rect 367928 300568 367980 300620
rect 509700 300568 509752 300620
rect 370872 300500 370924 300552
rect 513656 300500 513708 300552
rect 370964 300432 371016 300484
rect 514852 300432 514904 300484
rect 368112 300364 368164 300416
rect 513564 300364 513616 300416
rect 368020 300296 368072 300348
rect 516508 300296 516560 300348
rect 361028 300228 361080 300280
rect 512000 300228 512052 300280
rect 365352 300160 365404 300212
rect 516324 300160 516376 300212
rect 365260 300092 365312 300144
rect 517520 300092 517572 300144
rect 373448 300024 373500 300076
rect 509976 300024 510028 300076
rect 373540 299956 373592 300008
rect 510344 299956 510396 300008
rect 466092 299888 466144 299940
rect 551284 299888 551336 299940
rect 461584 299412 461636 299464
rect 580172 299412 580224 299464
rect 403624 298800 403676 298852
rect 502800 298800 502852 298852
rect 381636 298732 381688 298784
rect 485688 298732 485740 298784
rect 454960 298052 455012 298104
rect 566464 298052 566516 298104
rect 382924 297984 382976 298036
rect 519360 297984 519412 298036
rect 370596 297916 370648 297968
rect 518072 297916 518124 297968
rect 369216 297848 369268 297900
rect 518256 297848 518308 297900
rect 361120 297780 361172 297832
rect 512184 297780 512236 297832
rect 363972 297712 364024 297764
rect 515312 297712 515364 297764
rect 366548 297644 366600 297696
rect 518348 297644 518400 297696
rect 365076 297576 365128 297628
rect 516876 297576 516928 297628
rect 362408 297508 362460 297560
rect 515588 297508 515640 297560
rect 366456 297440 366508 297492
rect 519728 297440 519780 297492
rect 362500 297372 362552 297424
rect 516232 297372 516284 297424
rect 454776 295944 454828 295996
rect 573364 295944 573416 295996
rect 435364 295332 435416 295384
rect 440884 295332 440936 295384
rect 469864 295332 469916 295384
rect 471244 295332 471296 295384
rect 374644 295264 374696 295316
rect 507584 295264 507636 295316
rect 379152 295196 379204 295248
rect 514208 295196 514260 295248
rect 372068 295128 372120 295180
rect 509792 295128 509844 295180
rect 371976 295060 372028 295112
rect 510712 295060 510764 295112
rect 375104 294992 375156 295044
rect 517612 294992 517664 295044
rect 375012 294924 375064 294976
rect 517704 294924 517756 294976
rect 377588 294856 377640 294908
rect 520556 294856 520608 294908
rect 373356 294788 373408 294840
rect 517980 294788 518032 294840
rect 372344 294720 372396 294772
rect 519176 294720 519228 294772
rect 371884 294652 371936 294704
rect 518992 294652 519044 294704
rect 369400 294584 369452 294636
rect 516692 294584 516744 294636
rect 374920 294516 374972 294568
rect 507676 294516 507728 294568
rect 376208 294448 376260 294500
rect 507768 294448 507820 294500
rect 455052 294380 455104 294432
rect 570604 294380 570656 294432
rect 361764 293904 361816 293956
rect 436836 293904 436888 293956
rect 476856 293224 476908 293276
rect 558184 293224 558236 293276
rect 3424 292544 3476 292596
rect 4896 292544 4948 292596
rect 383476 292476 383528 292528
rect 507492 292476 507544 292528
rect 386052 292408 386104 292460
rect 520280 292408 520332 292460
rect 380440 292340 380492 292392
rect 514760 292340 514812 292392
rect 381360 292272 381412 292324
rect 516968 292272 517020 292324
rect 377772 292204 377824 292256
rect 514116 292204 514168 292256
rect 383384 292136 383436 292188
rect 520372 292136 520424 292188
rect 380532 292068 380584 292120
rect 520464 292068 520516 292120
rect 369124 292000 369176 292052
rect 516784 292000 516836 292052
rect 366364 291932 366416 291984
rect 519268 291932 519320 291984
rect 363880 291864 363932 291916
rect 520740 291864 520792 291916
rect 361212 291796 361264 291848
rect 519452 291796 519504 291848
rect 385868 291728 385920 291780
rect 507400 291728 507452 291780
rect 456156 291660 456208 291712
rect 572076 291660 572128 291712
rect 454960 290504 455012 290556
rect 485872 290504 485924 290556
rect 476028 290436 476080 290488
rect 569224 290436 569276 290488
rect 374828 289756 374880 289808
rect 507124 289756 507176 289808
rect 383200 289688 383252 289740
rect 517796 289688 517848 289740
rect 385960 289620 386012 289672
rect 521844 289620 521896 289672
rect 380348 289552 380400 289604
rect 516600 289552 516652 289604
rect 382188 289484 382240 289536
rect 518900 289484 518952 289536
rect 377496 289416 377548 289468
rect 514944 289416 514996 289468
rect 377680 289348 377732 289400
rect 519084 289348 519136 289400
rect 380256 289280 380308 289332
rect 523316 289280 523368 289332
rect 379060 289212 379112 289264
rect 523224 289212 523276 289264
rect 376116 289144 376168 289196
rect 521752 289144 521804 289196
rect 372252 289076 372304 289128
rect 520648 289076 520700 289128
rect 383292 289008 383344 289060
rect 507216 289008 507268 289060
rect 384672 288940 384724 288992
rect 507308 288940 507360 288992
rect 450360 288872 450412 288924
rect 455144 288872 455196 288924
rect 455328 288872 455380 288924
rect 574744 288872 574796 288924
rect 502248 287716 502300 287768
rect 538956 287716 539008 287768
rect 451188 287648 451240 287700
rect 505008 287648 505060 287700
rect 452108 286628 452160 286680
rect 487896 286628 487948 286680
rect 378784 286560 378836 286612
rect 475200 286560 475252 286612
rect 486516 286560 486568 286612
rect 531320 286560 531372 286612
rect 464988 286492 465040 286544
rect 571984 286492 572036 286544
rect 372160 286424 372212 286476
rect 523040 286424 523092 286476
rect 369308 286356 369360 286408
rect 521660 286356 521712 286408
rect 366640 286288 366692 286340
rect 523132 286288 523184 286340
rect 455052 284996 455104 285048
rect 494520 284996 494572 285048
rect 449808 284928 449860 284980
rect 536840 284928 536892 284980
rect 453580 283636 453632 283688
rect 493968 283636 494020 283688
rect 501420 283636 501472 283688
rect 540244 283636 540296 283688
rect 477224 283568 477276 283620
rect 580264 283568 580316 283620
rect 361764 282820 361816 282872
rect 439688 282820 439740 282872
rect 459284 282140 459336 282192
rect 492312 282140 492364 282192
rect 432604 282072 432656 282124
rect 435364 282072 435416 282124
rect 452384 280848 452436 280900
rect 493140 280848 493192 280900
rect 500868 280848 500920 280900
rect 540152 280848 540204 280900
rect 458088 280780 458140 280832
rect 505284 280780 505336 280832
rect 453672 279420 453724 279472
rect 493692 279420 493744 279472
rect 471980 279012 472032 279064
rect 475384 279012 475436 279064
rect 457628 277992 457680 278044
rect 493416 277992 493468 278044
rect 499212 277992 499264 278044
rect 541440 277992 541492 278044
rect 467104 277380 467156 277432
rect 472624 277380 472676 277432
rect 466460 276836 466512 276888
rect 471980 276836 472032 276888
rect 456432 276700 456484 276752
rect 492036 276700 492088 276752
rect 375840 276632 375892 276684
rect 485412 276632 485464 276684
rect 497740 276632 497792 276684
rect 541348 276632 541400 276684
rect 453488 275340 453540 275392
rect 488172 275340 488224 275392
rect 500500 275340 500552 275392
rect 540336 275340 540388 275392
rect 454868 275272 454920 275324
rect 491208 275272 491260 275324
rect 497832 275272 497884 275324
rect 541256 275272 541308 275324
rect 429200 274592 429252 274644
rect 432604 274592 432656 274644
rect 459192 273980 459244 274032
rect 487344 273980 487396 274032
rect 498936 273980 498988 274032
rect 540060 273980 540112 274032
rect 456340 273912 456392 273964
rect 490932 273912 490984 273964
rect 497556 273912 497608 273964
rect 541164 273912 541216 273964
rect 462228 273232 462280 273284
rect 466460 273232 466512 273284
rect 454776 272552 454828 272604
rect 487620 272552 487672 272604
rect 498384 272552 498436 272604
rect 539968 272552 540020 272604
rect 456248 272484 456300 272536
rect 490380 272484 490432 272536
rect 496176 272484 496228 272536
rect 543004 272484 543056 272536
rect 361764 271804 361816 271856
rect 438124 271804 438176 271856
rect 452292 271192 452344 271244
rect 489828 271192 489880 271244
rect 495072 271192 495124 271244
rect 542820 271192 542872 271244
rect 466644 271124 466696 271176
rect 580356 271124 580408 271176
rect 456524 270920 456576 270972
rect 462228 270920 462280 270972
rect 465816 269832 465868 269884
rect 555424 269832 555476 269884
rect 450452 269764 450504 269816
rect 457812 269764 457864 269816
rect 466368 269764 466420 269816
rect 580264 269764 580316 269816
rect 427084 269016 427136 269068
rect 429200 269016 429252 269068
rect 449900 268540 449952 268592
rect 469864 268540 469916 268592
rect 442264 268472 442316 268524
rect 467104 268472 467156 268524
rect 486884 268472 486936 268524
rect 531228 268472 531280 268524
rect 456156 268404 456208 268456
rect 489276 268404 489328 268456
rect 495348 268404 495400 268456
rect 542912 268404 542964 268456
rect 450912 268336 450964 268388
rect 504732 268336 504784 268388
rect 443184 266976 443236 267028
rect 456524 266976 456576 267028
rect 449164 263508 449216 263560
rect 456800 263508 456852 263560
rect 438124 261808 438176 261860
rect 443184 261808 443236 261860
rect 361764 260788 361816 260840
rect 399484 260788 399536 260840
rect 447784 260788 447836 260840
rect 449808 260788 449860 260840
rect 431316 258680 431368 258732
rect 455236 258680 455288 258732
rect 3976 253920 4028 253972
rect 5080 253920 5132 253972
rect 421564 250452 421616 250504
rect 427084 250452 427136 250504
rect 361764 249704 361816 249756
rect 443736 249704 443788 249756
rect 447140 249704 447192 249756
rect 456800 249704 456852 249756
rect 446404 248888 446456 248940
rect 447140 248888 447192 248940
rect 443736 245624 443788 245676
rect 447784 245624 447836 245676
rect 572076 245556 572128 245608
rect 580172 245556 580224 245608
rect 425704 244264 425756 244316
rect 431316 244264 431368 244316
rect 3792 243924 3844 243976
rect 4988 243924 5040 243976
rect 418528 238960 418580 239012
rect 421564 238960 421616 239012
rect 361764 238688 361816 238740
rect 439596 238688 439648 238740
rect 406384 236648 406436 236700
rect 418528 236648 418580 236700
rect 558184 233180 558236 233232
rect 580172 233180 580224 233232
rect 422944 232908 422996 232960
rect 425704 232908 425756 232960
rect 361764 227672 361816 227724
rect 443644 227672 443696 227724
rect 439596 224068 439648 224120
rect 443736 224068 443788 224120
rect 3884 222096 3936 222148
rect 5172 222096 5224 222148
rect 455144 222096 455196 222148
rect 457812 222096 457864 222148
rect 439688 218016 439740 218068
rect 442264 218016 442316 218068
rect 361672 216316 361724 216368
rect 364064 216316 364116 216368
rect 432604 213868 432656 213920
rect 438124 213868 438176 213920
rect 423036 209040 423088 209092
rect 432604 209040 432656 209092
rect 457720 207884 457772 207936
rect 459560 207884 459612 207936
rect 576124 206932 576176 206984
rect 579804 206932 579856 206984
rect 361764 205572 361816 205624
rect 436744 205572 436796 205624
rect 460572 201084 460624 201136
rect 462412 201084 462464 201136
rect 460756 200676 460808 200728
rect 462320 200676 462372 200728
rect 459468 200132 459520 200184
rect 460940 200132 460992 200184
rect 448244 199384 448296 199436
rect 461584 199384 461636 199436
rect 404084 197344 404136 197396
rect 406384 197344 406436 197396
rect 438032 197344 438084 197396
rect 439596 197344 439648 197396
rect 429200 195236 429252 195288
rect 439688 195236 439740 195288
rect 361764 194488 361816 194540
rect 431224 194488 431276 194540
rect 417424 194284 417476 194336
rect 422944 194284 422996 194336
rect 547144 193128 547196 193180
rect 580172 193128 580224 193180
rect 418068 192448 418120 192500
rect 429200 192448 429252 192500
rect 419540 191836 419592 191888
rect 423036 191836 423088 191888
rect 436376 191496 436428 191548
rect 438032 191496 438084 191548
rect 394700 191088 394752 191140
rect 404084 191088 404136 191140
rect 395344 189728 395396 189780
rect 418068 189728 418120 189780
rect 433064 187688 433116 187740
rect 436376 187688 436428 187740
rect 414664 186328 414716 186380
rect 417424 186328 417476 186380
rect 391204 185376 391256 185428
rect 394700 185376 394752 185428
rect 413928 183608 413980 183660
rect 419540 183608 419592 183660
rect 361764 183472 361816 183524
rect 447600 183472 447652 183524
rect 448152 183472 448204 183524
rect 447600 182792 447652 182844
rect 528560 182792 528612 182844
rect 430580 182180 430632 182232
rect 433064 182180 433116 182232
rect 400588 181432 400640 181484
rect 413928 181432 413980 181484
rect 551284 179324 551336 179376
rect 580172 179324 580224 179376
rect 398104 176672 398156 176724
rect 400588 176672 400640 176724
rect 422944 176604 422996 176656
rect 430580 176672 430632 176724
rect 361764 172456 361816 172508
rect 447140 172456 447192 172508
rect 447140 171776 447192 171828
rect 448336 171776 448388 171828
rect 524420 171776 524472 171828
rect 391296 171096 391348 171148
rect 395344 171096 395396 171148
rect 420184 169736 420236 169788
rect 422944 169736 422996 169788
rect 533436 166948 533488 167000
rect 580172 166948 580224 167000
rect 388536 166268 388588 166320
rect 391204 166268 391256 166320
rect 388444 164840 388496 164892
rect 398104 164840 398156 164892
rect 448428 164160 448480 164212
rect 449348 164160 449400 164212
rect 438584 163616 438636 163668
rect 439504 163616 439556 163668
rect 445208 163616 445260 163668
rect 446404 163616 446456 163668
rect 407028 162868 407080 162920
rect 414664 162868 414716 162920
rect 456800 162256 456852 162308
rect 457812 162256 457864 162308
rect 485780 162256 485832 162308
rect 418712 162188 418764 162240
rect 457996 162188 458048 162240
rect 415124 162120 415176 162172
rect 456800 162120 456852 162172
rect 489920 162120 489972 162172
rect 375196 161508 375248 161560
rect 418712 161508 418764 161560
rect 445208 161508 445260 161560
rect 451004 161508 451056 161560
rect 412088 161440 412140 161492
rect 459560 161440 459612 161492
rect 460204 161440 460256 161492
rect 361764 161372 361816 161424
rect 448336 161372 448388 161424
rect 359464 160692 359516 160744
rect 388536 160692 388588 160744
rect 448336 160692 448388 160744
rect 521660 160692 521712 160744
rect 425336 160488 425388 160540
rect 425888 160488 425940 160540
rect 496820 160488 496872 160540
rect 428648 160420 428700 160472
rect 500960 160420 501012 160472
rect 421840 160352 421892 160404
rect 494060 160352 494112 160404
rect 435272 160284 435324 160336
rect 436008 160284 436060 160336
rect 509240 160284 509292 160336
rect 431776 160216 431828 160268
rect 505100 160216 505152 160268
rect 386144 160148 386196 160200
rect 415124 160148 415176 160200
rect 438584 160148 438636 160200
rect 513380 160148 513432 160200
rect 387800 160080 387852 160132
rect 391296 160080 391348 160132
rect 409512 160080 409564 160132
rect 441574 160080 441626 160132
rect 442908 160080 442960 160132
rect 517520 160080 517572 160132
rect 409880 159740 409932 159792
rect 420184 159740 420236 159792
rect 409144 159672 409196 159724
rect 428004 159672 428056 159724
rect 409236 159604 409288 159656
rect 431316 159604 431368 159656
rect 409328 159536 409380 159588
rect 434812 159536 434864 159588
rect 409420 159468 409472 159520
rect 437940 159468 437992 159520
rect 384212 159400 384264 159452
rect 421380 159400 421432 159452
rect 386236 159332 386288 159384
rect 425152 159332 425204 159384
rect 451740 158652 451792 158704
rect 454960 158652 455012 158704
rect 361580 157972 361632 158024
rect 387800 157972 387852 158024
rect 398840 157972 398892 158024
rect 409880 157972 409932 158024
rect 451740 157292 451792 157344
rect 455052 157292 455104 157344
rect 402244 155184 402296 155236
rect 407028 155184 407080 155236
rect 452476 154436 452528 154488
rect 453580 154436 453632 154488
rect 389272 153824 389324 153876
rect 398748 153824 398800 153876
rect 537484 153144 537536 153196
rect 580172 153144 580224 153196
rect 452476 152940 452528 152992
rect 453672 152940 453724 152992
rect 452568 151444 452620 151496
rect 457628 151444 457680 151496
rect 386512 150560 386564 150612
rect 389272 150560 389324 150612
rect 361764 150356 361816 150408
rect 409512 150356 409564 150408
rect 371240 149744 371292 149796
rect 386512 149744 386564 149796
rect 368296 149676 368348 149728
rect 388444 149676 388496 149728
rect 365720 147636 365772 147688
rect 371240 147636 371292 147688
rect 452568 147364 452620 147416
rect 459100 147364 459152 147416
rect 393964 146956 394016 147008
rect 402244 146956 402296 147008
rect 451832 146208 451884 146260
rect 459284 146208 459336 146260
rect 364340 144848 364392 144900
rect 368296 144848 368348 144900
rect 451556 144780 451608 144832
rect 456432 144780 456484 144832
rect 362960 143556 363012 143608
rect 365628 143556 365680 143608
rect 460204 143488 460256 143540
rect 460848 143488 460900 143540
rect 452568 143420 452620 143472
rect 457444 143420 457496 143472
rect 460848 142196 460900 142248
rect 481916 142196 481968 142248
rect 451004 142128 451056 142180
rect 533988 142128 534040 142180
rect 540428 142128 540480 142180
rect 452568 141924 452620 141976
rect 459008 141924 459060 141976
rect 452568 140700 452620 140752
rect 454868 140700 454920 140752
rect 359648 140020 359700 140072
rect 393964 140020 394016 140072
rect 533344 140020 533396 140072
rect 542544 140020 542596 140072
rect 359556 139544 359608 139596
rect 364340 139544 364392 139596
rect 361764 139340 361816 139392
rect 409420 139340 409472 139392
rect 555424 139340 555476 139392
rect 580172 139340 580224 139392
rect 451556 139204 451608 139256
rect 456340 139204 456392 139256
rect 452568 137844 452620 137896
rect 457536 137844 457588 137896
rect 538956 136552 539008 136604
rect 539508 136552 539560 136604
rect 451556 136484 451608 136536
rect 456248 136484 456300 136536
rect 452016 135124 452068 135176
rect 458916 135124 458968 135176
rect 452292 132404 452344 132456
rect 453396 132404 453448 132456
rect 361396 131112 361448 131164
rect 362592 131112 362644 131164
rect 452568 131044 452620 131096
rect 456156 131044 456208 131096
rect 452108 129684 452160 129736
rect 453304 129684 453356 129736
rect 361764 128256 361816 128308
rect 409328 128256 409380 128308
rect 452568 126896 452620 126948
rect 458824 126896 458876 126948
rect 574744 126896 574796 126948
rect 580172 126896 580224 126948
rect 451740 126760 451792 126812
rect 453488 126760 453540 126812
rect 451740 123088 451792 123140
rect 454776 123088 454828 123140
rect 451924 122000 451976 122052
rect 459192 122000 459244 122052
rect 384948 119348 385000 119400
rect 456064 119348 456116 119400
rect 361764 117240 361816 117292
rect 409236 117240 409288 117292
rect 569224 113092 569276 113144
rect 579804 113092 579856 113144
rect 402152 107584 402204 107636
rect 403624 107584 403676 107636
rect 439136 107244 439188 107296
rect 450820 107244 450872 107296
rect 432972 107176 433024 107228
rect 450544 107176 450596 107228
rect 426808 107108 426860 107160
rect 450728 107108 450780 107160
rect 420644 107040 420696 107092
rect 450636 107040 450688 107092
rect 414480 106972 414532 107024
rect 454684 106972 454736 107024
rect 389824 106904 389876 106956
rect 451004 106904 451056 106956
rect 445300 106496 445352 106548
rect 450912 106496 450964 106548
rect 361764 106224 361816 106276
rect 409144 106224 409196 106276
rect 559564 100648 559616 100700
rect 580172 100648 580224 100700
rect 3608 98608 3660 98660
rect 20904 98608 20956 98660
rect 361764 95140 361816 95192
rect 386236 95140 386288 95192
rect 570604 86912 570656 86964
rect 580172 86912 580224 86964
rect 3700 86232 3752 86284
rect 20904 86232 20956 86284
rect 361764 84124 361816 84176
rect 384212 84124 384264 84176
rect 361764 73108 361816 73160
rect 375196 73108 375248 73160
rect 544384 73108 544436 73160
rect 580172 73108 580224 73160
rect 5080 71680 5132 71732
rect 5540 71680 5592 71732
rect 3608 70388 3660 70440
rect 19984 70388 20036 70440
rect 5540 70320 5592 70372
rect 7564 70320 7616 70372
rect 361764 62024 361816 62076
rect 386144 62024 386196 62076
rect 7564 60732 7616 60784
rect 10048 60664 10100 60716
rect 548524 60664 548576 60716
rect 580172 60664 580224 60716
rect 4804 59304 4856 59356
rect 5816 59304 5868 59356
rect 3608 57944 3660 57996
rect 20076 57944 20128 57996
rect 5816 57196 5868 57248
rect 9772 57196 9824 57248
rect 4896 56516 4948 56568
rect 7288 56516 7340 56568
rect 10048 56516 10100 56568
rect 12348 56516 12400 56568
rect 9772 56108 9824 56160
rect 12808 56108 12860 56160
rect 5540 54476 5592 54528
rect 12256 54476 12308 54528
rect 7288 54068 7340 54120
rect 11980 54068 12032 54120
rect 12348 53388 12400 53440
rect 15200 53388 15252 53440
rect 11980 52436 12032 52488
rect 19248 52368 19300 52420
rect 361764 51076 361816 51128
rect 386144 51076 386196 51128
rect 540612 51076 540664 51128
rect 543740 51076 543792 51128
rect 4988 50328 5040 50380
rect 11704 50328 11756 50380
rect 12808 50328 12860 50380
rect 20628 50328 20680 50380
rect 15200 49716 15252 49768
rect 18972 49648 19024 49700
rect 18972 47812 19024 47864
rect 20904 47812 20956 47864
rect 3056 46996 3108 47048
rect 384764 46996 384816 47048
rect 3700 46860 3752 46912
rect 384580 46860 384632 46912
rect 573364 46860 573416 46912
rect 580172 46860 580224 46912
rect 3240 46792 3292 46844
rect 381912 46792 381964 46844
rect 3332 46724 3384 46776
rect 382004 46724 382056 46776
rect 3976 46656 4028 46708
rect 378968 46656 379020 46708
rect 3884 46588 3936 46640
rect 378876 46588 378928 46640
rect 3792 46520 3844 46572
rect 378600 46520 378652 46572
rect 3424 46452 3476 46504
rect 375932 46452 375984 46504
rect 19984 46384 20036 46436
rect 384396 46384 384448 46436
rect 20076 46316 20128 46368
rect 382096 46316 382148 46368
rect 21456 46248 21508 46300
rect 376668 46248 376720 46300
rect 21364 46180 21416 46232
rect 373632 46180 373684 46232
rect 12440 46112 12492 46164
rect 359464 46112 359516 46164
rect 20904 46044 20956 46096
rect 359648 46044 359700 46096
rect 4068 45500 4120 45552
rect 381820 45500 381872 45552
rect 3516 45432 3568 45484
rect 376024 45432 376076 45484
rect 3424 45364 3476 45416
rect 375840 45364 375892 45416
rect 20904 45296 20956 45348
rect 361396 45296 361448 45348
rect 65524 45228 65576 45280
rect 376300 45228 376352 45280
rect 62028 45160 62080 45212
rect 376392 45160 376444 45212
rect 58440 45092 58492 45144
rect 379244 45092 379296 45144
rect 54944 45024 54996 45076
rect 379428 45024 379480 45076
rect 51356 44956 51408 45008
rect 378692 44956 378744 45008
rect 47860 44888 47912 44940
rect 379336 44888 379388 44940
rect 7656 44820 7708 44872
rect 381452 44820 381504 44872
rect 69112 44752 69164 44804
rect 376484 44752 376536 44804
rect 72608 44684 72660 44736
rect 376576 44684 376628 44736
rect 76196 44616 76248 44668
rect 373724 44616 373776 44668
rect 111616 42712 111668 42764
rect 365260 42712 365312 42764
rect 108120 42644 108172 42696
rect 367928 42644 367980 42696
rect 104532 42576 104584 42628
rect 368020 42576 368072 42628
rect 101036 42508 101088 42560
rect 367836 42508 367888 42560
rect 97448 42440 97500 42492
rect 368112 42440 368164 42492
rect 93952 42372 94004 42424
rect 370964 42372 371016 42424
rect 90364 42304 90416 42356
rect 370872 42304 370924 42356
rect 86868 42236 86920 42288
rect 370780 42236 370832 42288
rect 83280 42168 83332 42220
rect 370688 42168 370740 42220
rect 79692 42100 79744 42152
rect 373448 42100 373500 42152
rect 12348 42032 12400 42084
rect 373540 42032 373592 42084
rect 115204 41964 115256 42016
rect 365352 41964 365404 42016
rect 461584 41352 461636 41404
rect 536840 41352 536892 41404
rect 118792 39992 118844 40044
rect 362500 39992 362552 40044
rect 63224 39924 63276 39976
rect 372344 39924 372396 39976
rect 59636 39856 59688 39908
rect 369400 39856 369452 39908
rect 56048 39788 56100 39840
rect 370596 39788 370648 39840
rect 52552 39720 52604 39772
rect 369216 39720 369268 39772
rect 48964 39652 49016 39704
rect 366548 39652 366600 39704
rect 40684 39584 40736 39636
rect 366456 39584 366508 39636
rect 37188 39516 37240 39568
rect 363972 39516 364024 39568
rect 33600 39448 33652 39500
rect 362408 39448 362460 39500
rect 26516 39380 26568 39432
rect 365168 39380 365220 39432
rect 4068 39312 4120 39364
rect 368204 39312 368256 39364
rect 122288 39244 122340 39296
rect 362316 39244 362368 39296
rect 102232 37204 102284 37256
rect 377772 37204 377824 37256
rect 98644 37136 98696 37188
rect 379152 37136 379204 37188
rect 95148 37068 95200 37120
rect 377588 37068 377640 37120
rect 91560 37000 91612 37052
rect 375104 37000 375156 37052
rect 87972 36932 88024 36984
rect 375012 36932 375064 36984
rect 84476 36864 84528 36916
rect 376208 36864 376260 36916
rect 80888 36796 80940 36848
rect 374920 36796 374972 36848
rect 77392 36728 77444 36780
rect 372068 36728 372120 36780
rect 73804 36660 73856 36712
rect 373356 36660 373408 36712
rect 70308 36592 70360 36644
rect 371976 36592 372028 36644
rect 66720 36524 66772 36576
rect 371884 36524 371936 36576
rect 105728 36456 105780 36508
rect 380532 36456 380584 36508
rect 119896 34416 119948 34468
rect 386052 34416 386104 34468
rect 116400 34348 116452 34400
rect 383384 34348 383436 34400
rect 112812 34280 112864 34332
rect 380440 34280 380492 34332
rect 109316 34212 109368 34264
rect 381360 34212 381412 34264
rect 45468 34144 45520 34196
rect 372252 34144 372304 34196
rect 41880 34076 41932 34128
rect 369124 34076 369176 34128
rect 50160 34008 50212 34060
rect 377680 34008 377732 34060
rect 34796 33940 34848 33992
rect 363880 33940 363932 33992
rect 31300 33872 31352 33924
rect 361212 33872 361264 33924
rect 23020 33804 23072 33856
rect 384856 33804 384908 33856
rect 18236 33736 18288 33788
rect 383476 33736 383528 33788
rect 123484 33668 123536 33720
rect 385684 33668 385736 33720
rect 2872 33056 2924 33108
rect 383108 33056 383160 33108
rect 562324 33056 562376 33108
rect 580172 33056 580224 33108
rect 99840 31696 99892 31748
rect 366640 31696 366692 31748
rect 386144 31696 386196 31748
rect 460204 31696 460256 31748
rect 96252 31628 96304 31680
rect 376116 31628 376168 31680
rect 92756 31560 92808 31612
rect 379060 31560 379112 31612
rect 85672 31492 85724 31544
rect 382188 31492 382240 31544
rect 78588 31424 78640 31476
rect 385960 31424 386012 31476
rect 71504 31356 71556 31408
rect 383200 31356 383252 31408
rect 67916 31288 67968 31340
rect 380256 31288 380308 31340
rect 64328 31220 64380 31272
rect 377496 31220 377548 31272
rect 60832 31152 60884 31204
rect 383292 31152 383344 31204
rect 57244 31084 57296 31136
rect 380348 31084 380400 31136
rect 14740 31016 14792 31068
rect 384672 31016 384724 31068
rect 106924 30948 106976 31000
rect 369308 30948 369360 31000
rect 124680 28908 124732 28960
rect 380164 28908 380216 28960
rect 117596 28840 117648 28892
rect 373264 28840 373316 28892
rect 121092 28772 121144 28824
rect 377404 28772 377456 28824
rect 114008 28704 114060 28756
rect 372160 28704 372212 28756
rect 109684 28636 109736 28688
rect 384948 28636 385000 28688
rect 28908 28568 28960 28620
rect 383016 28568 383068 28620
rect 19432 28500 19484 28552
rect 374736 28500 374788 28552
rect 43076 28432 43128 28484
rect 462320 28432 462372 28484
rect 35992 28364 36044 28416
rect 461032 28364 461084 28416
rect 32404 28296 32456 28348
rect 462412 28296 462464 28348
rect 5264 28228 5316 28280
rect 460940 28228 460992 28280
rect 3424 20612 3476 20664
rect 378784 20612 378836 20664
rect 571984 20612 572036 20664
rect 579988 20612 580040 20664
rect 3424 6808 3476 6860
rect 381636 6808 381688 6860
rect 566464 6808 566516 6860
rect 580172 6808 580224 6860
rect 82084 4088 82136 4140
rect 370504 4088 370556 4140
rect 75000 4020 75052 4072
rect 367744 4020 367796 4072
rect 53748 3952 53800 4004
rect 364984 3952 365036 4004
rect 46664 3884 46716 3936
rect 363696 3884 363748 3936
rect 39580 3816 39632 3868
rect 360936 3816 360988 3868
rect 38384 3748 38436 3800
rect 366364 3748 366416 3800
rect 30104 3680 30156 3732
rect 363604 3680 363656 3732
rect 44272 3612 44324 3664
rect 382924 3612 382976 3664
rect 21824 3544 21876 3596
rect 363788 3544 363840 3596
rect 27712 3476 27764 3528
rect 385868 3476 385920 3528
rect 24216 3408 24268 3460
rect 385776 3408 385828 3460
rect 89168 3340 89220 3392
rect 361120 3340 361172 3392
rect 103336 3272 103388 3324
rect 361028 3272 361080 3324
rect 6460 3204 6512 3256
rect 109684 3204 109736 3256
rect 110512 3204 110564 3256
rect 360844 3204 360896 3256
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 8128 700330 8156 703520
rect 8116 700324 8168 700330
rect 8116 700266 8168 700272
rect 24320 686497 24348 703520
rect 40512 700369 40540 703520
rect 40498 700360 40554 700369
rect 40498 700295 40554 700304
rect 24306 686488 24362 686497
rect 24306 686423 24362 686432
rect 72988 685166 73016 703520
rect 89180 685234 89208 703520
rect 105464 700398 105492 703520
rect 105452 700392 105504 700398
rect 105452 700334 105504 700340
rect 137848 685302 137876 703520
rect 154132 700466 154160 703520
rect 170324 700534 170352 703520
rect 170312 700528 170364 700534
rect 202800 700505 202828 703520
rect 170312 700470 170364 700476
rect 202786 700496 202842 700505
rect 154120 700460 154172 700466
rect 202786 700431 202842 700440
rect 154120 700402 154172 700408
rect 218992 692102 219020 703520
rect 235184 700602 235212 703520
rect 267660 700670 267688 703520
rect 267648 700664 267700 700670
rect 267648 700606 267700 700612
rect 235172 700596 235224 700602
rect 235172 700538 235224 700544
rect 218980 692096 219032 692102
rect 218980 692038 219032 692044
rect 283852 687954 283880 703520
rect 300136 689353 300164 703520
rect 332520 700738 332548 703520
rect 332508 700732 332560 700738
rect 332508 700674 332560 700680
rect 300122 689344 300178 689353
rect 300122 689279 300178 689288
rect 283840 687948 283892 687954
rect 283840 687890 283892 687896
rect 348804 686526 348832 703520
rect 364996 700806 365024 703520
rect 397472 700874 397500 703520
rect 397460 700868 397512 700874
rect 397460 700810 397512 700816
rect 364984 700800 365036 700806
rect 364984 700742 365036 700748
rect 348792 686520 348844 686526
rect 348792 686462 348844 686468
rect 137836 685296 137888 685302
rect 137836 685238 137888 685244
rect 89168 685228 89220 685234
rect 89168 685170 89220 685176
rect 72976 685160 73028 685166
rect 72976 685102 73028 685108
rect 3884 684548 3936 684554
rect 3884 684490 3936 684496
rect 3238 684312 3294 684321
rect 3238 684247 3294 684256
rect 3252 683194 3280 684247
rect 3516 683664 3568 683670
rect 3516 683606 3568 683612
rect 3332 683596 3384 683602
rect 3332 683538 3384 683544
rect 3240 683188 3292 683194
rect 3240 683130 3292 683136
rect 3240 682712 3292 682718
rect 3240 682654 3292 682660
rect 3148 658232 3200 658238
rect 3146 658200 3148 658209
rect 3200 658200 3202 658209
rect 3146 658135 3202 658144
rect 3252 580009 3280 682654
rect 3238 580000 3294 580009
rect 3238 579935 3294 579944
rect 3344 566953 3372 683538
rect 3424 683460 3476 683466
rect 3424 683402 3476 683408
rect 3330 566944 3386 566953
rect 3330 566879 3386 566888
rect 3436 449585 3464 683402
rect 3528 462641 3556 683606
rect 3700 683528 3752 683534
rect 3700 683470 3752 683476
rect 3608 683392 3660 683398
rect 3608 683334 3660 683340
rect 3620 475697 3648 683334
rect 3712 632097 3740 683470
rect 3792 683324 3844 683330
rect 3792 683266 3844 683272
rect 3698 632088 3754 632097
rect 3698 632023 3754 632032
rect 3700 631372 3752 631378
rect 3700 631314 3752 631320
rect 3606 475688 3662 475697
rect 3606 475623 3662 475632
rect 3514 462632 3570 462641
rect 3514 462567 3570 462576
rect 3422 449576 3478 449585
rect 3422 449511 3478 449520
rect 3712 423609 3740 631314
rect 3804 501809 3832 683266
rect 3896 514865 3924 684490
rect 24124 683936 24176 683942
rect 24124 683878 24176 683884
rect 359464 683936 359516 683942
rect 359464 683878 359516 683884
rect 19984 683868 20036 683874
rect 19984 683810 20036 683816
rect 4068 683732 4120 683738
rect 4068 683674 4120 683680
rect 3976 683256 4028 683262
rect 3976 683198 4028 683204
rect 4080 683210 4108 683674
rect 3988 527921 4016 683198
rect 4080 683182 4200 683210
rect 4172 683074 4200 683182
rect 4080 683046 4200 683074
rect 4080 553897 4108 683046
rect 19248 682780 19300 682786
rect 19248 682722 19300 682728
rect 19260 680406 19288 682722
rect 17224 680400 17276 680406
rect 17224 680342 17276 680348
rect 19248 680400 19300 680406
rect 19248 680342 19300 680348
rect 17236 661094 17264 680342
rect 17224 661088 17276 661094
rect 17224 661030 17276 661036
rect 14188 661020 14240 661026
rect 14188 660962 14240 660968
rect 14200 656674 14228 660962
rect 19996 658238 20024 683810
rect 21364 683800 21416 683806
rect 21364 683742 21416 683748
rect 19984 658232 20036 658238
rect 19984 658174 20036 658180
rect 11704 656668 11756 656674
rect 11704 656610 11756 656616
rect 14188 656668 14240 656674
rect 14188 656610 14240 656616
rect 11716 645862 11744 656610
rect 10600 645856 10652 645862
rect 10600 645798 10652 645804
rect 11704 645856 11756 645862
rect 11704 645798 11756 645804
rect 10612 643754 10640 645798
rect 5540 643748 5592 643754
rect 5540 643690 5592 643696
rect 10600 643748 10652 643754
rect 10600 643690 10652 643696
rect 5552 640354 5580 643690
rect 4804 640348 4856 640354
rect 4804 640290 4856 640296
rect 5540 640348 5592 640354
rect 5540 640290 5592 640296
rect 4066 553888 4122 553897
rect 4066 553823 4122 553832
rect 3974 527912 4030 527921
rect 3974 527847 4030 527856
rect 3882 514856 3938 514865
rect 4816 514826 4844 640290
rect 21376 634814 21404 683742
rect 24136 682786 24164 683878
rect 24124 682780 24176 682786
rect 24124 682722 24176 682728
rect 20916 634786 21404 634814
rect 20916 631378 20944 634786
rect 20904 631372 20956 631378
rect 20904 631314 20956 631320
rect 359476 561678 359504 683878
rect 361764 679040 361816 679046
rect 361762 679008 361764 679017
rect 387064 679040 387116 679046
rect 361816 679008 361818 679017
rect 387064 678982 387116 678988
rect 361762 678943 361818 678952
rect 361762 667992 361818 668001
rect 361762 667927 361764 667936
rect 361816 667927 361818 667936
rect 382924 667956 382976 667962
rect 361764 667898 361816 667904
rect 382924 667898 382976 667904
rect 361762 656976 361818 656985
rect 361762 656911 361764 656920
rect 361816 656911 361818 656920
rect 381544 656940 381596 656946
rect 361764 656882 361816 656888
rect 381544 656882 381596 656888
rect 361762 645960 361818 645969
rect 361762 645895 361764 645904
rect 361816 645895 361818 645904
rect 378784 645924 378836 645930
rect 361764 645866 361816 645872
rect 378784 645866 378836 645872
rect 361578 634944 361634 634953
rect 361578 634879 361634 634888
rect 361592 634846 361620 634879
rect 361580 634840 361632 634846
rect 361580 634782 361632 634788
rect 361578 623928 361634 623937
rect 361578 623863 361634 623872
rect 361592 623830 361620 623863
rect 361580 623824 361632 623830
rect 361580 623766 361632 623772
rect 376024 623824 376076 623830
rect 376024 623766 376076 623772
rect 361578 612912 361634 612921
rect 361578 612847 361634 612856
rect 361592 612814 361620 612847
rect 361580 612808 361632 612814
rect 361580 612750 361632 612756
rect 361762 601896 361818 601905
rect 361762 601831 361818 601840
rect 361776 601730 361804 601831
rect 361764 601724 361816 601730
rect 361764 601666 361816 601672
rect 374644 601724 374696 601730
rect 374644 601666 374696 601672
rect 361762 590880 361818 590889
rect 361762 590815 361818 590824
rect 361776 590714 361804 590815
rect 361764 590708 361816 590714
rect 361764 590650 361816 590656
rect 361762 579864 361818 579873
rect 361762 579799 361818 579808
rect 361776 579698 361804 579799
rect 361764 579692 361816 579698
rect 361764 579634 361816 579640
rect 371884 579692 371936 579698
rect 371884 579634 371936 579640
rect 361578 568848 361634 568857
rect 361578 568783 361580 568792
rect 361632 568783 361634 568792
rect 363604 568812 363656 568818
rect 361580 568754 361632 568760
rect 363604 568754 363656 568760
rect 359464 561672 359516 561678
rect 359464 561614 359516 561620
rect 362224 561672 362276 561678
rect 362224 561614 362276 561620
rect 361670 557832 361726 557841
rect 361670 557767 361726 557776
rect 361684 557598 361712 557767
rect 361672 557592 361724 557598
rect 361672 557534 361724 557540
rect 362236 551342 362264 561614
rect 362224 551336 362276 551342
rect 362224 551278 362276 551284
rect 361762 546816 361818 546825
rect 361762 546751 361818 546760
rect 361776 546514 361804 546751
rect 361764 546508 361816 546514
rect 361764 546450 361816 546456
rect 361578 535800 361634 535809
rect 361578 535735 361634 535744
rect 361592 535498 361620 535735
rect 361580 535492 361632 535498
rect 361580 535434 361632 535440
rect 361578 524784 361634 524793
rect 361578 524719 361580 524728
rect 361632 524719 361634 524728
rect 361580 524690 361632 524696
rect 3882 514791 3938 514800
rect 3976 514820 4028 514826
rect 3976 514762 4028 514768
rect 4804 514820 4856 514826
rect 4804 514762 4856 514768
rect 3790 501800 3846 501809
rect 3790 501735 3846 501744
rect 3698 423600 3754 423609
rect 3698 423535 3754 423544
rect 3988 410553 4016 514762
rect 361762 513768 361818 513777
rect 361762 513703 361818 513712
rect 361776 513398 361804 513703
rect 361764 513392 361816 513398
rect 361764 513334 361816 513340
rect 361762 502752 361818 502761
rect 361762 502687 361818 502696
rect 361776 502382 361804 502687
rect 361764 502376 361816 502382
rect 361764 502318 361816 502324
rect 361762 491736 361818 491745
rect 361762 491671 361818 491680
rect 361776 491366 361804 491671
rect 361764 491360 361816 491366
rect 361764 491302 361816 491308
rect 361762 480720 361818 480729
rect 361762 480655 361818 480664
rect 361776 480282 361804 480655
rect 361764 480276 361816 480282
rect 361764 480218 361816 480224
rect 361762 469704 361818 469713
rect 361762 469639 361818 469648
rect 361776 469266 361804 469639
rect 361764 469260 361816 469266
rect 361764 469202 361816 469208
rect 361762 458688 361818 458697
rect 361762 458623 361818 458632
rect 361776 458250 361804 458623
rect 361764 458244 361816 458250
rect 361764 458186 361816 458192
rect 362222 447672 362278 447681
rect 362222 447607 362278 447616
rect 361762 436656 361818 436665
rect 361762 436591 361818 436600
rect 361776 436150 361804 436591
rect 361764 436144 361816 436150
rect 361764 436086 361816 436092
rect 362236 416090 362264 447607
rect 362314 425640 362370 425649
rect 362314 425575 362370 425584
rect 362328 418810 362356 425575
rect 362316 418804 362368 418810
rect 362316 418746 362368 418752
rect 362224 416084 362276 416090
rect 362224 416026 362276 416032
rect 361578 414624 361634 414633
rect 361578 414559 361634 414568
rect 361592 414050 361620 414559
rect 361580 414044 361632 414050
rect 361580 413986 361632 413992
rect 3974 410544 4030 410553
rect 3974 410479 4030 410488
rect 361578 403608 361634 403617
rect 361578 403543 361634 403552
rect 361592 403034 361620 403543
rect 361580 403028 361632 403034
rect 361580 402970 361632 402976
rect 3790 397488 3846 397497
rect 3790 397423 3846 397432
rect 3514 358456 3570 358465
rect 3514 358391 3570 358400
rect 3422 345400 3478 345409
rect 3422 345335 3478 345344
rect 3436 292602 3464 345335
rect 3528 307766 3556 358391
rect 3516 307760 3568 307766
rect 3516 307702 3568 307708
rect 3606 306232 3662 306241
rect 3606 306167 3662 306176
rect 3424 292596 3476 292602
rect 3424 292538 3476 292544
rect 3422 267200 3478 267209
rect 3422 267135 3478 267144
rect 3330 162888 3386 162897
rect 3330 162823 3386 162832
rect 3238 149832 3294 149841
rect 3238 149767 3294 149776
rect 3054 98696 3110 98705
rect 3054 98631 3110 98640
rect 3068 47054 3096 98631
rect 3056 47048 3108 47054
rect 3056 46990 3108 46996
rect 3252 46850 3280 149767
rect 3240 46844 3292 46850
rect 3240 46786 3292 46792
rect 3344 46782 3372 162823
rect 3332 46776 3384 46782
rect 3332 46718 3384 46724
rect 3436 46510 3464 267135
rect 3514 254144 3570 254153
rect 3514 254079 3570 254088
rect 3424 46504 3476 46510
rect 3424 46446 3476 46452
rect 3422 45520 3478 45529
rect 3528 45490 3556 254079
rect 3620 98666 3648 306167
rect 3698 293176 3754 293185
rect 3698 293111 3754 293120
rect 3608 98660 3660 98666
rect 3608 98602 3660 98608
rect 3712 86290 3740 293111
rect 3804 243982 3832 397423
rect 361578 392592 361634 392601
rect 361578 392527 361634 392536
rect 361592 392018 361620 392527
rect 361580 392012 361632 392018
rect 361580 391954 361632 391960
rect 361578 381576 361634 381585
rect 361578 381511 361634 381520
rect 361592 380934 361620 381511
rect 361580 380928 361632 380934
rect 361580 380870 361632 380876
rect 363616 378146 363644 568754
rect 370504 557592 370556 557598
rect 370504 557534 370556 557540
rect 369124 551336 369176 551342
rect 369124 551278 369176 551284
rect 367744 546508 367796 546514
rect 367744 546450 367796 546456
rect 363696 535492 363748 535498
rect 363696 535434 363748 535440
rect 363604 378140 363656 378146
rect 363604 378082 363656 378088
rect 363708 375358 363736 535434
rect 363788 524748 363840 524754
rect 363788 524690 363840 524696
rect 363696 375352 363748 375358
rect 363696 375294 363748 375300
rect 363800 375290 363828 524690
rect 367756 376718 367784 546450
rect 369136 522306 369164 551278
rect 369124 522300 369176 522306
rect 369124 522242 369176 522248
rect 367744 376712 367796 376718
rect 367744 376654 367796 376660
rect 370516 376650 370544 557534
rect 371896 378078 371924 579634
rect 373264 386436 373316 386442
rect 373264 386378 373316 386384
rect 371884 378072 371936 378078
rect 371884 378014 371936 378020
rect 370504 376644 370556 376650
rect 370504 376586 370556 376592
rect 363788 375284 363840 375290
rect 363788 375226 363840 375232
rect 3882 371376 3938 371385
rect 3882 371311 3938 371320
rect 3792 243976 3844 243982
rect 3792 243918 3844 243924
rect 3790 241088 3846 241097
rect 3790 241023 3846 241032
rect 3700 86284 3752 86290
rect 3700 86226 3752 86232
rect 3698 84688 3754 84697
rect 3698 84623 3754 84632
rect 3606 71632 3662 71641
rect 3606 71567 3662 71576
rect 3620 70446 3648 71567
rect 3608 70440 3660 70446
rect 3608 70382 3660 70388
rect 3606 58576 3662 58585
rect 3606 58511 3662 58520
rect 3620 58002 3648 58511
rect 3608 57996 3660 58002
rect 3608 57938 3660 57944
rect 3712 46918 3740 84623
rect 3700 46912 3752 46918
rect 3700 46854 3752 46860
rect 3804 46578 3832 241023
rect 3896 222154 3924 371311
rect 361578 370560 361634 370569
rect 361578 370495 361634 370504
rect 361592 369918 361620 370495
rect 361580 369912 361632 369918
rect 361580 369854 361632 369860
rect 362222 359544 362278 359553
rect 362222 359479 362278 359488
rect 361762 348528 361818 348537
rect 361762 348463 361818 348472
rect 361776 347818 361804 348463
rect 361764 347812 361816 347818
rect 361764 347754 361816 347760
rect 362236 347750 362264 359479
rect 362224 347744 362276 347750
rect 362224 347686 362276 347692
rect 361764 340944 361816 340950
rect 361764 340886 361816 340892
rect 361776 337521 361804 340886
rect 361762 337512 361818 337521
rect 361762 337447 361818 337456
rect 362224 336048 362276 336054
rect 362224 335990 362276 335996
rect 362236 326505 362264 335990
rect 364064 334008 364116 334014
rect 364064 333950 364116 333956
rect 362222 326496 362278 326505
rect 362222 326431 362278 326440
rect 3974 319288 4030 319297
rect 3974 319223 4030 319232
rect 3988 253978 4016 319223
rect 361764 315988 361816 315994
rect 361764 315930 361816 315936
rect 361776 315489 361804 315930
rect 361762 315480 361818 315489
rect 361762 315415 361818 315424
rect 4804 307760 4856 307766
rect 4804 307702 4856 307708
rect 3976 253972 4028 253978
rect 3976 253914 4028 253920
rect 3884 222148 3936 222154
rect 3884 222090 3936 222096
rect 3882 214976 3938 214985
rect 3882 214911 3938 214920
rect 3896 46646 3924 214911
rect 3974 201920 4030 201929
rect 3974 201855 4030 201864
rect 3988 46714 4016 201855
rect 4066 188864 4122 188873
rect 4066 188799 4122 188808
rect 3976 46708 4028 46714
rect 3976 46650 4028 46656
rect 3884 46640 3936 46646
rect 3884 46582 3936 46588
rect 3792 46572 3844 46578
rect 3792 46514 3844 46520
rect 4080 45558 4108 188799
rect 4816 59362 4844 307702
rect 360842 305688 360898 305697
rect 360842 305623 360898 305632
rect 362316 305652 362368 305658
rect 4896 292596 4948 292602
rect 4896 292538 4948 292544
rect 4804 59356 4856 59362
rect 4804 59298 4856 59304
rect 4908 56574 4936 292538
rect 5080 253972 5132 253978
rect 5080 253914 5132 253920
rect 4988 243976 5040 243982
rect 4988 243918 5040 243924
rect 4896 56568 4948 56574
rect 4896 56510 4948 56516
rect 5000 50386 5028 243918
rect 5092 71738 5120 253914
rect 5172 222148 5224 222154
rect 5172 222090 5224 222096
rect 5080 71732 5132 71738
rect 5080 71674 5132 71680
rect 5184 55214 5212 222090
rect 359464 160744 359516 160750
rect 359464 160686 359516 160692
rect 20904 98660 20956 98666
rect 20904 98602 20956 98608
rect 20916 93854 20944 98602
rect 20916 93826 21404 93854
rect 20904 86284 20956 86290
rect 20904 86226 20956 86232
rect 20916 73681 20944 86226
rect 21376 77294 21404 93826
rect 21284 77266 21404 77294
rect 20902 73672 20958 73681
rect 20902 73607 20958 73616
rect 5540 71732 5592 71738
rect 5540 71674 5592 71680
rect 5552 70378 5580 71674
rect 19984 70440 20036 70446
rect 19984 70382 20036 70388
rect 5540 70372 5592 70378
rect 5540 70314 5592 70320
rect 7564 70372 7616 70378
rect 7564 70314 7616 70320
rect 7576 60790 7604 70314
rect 7564 60784 7616 60790
rect 7564 60726 7616 60732
rect 10048 60716 10100 60722
rect 10048 60658 10100 60664
rect 5816 59356 5868 59362
rect 5816 59298 5868 59304
rect 5828 57254 5856 59298
rect 5816 57248 5868 57254
rect 5816 57190 5868 57196
rect 9772 57248 9824 57254
rect 9772 57190 9824 57196
rect 7288 56568 7340 56574
rect 7288 56510 7340 56516
rect 5184 55186 5580 55214
rect 5552 54534 5580 55186
rect 5540 54528 5592 54534
rect 5540 54470 5592 54476
rect 7300 54126 7328 56510
rect 9784 56166 9812 57190
rect 10060 56574 10088 60658
rect 10048 56568 10100 56574
rect 10048 56510 10100 56516
rect 12348 56568 12400 56574
rect 12348 56510 12400 56516
rect 9772 56160 9824 56166
rect 9772 56102 9824 56108
rect 12256 54528 12308 54534
rect 12256 54470 12308 54476
rect 7288 54120 7340 54126
rect 7288 54062 7340 54068
rect 11980 54120 12032 54126
rect 11980 54062 12032 54068
rect 11992 52494 12020 54062
rect 11980 52488 12032 52494
rect 11980 52430 12032 52436
rect 12268 52442 12296 54470
rect 12360 53446 12388 56510
rect 12808 56160 12860 56166
rect 12808 56102 12860 56108
rect 12348 53440 12400 53446
rect 12348 53382 12400 53388
rect 12268 52414 12480 52442
rect 4988 50380 5040 50386
rect 4988 50322 5040 50328
rect 11704 50380 11756 50386
rect 11704 50322 11756 50328
rect 11716 48929 11744 50322
rect 11702 48920 11758 48929
rect 11702 48855 11758 48864
rect 12452 46170 12480 52414
rect 12820 50386 12848 56102
rect 15200 53440 15252 53446
rect 15200 53382 15252 53388
rect 12808 50380 12860 50386
rect 12808 50322 12860 50328
rect 15212 49774 15240 53382
rect 19248 52420 19300 52426
rect 19248 52362 19300 52368
rect 15200 49768 15252 49774
rect 15200 49710 15252 49716
rect 18972 49700 19024 49706
rect 18972 49642 19024 49648
rect 18984 47870 19012 49642
rect 19260 49609 19288 52362
rect 19246 49600 19302 49609
rect 19246 49535 19302 49544
rect 18972 47864 19024 47870
rect 18972 47806 19024 47812
rect 19996 46442 20024 70382
rect 21284 67634 21312 77266
rect 21454 73672 21510 73681
rect 21454 73607 21510 73616
rect 21284 67606 21404 67634
rect 20076 57996 20128 58002
rect 20076 57938 20128 57944
rect 19984 46436 20036 46442
rect 19984 46378 20036 46384
rect 20088 46374 20116 57938
rect 20628 50380 20680 50386
rect 20628 50322 20680 50328
rect 20640 48226 20668 50322
rect 20640 48198 20760 48226
rect 20076 46368 20128 46374
rect 20076 46310 20128 46316
rect 12440 46164 12492 46170
rect 12440 46106 12492 46112
rect 4068 45552 4120 45558
rect 20732 45554 20760 48198
rect 20904 47864 20956 47870
rect 20904 47806 20956 47812
rect 20916 46102 20944 47806
rect 21376 46238 21404 67606
rect 21468 46306 21496 73607
rect 21456 46300 21508 46306
rect 21456 46242 21508 46248
rect 21364 46232 21416 46238
rect 21364 46174 21416 46180
rect 359476 46170 359504 160686
rect 359648 140072 359700 140078
rect 359648 140014 359700 140020
rect 359556 139596 359608 139602
rect 359556 139538 359608 139544
rect 359568 46481 359596 139538
rect 359554 46472 359610 46481
rect 359554 46407 359610 46416
rect 359464 46164 359516 46170
rect 359464 46106 359516 46112
rect 359660 46102 359688 140014
rect 20904 46096 20956 46102
rect 20904 46038 20956 46044
rect 359648 46096 359700 46102
rect 359648 46038 359700 46044
rect 20732 45526 20944 45554
rect 4068 45494 4120 45500
rect 3422 45455 3478 45464
rect 3516 45484 3568 45490
rect 3436 45422 3464 45455
rect 3516 45426 3568 45432
rect 3424 45416 3476 45422
rect 3424 45358 3476 45364
rect 20916 45354 20944 45526
rect 20904 45348 20956 45354
rect 20904 45290 20956 45296
rect 65524 45280 65576 45286
rect 65524 45222 65576 45228
rect 62028 45212 62080 45218
rect 62028 45154 62080 45160
rect 58440 45144 58492 45150
rect 58440 45086 58492 45092
rect 54944 45076 54996 45082
rect 54944 45018 54996 45024
rect 51356 45008 51408 45014
rect 51356 44950 51408 44956
rect 47860 44940 47912 44946
rect 47860 44882 47912 44888
rect 7656 44872 7708 44878
rect 7656 44814 7708 44820
rect 4068 39364 4120 39370
rect 4068 39306 4120 39312
rect 2872 33108 2924 33114
rect 2872 33050 2924 33056
rect 2884 32473 2912 33050
rect 2870 32464 2926 32473
rect 2870 32399 2926 32408
rect 3424 20664 3476 20670
rect 3424 20606 3476 20612
rect 3436 19417 3464 20606
rect 3422 19408 3478 19417
rect 3422 19343 3478 19352
rect 3424 6860 3476 6866
rect 3424 6802 3476 6808
rect 3436 6497 3464 6802
rect 3422 6488 3478 6497
rect 3422 6423 3478 6432
rect 2870 3632 2926 3641
rect 2870 3567 2926 3576
rect 1674 3496 1730 3505
rect 1674 3431 1730 3440
rect 570 3360 626 3369
rect 570 3295 626 3304
rect 584 480 612 3295
rect 1688 480 1716 3431
rect 2884 480 2912 3567
rect 4080 480 4108 39306
rect 5264 28280 5316 28286
rect 5264 28222 5316 28228
rect 5276 480 5304 28222
rect 6460 3256 6512 3262
rect 6460 3198 6512 3204
rect 6472 480 6500 3198
rect 7668 480 7696 44814
rect 12348 42084 12400 42090
rect 12348 42026 12400 42032
rect 8758 4040 8814 4049
rect 8758 3975 8814 3984
rect 8772 480 8800 3975
rect 9954 3768 10010 3777
rect 9954 3703 10010 3712
rect 9968 480 9996 3703
rect 12360 480 12388 42026
rect 40684 39636 40736 39642
rect 40684 39578 40736 39584
rect 37188 39568 37240 39574
rect 37188 39510 37240 39516
rect 33600 39500 33652 39506
rect 33600 39442 33652 39448
rect 26516 39432 26568 39438
rect 26516 39374 26568 39380
rect 23020 33856 23072 33862
rect 23020 33798 23072 33804
rect 18236 33788 18288 33794
rect 18236 33730 18288 33736
rect 14740 31068 14792 31074
rect 14740 31010 14792 31016
rect 13542 3904 13598 3913
rect 13542 3839 13598 3848
rect 13556 480 13584 3839
rect 14752 480 14780 31010
rect 17038 3224 17094 3233
rect 17038 3159 17094 3168
rect 17052 480 17080 3159
rect 18248 480 18276 33730
rect 19432 28552 19484 28558
rect 19432 28494 19484 28500
rect 19444 480 19472 28494
rect 21824 3596 21876 3602
rect 21824 3538 21876 3544
rect 21836 480 21864 3538
rect 23032 480 23060 33798
rect 24216 3460 24268 3466
rect 24216 3402 24268 3408
rect 24228 480 24256 3402
rect 26528 480 26556 39374
rect 31300 33924 31352 33930
rect 31300 33866 31352 33872
rect 28908 28620 28960 28626
rect 28908 28562 28960 28568
rect 27712 3528 27764 3534
rect 27712 3470 27764 3476
rect 27724 480 27752 3470
rect 28920 480 28948 28562
rect 30104 3732 30156 3738
rect 30104 3674 30156 3680
rect 30116 480 30144 3674
rect 31312 480 31340 33866
rect 32404 28348 32456 28354
rect 32404 28290 32456 28296
rect 32416 480 32444 28290
rect 33612 480 33640 39442
rect 34796 33992 34848 33998
rect 34796 33934 34848 33940
rect 34808 480 34836 33934
rect 35992 28416 36044 28422
rect 35992 28358 36044 28364
rect 36004 480 36032 28358
rect 37200 480 37228 39510
rect 39580 3868 39632 3874
rect 39580 3810 39632 3816
rect 38384 3800 38436 3806
rect 38384 3742 38436 3748
rect 38396 480 38424 3742
rect 39592 480 39620 3810
rect 40696 480 40724 39578
rect 45468 34196 45520 34202
rect 45468 34138 45520 34144
rect 41880 34128 41932 34134
rect 41880 34070 41932 34076
rect 41892 480 41920 34070
rect 43076 28484 43128 28490
rect 43076 28426 43128 28432
rect 43088 480 43116 28426
rect 44272 3664 44324 3670
rect 44272 3606 44324 3612
rect 44284 480 44312 3606
rect 45480 480 45508 34138
rect 46664 3936 46716 3942
rect 46664 3878 46716 3884
rect 46676 480 46704 3878
rect 47872 480 47900 44882
rect 48964 39704 49016 39710
rect 48964 39646 49016 39652
rect 48976 480 49004 39646
rect 50160 34060 50212 34066
rect 50160 34002 50212 34008
rect 50172 480 50200 34002
rect 51368 480 51396 44950
rect 52552 39772 52604 39778
rect 52552 39714 52604 39720
rect 52564 480 52592 39714
rect 53748 4004 53800 4010
rect 53748 3946 53800 3952
rect 53760 480 53788 3946
rect 54956 480 54984 45018
rect 56048 39840 56100 39846
rect 56048 39782 56100 39788
rect 56060 480 56088 39782
rect 57244 31136 57296 31142
rect 57244 31078 57296 31084
rect 57256 480 57284 31078
rect 58452 480 58480 45086
rect 59636 39908 59688 39914
rect 59636 39850 59688 39856
rect 59648 480 59676 39850
rect 60832 31204 60884 31210
rect 60832 31146 60884 31152
rect 60844 480 60872 31146
rect 62040 480 62068 45154
rect 63224 39976 63276 39982
rect 63224 39918 63276 39924
rect 63236 480 63264 39918
rect 64328 31272 64380 31278
rect 64328 31214 64380 31220
rect 64340 480 64368 31214
rect 65536 480 65564 45222
rect 69112 44804 69164 44810
rect 69112 44746 69164 44752
rect 66720 36576 66772 36582
rect 66720 36518 66772 36524
rect 66732 480 66760 36518
rect 67916 31340 67968 31346
rect 67916 31282 67968 31288
rect 67928 480 67956 31282
rect 69124 480 69152 44746
rect 72608 44736 72660 44742
rect 72608 44678 72660 44684
rect 70308 36644 70360 36650
rect 70308 36586 70360 36592
rect 70320 480 70348 36586
rect 71504 31408 71556 31414
rect 71504 31350 71556 31356
rect 71516 480 71544 31350
rect 72620 480 72648 44678
rect 76196 44668 76248 44674
rect 76196 44610 76248 44616
rect 73804 36712 73856 36718
rect 73804 36654 73856 36660
rect 73816 480 73844 36654
rect 75000 4072 75052 4078
rect 75000 4014 75052 4020
rect 75012 480 75040 4014
rect 76208 480 76236 44610
rect 111616 42764 111668 42770
rect 111616 42706 111668 42712
rect 108120 42696 108172 42702
rect 108120 42638 108172 42644
rect 104532 42628 104584 42634
rect 104532 42570 104584 42576
rect 101036 42560 101088 42566
rect 101036 42502 101088 42508
rect 97448 42492 97500 42498
rect 97448 42434 97500 42440
rect 93952 42424 94004 42430
rect 93952 42366 94004 42372
rect 90364 42356 90416 42362
rect 90364 42298 90416 42304
rect 86868 42288 86920 42294
rect 86868 42230 86920 42236
rect 83280 42220 83332 42226
rect 83280 42162 83332 42168
rect 79692 42152 79744 42158
rect 79692 42094 79744 42100
rect 77392 36780 77444 36786
rect 77392 36722 77444 36728
rect 77404 480 77432 36722
rect 78588 31476 78640 31482
rect 78588 31418 78640 31424
rect 78600 480 78628 31418
rect 79704 480 79732 42094
rect 80888 36848 80940 36854
rect 80888 36790 80940 36796
rect 80900 480 80928 36790
rect 82084 4140 82136 4146
rect 82084 4082 82136 4088
rect 82096 480 82124 4082
rect 83292 480 83320 42162
rect 84476 36916 84528 36922
rect 84476 36858 84528 36864
rect 84488 480 84516 36858
rect 85672 31544 85724 31550
rect 85672 31486 85724 31492
rect 85684 480 85712 31486
rect 86880 480 86908 42230
rect 87972 36984 88024 36990
rect 87972 36926 88024 36932
rect 87984 480 88012 36926
rect 89168 3392 89220 3398
rect 89168 3334 89220 3340
rect 89180 480 89208 3334
rect 90376 480 90404 42298
rect 91560 37052 91612 37058
rect 91560 36994 91612 37000
rect 91572 480 91600 36994
rect 92756 31612 92808 31618
rect 92756 31554 92808 31560
rect 92768 480 92796 31554
rect 93964 480 93992 42366
rect 95148 37120 95200 37126
rect 95148 37062 95200 37068
rect 95160 480 95188 37062
rect 96252 31680 96304 31686
rect 96252 31622 96304 31628
rect 96264 480 96292 31622
rect 97460 480 97488 42434
rect 98644 37188 98696 37194
rect 98644 37130 98696 37136
rect 98656 480 98684 37130
rect 99840 31748 99892 31754
rect 99840 31690 99892 31696
rect 99852 480 99880 31690
rect 101048 480 101076 42502
rect 102232 37256 102284 37262
rect 102232 37198 102284 37204
rect 102244 480 102272 37198
rect 103336 3324 103388 3330
rect 103336 3266 103388 3272
rect 103348 480 103376 3266
rect 104544 480 104572 42570
rect 105728 36508 105780 36514
rect 105728 36450 105780 36456
rect 105740 480 105768 36450
rect 106924 31000 106976 31006
rect 106924 30942 106976 30948
rect 106936 480 106964 30942
rect 108132 480 108160 42638
rect 109316 34264 109368 34270
rect 109316 34206 109368 34212
rect 109328 480 109356 34206
rect 109684 28688 109736 28694
rect 109684 28630 109736 28636
rect 109696 3262 109724 28630
rect 109684 3256 109736 3262
rect 109684 3198 109736 3204
rect 110512 3256 110564 3262
rect 110512 3198 110564 3204
rect 110524 480 110552 3198
rect 111628 480 111656 42706
rect 115204 42016 115256 42022
rect 115204 41958 115256 41964
rect 112812 34332 112864 34338
rect 112812 34274 112864 34280
rect 112824 480 112852 34274
rect 114008 28756 114060 28762
rect 114008 28698 114060 28704
rect 114020 480 114048 28698
rect 115216 480 115244 41958
rect 118792 40044 118844 40050
rect 118792 39986 118844 39992
rect 116400 34400 116452 34406
rect 116400 34342 116452 34348
rect 116412 480 116440 34342
rect 117596 28892 117648 28898
rect 117596 28834 117648 28840
rect 117608 480 117636 28834
rect 118804 480 118832 39986
rect 122288 39296 122340 39302
rect 122288 39238 122340 39244
rect 119896 34468 119948 34474
rect 119896 34410 119948 34416
rect 119908 480 119936 34410
rect 121092 28824 121144 28830
rect 121092 28766 121144 28772
rect 121104 480 121132 28766
rect 122300 480 122328 39238
rect 123484 33720 123536 33726
rect 123484 33662 123536 33668
rect 123496 480 123524 33662
rect 124680 28960 124732 28966
rect 124680 28902 124732 28908
rect 124692 480 124720 28902
rect 360856 3262 360884 305623
rect 362316 305594 362368 305600
rect 361764 304972 361816 304978
rect 361764 304914 361816 304920
rect 361776 304473 361804 304914
rect 361762 304464 361818 304473
rect 361762 304399 361818 304408
rect 360936 304292 360988 304298
rect 360936 304234 360988 304240
rect 360948 3874 360976 304234
rect 362222 302832 362278 302841
rect 362222 302767 362278 302776
rect 361028 300280 361080 300286
rect 361028 300222 361080 300228
rect 360936 3868 360988 3874
rect 360936 3810 360988 3816
rect 361040 3330 361068 300222
rect 361120 297832 361172 297838
rect 361120 297774 361172 297780
rect 361132 3398 361160 297774
rect 361764 293956 361816 293962
rect 361764 293898 361816 293904
rect 361776 293457 361804 293898
rect 361762 293448 361818 293457
rect 361762 293383 361818 293392
rect 361212 291848 361264 291854
rect 361212 291790 361264 291796
rect 361224 33930 361252 291790
rect 361764 282872 361816 282878
rect 361764 282814 361816 282820
rect 361776 282441 361804 282814
rect 361762 282432 361818 282441
rect 361762 282367 361818 282376
rect 361764 271856 361816 271862
rect 361764 271798 361816 271804
rect 361776 271425 361804 271798
rect 361762 271416 361818 271425
rect 361762 271351 361818 271360
rect 361764 260840 361816 260846
rect 361764 260782 361816 260788
rect 361776 260409 361804 260782
rect 361762 260400 361818 260409
rect 361762 260335 361818 260344
rect 361764 249756 361816 249762
rect 361764 249698 361816 249704
rect 361776 249393 361804 249698
rect 361762 249384 361818 249393
rect 361762 249319 361818 249328
rect 361764 238740 361816 238746
rect 361764 238682 361816 238688
rect 361776 238377 361804 238682
rect 361762 238368 361818 238377
rect 361762 238303 361818 238312
rect 361764 227724 361816 227730
rect 361764 227666 361816 227672
rect 361776 227361 361804 227666
rect 361762 227352 361818 227361
rect 361762 227287 361818 227296
rect 361672 216368 361724 216374
rect 361670 216336 361672 216345
rect 361724 216336 361726 216345
rect 361670 216271 361726 216280
rect 361764 205624 361816 205630
rect 361764 205566 361816 205572
rect 361776 205329 361804 205566
rect 361762 205320 361818 205329
rect 361762 205255 361818 205264
rect 361764 194540 361816 194546
rect 361764 194482 361816 194488
rect 361776 194313 361804 194482
rect 361762 194304 361818 194313
rect 361762 194239 361818 194248
rect 361764 183524 361816 183530
rect 361764 183466 361816 183472
rect 361776 183297 361804 183466
rect 361762 183288 361818 183297
rect 361762 183223 361818 183232
rect 361764 172508 361816 172514
rect 361764 172450 361816 172456
rect 361776 172281 361804 172450
rect 361762 172272 361818 172281
rect 361762 172207 361818 172216
rect 361764 161424 361816 161430
rect 361764 161366 361816 161372
rect 361776 161265 361804 161366
rect 361762 161256 361818 161265
rect 361762 161191 361818 161200
rect 361580 158024 361632 158030
rect 361580 157966 361632 157972
rect 361592 154442 361620 157966
rect 361316 154414 361620 154442
rect 361316 46617 361344 154414
rect 361764 150408 361816 150414
rect 361764 150350 361816 150356
rect 361776 150249 361804 150350
rect 361762 150240 361818 150249
rect 361762 150175 361818 150184
rect 361764 139392 361816 139398
rect 361764 139334 361816 139340
rect 361776 139233 361804 139334
rect 361762 139224 361818 139233
rect 361762 139159 361818 139168
rect 361396 131164 361448 131170
rect 361396 131106 361448 131112
rect 361302 46608 361358 46617
rect 361302 46543 361358 46552
rect 361408 45354 361436 131106
rect 361764 128308 361816 128314
rect 361764 128250 361816 128256
rect 361776 128217 361804 128250
rect 361762 128208 361818 128217
rect 361762 128143 361818 128152
rect 361764 117292 361816 117298
rect 361764 117234 361816 117240
rect 361776 117201 361804 117234
rect 361762 117192 361818 117201
rect 361762 117127 361818 117136
rect 361764 106276 361816 106282
rect 361764 106218 361816 106224
rect 361776 106185 361804 106218
rect 361762 106176 361818 106185
rect 361762 106111 361818 106120
rect 361764 95192 361816 95198
rect 361762 95160 361764 95169
rect 361816 95160 361818 95169
rect 361762 95095 361818 95104
rect 361764 84176 361816 84182
rect 361762 84144 361764 84153
rect 361816 84144 361818 84153
rect 361762 84079 361818 84088
rect 361764 73160 361816 73166
rect 361762 73128 361764 73137
rect 361816 73128 361818 73137
rect 361762 73063 361818 73072
rect 361762 62112 361818 62121
rect 361762 62047 361764 62056
rect 361816 62047 361818 62056
rect 361764 62018 361816 62024
rect 361764 51128 361816 51134
rect 361762 51096 361764 51105
rect 361816 51096 361818 51105
rect 361762 51031 361818 51040
rect 361396 45348 361448 45354
rect 361396 45290 361448 45296
rect 361212 33924 361264 33930
rect 361212 33866 361264 33872
rect 362236 4049 362264 302767
rect 362328 39302 362356 305594
rect 363604 304360 363656 304366
rect 363604 304302 363656 304308
rect 362408 297560 362460 297566
rect 362408 297502 362460 297508
rect 362420 39506 362448 297502
rect 362500 297424 362552 297430
rect 362500 297366 362552 297372
rect 362512 40050 362540 297366
rect 362960 143608 363012 143614
rect 362960 143550 363012 143556
rect 362972 137306 363000 143550
rect 362604 137278 363000 137306
rect 362604 131170 362632 137278
rect 362592 131164 362644 131170
rect 362592 131106 362644 131112
rect 362500 40044 362552 40050
rect 362500 39986 362552 39992
rect 362408 39500 362460 39506
rect 362408 39442 362460 39448
rect 362316 39296 362368 39302
rect 362316 39238 362368 39244
rect 362222 4040 362278 4049
rect 362222 3975 362278 3984
rect 363616 3738 363644 304302
rect 363694 302968 363750 302977
rect 363694 302903 363750 302912
rect 363708 3942 363736 302903
rect 363972 297764 364024 297770
rect 363972 297706 364024 297712
rect 363786 297392 363842 297401
rect 363786 297327 363842 297336
rect 363696 3936 363748 3942
rect 363696 3878 363748 3884
rect 363604 3732 363656 3738
rect 363604 3674 363656 3680
rect 363800 3602 363828 297327
rect 363880 291916 363932 291922
rect 363880 291858 363932 291864
rect 363892 33998 363920 291858
rect 363984 39574 364012 297706
rect 364076 216374 364104 333950
rect 367834 305824 367890 305833
rect 367834 305759 367890 305768
rect 364984 302932 365036 302938
rect 364984 302874 365036 302880
rect 364064 216368 364116 216374
rect 364064 216310 364116 216316
rect 364340 144900 364392 144906
rect 364340 144842 364392 144848
rect 364352 139602 364380 144842
rect 364340 139596 364392 139602
rect 364340 139538 364392 139544
rect 363972 39568 364024 39574
rect 363972 39510 364024 39516
rect 363880 33992 363932 33998
rect 363880 33934 363932 33940
rect 364996 4010 365024 302874
rect 367744 301504 367796 301510
rect 367744 301446 367796 301452
rect 365352 300212 365404 300218
rect 365352 300154 365404 300160
rect 365260 300144 365312 300150
rect 365260 300086 365312 300092
rect 365166 297664 365222 297673
rect 365076 297628 365128 297634
rect 365166 297599 365222 297608
rect 365076 297570 365128 297576
rect 364984 4004 365036 4010
rect 364984 3946 365036 3952
rect 363788 3596 363840 3602
rect 363788 3538 363840 3544
rect 361120 3392 361172 3398
rect 361120 3334 361172 3340
rect 361028 3324 361080 3330
rect 361028 3266 361080 3272
rect 360844 3256 360896 3262
rect 365088 3233 365116 297570
rect 365180 39438 365208 297599
rect 365272 42770 365300 300086
rect 365260 42764 365312 42770
rect 365260 42706 365312 42712
rect 365364 42022 365392 300154
rect 366548 297696 366600 297702
rect 366548 297638 366600 297644
rect 366456 297492 366508 297498
rect 366456 297434 366508 297440
rect 366364 291984 366416 291990
rect 366364 291926 366416 291932
rect 365720 147688 365772 147694
rect 365720 147630 365772 147636
rect 365732 144922 365760 147630
rect 365640 144894 365760 144922
rect 365640 143614 365668 144894
rect 365628 143608 365680 143614
rect 365628 143550 365680 143556
rect 365352 42016 365404 42022
rect 365352 41958 365404 41964
rect 365168 39432 365220 39438
rect 365168 39374 365220 39380
rect 366376 3806 366404 291926
rect 366468 39642 366496 297434
rect 366560 39710 366588 297638
rect 366640 286340 366692 286346
rect 366640 286282 366692 286288
rect 366548 39704 366600 39710
rect 366548 39646 366600 39652
rect 366456 39636 366508 39642
rect 366456 39578 366508 39584
rect 366652 31754 366680 286282
rect 366640 31748 366692 31754
rect 366640 31690 366692 31696
rect 367756 4078 367784 301446
rect 367848 42566 367876 305759
rect 370504 301572 370556 301578
rect 370504 301514 370556 301520
rect 367928 300620 367980 300626
rect 367928 300562 367980 300568
rect 367940 42702 367968 300562
rect 368112 300416 368164 300422
rect 368112 300358 368164 300364
rect 368020 300348 368072 300354
rect 368020 300290 368072 300296
rect 367928 42696 367980 42702
rect 367928 42638 367980 42644
rect 368032 42634 368060 300290
rect 368020 42628 368072 42634
rect 368020 42570 368072 42576
rect 367836 42560 367888 42566
rect 367836 42502 367888 42508
rect 368124 42498 368152 300358
rect 369216 297900 369268 297906
rect 369216 297842 369268 297848
rect 368202 297528 368258 297537
rect 368202 297463 368258 297472
rect 368112 42492 368164 42498
rect 368112 42434 368164 42440
rect 368216 39370 368244 297463
rect 369124 292052 369176 292058
rect 369124 291994 369176 292000
rect 368296 149728 368348 149734
rect 368296 149670 368348 149676
rect 368308 144906 368336 149670
rect 368296 144900 368348 144906
rect 368296 144842 368348 144848
rect 368204 39364 368256 39370
rect 368204 39306 368256 39312
rect 369136 34134 369164 291994
rect 369228 39778 369256 297842
rect 369400 294636 369452 294642
rect 369400 294578 369452 294584
rect 369308 286408 369360 286414
rect 369308 286350 369360 286356
rect 369216 39772 369268 39778
rect 369216 39714 369268 39720
rect 369124 34128 369176 34134
rect 369124 34070 369176 34076
rect 369320 31006 369348 286350
rect 369412 39914 369440 294578
rect 369400 39908 369452 39914
rect 369400 39850 369452 39856
rect 369308 31000 369360 31006
rect 369308 30942 369360 30948
rect 370516 4146 370544 301514
rect 370780 300756 370832 300762
rect 370780 300698 370832 300704
rect 370688 300688 370740 300694
rect 370688 300630 370740 300636
rect 370596 297968 370648 297974
rect 370596 297910 370648 297916
rect 370608 39846 370636 297910
rect 370700 42226 370728 300630
rect 370792 42294 370820 300698
rect 370872 300552 370924 300558
rect 370872 300494 370924 300500
rect 370884 42362 370912 300494
rect 370964 300484 371016 300490
rect 370964 300426 371016 300432
rect 370976 42430 371004 300426
rect 372068 295180 372120 295186
rect 372068 295122 372120 295128
rect 371976 295112 372028 295118
rect 371976 295054 372028 295060
rect 371884 294704 371936 294710
rect 371884 294646 371936 294652
rect 371240 149796 371292 149802
rect 371240 149738 371292 149744
rect 371252 147694 371280 149738
rect 371240 147688 371292 147694
rect 371240 147630 371292 147636
rect 370964 42424 371016 42430
rect 370964 42366 371016 42372
rect 370872 42356 370924 42362
rect 370872 42298 370924 42304
rect 370780 42288 370832 42294
rect 370780 42230 370832 42236
rect 370688 42220 370740 42226
rect 370688 42162 370740 42168
rect 370596 39840 370648 39846
rect 370596 39782 370648 39788
rect 371896 36582 371924 294646
rect 371988 36650 372016 295054
rect 372080 36786 372108 295122
rect 372344 294772 372396 294778
rect 372344 294714 372396 294720
rect 372252 289128 372304 289134
rect 372252 289070 372304 289076
rect 372160 286476 372212 286482
rect 372160 286418 372212 286424
rect 372068 36780 372120 36786
rect 372068 36722 372120 36728
rect 371976 36644 372028 36650
rect 371976 36586 372028 36592
rect 371884 36576 371936 36582
rect 371884 36518 371936 36524
rect 372172 28762 372200 286418
rect 372264 34202 372292 289070
rect 372356 39982 372384 294714
rect 372344 39976 372396 39982
rect 372344 39918 372396 39924
rect 372252 34196 372304 34202
rect 372252 34138 372304 34144
rect 373276 28898 373304 386378
rect 374656 379506 374684 601666
rect 376036 380866 376064 623766
rect 377404 385416 377456 385422
rect 377404 385358 377456 385364
rect 376024 380860 376076 380866
rect 376024 380802 376076 380808
rect 374644 379500 374696 379506
rect 374644 379442 374696 379448
rect 374644 339516 374696 339522
rect 374644 339458 374696 339464
rect 374656 315994 374684 339458
rect 374644 315988 374696 315994
rect 374644 315930 374696 315936
rect 376668 303544 376720 303550
rect 376668 303486 376720 303492
rect 376576 303204 376628 303210
rect 376576 303146 376628 303152
rect 376392 303136 376444 303142
rect 376392 303078 376444 303084
rect 376300 303000 376352 303006
rect 376300 302942 376352 302948
rect 373632 302864 373684 302870
rect 373632 302806 373684 302812
rect 373448 300076 373500 300082
rect 373448 300018 373500 300024
rect 373356 294840 373408 294846
rect 373356 294782 373408 294788
rect 373368 36718 373396 294782
rect 373460 42158 373488 300018
rect 373540 300008 373592 300014
rect 373540 299950 373592 299956
rect 373448 42152 373500 42158
rect 373448 42094 373500 42100
rect 373552 42090 373580 299950
rect 373644 46238 373672 302806
rect 376024 302796 376076 302802
rect 376024 302738 376076 302744
rect 375932 302728 375984 302734
rect 375932 302670 375984 302676
rect 373724 300824 373776 300830
rect 373724 300766 373776 300772
rect 373632 46232 373684 46238
rect 373632 46174 373684 46180
rect 373736 44674 373764 300766
rect 374644 295316 374696 295322
rect 374644 295258 374696 295264
rect 373724 44668 373776 44674
rect 373724 44610 373776 44616
rect 373540 42084 373592 42090
rect 373540 42026 373592 42032
rect 373356 36712 373408 36718
rect 373356 36654 373408 36660
rect 373264 28892 373316 28898
rect 373264 28834 373316 28840
rect 372160 28756 372212 28762
rect 372160 28698 372212 28704
rect 370504 4140 370556 4146
rect 370504 4082 370556 4088
rect 367744 4072 367796 4078
rect 367744 4014 367796 4020
rect 374656 3913 374684 295258
rect 375104 295044 375156 295050
rect 375104 294986 375156 294992
rect 375012 294976 375064 294982
rect 375012 294918 375064 294924
rect 374920 294568 374972 294574
rect 374920 294510 374972 294516
rect 374828 289808 374880 289814
rect 374828 289750 374880 289756
rect 374734 286376 374790 286385
rect 374734 286311 374790 286320
rect 374748 28558 374776 286311
rect 374736 28552 374788 28558
rect 374736 28494 374788 28500
rect 374642 3904 374698 3913
rect 374642 3839 374698 3848
rect 366364 3800 366416 3806
rect 374840 3777 374868 289750
rect 374932 36854 374960 294510
rect 375024 36990 375052 294918
rect 375116 37058 375144 294986
rect 375840 276684 375892 276690
rect 375840 276626 375892 276632
rect 375196 161560 375248 161566
rect 375196 161502 375248 161508
rect 375208 73166 375236 161502
rect 375196 73160 375248 73166
rect 375196 73102 375248 73108
rect 375852 45422 375880 276626
rect 375944 46510 375972 302670
rect 375932 46504 375984 46510
rect 375932 46446 375984 46452
rect 376036 45490 376064 302738
rect 376208 294500 376260 294506
rect 376208 294442 376260 294448
rect 376116 289196 376168 289202
rect 376116 289138 376168 289144
rect 376024 45484 376076 45490
rect 376024 45426 376076 45432
rect 375840 45416 375892 45422
rect 375840 45358 375892 45364
rect 375104 37052 375156 37058
rect 375104 36994 375156 37000
rect 375012 36984 375064 36990
rect 375012 36926 375064 36932
rect 374920 36848 374972 36854
rect 374920 36790 374972 36796
rect 376128 31686 376156 289138
rect 376220 36922 376248 294442
rect 376312 45286 376340 302942
rect 376300 45280 376352 45286
rect 376300 45222 376352 45228
rect 376404 45218 376432 303078
rect 376484 303068 376536 303074
rect 376484 303010 376536 303016
rect 376392 45212 376444 45218
rect 376392 45154 376444 45160
rect 376496 44810 376524 303010
rect 376484 44804 376536 44810
rect 376484 44746 376536 44752
rect 376588 44742 376616 303146
rect 376680 46306 376708 303486
rect 376668 46300 376720 46306
rect 376668 46242 376720 46248
rect 376576 44736 376628 44742
rect 376576 44678 376628 44684
rect 376208 36916 376260 36922
rect 376208 36858 376260 36864
rect 376116 31680 376168 31686
rect 376116 31622 376168 31628
rect 377416 28830 377444 385358
rect 378796 382226 378824 645866
rect 378876 522300 378928 522306
rect 378876 522242 378928 522248
rect 378888 508502 378916 522242
rect 378876 508496 378928 508502
rect 378876 508438 378928 508444
rect 381268 508496 381320 508502
rect 381268 508438 381320 508444
rect 381280 501634 381308 508438
rect 381268 501628 381320 501634
rect 381268 501570 381320 501576
rect 380164 386504 380216 386510
rect 380164 386446 380216 386452
rect 378784 382220 378836 382226
rect 378784 382162 378836 382168
rect 378876 306196 378928 306202
rect 378876 306138 378928 306144
rect 378600 303612 378652 303618
rect 378600 303554 378652 303560
rect 377588 294908 377640 294914
rect 377588 294850 377640 294856
rect 377496 289468 377548 289474
rect 377496 289410 377548 289416
rect 377508 31278 377536 289410
rect 377600 37126 377628 294850
rect 377772 292256 377824 292262
rect 377772 292198 377824 292204
rect 377680 289400 377732 289406
rect 377680 289342 377732 289348
rect 377588 37120 377640 37126
rect 377588 37062 377640 37068
rect 377692 34066 377720 289342
rect 377784 37262 377812 292198
rect 378612 46578 378640 303554
rect 378692 303408 378744 303414
rect 378692 303350 378744 303356
rect 378600 46572 378652 46578
rect 378600 46514 378652 46520
rect 378704 45014 378732 303350
rect 378784 286612 378836 286618
rect 378784 286554 378836 286560
rect 378692 45008 378744 45014
rect 378692 44950 378744 44956
rect 377772 37256 377824 37262
rect 377772 37198 377824 37204
rect 377680 34060 377732 34066
rect 377680 34002 377732 34008
rect 377496 31272 377548 31278
rect 377496 31214 377548 31220
rect 377404 28824 377456 28830
rect 377404 28766 377456 28772
rect 378796 20670 378824 286554
rect 378888 46646 378916 306138
rect 378968 305924 379020 305930
rect 378968 305866 379020 305872
rect 378980 46714 379008 305866
rect 379336 303476 379388 303482
rect 379336 303418 379388 303424
rect 379244 303340 379296 303346
rect 379244 303282 379296 303288
rect 379152 295248 379204 295254
rect 379152 295190 379204 295196
rect 379060 289264 379112 289270
rect 379060 289206 379112 289212
rect 378968 46708 379020 46714
rect 378968 46650 379020 46656
rect 378876 46640 378928 46646
rect 378876 46582 378928 46588
rect 379072 31618 379100 289206
rect 379164 37194 379192 295190
rect 379256 45150 379284 303282
rect 379244 45144 379296 45150
rect 379244 45086 379296 45092
rect 379348 44946 379376 303418
rect 379428 303272 379480 303278
rect 379428 303214 379480 303220
rect 379440 45082 379468 303214
rect 379428 45076 379480 45082
rect 379428 45018 379480 45024
rect 379336 44940 379388 44946
rect 379336 44882 379388 44888
rect 379152 37188 379204 37194
rect 379152 37130 379204 37136
rect 379060 31612 379112 31618
rect 379060 31554 379112 31560
rect 380176 28966 380204 386446
rect 381556 383654 381584 656882
rect 381544 383648 381596 383654
rect 381544 383590 381596 383596
rect 382936 383586 382964 667898
rect 385776 458244 385828 458250
rect 385776 458186 385828 458192
rect 385684 386572 385736 386578
rect 385684 386514 385736 386520
rect 382924 383580 382976 383586
rect 382924 383522 382976 383528
rect 383016 307080 383068 307086
rect 383016 307022 383068 307028
rect 382004 306264 382056 306270
rect 382004 306206 382056 306212
rect 381542 306096 381598 306105
rect 381542 306031 381598 306040
rect 381912 306060 381964 306066
rect 381450 303104 381506 303113
rect 381450 303039 381506 303048
rect 380440 292392 380492 292398
rect 380440 292334 380492 292340
rect 380348 289604 380400 289610
rect 380348 289546 380400 289552
rect 380256 289332 380308 289338
rect 380256 289274 380308 289280
rect 380268 31346 380296 289274
rect 380256 31340 380308 31346
rect 380256 31282 380308 31288
rect 380360 31142 380388 289546
rect 380452 34338 380480 292334
rect 381360 292324 381412 292330
rect 381360 292266 381412 292272
rect 380532 292120 380584 292126
rect 380532 292062 380584 292068
rect 380544 36514 380572 292062
rect 380532 36508 380584 36514
rect 380532 36450 380584 36456
rect 380440 34332 380492 34338
rect 380440 34274 380492 34280
rect 381372 34270 381400 292266
rect 381464 44878 381492 303039
rect 381452 44872 381504 44878
rect 381452 44814 381504 44820
rect 381360 34264 381412 34270
rect 381360 34206 381412 34212
rect 380348 31136 380400 31142
rect 380348 31078 380400 31084
rect 380164 28960 380216 28966
rect 380164 28902 380216 28908
rect 378784 20664 378836 20670
rect 378784 20606 378836 20612
rect 366364 3742 366416 3748
rect 374826 3768 374882 3777
rect 374826 3703 374882 3712
rect 381556 3641 381584 306031
rect 381912 306002 381964 306008
rect 381726 305960 381782 305969
rect 381726 305895 381782 305904
rect 381636 298784 381688 298790
rect 381636 298726 381688 298732
rect 381648 6866 381676 298726
rect 381636 6860 381688 6866
rect 381636 6802 381688 6808
rect 381542 3632 381598 3641
rect 381542 3567 381598 3576
rect 381740 3505 381768 305895
rect 381820 305720 381872 305726
rect 381820 305662 381872 305668
rect 381832 45558 381860 305662
rect 381924 46850 381952 306002
rect 381912 46844 381964 46850
rect 381912 46786 381964 46792
rect 382016 46782 382044 306206
rect 382096 305992 382148 305998
rect 382096 305934 382148 305940
rect 382004 46776 382056 46782
rect 382004 46718 382056 46724
rect 382108 46374 382136 305934
rect 382924 298036 382976 298042
rect 382924 297978 382976 297984
rect 382188 289536 382240 289542
rect 382188 289478 382240 289484
rect 382096 46368 382148 46374
rect 382096 46310 382148 46316
rect 381820 45552 381872 45558
rect 381820 45494 381872 45500
rect 382200 31550 382228 289478
rect 382188 31544 382240 31550
rect 382188 31486 382240 31492
rect 382936 3670 382964 297978
rect 383028 28626 383056 307022
rect 383108 306332 383160 306338
rect 383108 306274 383160 306280
rect 383120 33114 383148 306274
rect 384488 306128 384540 306134
rect 384488 306070 384540 306076
rect 384396 305584 384448 305590
rect 384396 305526 384448 305532
rect 384304 305516 384356 305522
rect 384304 305458 384356 305464
rect 383476 292528 383528 292534
rect 383476 292470 383528 292476
rect 383384 292188 383436 292194
rect 383384 292130 383436 292136
rect 383200 289740 383252 289746
rect 383200 289682 383252 289688
rect 383108 33108 383160 33114
rect 383108 33050 383160 33056
rect 383212 31414 383240 289682
rect 383292 289060 383344 289066
rect 383292 289002 383344 289008
rect 383200 31408 383252 31414
rect 383200 31350 383252 31356
rect 383304 31210 383332 289002
rect 383396 34406 383424 292130
rect 383384 34400 383436 34406
rect 383384 34342 383436 34348
rect 383488 33794 383516 292470
rect 384212 159452 384264 159458
rect 384212 159394 384264 159400
rect 384224 84182 384252 159394
rect 384212 84176 384264 84182
rect 384212 84118 384264 84124
rect 384316 46753 384344 305458
rect 384302 46744 384358 46753
rect 384302 46679 384358 46688
rect 384408 46442 384436 305526
rect 384500 46889 384528 306070
rect 384764 305856 384816 305862
rect 384764 305798 384816 305804
rect 384580 305788 384632 305794
rect 384580 305730 384632 305736
rect 384592 46918 384620 305730
rect 384672 288992 384724 288998
rect 384672 288934 384724 288940
rect 384580 46912 384632 46918
rect 384486 46880 384542 46889
rect 384580 46854 384632 46860
rect 384486 46815 384542 46824
rect 384396 46436 384448 46442
rect 384396 46378 384448 46384
rect 383476 33788 383528 33794
rect 383476 33730 383528 33736
rect 383292 31204 383344 31210
rect 383292 31146 383344 31152
rect 384684 31074 384712 288934
rect 384776 47054 384804 305798
rect 384854 291816 384910 291825
rect 384854 291751 384910 291760
rect 384764 47048 384816 47054
rect 384764 46990 384816 46996
rect 384868 33862 384896 291751
rect 384948 119400 385000 119406
rect 384948 119342 385000 119348
rect 384856 33856 384908 33862
rect 384856 33798 384908 33804
rect 384672 31068 384724 31074
rect 384672 31010 384724 31016
rect 384960 28694 384988 119342
rect 385696 33726 385724 386514
rect 385788 371210 385816 458186
rect 387076 385014 387104 678982
rect 403624 634840 403676 634846
rect 403624 634782 403676 634788
rect 387340 501628 387392 501634
rect 387340 501570 387392 501576
rect 387352 498166 387380 501570
rect 387340 498160 387392 498166
rect 387340 498102 387392 498108
rect 393964 498160 394016 498166
rect 393964 498102 394016 498108
rect 393976 466342 394004 498102
rect 393964 466336 394016 466342
rect 393964 466278 394016 466284
rect 398104 466336 398156 466342
rect 398104 466278 398156 466284
rect 398116 416158 398144 466278
rect 398104 416152 398156 416158
rect 398104 416094 398156 416100
rect 387064 385008 387116 385014
rect 387064 384950 387116 384956
rect 403636 382158 403664 634782
rect 406384 612808 406436 612814
rect 406384 612750 406436 612756
rect 403624 382152 403676 382158
rect 403624 382094 403676 382100
rect 406396 380798 406424 612750
rect 407764 590708 407816 590714
rect 407764 590650 407816 590656
rect 406384 380792 406436 380798
rect 406384 380734 406436 380740
rect 407776 379438 407804 590650
rect 410524 513392 410576 513398
rect 410524 513334 410576 513340
rect 409144 416152 409196 416158
rect 409144 416094 409196 416100
rect 407764 379432 407816 379438
rect 407764 379374 407816 379380
rect 385776 371204 385828 371210
rect 385776 371146 385828 371152
rect 409156 363662 409184 416094
rect 410536 373998 410564 513334
rect 411904 502376 411956 502382
rect 411904 502318 411956 502324
rect 410524 373992 410576 373998
rect 410524 373934 410576 373940
rect 411916 373930 411944 502318
rect 411904 373924 411956 373930
rect 411904 373866 411956 373872
rect 409880 369912 409932 369918
rect 409880 369854 409932 369860
rect 409892 365702 409920 369854
rect 409880 365696 409932 365702
rect 409880 365638 409932 365644
rect 409144 363656 409196 363662
rect 409144 363598 409196 363604
rect 395988 351960 396040 351966
rect 395988 351902 396040 351908
rect 385776 304428 385828 304434
rect 385776 304370 385828 304376
rect 385684 33720 385736 33726
rect 385684 33662 385736 33668
rect 384948 28688 385000 28694
rect 384948 28630 385000 28636
rect 383016 28620 383068 28626
rect 383016 28562 383068 28568
rect 382924 3664 382976 3670
rect 382924 3606 382976 3612
rect 381726 3496 381782 3505
rect 385788 3466 385816 304370
rect 386052 292460 386104 292466
rect 386052 292402 386104 292408
rect 385868 291780 385920 291786
rect 385868 291722 385920 291728
rect 385880 3534 385908 291722
rect 385960 289672 386012 289678
rect 385960 289614 386012 289620
rect 385972 31482 386000 289614
rect 386064 34474 386092 292402
rect 394700 191140 394752 191146
rect 394700 191082 394752 191088
rect 394712 185434 394740 191082
rect 395344 189780 395396 189786
rect 395344 189722 395396 189728
rect 391204 185428 391256 185434
rect 391204 185370 391256 185376
rect 394700 185428 394752 185434
rect 394700 185370 394752 185376
rect 391216 166326 391244 185370
rect 395356 171154 395384 189722
rect 391296 171148 391348 171154
rect 391296 171090 391348 171096
rect 395344 171148 395396 171154
rect 395344 171090 395396 171096
rect 388536 166320 388588 166326
rect 388536 166262 388588 166268
rect 391204 166320 391256 166326
rect 391204 166262 391256 166268
rect 388444 164892 388496 164898
rect 388444 164834 388496 164840
rect 386144 160200 386196 160206
rect 386144 160142 386196 160148
rect 386156 62082 386184 160142
rect 387800 160132 387852 160138
rect 387800 160074 387852 160080
rect 386236 159384 386288 159390
rect 386236 159326 386288 159332
rect 386248 95198 386276 159326
rect 387812 158030 387840 160074
rect 387800 158024 387852 158030
rect 387800 157966 387852 157972
rect 386512 150612 386564 150618
rect 386512 150554 386564 150560
rect 386524 149802 386552 150554
rect 386512 149796 386564 149802
rect 386512 149738 386564 149744
rect 388456 149734 388484 164834
rect 388548 160750 388576 166262
rect 388536 160744 388588 160750
rect 388536 160686 388588 160692
rect 391308 160138 391336 171090
rect 391296 160132 391348 160138
rect 391296 160074 391348 160080
rect 389272 153876 389324 153882
rect 389272 153818 389324 153824
rect 389284 150618 389312 153818
rect 389272 150612 389324 150618
rect 389272 150554 389324 150560
rect 388444 149728 388496 149734
rect 388444 149670 388496 149676
rect 393964 147008 394016 147014
rect 393964 146950 394016 146956
rect 393976 140078 394004 146950
rect 393964 140072 394016 140078
rect 393964 140014 394016 140020
rect 389824 106956 389876 106962
rect 389824 106898 389876 106904
rect 389836 104938 389864 106898
rect 396000 104938 396028 351902
rect 407028 350600 407080 350606
rect 407028 350542 407080 350548
rect 402244 347812 402296 347818
rect 402244 347754 402296 347760
rect 402256 337414 402284 347754
rect 402244 337408 402296 337414
rect 402244 337350 402296 337356
rect 399484 336116 399536 336122
rect 399484 336058 399536 336064
rect 399496 260846 399524 336058
rect 402256 334914 402284 337350
rect 407040 335354 407068 350542
rect 413100 336864 413152 336870
rect 413100 336806 413152 336812
rect 409420 336796 409472 336802
rect 409420 336738 409472 336744
rect 406120 335326 407068 335354
rect 406120 334914 406148 335326
rect 402086 334886 402284 334914
rect 405766 334886 406148 334914
rect 409432 334900 409460 336738
rect 413112 334900 413140 336806
rect 413664 336190 413692 703520
rect 429856 700641 429884 703520
rect 444104 700868 444156 700874
rect 444104 700810 444156 700816
rect 429842 700632 429898 700641
rect 429842 700567 429898 700576
rect 418804 700324 418856 700330
rect 418804 700266 418856 700272
rect 416044 685228 416096 685234
rect 416044 685170 416096 685176
rect 414664 491360 414716 491366
rect 414664 491302 414716 491308
rect 414676 372570 414704 491302
rect 414664 372564 414716 372570
rect 414664 372506 414716 372512
rect 416056 336258 416084 685170
rect 417424 469260 417476 469266
rect 417424 469202 417476 469208
rect 417436 371142 417464 469202
rect 417424 371136 417476 371142
rect 417424 371078 417476 371084
rect 416136 363656 416188 363662
rect 416136 363598 416188 363604
rect 416148 346458 416176 363598
rect 416136 346452 416188 346458
rect 416136 346394 416188 346400
rect 416780 336932 416832 336938
rect 416780 336874 416832 336880
rect 416044 336252 416096 336258
rect 416044 336194 416096 336200
rect 413652 336184 413704 336190
rect 413652 336126 413704 336132
rect 416792 334900 416820 336874
rect 418816 336326 418844 700266
rect 418896 685160 418948 685166
rect 418896 685102 418948 685108
rect 418908 336394 418936 685102
rect 418988 683868 419040 683874
rect 418988 683810 419040 683816
rect 419000 336462 419028 683810
rect 420644 683800 420696 683806
rect 420644 683742 420696 683748
rect 420184 683732 420236 683738
rect 420184 683674 420236 683680
rect 420090 682816 420146 682825
rect 420090 682751 420146 682760
rect 419080 480276 419132 480282
rect 419080 480218 419132 480224
rect 419092 372502 419120 480218
rect 419172 436144 419224 436150
rect 419172 436086 419224 436092
rect 419080 372496 419132 372502
rect 419080 372438 419132 372444
rect 419184 369850 419212 436086
rect 419172 369844 419224 369850
rect 419172 369786 419224 369792
rect 418988 336456 419040 336462
rect 418988 336398 419040 336404
rect 418896 336388 418948 336394
rect 418896 336330 418948 336336
rect 418804 336320 418856 336326
rect 418804 336262 418856 336268
rect 420104 334626 420132 682751
rect 420196 335034 420224 683674
rect 420368 683664 420420 683670
rect 420368 683606 420420 683612
rect 420276 683596 420328 683602
rect 420276 683538 420328 683544
rect 420184 335028 420236 335034
rect 420184 334970 420236 334976
rect 420288 334830 420316 683538
rect 420276 334824 420328 334830
rect 420276 334766 420328 334772
rect 420276 334688 420328 334694
rect 420380 334642 420408 683606
rect 420552 683460 420604 683466
rect 420552 683402 420604 683408
rect 420564 335102 420592 683402
rect 420552 335096 420604 335102
rect 420552 335038 420604 335044
rect 420656 334898 420684 683742
rect 420736 683528 420788 683534
rect 420736 683470 420788 683476
rect 420644 334892 420696 334898
rect 420644 334834 420696 334840
rect 420748 334762 420776 683470
rect 420828 683392 420880 683398
rect 420828 683334 420880 683340
rect 420840 334966 420868 683334
rect 422484 447364 422536 447370
rect 422484 447306 422536 447312
rect 422496 444924 422524 447306
rect 437388 447296 437440 447302
rect 437388 447238 437440 447244
rect 432420 447228 432472 447234
rect 432420 447170 432472 447176
rect 432432 444924 432460 447170
rect 437400 444924 437428 447238
rect 427728 444440 427780 444446
rect 427478 444388 427728 444394
rect 427478 444382 427780 444388
rect 427478 444366 427768 444382
rect 442382 444378 442672 444394
rect 442382 444372 442684 444378
rect 442382 444366 442632 444372
rect 442632 444314 442684 444320
rect 421484 417586 421512 420036
rect 422128 417654 422156 420036
rect 422786 420022 423168 420050
rect 423430 420022 423536 420050
rect 422116 417648 422168 417654
rect 422116 417590 422168 417596
rect 421472 417580 421524 417586
rect 421472 417522 421524 417528
rect 423140 416022 423168 420022
rect 423128 416016 423180 416022
rect 423128 415958 423180 415964
rect 423508 391270 423536 420022
rect 424060 417518 424088 420036
rect 424704 417722 424732 420036
rect 425348 417790 425376 420036
rect 425336 417784 425388 417790
rect 425336 417726 425388 417732
rect 424692 417716 424744 417722
rect 424692 417658 424744 417664
rect 424048 417512 424100 417518
rect 424048 417454 424100 417460
rect 425992 417450 426020 420036
rect 442264 418804 442316 418810
rect 442264 418746 442316 418752
rect 425980 417444 426032 417450
rect 425980 417386 426032 417392
rect 436744 416084 436796 416090
rect 436744 416026 436796 416032
rect 423588 416016 423640 416022
rect 423588 415958 423640 415964
rect 423496 391264 423548 391270
rect 423496 391206 423548 391212
rect 423600 389842 423628 415958
rect 423588 389836 423640 389842
rect 423588 389778 423640 389784
rect 436756 369782 436784 416026
rect 439504 403028 439556 403034
rect 439504 402970 439556 402976
rect 436744 369776 436796 369782
rect 436744 369718 436796 369724
rect 439516 367062 439544 402970
rect 441528 387116 441580 387122
rect 441528 387058 441580 387064
rect 439504 367056 439556 367062
rect 439504 366998 439556 367004
rect 432696 363044 432748 363050
rect 432696 362986 432748 362992
rect 432604 361616 432656 361622
rect 432604 361558 432656 361564
rect 423680 346452 423732 346458
rect 423680 346394 423732 346400
rect 423692 341630 423720 346394
rect 423680 341624 423732 341630
rect 423680 341566 423732 341572
rect 429844 341624 429896 341630
rect 429844 341566 429896 341572
rect 427818 337104 427874 337113
rect 427818 337039 427874 337048
rect 420828 334960 420880 334966
rect 420828 334902 420880 334908
rect 420736 334756 420788 334762
rect 420736 334698 420788 334704
rect 420328 334636 420408 334642
rect 420276 334630 420408 334636
rect 420092 334620 420144 334626
rect 420288 334614 420408 334630
rect 427832 334642 427860 337039
rect 427832 334628 427952 334642
rect 427846 334614 427952 334628
rect 420092 334562 420144 334568
rect 427924 334506 427952 334614
rect 428094 334520 428150 334529
rect 427846 334478 428094 334506
rect 428094 334455 428150 334464
rect 420458 334384 420514 334393
rect 420458 334319 420514 334328
rect 424138 334384 424194 334393
rect 424138 334319 424194 334328
rect 429856 322250 429884 341566
rect 431224 332648 431276 332654
rect 431224 332590 431276 332596
rect 429844 322244 429896 322250
rect 429844 322186 429896 322192
rect 408408 301640 408460 301646
rect 408408 301582 408460 301588
rect 403624 298852 403676 298858
rect 403624 298794 403676 298800
rect 399484 260840 399536 260846
rect 399484 260782 399536 260788
rect 400588 181484 400640 181490
rect 400588 181426 400640 181432
rect 400600 176730 400628 181426
rect 398104 176724 398156 176730
rect 398104 176666 398156 176672
rect 400588 176724 400640 176730
rect 400588 176666 400640 176672
rect 398116 164898 398144 176666
rect 398104 164892 398156 164898
rect 398104 164834 398156 164840
rect 398840 158024 398892 158030
rect 398840 157966 398892 157972
rect 398852 156074 398880 157966
rect 398760 156046 398880 156074
rect 398760 153882 398788 156046
rect 402244 155236 402296 155242
rect 402244 155178 402296 155184
rect 398748 153876 398800 153882
rect 398748 153818 398800 153824
rect 402256 147014 402284 155178
rect 402244 147008 402296 147014
rect 402244 146950 402296 146956
rect 403636 107642 403664 298794
rect 406384 236700 406436 236706
rect 406384 236642 406436 236648
rect 406396 197402 406424 236642
rect 404084 197396 404136 197402
rect 404084 197338 404136 197344
rect 406384 197396 406436 197402
rect 406384 197338 406436 197344
rect 404096 191146 404124 197338
rect 404084 191140 404136 191146
rect 404084 191082 404136 191088
rect 407028 162920 407080 162926
rect 407028 162862 407080 162868
rect 407040 155242 407068 162862
rect 407028 155236 407080 155242
rect 407028 155178 407080 155184
rect 402152 107636 402204 107642
rect 402152 107578 402204 107584
rect 403624 107636 403676 107642
rect 403624 107578 403676 107584
rect 402164 104938 402192 107578
rect 408420 104938 408448 301582
rect 429200 274644 429252 274650
rect 429200 274586 429252 274592
rect 429212 269074 429240 274586
rect 427084 269068 427136 269074
rect 427084 269010 427136 269016
rect 429200 269068 429252 269074
rect 429200 269010 429252 269016
rect 427096 250510 427124 269010
rect 421564 250504 421616 250510
rect 421564 250446 421616 250452
rect 427084 250504 427136 250510
rect 427084 250446 427136 250452
rect 421576 239018 421604 250446
rect 425704 244316 425756 244322
rect 425704 244258 425756 244264
rect 418528 239012 418580 239018
rect 418528 238954 418580 238960
rect 421564 239012 421616 239018
rect 421564 238954 421616 238960
rect 418540 236706 418568 238954
rect 418528 236700 418580 236706
rect 418528 236642 418580 236648
rect 425716 232966 425744 244258
rect 422944 232960 422996 232966
rect 422944 232902 422996 232908
rect 425704 232960 425756 232966
rect 425704 232902 425756 232908
rect 422956 194342 422984 232902
rect 423036 209092 423088 209098
rect 423036 209034 423088 209040
rect 417424 194336 417476 194342
rect 417424 194278 417476 194284
rect 422944 194336 422996 194342
rect 422944 194278 422996 194284
rect 417436 186386 417464 194278
rect 418068 192500 418120 192506
rect 418068 192442 418120 192448
rect 418080 189786 418108 192442
rect 423048 191894 423076 209034
rect 429200 195288 429252 195294
rect 429200 195230 429252 195236
rect 429212 192506 429240 195230
rect 431236 194546 431264 332590
rect 431868 327140 431920 327146
rect 431868 327082 431920 327088
rect 431316 258732 431368 258738
rect 431316 258674 431368 258680
rect 431328 244322 431356 258674
rect 431316 244316 431368 244322
rect 431316 244258 431368 244264
rect 431224 194540 431276 194546
rect 431224 194482 431276 194488
rect 429200 192500 429252 192506
rect 429200 192442 429252 192448
rect 419540 191888 419592 191894
rect 419540 191830 419592 191836
rect 423036 191888 423088 191894
rect 423036 191830 423088 191836
rect 418068 189780 418120 189786
rect 418068 189722 418120 189728
rect 414664 186380 414716 186386
rect 414664 186322 414716 186328
rect 417424 186380 417476 186386
rect 417424 186322 417476 186328
rect 413928 183660 413980 183666
rect 413928 183602 413980 183608
rect 413940 181490 413968 183602
rect 413928 181484 413980 181490
rect 413928 181426 413980 181432
rect 414676 162926 414704 186322
rect 419552 183666 419580 191830
rect 419540 183660 419592 183666
rect 419540 183602 419592 183608
rect 430580 182232 430632 182238
rect 430580 182174 430632 182180
rect 430592 176730 430620 182174
rect 430580 176724 430632 176730
rect 430580 176666 430632 176672
rect 422944 176656 422996 176662
rect 422944 176598 422996 176604
rect 422956 169794 422984 176598
rect 420184 169788 420236 169794
rect 420184 169730 420236 169736
rect 422944 169788 422996 169794
rect 422944 169730 422996 169736
rect 414664 162920 414716 162926
rect 414664 162862 414716 162868
rect 418712 162240 418764 162246
rect 418712 162182 418764 162188
rect 415124 162172 415176 162178
rect 415124 162114 415176 162120
rect 412088 161492 412140 161498
rect 412088 161434 412140 161440
rect 409512 160132 409564 160138
rect 409512 160074 409564 160080
rect 409144 159724 409196 159730
rect 409144 159666 409196 159672
rect 409156 106282 409184 159666
rect 409236 159656 409288 159662
rect 409236 159598 409288 159604
rect 409248 117298 409276 159598
rect 409328 159588 409380 159594
rect 409328 159530 409380 159536
rect 409340 128314 409368 159530
rect 409420 159520 409472 159526
rect 409420 159462 409472 159468
rect 409432 139398 409460 159462
rect 409524 150414 409552 160074
rect 412100 159882 412128 161434
rect 415136 160206 415164 162114
rect 418724 161566 418752 162182
rect 418712 161560 418764 161566
rect 418712 161502 418764 161508
rect 415124 160200 415176 160206
rect 411792 159854 412128 159882
rect 415090 160148 415124 160154
rect 415090 160142 415176 160148
rect 415090 160126 415164 160142
rect 415090 159868 415118 160126
rect 418724 159882 418752 161502
rect 418416 159854 418752 159882
rect 420196 159798 420224 169730
rect 421838 162752 421894 162761
rect 421838 162687 421894 162696
rect 425886 162752 425942 162761
rect 425886 162687 425942 162696
rect 428646 162752 428702 162761
rect 428646 162687 428702 162696
rect 421852 160410 421880 162687
rect 425900 160546 425928 162687
rect 425336 160540 425388 160546
rect 425336 160482 425388 160488
rect 425888 160540 425940 160546
rect 425888 160482 425940 160488
rect 421840 160404 421892 160410
rect 421840 160346 421892 160352
rect 409880 159792 409932 159798
rect 409880 159734 409932 159740
rect 420184 159792 420236 159798
rect 420184 159734 420236 159740
rect 409892 158030 409920 159734
rect 421380 159452 421432 159458
rect 421380 159394 421432 159400
rect 421392 159338 421420 159394
rect 421852 159338 421880 160346
rect 425348 159882 425376 160482
rect 428660 160478 428688 162687
rect 431880 161474 431908 327082
rect 432616 325553 432644 361558
rect 432708 329225 432736 362986
rect 432788 362976 432840 362982
rect 432788 362918 432840 362924
rect 432800 332897 432828 362918
rect 436928 360256 436980 360262
rect 436928 360198 436980 360204
rect 435364 358828 435416 358834
rect 435364 358770 435416 358776
rect 432786 332888 432842 332897
rect 432786 332823 432842 332832
rect 432788 331900 432840 331906
rect 432788 331842 432840 331848
rect 432694 329216 432750 329225
rect 432694 329151 432750 329160
rect 432602 325544 432658 325553
rect 432602 325479 432658 325488
rect 432696 324964 432748 324970
rect 432696 324906 432748 324912
rect 432604 322992 432656 322998
rect 432604 322934 432656 322940
rect 432052 318572 432104 318578
rect 432052 318514 432104 318520
rect 432064 310865 432092 318514
rect 432616 314537 432644 322934
rect 432708 318209 432736 324906
rect 432800 321881 432828 331842
rect 432786 321872 432842 321881
rect 432786 321807 432842 321816
rect 435376 318578 435404 358770
rect 435456 339584 435508 339590
rect 435456 339526 435508 339532
rect 435364 318572 435416 318578
rect 435364 318514 435416 318520
rect 432694 318200 432750 318209
rect 432694 318135 432750 318144
rect 432602 314528 432658 314537
rect 432602 314463 432658 314472
rect 432696 313948 432748 313954
rect 432696 313890 432748 313896
rect 432050 310856 432106 310865
rect 432050 310791 432106 310800
rect 432708 307193 432736 313890
rect 432694 307184 432750 307193
rect 432694 307119 432750 307128
rect 435468 304978 435496 339526
rect 436836 338156 436888 338162
rect 436836 338098 436888 338104
rect 436744 332716 436796 332722
rect 436744 332658 436796 332664
rect 436008 328500 436060 328506
rect 436008 328442 436060 328448
rect 435456 304972 435508 304978
rect 435456 304914 435508 304920
rect 435364 295384 435416 295390
rect 435364 295326 435416 295332
rect 435376 282130 435404 295326
rect 432604 282124 432656 282130
rect 432604 282066 432656 282072
rect 435364 282124 435416 282130
rect 435364 282066 435416 282072
rect 432616 274650 432644 282066
rect 432604 274644 432656 274650
rect 432604 274586 432656 274592
rect 432604 213920 432656 213926
rect 432604 213862 432656 213868
rect 432616 209098 432644 213862
rect 432604 209092 432656 209098
rect 432604 209034 432656 209040
rect 433064 187740 433116 187746
rect 433064 187682 433116 187688
rect 433076 182238 433104 187682
rect 433064 182232 433116 182238
rect 433064 182174 433116 182180
rect 431788 161446 431908 161474
rect 428648 160472 428700 160478
rect 428648 160414 428700 160420
rect 425040 159854 425376 159882
rect 425164 159390 425192 159854
rect 428660 159746 428688 160414
rect 431788 160274 431816 161446
rect 436020 160342 436048 328442
rect 436756 205630 436784 332658
rect 436848 293962 436876 338098
rect 436940 322998 436968 360198
rect 438860 341012 438912 341018
rect 438860 340954 438912 340960
rect 438124 336524 438176 336530
rect 438124 336466 438176 336472
rect 436928 322992 436980 322998
rect 436928 322934 436980 322940
rect 436836 293956 436888 293962
rect 436836 293898 436888 293904
rect 438136 271862 438164 336466
rect 438872 336054 438900 340954
rect 439688 338224 439740 338230
rect 439688 338166 439740 338172
rect 438860 336048 438912 336054
rect 438860 335990 438912 335996
rect 439596 335368 439648 335374
rect 439596 335310 439648 335316
rect 439504 329112 439556 329118
rect 439504 329054 439556 329060
rect 438124 271856 438176 271862
rect 438124 271798 438176 271804
rect 438124 261860 438176 261866
rect 438124 261802 438176 261808
rect 438136 213926 438164 261802
rect 438124 213920 438176 213926
rect 438124 213862 438176 213868
rect 436744 205624 436796 205630
rect 436744 205566 436796 205572
rect 438032 197396 438084 197402
rect 438032 197338 438084 197344
rect 438044 191554 438072 197338
rect 436376 191548 436428 191554
rect 436376 191490 436428 191496
rect 438032 191548 438084 191554
rect 438032 191490 438084 191496
rect 436388 187746 436416 191490
rect 436376 187740 436428 187746
rect 436376 187682 436428 187688
rect 439516 163674 439544 329054
rect 439608 238746 439636 335310
rect 439700 282878 439728 338166
rect 439964 336252 440016 336258
rect 439964 336194 440016 336200
rect 439780 335096 439832 335102
rect 439780 335038 439832 335044
rect 439792 318646 439820 335038
rect 439872 335028 439924 335034
rect 439872 334970 439924 334976
rect 439884 319258 439912 334970
rect 439976 322697 440004 336194
rect 439962 322688 440018 322697
rect 439962 322623 440018 322632
rect 441540 320550 441568 387058
rect 442276 368422 442304 418746
rect 443644 414044 443696 414050
rect 443644 413986 443696 413992
rect 443656 368490 443684 413986
rect 443736 392012 443788 392018
rect 443736 391954 443788 391960
rect 443644 368484 443696 368490
rect 443644 368426 443696 368432
rect 442264 368416 442316 368422
rect 442264 368358 442316 368364
rect 443748 366994 443776 391954
rect 443828 380928 443880 380934
rect 443828 380870 443880 380876
rect 443736 366988 443788 366994
rect 443736 366930 443788 366936
rect 443840 365634 443868 380870
rect 443828 365628 443880 365634
rect 443828 365570 443880 365576
rect 443920 361684 443972 361690
rect 443920 361626 443972 361632
rect 442264 360324 442316 360330
rect 442264 360266 442316 360272
rect 442276 324970 442304 360266
rect 443828 358896 443880 358902
rect 443828 358838 443880 358844
rect 442356 336456 442408 336462
rect 442356 336398 442408 336404
rect 442264 324964 442316 324970
rect 442264 324906 442316 324912
rect 441528 320544 441580 320550
rect 441528 320486 441580 320492
rect 439872 319252 439924 319258
rect 439872 319194 439924 319200
rect 439780 318640 439832 318646
rect 439780 318582 439832 318588
rect 442368 318578 442396 336398
rect 442448 336388 442500 336394
rect 442448 336330 442500 336336
rect 442460 320113 442488 336330
rect 442724 336320 442776 336326
rect 442724 336262 442776 336268
rect 442540 334960 442592 334966
rect 442540 334902 442592 334908
rect 442446 320104 442502 320113
rect 442446 320039 442502 320048
rect 442552 320006 442580 334902
rect 442632 334892 442684 334898
rect 442632 334834 442684 334840
rect 442644 320074 442672 334834
rect 442736 321201 442764 336262
rect 443736 335708 443788 335714
rect 443736 335650 443788 335656
rect 442816 334824 442868 334830
rect 442816 334766 442868 334772
rect 442828 321910 442856 334766
rect 443644 334076 443696 334082
rect 443644 334018 443696 334024
rect 442908 330132 442960 330138
rect 442908 330074 442960 330080
rect 442816 321904 442868 321910
rect 442816 321846 442868 321852
rect 442722 321192 442778 321201
rect 442722 321127 442778 321136
rect 442632 320068 442684 320074
rect 442632 320010 442684 320016
rect 442540 320000 442592 320006
rect 442540 319942 442592 319948
rect 442356 318572 442408 318578
rect 442356 318514 442408 318520
rect 440884 311160 440936 311166
rect 440884 311102 440936 311108
rect 440896 295390 440924 311102
rect 440884 295384 440936 295390
rect 440884 295326 440936 295332
rect 439688 282872 439740 282878
rect 439688 282814 439740 282820
rect 442264 268524 442316 268530
rect 442264 268466 442316 268472
rect 439596 238740 439648 238746
rect 439596 238682 439648 238688
rect 439596 224120 439648 224126
rect 439596 224062 439648 224068
rect 439608 197402 439636 224062
rect 442276 218074 442304 268466
rect 439688 218068 439740 218074
rect 439688 218010 439740 218016
rect 442264 218068 442316 218074
rect 442264 218010 442316 218016
rect 439596 197396 439648 197402
rect 439596 197338 439648 197344
rect 439700 195294 439728 218010
rect 439688 195288 439740 195294
rect 439688 195230 439740 195236
rect 438584 163668 438636 163674
rect 438584 163610 438636 163616
rect 439504 163668 439556 163674
rect 439504 163610 439556 163616
rect 435272 160336 435324 160342
rect 435272 160278 435324 160284
rect 436008 160336 436060 160342
rect 436008 160278 436060 160284
rect 431776 160268 431828 160274
rect 431776 160210 431828 160216
rect 428016 159730 428688 159746
rect 428004 159724 428688 159730
rect 428056 159718 428688 159724
rect 428004 159666 428056 159672
rect 431316 159656 431368 159662
rect 431316 159598 431368 159604
rect 431328 159474 431356 159598
rect 431788 159474 431816 160210
rect 435284 159882 435312 160278
rect 438596 160206 438624 163610
rect 438584 160200 438636 160206
rect 438584 160142 438636 160148
rect 434824 159854 435312 159882
rect 434824 159594 434852 159854
rect 434812 159588 434864 159594
rect 434812 159530 434864 159536
rect 431328 159446 431816 159474
rect 437940 159520 437992 159526
rect 438596 159474 438624 160142
rect 442920 160138 442948 330074
rect 443184 267028 443236 267034
rect 443184 266970 443236 266976
rect 443196 261866 443224 266970
rect 443184 261860 443236 261866
rect 443184 261802 443236 261808
rect 443656 227730 443684 334018
rect 443748 249762 443776 335650
rect 443840 313954 443868 358838
rect 443932 331906 443960 361626
rect 444012 334756 444064 334762
rect 444012 334698 444064 334704
rect 443920 331900 443972 331906
rect 443920 331842 443972 331848
rect 444024 320686 444052 334698
rect 444116 321094 444144 700810
rect 446496 700800 446548 700806
rect 446496 700742 446548 700748
rect 445024 700732 445076 700738
rect 445024 700674 445076 700680
rect 444196 700392 444248 700398
rect 444196 700334 444248 700340
rect 444208 421977 444236 700334
rect 444288 423020 444340 423026
rect 444288 422962 444340 422968
rect 444194 421968 444250 421977
rect 444194 421903 444250 421912
rect 444104 321088 444156 321094
rect 444104 321030 444156 321036
rect 444012 320680 444064 320686
rect 444012 320622 444064 320628
rect 444300 319938 444328 422962
rect 444932 334688 444984 334694
rect 444932 334630 444984 334636
rect 444840 334620 444892 334626
rect 444840 334562 444892 334568
rect 444852 322833 444880 334562
rect 444838 322824 444894 322833
rect 444838 322759 444894 322768
rect 444288 319932 444340 319938
rect 444288 319874 444340 319880
rect 444944 318510 444972 334630
rect 445036 321026 445064 700674
rect 446404 700528 446456 700534
rect 446404 700470 446456 700476
rect 445116 700460 445168 700466
rect 445116 700402 445168 700408
rect 445024 321020 445076 321026
rect 445024 320962 445076 320968
rect 445128 320618 445156 700402
rect 445668 700392 445720 700398
rect 445668 700334 445720 700340
rect 445208 686520 445260 686526
rect 445208 686462 445260 686468
rect 445116 320612 445168 320618
rect 445116 320554 445168 320560
rect 445220 319598 445248 686462
rect 445576 684548 445628 684554
rect 445576 684490 445628 684496
rect 445300 683324 445352 683330
rect 445300 683266 445352 683272
rect 445208 319592 445260 319598
rect 445208 319534 445260 319540
rect 445312 319326 445340 683266
rect 445484 683256 445536 683262
rect 445484 683198 445536 683204
rect 445392 683188 445444 683194
rect 445392 683130 445444 683136
rect 445404 320754 445432 683130
rect 445496 320822 445524 683198
rect 445588 321774 445616 684490
rect 445576 321768 445628 321774
rect 445576 321710 445628 321716
rect 445484 320816 445536 320822
rect 445484 320758 445536 320764
rect 445392 320748 445444 320754
rect 445392 320690 445444 320696
rect 445300 319320 445352 319326
rect 445300 319262 445352 319268
rect 444932 318504 444984 318510
rect 444932 318446 444984 318452
rect 445680 318442 445708 700334
rect 446312 444440 446364 444446
rect 446312 444382 446364 444388
rect 446220 444372 446272 444378
rect 446220 444314 446272 444320
rect 446232 352714 446260 444314
rect 446220 352708 446272 352714
rect 446220 352650 446272 352656
rect 446324 344758 446352 444382
rect 446312 344752 446364 344758
rect 446312 344694 446364 344700
rect 446416 321366 446444 700470
rect 446508 321502 446536 700742
rect 449256 700664 449308 700670
rect 449256 700606 449308 700612
rect 449164 700596 449216 700602
rect 449164 700538 449216 700544
rect 447876 700324 447928 700330
rect 447876 700266 447928 700272
rect 446588 692096 446640 692102
rect 446588 692038 446640 692044
rect 446496 321496 446548 321502
rect 446496 321438 446548 321444
rect 446404 321360 446456 321366
rect 446404 321302 446456 321308
rect 446600 319734 446628 692038
rect 446680 687948 446732 687954
rect 446680 687890 446732 687896
rect 446692 319802 446720 687890
rect 446772 685296 446824 685302
rect 446772 685238 446824 685244
rect 446680 319796 446732 319802
rect 446680 319738 446732 319744
rect 446588 319728 446640 319734
rect 446588 319670 446640 319676
rect 446784 319190 446812 685238
rect 446862 683360 446918 683369
rect 446862 683295 446918 683304
rect 446876 319530 446904 683295
rect 447046 683224 447102 683233
rect 447046 683159 447102 683168
rect 446956 682712 447008 682718
rect 446956 682654 447008 682660
rect 446968 320958 446996 682654
rect 447060 322561 447088 683159
rect 447784 669996 447836 670002
rect 447784 669938 447836 669944
rect 447324 447976 447376 447982
rect 447324 447918 447376 447924
rect 447232 447908 447284 447914
rect 447232 447850 447284 447856
rect 447140 447840 447192 447846
rect 447140 447782 447192 447788
rect 447152 447302 447180 447782
rect 447244 447370 447272 447850
rect 447232 447364 447284 447370
rect 447232 447306 447284 447312
rect 447140 447296 447192 447302
rect 447140 447238 447192 447244
rect 447336 447234 447364 447918
rect 447324 447228 447376 447234
rect 447324 447170 447376 447176
rect 447416 388476 447468 388482
rect 447416 388418 447468 388424
rect 447140 385008 447192 385014
rect 447140 384950 447192 384956
rect 447152 383897 447180 384950
rect 447138 383888 447194 383897
rect 447138 383823 447194 383832
rect 447232 383648 447284 383654
rect 447232 383590 447284 383596
rect 447140 383580 447192 383586
rect 447140 383522 447192 383528
rect 447152 383217 447180 383522
rect 447138 383208 447194 383217
rect 447138 383143 447194 383152
rect 447244 382537 447272 383590
rect 447230 382528 447286 382537
rect 447230 382463 447286 382472
rect 447140 382220 447192 382226
rect 447140 382162 447192 382168
rect 447152 381857 447180 382162
rect 447232 382152 447284 382158
rect 447232 382094 447284 382100
rect 447138 381848 447194 381857
rect 447138 381783 447194 381792
rect 447244 381177 447272 382094
rect 447230 381168 447286 381177
rect 447230 381103 447286 381112
rect 447140 380860 447192 380866
rect 447140 380802 447192 380808
rect 447152 380497 447180 380802
rect 447232 380792 447284 380798
rect 447232 380734 447284 380740
rect 447138 380488 447194 380497
rect 447138 380423 447194 380432
rect 447244 379817 447272 380734
rect 447230 379808 447286 379817
rect 447230 379743 447286 379752
rect 447140 379500 447192 379506
rect 447140 379442 447192 379448
rect 447152 379137 447180 379442
rect 447232 379432 447284 379438
rect 447232 379374 447284 379380
rect 447138 379128 447194 379137
rect 447138 379063 447194 379072
rect 447244 378457 447272 379374
rect 447230 378448 447286 378457
rect 447230 378383 447286 378392
rect 447232 378140 447284 378146
rect 447232 378082 447284 378088
rect 447140 378072 447192 378078
rect 447140 378014 447192 378020
rect 447152 377777 447180 378014
rect 447138 377768 447194 377777
rect 447138 377703 447194 377712
rect 447244 377097 447272 378082
rect 447230 377088 447286 377097
rect 447230 377023 447286 377032
rect 447232 376712 447284 376718
rect 447232 376654 447284 376660
rect 447140 376644 447192 376650
rect 447140 376586 447192 376592
rect 447152 376417 447180 376586
rect 447138 376408 447194 376417
rect 447138 376343 447194 376352
rect 447244 375737 447272 376654
rect 447230 375728 447286 375737
rect 447230 375663 447286 375672
rect 447140 375352 447192 375358
rect 447140 375294 447192 375300
rect 447152 375057 447180 375294
rect 447232 375284 447284 375290
rect 447232 375226 447284 375232
rect 447138 375048 447194 375057
rect 447138 374983 447194 374992
rect 447244 374377 447272 375226
rect 447230 374368 447286 374377
rect 447230 374303 447286 374312
rect 447140 373992 447192 373998
rect 447140 373934 447192 373940
rect 447152 373697 447180 373934
rect 447232 373924 447284 373930
rect 447232 373866 447284 373872
rect 447138 373688 447194 373697
rect 447138 373623 447194 373632
rect 447244 373017 447272 373866
rect 447230 373008 447286 373017
rect 447230 372943 447286 372952
rect 447140 372564 447192 372570
rect 447140 372506 447192 372512
rect 447152 372337 447180 372506
rect 447232 372496 447284 372502
rect 447232 372438 447284 372444
rect 447138 372328 447194 372337
rect 447138 372263 447194 372272
rect 447244 371657 447272 372438
rect 447230 371648 447286 371657
rect 447230 371583 447286 371592
rect 447232 371204 447284 371210
rect 447232 371146 447284 371152
rect 447140 371136 447192 371142
rect 447140 371078 447192 371084
rect 447152 370977 447180 371078
rect 447138 370968 447194 370977
rect 447138 370903 447194 370912
rect 447244 370297 447272 371146
rect 447230 370288 447286 370297
rect 447230 370223 447286 370232
rect 447232 369844 447284 369850
rect 447232 369786 447284 369792
rect 447140 369776 447192 369782
rect 447140 369718 447192 369724
rect 447152 369617 447180 369718
rect 447138 369608 447194 369617
rect 447138 369543 447194 369552
rect 447244 368937 447272 369786
rect 447230 368928 447286 368937
rect 447230 368863 447286 368872
rect 447140 368484 447192 368490
rect 447140 368426 447192 368432
rect 447152 367577 447180 368426
rect 447232 368416 447284 368422
rect 447232 368358 447284 368364
rect 447244 368257 447272 368358
rect 447230 368248 447286 368257
rect 447230 368183 447286 368192
rect 447138 367568 447194 367577
rect 447138 367503 447194 367512
rect 447140 367056 447192 367062
rect 447140 366998 447192 367004
rect 447152 366897 447180 366998
rect 447232 366988 447284 366994
rect 447232 366930 447284 366936
rect 447138 366888 447194 366897
rect 447138 366823 447194 366832
rect 447244 366217 447272 366930
rect 447230 366208 447286 366217
rect 447230 366143 447286 366152
rect 447140 365696 447192 365702
rect 447140 365638 447192 365644
rect 447152 364857 447180 365638
rect 447232 365628 447284 365634
rect 447232 365570 447284 365576
rect 447244 365537 447272 365570
rect 447230 365528 447286 365537
rect 447230 365463 447286 365472
rect 447138 364848 447194 364857
rect 447138 364783 447194 364792
rect 447230 364168 447286 364177
rect 447230 364103 447286 364112
rect 447138 363488 447194 363497
rect 447138 363423 447194 363432
rect 447152 363050 447180 363423
rect 447140 363044 447192 363050
rect 447140 362986 447192 362992
rect 447244 362982 447272 364103
rect 447232 362976 447284 362982
rect 447232 362918 447284 362924
rect 447138 362808 447194 362817
rect 447138 362743 447194 362752
rect 447152 361622 447180 362743
rect 447230 362128 447286 362137
rect 447230 362063 447286 362072
rect 447244 361690 447272 362063
rect 447232 361684 447284 361690
rect 447232 361626 447284 361632
rect 447140 361616 447192 361622
rect 447140 361558 447192 361564
rect 447230 361448 447286 361457
rect 447230 361383 447286 361392
rect 447138 360768 447194 360777
rect 447138 360703 447194 360712
rect 447152 360262 447180 360703
rect 447244 360330 447272 361383
rect 447232 360324 447284 360330
rect 447232 360266 447284 360272
rect 447140 360256 447192 360262
rect 447140 360198 447192 360204
rect 447138 360088 447194 360097
rect 447138 360023 447194 360032
rect 447152 358834 447180 360023
rect 447230 359408 447286 359417
rect 447230 359343 447286 359352
rect 447244 358902 447272 359343
rect 447232 358896 447284 358902
rect 447232 358838 447284 358844
rect 447140 358828 447192 358834
rect 447140 358770 447192 358776
rect 447428 356017 447456 388418
rect 447600 387320 447652 387326
rect 447600 387262 447652 387268
rect 447414 356008 447470 356017
rect 447414 355943 447470 355952
rect 447612 353977 447640 387262
rect 447692 387252 447744 387258
rect 447692 387194 447744 387200
rect 447704 354657 447732 387194
rect 447796 387122 447824 669938
rect 447888 423026 447916 700266
rect 448428 447908 448480 447914
rect 448428 447850 448480 447856
rect 448060 447840 448112 447846
rect 448060 447782 448112 447788
rect 447968 447228 448020 447234
rect 447968 447170 448020 447176
rect 447876 423020 447928 423026
rect 447876 422962 447928 422968
rect 447784 387116 447836 387122
rect 447784 387058 447836 387064
rect 447876 385688 447928 385694
rect 447876 385630 447928 385636
rect 447690 354648 447746 354657
rect 447690 354583 447746 354592
rect 447598 353968 447654 353977
rect 447598 353903 447654 353912
rect 447888 353297 447916 385630
rect 447874 353288 447930 353297
rect 447874 353223 447930 353232
rect 447784 352708 447836 352714
rect 447784 352650 447836 352656
rect 447140 351960 447192 351966
rect 447138 351928 447140 351937
rect 447192 351928 447194 351937
rect 447138 351863 447194 351872
rect 447140 350600 447192 350606
rect 447138 350568 447140 350577
rect 447192 350568 447194 350577
rect 447138 350503 447194 350512
rect 447598 349888 447654 349897
rect 447598 349823 447654 349832
rect 447140 347744 447192 347750
rect 447140 347686 447192 347692
rect 447152 347177 447180 347686
rect 447138 347168 447194 347177
rect 447138 347103 447194 347112
rect 447230 341728 447286 341737
rect 447230 341663 447286 341672
rect 447138 341048 447194 341057
rect 447138 340983 447140 340992
rect 447192 340983 447194 340992
rect 447140 340954 447192 340960
rect 447244 340950 447272 341663
rect 447232 340944 447284 340950
rect 447232 340886 447284 340892
rect 447230 340368 447286 340377
rect 447230 340303 447286 340312
rect 447138 339688 447194 339697
rect 447138 339623 447194 339632
rect 447152 339590 447180 339623
rect 447140 339584 447192 339590
rect 447140 339526 447192 339532
rect 447244 339522 447272 340303
rect 447232 339516 447284 339522
rect 447232 339458 447284 339464
rect 447230 339008 447286 339017
rect 447230 338943 447286 338952
rect 447138 338328 447194 338337
rect 447138 338263 447194 338272
rect 447152 338230 447180 338263
rect 447140 338224 447192 338230
rect 447140 338166 447192 338172
rect 447244 338162 447272 338943
rect 447232 338156 447284 338162
rect 447232 338098 447284 338104
rect 447138 337648 447194 337657
rect 447138 337583 447194 337592
rect 447152 336530 447180 337583
rect 447324 337408 447376 337414
rect 447324 337350 447376 337356
rect 447230 336968 447286 336977
rect 447230 336903 447286 336912
rect 447140 336524 447192 336530
rect 447140 336466 447192 336472
rect 447138 336288 447194 336297
rect 447138 336223 447194 336232
rect 447152 335714 447180 336223
rect 447244 336122 447272 336903
rect 447232 336116 447284 336122
rect 447232 336058 447284 336064
rect 447140 335708 447192 335714
rect 447140 335650 447192 335656
rect 447138 335608 447194 335617
rect 447138 335543 447194 335552
rect 447152 335374 447180 335543
rect 447140 335368 447192 335374
rect 447140 335310 447192 335316
rect 447230 334928 447286 334937
rect 447230 334863 447286 334872
rect 447138 334248 447194 334257
rect 447138 334183 447194 334192
rect 447152 334014 447180 334183
rect 447244 334082 447272 334863
rect 447232 334076 447284 334082
rect 447232 334018 447284 334024
rect 447140 334008 447192 334014
rect 447140 333950 447192 333956
rect 447230 333568 447286 333577
rect 447230 333503 447286 333512
rect 447138 332888 447194 332897
rect 447138 332823 447194 332832
rect 447152 332654 447180 332823
rect 447244 332722 447272 333503
rect 447232 332716 447284 332722
rect 447232 332658 447284 332664
rect 447140 332648 447192 332654
rect 447140 332590 447192 332596
rect 447138 330168 447194 330177
rect 447138 330103 447140 330112
rect 447192 330103 447194 330112
rect 447140 330074 447192 330080
rect 447138 329488 447194 329497
rect 447138 329423 447194 329432
rect 447152 329118 447180 329423
rect 447140 329112 447192 329118
rect 447140 329054 447192 329060
rect 447046 322552 447102 322561
rect 447046 322487 447102 322496
rect 446956 320952 447008 320958
rect 446956 320894 447008 320900
rect 446864 319524 446916 319530
rect 446864 319466 446916 319472
rect 446772 319184 446824 319190
rect 446772 319126 446824 319132
rect 445668 318436 445720 318442
rect 445668 318378 445720 318384
rect 447336 316034 447364 337350
rect 447612 318782 447640 349823
rect 447796 330857 447824 352650
rect 447782 330848 447838 330857
rect 447782 330783 447838 330792
rect 447980 329497 448008 447170
rect 448072 330177 448100 447782
rect 448244 392692 448296 392698
rect 448244 392634 448296 392640
rect 448152 386028 448204 386034
rect 448152 385970 448204 385976
rect 448164 352617 448192 385970
rect 448256 355337 448284 392634
rect 448440 386646 448468 447850
rect 448980 387184 449032 387190
rect 448980 387126 449032 387132
rect 448428 386640 448480 386646
rect 448428 386582 448480 386588
rect 448336 385552 448388 385558
rect 448336 385494 448388 385500
rect 448242 355328 448298 355337
rect 448242 355263 448298 355272
rect 448150 352608 448206 352617
rect 448150 352543 448206 352552
rect 448242 351248 448298 351257
rect 448242 351183 448298 351192
rect 448150 332208 448206 332217
rect 448150 332143 448206 332152
rect 448058 330168 448114 330177
rect 448058 330103 448114 330112
rect 447966 329488 448022 329497
rect 447966 329423 448022 329432
rect 447600 318776 447652 318782
rect 447600 318718 447652 318724
rect 447152 316006 447364 316034
rect 443828 313948 443880 313954
rect 443828 313890 443880 313896
rect 447152 249762 447180 316006
rect 447784 260840 447836 260846
rect 447784 260782 447836 260788
rect 443736 249756 443788 249762
rect 443736 249698 443788 249704
rect 447140 249756 447192 249762
rect 447140 249698 447192 249704
rect 447152 248946 447180 249698
rect 446404 248940 446456 248946
rect 446404 248882 446456 248888
rect 447140 248940 447192 248946
rect 447140 248882 447192 248888
rect 443736 245676 443788 245682
rect 443736 245618 443788 245624
rect 443644 227724 443696 227730
rect 443644 227666 443696 227672
rect 443748 224126 443776 245618
rect 443736 224120 443788 224126
rect 443736 224062 443788 224068
rect 446416 163674 446444 248882
rect 447796 245682 447824 260782
rect 447784 245676 447836 245682
rect 447784 245618 447836 245624
rect 448164 183530 448192 332143
rect 448256 199442 448284 351183
rect 448348 348537 448376 385494
rect 448334 348528 448390 348537
rect 448334 348463 448390 348472
rect 448336 344752 448388 344758
rect 448336 344694 448388 344700
rect 448348 344457 448376 344694
rect 448334 344448 448390 344457
rect 448334 344383 448390 344392
rect 448440 343097 448468 386582
rect 448992 358737 449020 387126
rect 449070 387016 449126 387025
rect 449070 386951 449126 386960
rect 448978 358728 449034 358737
rect 448978 358663 449034 358672
rect 449084 357377 449112 386951
rect 449070 357368 449126 357377
rect 449070 357303 449126 357312
rect 448426 343088 448482 343097
rect 448426 343023 448482 343032
rect 448440 337414 448468 343023
rect 448428 337408 448480 337414
rect 448428 337350 448480 337356
rect 448334 331528 448390 331537
rect 448334 331463 448390 331472
rect 448244 199436 448296 199442
rect 448244 199378 448296 199384
rect 447600 183524 447652 183530
rect 447600 183466 447652 183472
rect 448152 183524 448204 183530
rect 448152 183466 448204 183472
rect 447612 182850 447640 183466
rect 447600 182844 447652 182850
rect 447600 182786 447652 182792
rect 447140 172508 447192 172514
rect 447140 172450 447192 172456
rect 447152 171834 447180 172450
rect 448348 171834 448376 331463
rect 448426 330848 448482 330857
rect 448426 330783 448482 330792
rect 447140 171828 447192 171834
rect 447140 171770 447192 171776
rect 448336 171828 448388 171834
rect 448336 171770 448388 171776
rect 448440 171134 448468 330783
rect 448520 322244 448572 322250
rect 448520 322186 448572 322192
rect 448532 319666 448560 322186
rect 449176 321434 449204 700538
rect 449268 321842 449296 700606
rect 462332 670002 462360 703520
rect 478524 700398 478552 703520
rect 478512 700392 478564 700398
rect 478512 700334 478564 700340
rect 494808 700330 494836 703520
rect 494796 700324 494848 700330
rect 494796 700266 494848 700272
rect 527192 699825 527220 703520
rect 543476 700369 543504 703520
rect 543462 700360 543518 700369
rect 543462 700295 543518 700304
rect 559668 699825 559696 703520
rect 527178 699816 527234 699825
rect 527178 699751 527234 699760
rect 559654 699816 559710 699825
rect 559654 699751 559710 699760
rect 580170 697232 580226 697241
rect 580170 697167 580226 697176
rect 580184 696998 580212 697167
rect 571984 696992 572036 696998
rect 571984 696934 572036 696940
rect 580172 696992 580224 696998
rect 580172 696934 580224 696940
rect 570604 670744 570656 670750
rect 570604 670686 570656 670692
rect 462320 669996 462372 670002
rect 462320 669938 462372 669944
rect 460202 668128 460258 668137
rect 460202 668063 460258 668072
rect 458086 659968 458142 659977
rect 458086 659903 458142 659912
rect 457810 657520 457866 657529
rect 457810 657455 457866 657464
rect 457718 652896 457774 652905
rect 457718 652831 457774 652840
rect 457626 650176 457682 650185
rect 457626 650111 457682 650120
rect 457534 645960 457590 645969
rect 457534 645895 457590 645904
rect 457442 643240 457498 643249
rect 457442 643175 457498 643184
rect 457350 623928 457406 623937
rect 457350 623863 457406 623872
rect 457258 621072 457314 621081
rect 457258 621007 457314 621016
rect 450544 596828 450596 596834
rect 450544 596770 450596 596776
rect 449808 518220 449860 518226
rect 449808 518162 449860 518168
rect 449820 503509 449848 518162
rect 450360 517540 450412 517546
rect 450360 517482 450412 517488
rect 449992 516792 450044 516798
rect 449992 516734 450044 516740
rect 450004 507657 450032 516734
rect 450372 510241 450400 517482
rect 450450 516896 450506 516905
rect 450450 516831 450506 516840
rect 450464 514729 450492 516831
rect 450450 514720 450506 514729
rect 450450 514655 450506 514664
rect 450556 512417 450584 596770
rect 457272 592686 457300 621007
rect 457364 596222 457392 623863
rect 457456 599622 457484 643175
rect 457444 599616 457496 599622
rect 457444 599558 457496 599564
rect 457548 598262 457576 645895
rect 457640 600642 457668 650111
rect 457628 600636 457680 600642
rect 457628 600578 457680 600584
rect 457732 600302 457760 652831
rect 457720 600296 457772 600302
rect 457720 600238 457772 600244
rect 457536 598256 457588 598262
rect 457536 598198 457588 598204
rect 457352 596216 457404 596222
rect 457352 596158 457404 596164
rect 457824 595474 457852 657455
rect 457994 635488 458050 635497
rect 457994 635423 458050 635432
rect 457902 618352 457958 618361
rect 457902 618287 457958 618296
rect 457812 595468 457864 595474
rect 457812 595410 457864 595416
rect 457260 592680 457312 592686
rect 457260 592622 457312 592628
rect 457916 520946 457944 618287
rect 457904 520940 457956 520946
rect 457904 520882 457956 520888
rect 458008 518294 458036 635423
rect 458100 519586 458128 659903
rect 459374 647728 459430 647737
rect 459374 647663 459430 647672
rect 459282 640384 459338 640393
rect 459282 640319 459338 640328
rect 459190 637936 459246 637945
rect 459190 637871 459246 637880
rect 459098 633448 459154 633457
rect 459098 633383 459154 633392
rect 459006 630728 459062 630737
rect 459006 630663 459062 630672
rect 458822 616040 458878 616049
rect 458822 615975 458878 615984
rect 458730 611416 458786 611425
rect 458730 611351 458786 611360
rect 458638 608696 458694 608705
rect 458638 608631 458694 608640
rect 458652 599758 458680 608631
rect 458640 599752 458692 599758
rect 458640 599694 458692 599700
rect 458744 598398 458772 611351
rect 458836 599690 458864 615975
rect 458914 614136 458970 614145
rect 458914 614071 458970 614080
rect 458824 599684 458876 599690
rect 458824 599626 458876 599632
rect 458732 598392 458784 598398
rect 458732 598334 458784 598340
rect 458928 596902 458956 614071
rect 458916 596896 458968 596902
rect 458916 596838 458968 596844
rect 459020 595649 459048 630663
rect 459112 598233 459140 633383
rect 459204 599593 459232 637871
rect 459190 599584 459246 599593
rect 459190 599519 459246 599528
rect 459098 598224 459154 598233
rect 459098 598159 459154 598168
rect 459006 595640 459062 595649
rect 459006 595575 459062 595584
rect 459296 589937 459324 640319
rect 459388 591297 459416 647663
rect 459466 628144 459522 628153
rect 459466 628079 459522 628088
rect 459374 591288 459430 591297
rect 459374 591223 459430 591232
rect 459282 589928 459338 589937
rect 459282 589863 459338 589872
rect 459480 544406 459508 628079
rect 460110 625832 460166 625841
rect 460110 625767 460166 625776
rect 460018 606384 460074 606393
rect 460018 606319 460074 606328
rect 459926 603664 459982 603673
rect 459926 603599 459982 603608
rect 459834 601896 459890 601905
rect 459834 601831 459890 601840
rect 459468 544400 459520 544406
rect 459468 544342 459520 544348
rect 458088 519580 458140 519586
rect 458088 519522 458140 519528
rect 459848 518430 459876 601831
rect 459940 597038 459968 603599
rect 460032 599894 460060 606319
rect 460020 599888 460072 599894
rect 460020 599830 460072 599836
rect 460124 598330 460152 625767
rect 460112 598324 460164 598330
rect 460112 598266 460164 598272
rect 459928 597032 459980 597038
rect 459928 596974 459980 596980
rect 460216 594454 460244 668063
rect 569224 616888 569276 616894
rect 569224 616830 569276 616836
rect 461584 600636 461636 600642
rect 461584 600578 461636 600584
rect 460204 594448 460256 594454
rect 460204 594390 460256 594396
rect 459836 518424 459888 518430
rect 459836 518366 459888 518372
rect 457996 518288 458048 518294
rect 457996 518230 458048 518236
rect 450636 516860 450688 516866
rect 450636 516802 450688 516808
rect 450542 512408 450598 512417
rect 450542 512343 450598 512352
rect 450358 510232 450414 510241
rect 450358 510167 450414 510176
rect 450372 509234 450400 510167
rect 450372 509206 450492 509234
rect 449990 507648 450046 507657
rect 449990 507583 450046 507592
rect 449806 503500 449862 503509
rect 449806 503435 449862 503444
rect 449808 464364 449860 464370
rect 449808 464306 449860 464312
rect 449716 461100 449768 461106
rect 449716 461042 449768 461048
rect 449624 454776 449676 454782
rect 449624 454718 449676 454724
rect 449532 454708 449584 454714
rect 449532 454650 449584 454656
rect 449440 387116 449492 387122
rect 449440 387058 449492 387064
rect 449348 385484 449400 385490
rect 449348 385426 449400 385432
rect 449360 347857 449388 385426
rect 449346 347848 449402 347857
rect 449346 347783 449402 347792
rect 449346 343768 449402 343777
rect 449346 343703 449402 343712
rect 449256 321836 449308 321842
rect 449256 321778 449308 321784
rect 449164 321428 449216 321434
rect 449164 321370 449216 321376
rect 448520 319660 448572 319666
rect 448520 319602 448572 319608
rect 449164 318776 449216 318782
rect 449164 318718 449216 318724
rect 448520 314152 448572 314158
rect 448520 314094 448572 314100
rect 448532 311166 448560 314094
rect 448520 311160 448572 311166
rect 448520 311102 448572 311108
rect 449176 263566 449204 318718
rect 449164 263560 449216 263566
rect 449164 263502 449216 263508
rect 448348 171106 448468 171134
rect 445208 163668 445260 163674
rect 445208 163610 445260 163616
rect 446404 163668 446456 163674
rect 446404 163610 446456 163616
rect 445220 161566 445248 163610
rect 445208 161560 445260 161566
rect 445208 161502 445260 161508
rect 441574 160132 441626 160138
rect 441574 160074 441626 160080
rect 442908 160132 442960 160138
rect 442908 160074 442960 160080
rect 441586 159868 441614 160074
rect 445220 159882 445248 161502
rect 448348 161430 448376 171106
rect 449360 164218 449388 343703
rect 449452 342417 449480 387058
rect 449544 358057 449572 454650
rect 449530 358048 449586 358057
rect 449530 357983 449586 357992
rect 449636 356697 449664 454718
rect 449622 356688 449678 356697
rect 449622 356623 449678 356632
rect 449728 346497 449756 461042
rect 449714 346488 449770 346497
rect 449714 346423 449770 346432
rect 449820 345817 449848 464306
rect 449806 345808 449862 345817
rect 449806 345743 449862 345752
rect 449806 345128 449862 345137
rect 449806 345063 449862 345072
rect 449438 342408 449494 342417
rect 449438 342343 449494 342352
rect 449440 336184 449492 336190
rect 449440 336126 449492 336132
rect 449452 319462 449480 336126
rect 449440 319456 449492 319462
rect 449440 319398 449492 319404
rect 449820 284986 449848 345063
rect 450004 333985 450032 507583
rect 450082 505472 450138 505481
rect 450082 505407 450138 505416
rect 450096 337482 450124 505407
rect 450174 503296 450230 503305
rect 450174 503231 450230 503240
rect 450084 337476 450136 337482
rect 450084 337418 450136 337424
rect 450188 336870 450216 503231
rect 450266 338056 450322 338065
rect 450266 337991 450322 338000
rect 450280 337113 450308 337991
rect 450360 337476 450412 337482
rect 450360 337418 450412 337424
rect 450266 337104 450322 337113
rect 450266 337039 450322 337048
rect 450176 336864 450228 336870
rect 450176 336806 450228 336812
rect 449990 333976 450046 333985
rect 449990 333911 450046 333920
rect 449898 328536 449954 328545
rect 449898 328471 449900 328480
rect 449952 328471 449954 328480
rect 449900 328442 449952 328448
rect 449898 327856 449954 327865
rect 449898 327791 449954 327800
rect 449912 327146 449940 327791
rect 449900 327140 449952 327146
rect 449900 327082 449952 327088
rect 450004 326233 450032 333911
rect 450084 330540 450136 330546
rect 450084 330482 450136 330488
rect 449990 326224 450046 326233
rect 449990 326159 450046 326168
rect 450096 324193 450124 330482
rect 450188 324442 450216 336806
rect 450280 327593 450308 337039
rect 450372 336938 450400 337418
rect 450360 336932 450412 336938
rect 450360 336874 450412 336880
rect 450266 327584 450322 327593
rect 450266 327519 450322 327528
rect 450372 325694 450400 336874
rect 450464 334393 450492 509206
rect 450556 462398 450584 512343
rect 450648 505481 450676 516802
rect 450634 505472 450690 505481
rect 450634 505407 450690 505416
rect 450648 500126 450754 500154
rect 451936 500126 452226 500154
rect 450544 462392 450596 462398
rect 450544 462334 450596 462340
rect 450556 338065 450584 462334
rect 450648 402974 450676 500126
rect 450648 402946 450860 402974
rect 450728 387388 450780 387394
rect 450728 387330 450780 387336
rect 450542 338056 450598 338065
rect 450542 337991 450598 338000
rect 450740 336802 450768 387330
rect 450832 385900 450860 402946
rect 451936 385914 451964 500126
rect 453304 497548 453356 497554
rect 453304 497490 453356 497496
rect 452568 496868 452620 496874
rect 452568 496810 452620 496816
rect 452016 455456 452068 455462
rect 452016 455398 452068 455404
rect 451582 385886 451964 385914
rect 452028 385558 452056 455398
rect 452580 385914 452608 496810
rect 453028 389156 453080 389162
rect 453028 389098 453080 389104
rect 452318 385886 452608 385914
rect 453040 385900 453068 389098
rect 453316 386034 453344 497490
rect 453684 496874 453712 500140
rect 454052 500126 455170 500154
rect 453672 496868 453724 496874
rect 453672 496810 453724 496816
rect 453948 496868 454000 496874
rect 453948 496810 454000 496816
rect 453304 386028 453356 386034
rect 453304 385970 453356 385976
rect 453960 385914 453988 496810
rect 454052 389162 454080 500126
rect 455328 497072 455380 497078
rect 455328 497014 455380 497020
rect 455144 496936 455196 496942
rect 455144 496878 455196 496884
rect 455156 393314 455184 496878
rect 455340 393314 455368 497014
rect 456524 497004 456576 497010
rect 456524 496946 456576 496952
rect 456536 393314 456564 496946
rect 456628 496874 456656 500140
rect 457628 497684 457680 497690
rect 457628 497626 457680 497632
rect 457444 497616 457496 497622
rect 457444 497558 457496 497564
rect 456616 496868 456668 496874
rect 456616 496810 456668 496816
rect 454880 393286 455184 393314
rect 455248 393286 455368 393314
rect 456352 393286 456564 393314
rect 454040 389156 454092 389162
rect 454040 389098 454092 389104
rect 454880 385914 454908 393286
rect 453790 385886 453988 385914
rect 454526 385886 454908 385914
rect 455248 385900 455276 393286
rect 456352 385914 456380 393286
rect 456708 389156 456760 389162
rect 456708 389098 456760 389104
rect 455998 385886 456380 385914
rect 456720 385900 456748 389098
rect 457456 387326 457484 497558
rect 457536 427100 457588 427106
rect 457536 427042 457588 427048
rect 457548 389162 457576 427042
rect 457536 389156 457588 389162
rect 457536 389098 457588 389104
rect 457444 387320 457496 387326
rect 457444 387262 457496 387268
rect 457640 386186 457668 497626
rect 458100 496942 458128 500140
rect 458824 497480 458876 497486
rect 458824 497422 458876 497428
rect 458088 496936 458140 496942
rect 458088 496878 458140 496884
rect 458088 429956 458140 429962
rect 458088 429898 458140 429904
rect 458100 393314 458128 429898
rect 457364 386158 457668 386186
rect 457824 393286 458128 393314
rect 457364 385694 457392 386158
rect 457824 385914 457852 393286
rect 458180 392760 458232 392766
rect 458180 392702 458232 392708
rect 457470 385886 457852 385914
rect 458192 385900 458220 392702
rect 458836 388482 458864 497422
rect 459572 497078 459600 500140
rect 459560 497072 459612 497078
rect 459560 497014 459612 497020
rect 461044 497010 461072 500140
rect 461032 497004 461084 497010
rect 461032 496946 461084 496952
rect 458916 460964 458968 460970
rect 458916 460906 458968 460912
rect 458928 447982 458956 460906
rect 460204 455524 460256 455530
rect 460204 455466 460256 455472
rect 458916 447976 458968 447982
rect 458916 447918 458968 447924
rect 459468 429888 459520 429894
rect 459468 429830 459520 429836
rect 459480 393314 459508 429830
rect 459296 393286 459508 393314
rect 458824 388476 458876 388482
rect 458824 388418 458876 388424
rect 459296 385914 459324 393286
rect 459652 388204 459704 388210
rect 459652 388146 459704 388152
rect 458942 385886 459324 385914
rect 459664 385900 459692 388146
rect 460216 387394 460244 455466
rect 461124 392624 461176 392630
rect 461124 392566 461176 392572
rect 460388 389156 460440 389162
rect 460388 389098 460440 389104
rect 460204 387388 460256 387394
rect 460204 387330 460256 387336
rect 460400 385900 460428 389098
rect 461136 385900 461164 392566
rect 461596 388550 461624 600578
rect 461676 600296 461728 600302
rect 461676 600238 461728 600244
rect 461688 388618 461716 600238
rect 463068 600086 463266 600114
rect 469614 600086 470088 600114
rect 475962 600086 476068 600114
rect 461766 597680 461822 597689
rect 461766 597615 461822 597624
rect 461676 388612 461728 388618
rect 461676 388554 461728 388560
rect 461584 388544 461636 388550
rect 461584 388486 461636 388492
rect 461780 388482 461808 597615
rect 462964 596216 463016 596222
rect 462964 596158 463016 596164
rect 462320 594448 462372 594454
rect 462320 594390 462372 594396
rect 461860 461032 461912 461038
rect 461860 460974 461912 460980
rect 461872 447846 461900 460974
rect 461952 454096 462004 454102
rect 461952 454038 462004 454044
rect 461964 447914 461992 454038
rect 461952 447908 462004 447914
rect 461952 447850 462004 447856
rect 461860 447840 461912 447846
rect 461860 447782 461912 447788
rect 462228 395344 462280 395350
rect 462228 395286 462280 395292
rect 461768 388476 461820 388482
rect 461768 388418 461820 388424
rect 462240 385914 462268 395286
rect 461886 385886 462268 385914
rect 462332 385914 462360 594390
rect 462412 518424 462464 518430
rect 462412 518366 462464 518372
rect 462424 402974 462452 518366
rect 462424 402946 462544 402974
rect 462516 386186 462544 402946
rect 462596 393984 462648 393990
rect 462596 393926 462648 393932
rect 462608 389162 462636 393926
rect 462780 389904 462832 389910
rect 462780 389846 462832 389852
rect 462596 389156 462648 389162
rect 462596 389098 462648 389104
rect 462792 388210 462820 389846
rect 462976 388414 463004 596158
rect 463068 501129 463096 600086
rect 463700 599888 463752 599894
rect 463700 599830 463752 599836
rect 463054 501120 463110 501129
rect 463054 501055 463110 501064
rect 463712 389298 463740 599830
rect 465080 599752 465132 599758
rect 465080 599694 465132 599700
rect 463792 597032 463844 597038
rect 463792 596974 463844 596980
rect 463700 389292 463752 389298
rect 463700 389234 463752 389240
rect 462964 388408 463016 388414
rect 462964 388350 463016 388356
rect 462780 388204 462832 388210
rect 462780 388146 462832 388152
rect 462516 386158 462912 386186
rect 462884 385914 462912 386158
rect 463804 385914 463832 596974
rect 464344 520328 464396 520334
rect 464344 520270 464396 520276
rect 464356 388385 464384 520270
rect 464436 497752 464488 497758
rect 464436 497694 464488 497700
rect 464448 392698 464476 497694
rect 464436 392692 464488 392698
rect 464436 392634 464488 392640
rect 464436 389292 464488 389298
rect 464436 389234 464488 389240
rect 464342 388376 464398 388385
rect 464342 388311 464398 388320
rect 464448 385914 464476 389234
rect 465092 385914 465120 599694
rect 466460 599684 466512 599690
rect 466460 599626 466512 599632
rect 465172 598392 465224 598398
rect 465172 598334 465224 598340
rect 465184 402974 465212 598334
rect 465724 592680 465776 592686
rect 465724 592622 465776 592628
rect 465184 402946 465672 402974
rect 465644 386050 465672 402946
rect 465736 388686 465764 592622
rect 465816 519580 465868 519586
rect 465816 519522 465868 519528
rect 465828 388958 465856 519522
rect 466472 389298 466500 599626
rect 469864 599616 469916 599622
rect 469864 599558 469916 599564
rect 468484 598256 468536 598262
rect 468484 598198 468536 598204
rect 466552 596896 466604 596902
rect 466552 596838 466604 596844
rect 466460 389292 466512 389298
rect 466460 389234 466512 389240
rect 465816 388952 465868 388958
rect 465816 388894 465868 388900
rect 465724 388680 465776 388686
rect 465724 388622 465776 388628
rect 465644 386022 465856 386050
rect 465828 385914 465856 386022
rect 466564 385914 466592 596838
rect 467932 520940 467984 520946
rect 467932 520882 467984 520888
rect 467102 518120 467158 518129
rect 467102 518055 467158 518064
rect 467116 388754 467144 518055
rect 467944 402974 467972 520882
rect 467944 402946 468064 402974
rect 467380 389292 467432 389298
rect 467380 389234 467432 389240
rect 467104 388748 467156 388754
rect 467104 388690 467156 388696
rect 467392 385914 467420 389234
rect 468036 385914 468064 402946
rect 468496 388890 468524 598198
rect 468576 595468 468628 595474
rect 468576 595410 468628 595416
rect 468484 388884 468536 388890
rect 468484 388826 468536 388832
rect 468588 388822 468616 595410
rect 468668 497820 468720 497826
rect 468668 497762 468720 497768
rect 468576 388816 468628 388822
rect 468576 388758 468628 388764
rect 468680 387258 468708 497762
rect 469876 388958 469904 599558
rect 469956 518288 470008 518294
rect 469956 518230 470008 518236
rect 469968 389026 469996 518230
rect 470060 518226 470088 600086
rect 470600 598324 470652 598330
rect 470600 598266 470652 598272
rect 470048 518220 470100 518226
rect 470048 518162 470100 518168
rect 469956 389020 470008 389026
rect 469956 388962 470008 388968
rect 469404 388952 469456 388958
rect 469404 388894 469456 388900
rect 469864 388952 469916 388958
rect 469864 388894 469916 388900
rect 469416 388754 469444 388894
rect 469404 388748 469456 388754
rect 469404 388690 469456 388696
rect 469220 388680 469272 388686
rect 469220 388622 469272 388628
rect 468668 387252 468720 387258
rect 468668 387194 468720 387200
rect 462332 385886 462622 385914
rect 462884 385886 463358 385914
rect 463804 385886 464094 385914
rect 464448 385886 464830 385914
rect 465092 385886 465566 385914
rect 465828 385886 466302 385914
rect 466564 385886 467038 385914
rect 467392 385886 467774 385914
rect 468036 385886 468510 385914
rect 469232 385900 469260 388622
rect 469956 388408 470008 388414
rect 469956 388350 470008 388356
rect 469968 385900 469996 388350
rect 470612 385914 470640 598266
rect 470876 544400 470928 544406
rect 470876 544342 470928 544348
rect 470888 402974 470916 544342
rect 476040 517614 476068 600086
rect 476028 517608 476080 517614
rect 476028 517550 476080 517556
rect 476040 516866 476068 517550
rect 482296 517478 482324 600100
rect 488644 598262 488672 600100
rect 488632 598256 488684 598262
rect 488632 598198 488684 598204
rect 494060 598256 494112 598262
rect 494060 598198 494112 598204
rect 482928 520940 482980 520946
rect 482928 520882 482980 520888
rect 482742 517576 482798 517585
rect 482940 517562 482968 520882
rect 488632 520328 488684 520334
rect 488632 520270 488684 520276
rect 488644 517970 488672 520270
rect 488644 517942 488980 517970
rect 482798 517534 483000 517562
rect 494072 517546 494100 598198
rect 494992 596834 495020 600100
rect 500972 600086 501354 600114
rect 507136 600086 507702 600114
rect 513392 600086 514050 600114
rect 520292 600086 520398 600114
rect 525812 600086 526746 600114
rect 494980 596828 495032 596834
rect 494980 596770 495032 596776
rect 494244 518220 494296 518226
rect 494244 518162 494296 518168
rect 494152 517608 494204 517614
rect 494152 517550 494204 517556
rect 494060 517540 494112 517546
rect 482742 517511 482798 517520
rect 494060 517482 494112 517488
rect 482284 517472 482336 517478
rect 482284 517414 482336 517420
rect 476028 516860 476080 516866
rect 476028 516802 476080 516808
rect 492128 516792 492180 516798
rect 492128 516734 492180 516740
rect 492140 512650 492168 516734
rect 494072 515545 494100 517482
rect 494058 515536 494114 515545
rect 494058 515471 494114 515480
rect 492128 512644 492180 512650
rect 492128 512586 492180 512592
rect 492140 512485 492168 512586
rect 492126 512476 492182 512485
rect 492126 512411 492182 512420
rect 494072 509930 494100 515471
rect 494060 509924 494112 509930
rect 494060 509866 494112 509872
rect 494164 508881 494192 517550
rect 494150 508872 494206 508881
rect 494150 508807 494206 508816
rect 494164 508570 494192 508807
rect 494152 508564 494204 508570
rect 494152 508506 494204 508512
rect 494256 505753 494284 518162
rect 500972 516905 501000 600086
rect 500958 516896 501014 516905
rect 500958 516831 501014 516840
rect 502246 516896 502302 516905
rect 502246 516831 502302 516840
rect 502260 514078 502288 516831
rect 507136 516769 507164 600086
rect 507122 516760 507178 516769
rect 507122 516695 507178 516704
rect 502248 514072 502300 514078
rect 502248 514014 502300 514020
rect 495072 505776 495124 505782
rect 494242 505744 494298 505753
rect 494242 505679 494298 505688
rect 495070 505744 495072 505753
rect 495124 505744 495126 505753
rect 495070 505679 495126 505688
rect 494702 501256 494758 501265
rect 494702 501191 494758 501200
rect 480272 500126 480608 500154
rect 481652 500126 481804 500154
rect 482664 500126 483000 500154
rect 483860 500126 484196 500154
rect 485056 500126 485392 500154
rect 486252 500126 486588 500154
rect 487172 500126 487784 500154
rect 488980 500126 489224 500154
rect 480272 497554 480300 500126
rect 481652 497690 481680 500126
rect 481640 497684 481692 497690
rect 481640 497626 481692 497632
rect 482664 497622 482692 500126
rect 483860 497826 483888 500126
rect 483848 497820 483900 497826
rect 483848 497762 483900 497768
rect 485056 497758 485084 500126
rect 485044 497752 485096 497758
rect 485044 497694 485096 497700
rect 482652 497616 482704 497622
rect 482652 497558 482704 497564
rect 480260 497548 480312 497554
rect 480260 497490 480312 497496
rect 486252 497486 486280 500126
rect 486240 497480 486292 497486
rect 486240 497422 486292 497428
rect 473726 462904 473782 462913
rect 473726 462839 473782 462848
rect 473740 454102 473768 462839
rect 480996 455456 481048 455462
rect 480996 455398 481048 455404
rect 473728 454096 473780 454102
rect 473728 454038 473780 454044
rect 473740 453900 473768 454038
rect 481008 453900 481036 455398
rect 487172 454782 487200 500126
rect 489196 496913 489224 500126
rect 489932 500126 490176 500154
rect 491312 500126 491372 500154
rect 489182 496904 489238 496913
rect 489182 496839 489238 496848
rect 488264 456068 488316 456074
rect 488264 456010 488316 456016
rect 488276 455530 488304 456010
rect 488264 455524 488316 455530
rect 488264 455466 488316 455472
rect 487160 454776 487212 454782
rect 487160 454718 487212 454724
rect 488276 453900 488304 455466
rect 489932 454714 489960 500126
rect 489920 454708 489972 454714
rect 489920 454650 489972 454656
rect 471624 427106 471652 432140
rect 474292 429962 474320 432140
rect 474280 429956 474332 429962
rect 474280 429898 474332 429904
rect 476960 429214 476988 432140
rect 479628 429894 479656 432140
rect 481652 432126 482310 432154
rect 484412 432126 484978 432154
rect 487172 432126 487646 432154
rect 489932 432126 490314 432154
rect 479616 429888 479668 429894
rect 479616 429830 479668 429836
rect 475384 429208 475436 429214
rect 475384 429150 475436 429156
rect 476948 429208 477000 429214
rect 476948 429150 477000 429156
rect 471612 427100 471664 427106
rect 471612 427042 471664 427048
rect 470888 402946 471008 402974
rect 470980 385914 471008 402946
rect 475396 392766 475424 429150
rect 475384 392760 475436 392766
rect 475384 392702 475436 392708
rect 481652 389910 481680 432126
rect 484308 423428 484360 423434
rect 484308 423370 484360 423376
rect 484216 421592 484268 421598
rect 484216 421534 484268 421540
rect 484228 393314 484256 421534
rect 483584 393286 484256 393314
rect 481640 389904 481692 389910
rect 481640 389846 481692 389852
rect 472162 389056 472218 389065
rect 474370 389056 474426 389065
rect 472162 388991 472218 389000
rect 473636 389020 473688 389026
rect 470612 385886 470718 385914
rect 470980 385886 471454 385914
rect 472176 385900 472204 388991
rect 474370 388991 474426 389000
rect 475106 389056 475162 389065
rect 475106 388991 475162 389000
rect 477314 389056 477370 389065
rect 477314 388991 477370 389000
rect 479522 389056 479578 389065
rect 479522 388991 479578 389000
rect 473636 388962 473688 388968
rect 472898 388920 472954 388929
rect 472898 388855 472954 388864
rect 472912 385900 472940 388855
rect 473648 385900 473676 388962
rect 474384 385900 474412 388991
rect 475120 385900 475148 388991
rect 475844 388952 475896 388958
rect 475844 388894 475896 388900
rect 475856 385900 475884 388894
rect 476580 388884 476632 388890
rect 476580 388826 476632 388832
rect 476592 385900 476620 388826
rect 477328 385900 477356 388991
rect 478788 388612 478840 388618
rect 478788 388554 478840 388560
rect 478052 388544 478104 388550
rect 478052 388486 478104 388492
rect 478064 385900 478092 388486
rect 478800 385900 478828 388554
rect 479536 385900 479564 388991
rect 480260 388816 480312 388822
rect 480260 388758 480312 388764
rect 480272 385900 480300 388758
rect 480996 388748 481048 388754
rect 480996 388690 481048 388696
rect 481008 385900 481036 388690
rect 481732 388680 481784 388686
rect 481732 388622 481784 388628
rect 481744 385900 481772 388622
rect 482468 388476 482520 388482
rect 482468 388418 482520 388424
rect 482480 385900 482508 388418
rect 483584 385914 483612 393286
rect 484320 385914 484348 423370
rect 484412 393990 484440 432126
rect 487068 423360 487120 423366
rect 487068 423302 487120 423308
rect 486976 416084 487028 416090
rect 486976 416026 487028 416032
rect 484400 393984 484452 393990
rect 484400 393926 484452 393932
rect 486988 393314 487016 416026
rect 486896 393286 487016 393314
rect 486424 389292 486476 389298
rect 486424 389234 486476 389240
rect 484676 388816 484728 388822
rect 484676 388758 484728 388764
rect 483230 385886 483612 385914
rect 483966 385886 484348 385914
rect 484688 385900 484716 388758
rect 485412 388612 485464 388618
rect 485412 388554 485464 388560
rect 485424 385900 485452 388554
rect 486436 385914 486464 389234
rect 486174 385886 486464 385914
rect 486896 385900 486924 393286
rect 487080 389298 487108 423302
rect 487172 392630 487200 432126
rect 488264 423292 488316 423298
rect 488264 423234 488316 423240
rect 488276 393314 488304 423234
rect 489644 423224 489696 423230
rect 489644 423166 489696 423172
rect 489656 393314 489684 423166
rect 489932 395350 489960 432126
rect 489920 395344 489972 395350
rect 489920 395286 489972 395292
rect 488000 393286 488304 393314
rect 489472 393286 489684 393314
rect 487160 392624 487212 392630
rect 487160 392566 487212 392572
rect 487068 389292 487120 389298
rect 487068 389234 487120 389240
rect 488000 385914 488028 393286
rect 488356 388476 488408 388482
rect 488356 388418 488408 388424
rect 487646 385886 488028 385914
rect 488368 385900 488396 388418
rect 489472 385914 489500 393286
rect 490564 392624 490616 392630
rect 490564 392566 490616 392572
rect 489828 388544 489880 388550
rect 489828 388486 489880 388492
rect 489118 385886 489500 385914
rect 489840 385900 489868 388486
rect 490576 385900 490604 392566
rect 491312 387190 491340 500126
rect 494716 462466 494744 501191
rect 494704 462460 494756 462466
rect 494704 462402 494756 462408
rect 494716 456074 494744 462402
rect 494704 456068 494756 456074
rect 494704 456010 494756 456016
rect 503628 424380 503680 424386
rect 503628 424322 503680 424328
rect 502984 423564 503036 423570
rect 502984 423506 503036 423512
rect 498108 423156 498160 423162
rect 498108 423098 498160 423104
rect 495348 420232 495400 420238
rect 495348 420174 495400 420180
rect 494612 398132 494664 398138
rect 494612 398074 494664 398080
rect 493968 396772 494020 396778
rect 493968 396714 494020 396720
rect 493140 395344 493192 395350
rect 493140 395286 493192 395292
rect 491668 393984 491720 393990
rect 491668 393926 491720 393932
rect 491300 387184 491352 387190
rect 491300 387126 491352 387132
rect 491680 385914 491708 393926
rect 492036 389904 492088 389910
rect 492036 389846 492088 389852
rect 491326 385886 491708 385914
rect 492048 385900 492076 389846
rect 493152 385914 493180 395286
rect 493980 385914 494008 396714
rect 494624 385914 494652 398074
rect 495360 385914 495388 420174
rect 497924 400920 497976 400926
rect 497924 400862 497976 400868
rect 496728 399492 496780 399498
rect 496728 399434 496780 399440
rect 495716 391332 495768 391338
rect 495716 391274 495768 391280
rect 492798 385886 493180 385914
rect 493534 385886 494008 385914
rect 494270 385886 494652 385914
rect 495006 385886 495388 385914
rect 495728 385900 495756 391274
rect 496740 385914 496768 399434
rect 497464 389292 497516 389298
rect 497464 389234 497516 389240
rect 497476 385914 497504 389234
rect 496478 385886 496768 385914
rect 497214 385886 497504 385914
rect 497936 385900 497964 400862
rect 498120 389298 498148 423098
rect 499304 423088 499356 423094
rect 499304 423030 499356 423036
rect 499316 393314 499344 423030
rect 500684 423020 500736 423026
rect 500684 422962 500736 422968
rect 500696 393314 500724 422962
rect 502248 422952 502300 422958
rect 502248 422894 502300 422900
rect 502260 393314 502288 422894
rect 499040 393286 499344 393314
rect 500512 393286 500724 393314
rect 501984 393286 502288 393314
rect 498108 389292 498160 389298
rect 498108 389234 498160 389240
rect 499040 385914 499068 393286
rect 499396 388680 499448 388686
rect 499396 388622 499448 388628
rect 498686 385886 499068 385914
rect 499408 385900 499436 388622
rect 500512 385914 500540 393286
rect 500868 388748 500920 388754
rect 500868 388690 500920 388696
rect 500158 385886 500540 385914
rect 500880 385900 500908 388690
rect 501984 385914 502012 393286
rect 502340 388952 502392 388958
rect 502340 388894 502392 388900
rect 501630 385886 502012 385914
rect 502352 385900 502380 388894
rect 502996 388822 503024 423506
rect 503640 393314 503668 424322
rect 507860 417784 507912 417790
rect 507860 417726 507912 417732
rect 506480 417716 506532 417722
rect 506480 417658 506532 417664
rect 503996 417648 504048 417654
rect 503996 417590 504048 417596
rect 503720 417580 503772 417586
rect 503720 417522 503772 417528
rect 503456 393286 503668 393314
rect 502984 388816 503036 388822
rect 502984 388758 503036 388764
rect 503456 385914 503484 393286
rect 503102 385886 503484 385914
rect 503732 385914 503760 417522
rect 504008 402974 504036 417590
rect 504008 402946 504128 402974
rect 504100 385914 504128 402946
rect 506020 391264 506072 391270
rect 506020 391206 506072 391212
rect 505284 389836 505336 389842
rect 505284 389778 505336 389784
rect 503732 385886 503838 385914
rect 504100 385886 504574 385914
rect 505296 385900 505324 389778
rect 506032 385900 506060 391206
rect 506492 389298 506520 417658
rect 506572 417512 506624 417518
rect 506572 417454 506624 417460
rect 506480 389292 506532 389298
rect 506480 389234 506532 389240
rect 506584 385914 506612 417454
rect 507124 389292 507176 389298
rect 507124 389234 507176 389240
rect 507136 385914 507164 389234
rect 507872 385914 507900 417726
rect 507952 417444 508004 417450
rect 507952 417386 508004 417392
rect 507964 402974 507992 417386
rect 511264 404388 511316 404394
rect 511264 404330 511316 404336
rect 507964 402946 508544 402974
rect 508516 385914 508544 402946
rect 506584 385886 506782 385914
rect 507136 385886 507518 385914
rect 507872 385886 508254 385914
rect 508516 385886 508990 385914
rect 457352 385688 457404 385694
rect 457352 385630 457404 385636
rect 452016 385552 452068 385558
rect 452016 385494 452068 385500
rect 509698 370152 509754 370161
rect 509698 370087 509754 370096
rect 450728 336796 450780 336802
rect 450728 336738 450780 336744
rect 450450 334384 450506 334393
rect 450450 334319 450506 334328
rect 450464 326913 450492 334319
rect 450740 330546 450768 336738
rect 450728 330540 450780 330546
rect 450728 330482 450780 330488
rect 450450 326904 450506 326913
rect 450450 326839 450506 326848
rect 509712 326346 509740 370087
rect 509882 360360 509938 360369
rect 509882 360295 509938 360304
rect 509792 349852 509844 349858
rect 509792 349794 509844 349800
rect 509804 326466 509832 349794
rect 509792 326460 509844 326466
rect 509792 326402 509844 326408
rect 509712 326318 509832 326346
rect 450372 325666 450492 325694
rect 450464 325553 450492 325666
rect 450450 325544 450506 325553
rect 450450 325479 450506 325488
rect 450358 324456 450414 324465
rect 450188 324414 450358 324442
rect 450358 324391 450414 324400
rect 450082 324184 450138 324193
rect 450082 324119 450138 324128
rect 450372 288930 450400 324391
rect 450360 288924 450412 288930
rect 450360 288866 450412 288872
rect 449808 284980 449860 284986
rect 449808 284922 449860 284928
rect 450464 269822 450492 325479
rect 450634 323776 450690 323785
rect 450634 323711 450690 323720
rect 450648 318102 450676 323711
rect 509698 322960 509754 322969
rect 509698 322895 509754 322904
rect 471058 322688 471114 322697
rect 471058 322623 471114 322632
rect 482374 322688 482430 322697
rect 482374 322623 482430 322632
rect 471886 322552 471942 322561
rect 471886 322487 471942 322496
rect 459190 322416 459246 322425
rect 459190 322351 459246 322360
rect 454558 321910 454586 322116
rect 454546 321904 454598 321910
rect 454546 321846 454598 321852
rect 450636 318096 450688 318102
rect 450636 318038 450688 318044
rect 453304 316872 453356 316878
rect 453304 316814 453356 316820
rect 450544 316736 450596 316742
rect 450544 316678 450596 316684
rect 450452 269816 450504 269822
rect 450452 269758 450504 269764
rect 449900 268592 449952 268598
rect 449900 268534 449952 268540
rect 449912 263650 449940 268534
rect 449820 263622 449940 263650
rect 449820 260846 449848 263622
rect 449808 260840 449860 260846
rect 449808 260782 449860 260788
rect 448428 164212 448480 164218
rect 448428 164154 448480 164160
rect 449348 164212 449400 164218
rect 449348 164154 449400 164160
rect 448336 161424 448388 161430
rect 448336 161366 448388 161372
rect 448348 160750 448376 161366
rect 448336 160744 448388 160750
rect 448336 160686 448388 160692
rect 448440 159882 448468 164154
rect 444912 159854 445248 159882
rect 448224 159854 448468 159882
rect 437992 159468 438624 159474
rect 437940 159462 438624 159468
rect 437952 159446 438624 159462
rect 421392 159310 421880 159338
rect 425152 159384 425204 159390
rect 425152 159326 425204 159332
rect 409880 158024 409932 158030
rect 409880 157966 409932 157972
rect 409512 150408 409564 150414
rect 409512 150350 409564 150356
rect 409420 139392 409472 139398
rect 409420 139334 409472 139340
rect 409328 128308 409380 128314
rect 409328 128250 409380 128256
rect 409236 117292 409288 117298
rect 409236 117234 409288 117240
rect 439136 107296 439188 107302
rect 439136 107238 439188 107244
rect 432972 107228 433024 107234
rect 432972 107170 433024 107176
rect 426808 107160 426860 107166
rect 426808 107102 426860 107108
rect 420644 107092 420696 107098
rect 420644 107034 420696 107040
rect 414480 107024 414532 107030
rect 414480 106966 414532 106972
rect 409144 106276 409196 106282
rect 409144 106218 409196 106224
rect 414492 104938 414520 106966
rect 420656 104938 420684 107034
rect 426820 104938 426848 107102
rect 432984 104938 433012 107170
rect 439148 104938 439176 107238
rect 450556 107234 450584 316678
rect 450636 315308 450688 315314
rect 450636 315250 450688 315256
rect 450544 107228 450596 107234
rect 450544 107170 450596 107176
rect 450648 107098 450676 315250
rect 452016 314084 452068 314090
rect 452016 314026 452068 314032
rect 450728 314016 450780 314022
rect 450728 313958 450780 313964
rect 450740 107166 450768 313958
rect 450820 311228 450872 311234
rect 450820 311170 450872 311176
rect 450832 107302 450860 311170
rect 451924 308508 451976 308514
rect 451924 308450 451976 308456
rect 451188 287700 451240 287706
rect 451188 287642 451240 287648
rect 450912 268388 450964 268394
rect 450912 268330 450964 268336
rect 450820 107296 450872 107302
rect 450820 107238 450872 107244
rect 450728 107160 450780 107166
rect 450728 107102 450780 107108
rect 450636 107092 450688 107098
rect 450636 107034 450688 107040
rect 450924 106554 450952 268330
rect 451004 161560 451056 161566
rect 451004 161502 451056 161508
rect 451016 142186 451044 161502
rect 451004 142180 451056 142186
rect 451004 142122 451056 142128
rect 451016 106962 451044 142122
rect 451004 106956 451056 106962
rect 451004 106898 451056 106904
rect 445300 106548 445352 106554
rect 445300 106490 445352 106496
rect 450912 106548 450964 106554
rect 450912 106490 450964 106496
rect 445312 104938 445340 106490
rect 451200 104938 451228 287642
rect 451740 158704 451792 158710
rect 451740 158646 451792 158652
rect 451752 158273 451780 158646
rect 451738 158264 451794 158273
rect 451738 158199 451794 158208
rect 451740 157344 451792 157350
rect 451740 157286 451792 157292
rect 451752 156913 451780 157286
rect 451738 156904 451794 156913
rect 451738 156839 451794 156848
rect 451832 146260 451884 146266
rect 451832 146202 451884 146208
rect 451844 146033 451872 146202
rect 451830 146024 451886 146033
rect 451830 145959 451886 145968
rect 451556 144832 451608 144838
rect 451556 144774 451608 144780
rect 451568 144673 451596 144774
rect 451554 144664 451610 144673
rect 451554 144599 451610 144608
rect 451556 139256 451608 139262
rect 451554 139224 451556 139233
rect 451608 139224 451610 139233
rect 451554 139159 451610 139168
rect 451556 136536 451608 136542
rect 451554 136504 451556 136513
rect 451608 136504 451610 136513
rect 451554 136439 451610 136448
rect 451936 128353 451964 308450
rect 452028 148753 452056 314026
rect 452200 311296 452252 311302
rect 452200 311238 452252 311244
rect 452108 286680 452160 286686
rect 452108 286622 452160 286628
rect 452014 148744 452070 148753
rect 452014 148679 452070 148688
rect 452016 135176 452068 135182
rect 452014 135144 452016 135153
rect 452068 135144 452070 135153
rect 452014 135079 452070 135088
rect 452120 132494 452148 286622
rect 452212 155553 452240 311238
rect 452384 280900 452436 280906
rect 452384 280842 452436 280848
rect 452292 271244 452344 271250
rect 452292 271186 452344 271192
rect 452198 155544 452254 155553
rect 452198 155479 452254 155488
rect 452304 133793 452332 271186
rect 452396 150113 452424 280842
rect 452476 154488 452528 154494
rect 452476 154430 452528 154436
rect 452488 154193 452516 154430
rect 452474 154184 452530 154193
rect 452474 154119 452530 154128
rect 452476 152992 452528 152998
rect 452476 152934 452528 152940
rect 452488 152833 452516 152934
rect 452474 152824 452530 152833
rect 452474 152759 452530 152768
rect 452568 151496 452620 151502
rect 452566 151464 452568 151473
rect 452620 151464 452622 151473
rect 452566 151399 452622 151408
rect 452382 150104 452438 150113
rect 452382 150039 452438 150048
rect 452568 147416 452620 147422
rect 452566 147384 452568 147393
rect 452620 147384 452622 147393
rect 452566 147319 452622 147328
rect 452568 143472 452620 143478
rect 452568 143414 452620 143420
rect 452580 143313 452608 143414
rect 452566 143304 452622 143313
rect 452566 143239 452622 143248
rect 452568 141976 452620 141982
rect 452566 141944 452568 141953
rect 452620 141944 452622 141953
rect 452566 141879 452622 141888
rect 452568 140752 452620 140758
rect 452568 140694 452620 140700
rect 452580 140593 452608 140694
rect 452566 140584 452622 140593
rect 452566 140519 452622 140528
rect 452568 137896 452620 137902
rect 452566 137864 452568 137873
rect 452620 137864 452622 137873
rect 452566 137799 452622 137808
rect 452290 133784 452346 133793
rect 452290 133719 452346 133728
rect 452028 132466 452148 132494
rect 451922 128344 451978 128353
rect 451922 128279 451978 128288
rect 451740 126812 451792 126818
rect 451740 126754 451792 126760
rect 451752 125633 451780 126754
rect 451738 125624 451794 125633
rect 451738 125559 451794 125568
rect 452028 124273 452056 132466
rect 452292 132456 452344 132462
rect 452290 132424 452292 132433
rect 452344 132424 452346 132433
rect 452290 132359 452346 132368
rect 452568 131096 452620 131102
rect 452566 131064 452568 131073
rect 452620 131064 452622 131073
rect 452566 130999 452622 131008
rect 453316 129742 453344 316814
rect 454684 316804 454736 316810
rect 454684 316746 454736 316752
rect 453396 315376 453448 315382
rect 453396 315318 453448 315324
rect 453408 132462 453436 315318
rect 453580 283688 453632 283694
rect 453580 283630 453632 283636
rect 453488 275392 453540 275398
rect 453488 275334 453540 275340
rect 453396 132456 453448 132462
rect 453396 132398 453448 132404
rect 452108 129736 452160 129742
rect 452106 129704 452108 129713
rect 453304 129736 453356 129742
rect 452160 129704 452162 129713
rect 453304 129678 453356 129684
rect 452106 129639 452162 129648
rect 452566 126984 452622 126993
rect 452566 126919 452568 126928
rect 452620 126919 452622 126928
rect 452568 126890 452620 126896
rect 453500 126818 453528 275334
rect 453592 154494 453620 283630
rect 453672 279472 453724 279478
rect 453672 279414 453724 279420
rect 453580 154488 453632 154494
rect 453580 154430 453632 154436
rect 453684 152998 453712 279414
rect 453672 152992 453724 152998
rect 453672 152934 453724 152940
rect 453488 126812 453540 126818
rect 453488 126754 453540 126760
rect 452014 124264 452070 124273
rect 452014 124199 452070 124208
rect 451740 123140 451792 123146
rect 451740 123082 451792 123088
rect 451752 122913 451780 123082
rect 451738 122904 451794 122913
rect 451738 122839 451794 122848
rect 451924 122052 451976 122058
rect 451924 121994 451976 122000
rect 451936 121553 451964 121994
rect 451922 121544 451978 121553
rect 451922 121479 451978 121488
rect 454696 107030 454724 316746
rect 454788 296002 454816 322116
rect 454960 321904 455012 321910
rect 454960 321846 455012 321852
rect 454972 298110 455000 321846
rect 454960 298104 455012 298110
rect 454960 298046 455012 298052
rect 454776 295996 454828 296002
rect 454776 295938 454828 295944
rect 455064 294438 455092 322116
rect 455236 313948 455288 313954
rect 455236 313890 455288 313896
rect 455052 294432 455104 294438
rect 455052 294374 455104 294380
rect 454960 290556 455012 290562
rect 454960 290498 455012 290504
rect 454868 275324 454920 275330
rect 454868 275266 454920 275272
rect 454776 272604 454828 272610
rect 454776 272546 454828 272552
rect 454788 123146 454816 272546
rect 454880 140758 454908 275266
rect 454972 158710 455000 290498
rect 455144 288924 455196 288930
rect 455144 288866 455196 288872
rect 455052 285048 455104 285054
rect 455052 284990 455104 284996
rect 454960 158704 455012 158710
rect 454960 158646 455012 158652
rect 455064 157350 455092 284990
rect 455156 222154 455184 288866
rect 455248 258738 455276 313890
rect 455340 288930 455368 322116
rect 455616 313886 455644 322116
rect 455604 313880 455656 313886
rect 455604 313822 455656 313828
rect 455892 307154 455920 322116
rect 456062 318064 456118 318073
rect 456062 317999 456118 318008
rect 455880 307148 455932 307154
rect 455880 307090 455932 307096
rect 455328 288924 455380 288930
rect 455328 288866 455380 288872
rect 455236 258732 455288 258738
rect 455236 258674 455288 258680
rect 455144 222148 455196 222154
rect 455144 222090 455196 222096
rect 455052 157344 455104 157350
rect 455052 157286 455104 157292
rect 454868 140752 454920 140758
rect 454868 140694 454920 140700
rect 454776 123140 454828 123146
rect 454776 123082 454828 123088
rect 456076 119406 456104 317999
rect 456168 291718 456196 322116
rect 456444 316062 456472 322116
rect 456720 321230 456748 322116
rect 456708 321224 456760 321230
rect 456708 321166 456760 321172
rect 456996 321162 457024 322116
rect 456984 321156 457036 321162
rect 456984 321098 457036 321104
rect 457272 318782 457300 322116
rect 457548 320890 457576 322116
rect 457824 321638 457852 322116
rect 457812 321632 457864 321638
rect 457812 321574 457864 321580
rect 457536 320884 457588 320890
rect 457536 320826 457588 320832
rect 457260 318776 457312 318782
rect 457260 318718 457312 318724
rect 458100 318714 458128 322116
rect 458376 321570 458404 322116
rect 458364 321564 458416 321570
rect 458364 321506 458416 321512
rect 458652 320657 458680 322116
rect 458638 320648 458694 320657
rect 458638 320583 458694 320592
rect 458928 319938 458956 322116
rect 459480 321502 459508 322116
rect 459468 321496 459520 321502
rect 459468 321438 459520 321444
rect 458916 319932 458968 319938
rect 458916 319874 458968 319880
rect 459756 319841 459784 322116
rect 460032 321366 460060 322116
rect 460020 321360 460072 321366
rect 460020 321302 460072 321308
rect 460308 321298 460336 322116
rect 460584 321473 460612 322116
rect 460570 321464 460626 321473
rect 460570 321399 460626 321408
rect 460860 321337 460888 322116
rect 460846 321328 460902 321337
rect 460296 321292 460348 321298
rect 460846 321263 460902 321272
rect 460296 321234 460348 321240
rect 461136 320754 461164 322116
rect 461124 320748 461176 320754
rect 461124 320690 461176 320696
rect 461412 320686 461440 322116
rect 461688 320958 461716 322116
rect 461676 320952 461728 320958
rect 461676 320894 461728 320900
rect 461964 320822 461992 322116
rect 461952 320816 462004 320822
rect 461952 320758 462004 320764
rect 461400 320680 461452 320686
rect 461400 320622 461452 320628
rect 462240 320006 462268 322116
rect 462516 320074 462544 322116
rect 462504 320068 462556 320074
rect 462504 320010 462556 320016
rect 462228 320000 462280 320006
rect 462228 319942 462280 319948
rect 459742 319832 459798 319841
rect 459742 319767 459798 319776
rect 458088 318708 458140 318714
rect 458088 318650 458140 318656
rect 460570 318336 460626 318345
rect 458916 318300 458968 318306
rect 460570 318271 460626 318280
rect 458916 318242 458968 318248
rect 457720 318096 457772 318102
rect 457720 318038 457772 318044
rect 456432 316056 456484 316062
rect 456432 315998 456484 316004
rect 457444 315444 457496 315450
rect 457444 315386 457496 315392
rect 456156 291712 456208 291718
rect 456156 291654 456208 291660
rect 456432 276752 456484 276758
rect 456432 276694 456484 276700
rect 456340 273964 456392 273970
rect 456340 273906 456392 273912
rect 456248 272536 456300 272542
rect 456248 272478 456300 272484
rect 456156 268456 456208 268462
rect 456156 268398 456208 268404
rect 456168 131102 456196 268398
rect 456260 136542 456288 272478
rect 456352 139262 456380 273906
rect 456444 144838 456472 276694
rect 456524 270972 456576 270978
rect 456524 270914 456576 270920
rect 456536 267034 456564 270914
rect 456524 267028 456576 267034
rect 456524 266970 456576 266976
rect 456800 263560 456852 263566
rect 456800 263502 456852 263508
rect 456812 262721 456840 263502
rect 456798 262712 456854 262721
rect 456798 262647 456854 262656
rect 456800 249756 456852 249762
rect 456800 249698 456852 249704
rect 456812 248849 456840 249698
rect 456798 248840 456854 248849
rect 456798 248775 456854 248784
rect 456800 162308 456852 162314
rect 456800 162250 456852 162256
rect 456812 162178 456840 162250
rect 456800 162172 456852 162178
rect 456800 162114 456852 162120
rect 456432 144832 456484 144838
rect 456432 144774 456484 144780
rect 457456 143478 457484 315386
rect 457536 305448 457588 305454
rect 457536 305390 457588 305396
rect 457444 143472 457496 143478
rect 457444 143414 457496 143420
rect 456340 139256 456392 139262
rect 456340 139198 456392 139204
rect 457548 137902 457576 305390
rect 457628 278044 457680 278050
rect 457628 277986 457680 277992
rect 457640 151502 457668 277986
rect 457732 207942 457760 318038
rect 458824 309868 458876 309874
rect 458824 309810 458876 309816
rect 458088 280832 458140 280838
rect 458088 280774 458140 280780
rect 457812 269816 457864 269822
rect 457812 269758 457864 269764
rect 457824 248414 457852 269758
rect 457824 248386 458036 248414
rect 458008 234977 458036 248386
rect 457994 234968 458050 234977
rect 457994 234903 458050 234912
rect 457812 222148 457864 222154
rect 457812 222090 457864 222096
rect 457824 221105 457852 222090
rect 457810 221096 457866 221105
rect 457810 221031 457866 221040
rect 457720 207936 457772 207942
rect 457720 207878 457772 207884
rect 457824 162314 457852 221031
rect 457812 162308 457864 162314
rect 457812 162250 457864 162256
rect 458008 162246 458036 234903
rect 457996 162240 458048 162246
rect 457996 162182 458048 162188
rect 457628 151496 457680 151502
rect 457628 151438 457680 151444
rect 457536 137896 457588 137902
rect 457536 137838 457588 137844
rect 456248 136536 456300 136542
rect 456248 136478 456300 136484
rect 456156 131096 456208 131102
rect 456156 131038 456208 131044
rect 456064 119400 456116 119406
rect 456064 119342 456116 119348
rect 458100 113174 458128 280774
rect 458836 126954 458864 309810
rect 458928 135182 458956 318242
rect 459100 318232 459152 318238
rect 459100 318174 459152 318180
rect 459466 318200 459522 318209
rect 459008 317008 459060 317014
rect 459008 316950 459060 316956
rect 459020 141982 459048 316950
rect 459112 147422 459140 318174
rect 459466 318135 459522 318144
rect 459284 282192 459336 282198
rect 459284 282134 459336 282140
rect 459192 274032 459244 274038
rect 459192 273974 459244 273980
rect 459100 147416 459152 147422
rect 459100 147358 459152 147364
rect 459008 141976 459060 141982
rect 459008 141918 459060 141924
rect 458916 135176 458968 135182
rect 458916 135118 458968 135124
rect 458824 126948 458876 126954
rect 458824 126890 458876 126896
rect 459204 122058 459232 273974
rect 459296 146266 459324 282134
rect 459480 200190 459508 318135
rect 459560 207936 459612 207942
rect 459560 207878 459612 207884
rect 459572 207233 459600 207878
rect 459558 207224 459614 207233
rect 459558 207159 459614 207168
rect 459468 200184 459520 200190
rect 459468 200126 459520 200132
rect 459572 161498 459600 207159
rect 460584 201142 460612 318271
rect 460756 318164 460808 318170
rect 460756 318106 460808 318112
rect 460664 318096 460716 318102
rect 460664 318038 460716 318044
rect 460572 201136 460624 201142
rect 460572 201078 460624 201084
rect 460676 200274 460704 318038
rect 460768 200734 460796 318106
rect 461584 316056 461636 316062
rect 461584 315998 461636 316004
rect 461596 299470 461624 315998
rect 462792 314158 462820 322116
rect 462780 314152 462832 314158
rect 462780 314094 462832 314100
rect 463068 313954 463096 322116
rect 463056 313948 463108 313954
rect 463056 313890 463108 313896
rect 463344 302734 463372 322116
rect 463620 306202 463648 322116
rect 463896 306270 463924 322116
rect 463884 306264 463936 306270
rect 463884 306206 463936 306212
rect 463608 306196 463660 306202
rect 463608 306138 463660 306144
rect 464172 305522 464200 322116
rect 464448 305590 464476 322116
rect 464724 306338 464752 322116
rect 464712 306332 464764 306338
rect 464712 306274 464764 306280
rect 464436 305584 464488 305590
rect 464436 305526 464488 305532
rect 464160 305516 464212 305522
rect 464160 305458 464212 305464
rect 463332 302728 463384 302734
rect 463332 302670 463384 302676
rect 461584 299464 461636 299470
rect 461584 299406 461636 299412
rect 465000 286550 465028 322116
rect 465276 308446 465304 322116
rect 465264 308440 465316 308446
rect 465264 308382 465316 308388
rect 465552 301714 465580 322116
rect 465540 301708 465592 301714
rect 465540 301650 465592 301656
rect 464988 286544 465040 286550
rect 464988 286486 465040 286492
rect 462228 273284 462280 273290
rect 462228 273226 462280 273232
rect 462240 270978 462268 273226
rect 462228 270972 462280 270978
rect 462228 270914 462280 270920
rect 465828 269890 465856 322116
rect 466104 299946 466132 322116
rect 466092 299940 466144 299946
rect 466092 299882 466144 299888
rect 465816 269884 465868 269890
rect 465816 269826 465868 269832
rect 466380 269822 466408 322116
rect 466460 276888 466512 276894
rect 466460 276830 466512 276836
rect 466472 273290 466500 276830
rect 466460 273284 466512 273290
rect 466460 273226 466512 273232
rect 466656 271182 466684 322116
rect 466932 313274 466960 322116
rect 467208 321366 467236 322116
rect 467196 321360 467248 321366
rect 467196 321302 467248 321308
rect 467484 319938 467512 322116
rect 467760 320006 467788 322116
rect 467748 320000 467800 320006
rect 467748 319942 467800 319948
rect 467472 319932 467524 319938
rect 467472 319874 467524 319880
rect 468036 319870 468064 322116
rect 468312 321910 468340 322116
rect 468300 321904 468352 321910
rect 468300 321846 468352 321852
rect 468588 320074 468616 322116
rect 468864 321434 468892 322116
rect 468852 321428 468904 321434
rect 468852 321370 468904 321376
rect 469140 321337 469168 322116
rect 469126 321328 469182 321337
rect 469126 321263 469182 321272
rect 468576 320068 468628 320074
rect 468576 320010 468628 320016
rect 468024 319864 468076 319870
rect 468024 319806 468076 319812
rect 469416 318442 469444 322116
rect 469692 319462 469720 322116
rect 469968 319598 469996 322116
rect 470244 319802 470272 322116
rect 470232 319796 470284 319802
rect 470232 319738 470284 319744
rect 470520 319734 470548 322116
rect 470796 320618 470824 322116
rect 470784 320612 470836 320618
rect 470784 320554 470836 320560
rect 471348 319977 471376 322116
rect 471334 319968 471390 319977
rect 471334 319903 471390 319912
rect 470508 319728 470560 319734
rect 470508 319670 470560 319676
rect 469956 319592 470008 319598
rect 469956 319534 470008 319540
rect 471624 319530 471652 322116
rect 472176 321994 472204 322116
rect 471796 321972 471848 321978
rect 471796 321914 471848 321920
rect 472084 321966 472204 321994
rect 471808 321858 471836 321914
rect 472084 321858 472112 321966
rect 471808 321830 472112 321858
rect 472452 321774 472480 322116
rect 472440 321768 472492 321774
rect 472440 321710 472492 321716
rect 471612 319524 471664 319530
rect 471612 319466 471664 319472
rect 469680 319456 469732 319462
rect 469680 319398 469732 319404
rect 472728 318510 472756 322116
rect 473004 319666 473032 322116
rect 472992 319660 473044 319666
rect 472992 319602 473044 319608
rect 472716 318504 472768 318510
rect 472716 318446 472768 318452
rect 469404 318436 469456 318442
rect 469404 318378 469456 318384
rect 466920 313268 466972 313274
rect 466920 313210 466972 313216
rect 472624 311364 472676 311370
rect 472624 311306 472676 311312
rect 471244 301096 471296 301102
rect 471244 301038 471296 301044
rect 471256 295390 471284 301038
rect 469864 295384 469916 295390
rect 469864 295326 469916 295332
rect 471244 295384 471296 295390
rect 471244 295326 471296 295332
rect 467104 277432 467156 277438
rect 467104 277374 467156 277380
rect 466644 271176 466696 271182
rect 466644 271118 466696 271124
rect 466368 269816 466420 269822
rect 466368 269758 466420 269764
rect 467116 268530 467144 277374
rect 469876 268598 469904 295326
rect 471980 279064 472032 279070
rect 471980 279006 472032 279012
rect 471992 276894 472020 279006
rect 472636 277438 472664 311306
rect 473280 301102 473308 322116
rect 473556 302870 473584 322116
rect 473544 302864 473596 302870
rect 473544 302806 473596 302812
rect 473832 302802 473860 322116
rect 474108 305930 474136 322116
rect 474384 306066 474412 322116
rect 474660 306134 474688 322116
rect 474648 306128 474700 306134
rect 474648 306070 474700 306076
rect 474372 306060 474424 306066
rect 474372 306002 474424 306008
rect 474936 305998 474964 322116
rect 474924 305992 474976 305998
rect 474924 305934 474976 305940
rect 474096 305924 474148 305930
rect 474096 305866 474148 305872
rect 473820 302796 473872 302802
rect 473820 302738 473872 302744
rect 473268 301096 473320 301102
rect 473268 301038 473320 301044
rect 475212 286618 475240 322116
rect 475488 305930 475516 322116
rect 475764 311166 475792 322116
rect 475752 311160 475804 311166
rect 475752 311102 475804 311108
rect 475476 305924 475528 305930
rect 475476 305866 475528 305872
rect 475384 303680 475436 303686
rect 475384 303622 475436 303628
rect 475200 286612 475252 286618
rect 475200 286554 475252 286560
rect 475396 279070 475424 303622
rect 476040 290494 476068 322116
rect 476316 309806 476344 322116
rect 476304 309800 476356 309806
rect 476304 309742 476356 309748
rect 476592 302870 476620 322116
rect 476580 302864 476632 302870
rect 476580 302806 476632 302812
rect 476868 293282 476896 322116
rect 477144 316034 477172 322116
rect 477420 321858 477448 322116
rect 477500 321904 477552 321910
rect 477420 321852 477500 321858
rect 477420 321846 477552 321852
rect 477420 321830 477540 321846
rect 477696 320958 477724 322116
rect 477972 321298 478000 322116
rect 477960 321292 478012 321298
rect 477960 321234 478012 321240
rect 477684 320952 477736 320958
rect 477684 320894 477736 320900
rect 478248 319598 478276 322116
rect 478524 319666 478552 322116
rect 478800 319802 478828 322116
rect 478788 319796 478840 319802
rect 478788 319738 478840 319744
rect 478512 319660 478564 319666
rect 478512 319602 478564 319608
rect 478236 319592 478288 319598
rect 478236 319534 478288 319540
rect 479076 319530 479104 322116
rect 479352 320142 479380 322116
rect 479340 320136 479392 320142
rect 479340 320078 479392 320084
rect 479628 319734 479656 322116
rect 479904 320550 479932 322116
rect 480180 321094 480208 322116
rect 480168 321088 480220 321094
rect 480168 321030 480220 321036
rect 480456 321026 480484 322116
rect 480732 321842 480760 322116
rect 480720 321836 480772 321842
rect 480720 321778 480772 321784
rect 481008 321065 481036 322116
rect 480994 321056 481050 321065
rect 480444 321020 480496 321026
rect 480994 320991 481050 321000
rect 480444 320962 480496 320968
rect 479892 320544 479944 320550
rect 479892 320486 479944 320492
rect 479616 319728 479668 319734
rect 479616 319670 479668 319676
rect 479064 319524 479116 319530
rect 479064 319466 479116 319472
rect 479524 319456 479576 319462
rect 479524 319398 479576 319404
rect 477144 316006 477264 316034
rect 476856 293276 476908 293282
rect 476856 293218 476908 293224
rect 476028 290488 476080 290494
rect 476028 290430 476080 290436
rect 477236 283626 477264 316006
rect 479536 303686 479564 319398
rect 481284 319190 481312 322116
rect 481560 320113 481588 322116
rect 481836 321201 481864 322116
rect 481822 321192 481878 321201
rect 481822 321127 481878 321136
rect 481546 320104 481602 320113
rect 481546 320039 481602 320048
rect 481272 319184 481324 319190
rect 481272 319126 481324 319132
rect 480904 319116 480956 319122
rect 480904 319058 480956 319064
rect 480916 311370 480944 319058
rect 482112 318578 482140 322116
rect 482664 319258 482692 322116
rect 482940 319326 482968 322116
rect 482928 319320 482980 319326
rect 482928 319262 482980 319268
rect 482652 319252 482704 319258
rect 482652 319194 482704 319200
rect 483216 318646 483244 322116
rect 483492 319462 483520 322116
rect 483480 319456 483532 319462
rect 483480 319398 483532 319404
rect 483768 319122 483796 322116
rect 483756 319116 483808 319122
rect 483756 319058 483808 319064
rect 483204 318640 483256 318646
rect 483204 318582 483256 318588
rect 482100 318572 482152 318578
rect 482100 318514 482152 318520
rect 480904 311364 480956 311370
rect 480904 311306 480956 311312
rect 479524 303680 479576 303686
rect 479524 303622 479576 303628
rect 484044 303550 484072 322116
rect 484320 303618 484348 322116
rect 484596 305726 484624 322116
rect 484872 305862 484900 322116
rect 484860 305856 484912 305862
rect 484860 305798 484912 305804
rect 485148 305794 485176 322116
rect 485136 305788 485188 305794
rect 485136 305730 485188 305736
rect 484584 305720 484636 305726
rect 484584 305662 484636 305668
rect 484308 303612 484360 303618
rect 484308 303554 484360 303560
rect 484032 303544 484084 303550
rect 484032 303486 484084 303492
rect 477224 283620 477276 283626
rect 477224 283562 477276 283568
rect 475384 279064 475436 279070
rect 475384 279006 475436 279012
rect 472624 277432 472676 277438
rect 472624 277374 472676 277380
rect 471980 276888 472032 276894
rect 471980 276830 472032 276836
rect 485424 276690 485452 322116
rect 485700 298790 485728 322116
rect 485872 319116 485924 319122
rect 485872 319058 485924 319064
rect 485688 298784 485740 298790
rect 485688 298726 485740 298732
rect 485884 290562 485912 319058
rect 485976 316946 486004 322116
rect 485964 316940 486016 316946
rect 485964 316882 486016 316888
rect 486252 304502 486280 322116
rect 486240 304496 486292 304502
rect 486240 304438 486292 304444
rect 485872 290556 485924 290562
rect 485872 290498 485924 290504
rect 486528 286618 486556 322116
rect 486804 316034 486832 322116
rect 487080 319122 487108 322116
rect 487068 319116 487120 319122
rect 487068 319058 487120 319064
rect 486804 316006 486924 316034
rect 486516 286612 486568 286618
rect 486516 286554 486568 286560
rect 485412 276684 485464 276690
rect 485412 276626 485464 276632
rect 469864 268592 469916 268598
rect 469864 268534 469916 268540
rect 486896 268530 486924 316006
rect 487356 274038 487384 322116
rect 487344 274032 487396 274038
rect 487344 273974 487396 273980
rect 487632 272610 487660 322116
rect 487908 286686 487936 322116
rect 487896 286680 487948 286686
rect 487896 286622 487948 286628
rect 488184 275398 488212 322116
rect 488460 309874 488488 322116
rect 488448 309868 488500 309874
rect 488448 309810 488500 309816
rect 488736 308514 488764 322116
rect 489012 316878 489040 322116
rect 489000 316872 489052 316878
rect 489000 316814 489052 316820
rect 488724 308508 488776 308514
rect 488724 308450 488776 308456
rect 488172 275392 488224 275398
rect 488172 275334 488224 275340
rect 487620 272604 487672 272610
rect 487620 272546 487672 272552
rect 467104 268524 467156 268530
rect 467104 268466 467156 268472
rect 486884 268524 486936 268530
rect 486884 268466 486936 268472
rect 489288 268462 489316 322116
rect 489564 315382 489592 322116
rect 489552 315376 489604 315382
rect 489552 315318 489604 315324
rect 489840 271250 489868 322116
rect 490116 318306 490144 322116
rect 490104 318300 490156 318306
rect 490104 318242 490156 318248
rect 490392 272542 490420 322116
rect 490668 305454 490696 322116
rect 490656 305448 490708 305454
rect 490656 305390 490708 305396
rect 490944 273970 490972 322116
rect 491220 275330 491248 322116
rect 491496 317014 491524 322116
rect 491484 317008 491536 317014
rect 491484 316950 491536 316956
rect 491772 315450 491800 322116
rect 491760 315444 491812 315450
rect 491760 315386 491812 315392
rect 492048 276758 492076 322116
rect 492324 282198 492352 322116
rect 492600 318238 492628 322116
rect 492588 318232 492640 318238
rect 492588 318174 492640 318180
rect 492876 314090 492904 322116
rect 492864 314084 492916 314090
rect 492864 314026 492916 314032
rect 492312 282192 492364 282198
rect 492312 282134 492364 282140
rect 493152 280906 493180 322116
rect 493140 280900 493192 280906
rect 493140 280842 493192 280848
rect 493428 278050 493456 322116
rect 493704 279478 493732 322116
rect 493980 283694 494008 322116
rect 494256 311302 494284 322116
rect 494244 311296 494296 311302
rect 494244 311238 494296 311244
rect 494532 285054 494560 322116
rect 494808 318238 494836 322116
rect 494796 318232 494848 318238
rect 494796 318174 494848 318180
rect 494520 285048 494572 285054
rect 494520 284990 494572 284996
rect 493968 283688 494020 283694
rect 493968 283630 494020 283636
rect 493692 279472 493744 279478
rect 493692 279414 493744 279420
rect 493416 278044 493468 278050
rect 493416 277986 493468 277992
rect 492036 276752 492088 276758
rect 492036 276694 492088 276700
rect 491208 275324 491260 275330
rect 491208 275266 491260 275272
rect 490932 273964 490984 273970
rect 490932 273906 490984 273912
rect 490380 272536 490432 272542
rect 490380 272478 490432 272484
rect 495084 271250 495112 322116
rect 489828 271244 489880 271250
rect 489828 271186 489880 271192
rect 495072 271244 495124 271250
rect 495072 271186 495124 271192
rect 495360 268462 495388 322116
rect 495636 316878 495664 322116
rect 495624 316872 495676 316878
rect 495624 316814 495676 316820
rect 495912 309874 495940 322116
rect 495900 309868 495952 309874
rect 495900 309810 495952 309816
rect 496188 272542 496216 322116
rect 496464 318306 496492 322116
rect 496452 318300 496504 318306
rect 496452 318242 496504 318248
rect 496740 316034 496768 322116
rect 496372 316006 496768 316034
rect 496372 312594 496400 316006
rect 496360 312588 496412 312594
rect 496360 312530 496412 312536
rect 497016 308514 497044 322116
rect 497292 319394 497320 322116
rect 497280 319388 497332 319394
rect 497280 319330 497332 319336
rect 497004 308508 497056 308514
rect 497004 308450 497056 308456
rect 497568 273970 497596 322116
rect 497740 317756 497792 317762
rect 497740 317698 497792 317704
rect 497752 276690 497780 317698
rect 497740 276684 497792 276690
rect 497740 276626 497792 276632
rect 497844 275330 497872 322116
rect 498120 317762 498148 322116
rect 498108 317756 498160 317762
rect 498108 317698 498160 317704
rect 497832 275324 497884 275330
rect 497832 275266 497884 275272
rect 497556 273964 497608 273970
rect 497556 273906 497608 273912
rect 498396 272610 498424 322116
rect 498672 317082 498700 322116
rect 498660 317076 498712 317082
rect 498660 317018 498712 317024
rect 498948 274038 498976 322116
rect 499224 319274 499252 322116
rect 499040 319246 499252 319274
rect 499040 316062 499068 319246
rect 499500 319002 499528 322116
rect 499132 318974 499528 319002
rect 499028 316056 499080 316062
rect 499028 315998 499080 316004
rect 499132 315382 499160 318974
rect 499776 317014 499804 322116
rect 499764 317008 499816 317014
rect 499764 316950 499816 316956
rect 499212 316056 499264 316062
rect 499212 315998 499264 316004
rect 499120 315376 499172 315382
rect 499120 315318 499172 315324
rect 499224 278050 499252 315998
rect 500052 312662 500080 322116
rect 500328 314090 500356 322116
rect 500604 316034 500632 322116
rect 500512 316006 500632 316034
rect 500316 314084 500368 314090
rect 500316 314026 500368 314032
rect 500040 312656 500092 312662
rect 500040 312598 500092 312604
rect 499212 278044 499264 278050
rect 499212 277986 499264 277992
rect 500512 275398 500540 316006
rect 500880 280906 500908 322116
rect 501156 315353 501184 322116
rect 501142 315344 501198 315353
rect 501142 315279 501198 315288
rect 501432 283694 501460 322116
rect 501708 313993 501736 322116
rect 501694 313984 501750 313993
rect 501694 313919 501750 313928
rect 501984 311302 502012 322116
rect 501972 311296 502024 311302
rect 501972 311238 502024 311244
rect 502260 287774 502288 322116
rect 502536 319462 502564 322116
rect 502524 319456 502576 319462
rect 502524 319398 502576 319404
rect 502708 319116 502760 319122
rect 502708 319058 502760 319064
rect 502720 315314 502748 319058
rect 502708 315308 502760 315314
rect 502708 315250 502760 315256
rect 502812 298858 502840 322116
rect 503088 301646 503116 322116
rect 503364 316810 503392 322116
rect 503640 319122 503668 322116
rect 503628 319116 503680 319122
rect 503628 319058 503680 319064
rect 503352 316804 503404 316810
rect 503352 316746 503404 316752
rect 503916 314022 503944 322116
rect 504192 316742 504220 322116
rect 504180 316736 504232 316742
rect 504180 316678 504232 316684
rect 503904 314016 503956 314022
rect 503904 313958 503956 313964
rect 504468 311234 504496 322116
rect 504456 311228 504508 311234
rect 504456 311170 504508 311176
rect 503076 301640 503128 301646
rect 503076 301582 503128 301588
rect 502800 298852 502852 298858
rect 502800 298794 502852 298800
rect 502248 287768 502300 287774
rect 502248 287710 502300 287716
rect 501420 283688 501472 283694
rect 501420 283630 501472 283636
rect 500868 280900 500920 280906
rect 500868 280842 500920 280848
rect 500500 275392 500552 275398
rect 500500 275334 500552 275340
rect 498936 274032 498988 274038
rect 498936 273974 498988 273980
rect 498384 272604 498436 272610
rect 498384 272546 498436 272552
rect 496176 272536 496228 272542
rect 496176 272478 496228 272484
rect 489276 268456 489328 268462
rect 489276 268398 489328 268404
rect 495348 268456 495400 268462
rect 495348 268398 495400 268404
rect 504744 268394 504772 322116
rect 505020 287706 505048 322116
rect 505008 287700 505060 287706
rect 505008 287642 505060 287648
rect 505296 280838 505324 322116
rect 507122 321872 507178 321881
rect 507122 321807 507178 321816
rect 507216 321836 507268 321842
rect 507136 289814 507164 321807
rect 507216 321778 507268 321784
rect 507124 289808 507176 289814
rect 507124 289750 507176 289756
rect 507228 289066 507256 321778
rect 507400 321768 507452 321774
rect 507400 321710 507452 321716
rect 507306 321600 507362 321609
rect 507306 321535 507362 321544
rect 507216 289060 507268 289066
rect 507216 289002 507268 289008
rect 507320 288998 507348 321535
rect 507412 291786 507440 321710
rect 509712 320793 509740 322895
rect 509698 320784 509754 320793
rect 509698 320719 509754 320728
rect 507676 320340 507728 320346
rect 507676 320282 507728 320288
rect 507582 320240 507638 320249
rect 507492 320204 507544 320210
rect 507582 320175 507638 320184
rect 507492 320146 507544 320152
rect 507504 292534 507532 320146
rect 507596 295322 507624 320175
rect 507584 295316 507636 295322
rect 507584 295258 507636 295264
rect 507688 294574 507716 320282
rect 507768 320272 507820 320278
rect 507768 320214 507820 320220
rect 507676 294568 507728 294574
rect 507676 294510 507728 294516
rect 507780 294506 507808 320214
rect 509804 316690 509832 326318
rect 509712 316662 509832 316690
rect 509712 300626 509740 316662
rect 509792 314220 509844 314226
rect 509792 314162 509844 314168
rect 509700 300620 509752 300626
rect 509700 300562 509752 300568
rect 509804 295186 509832 314162
rect 509896 300762 509924 360295
rect 511078 359680 511134 359689
rect 511078 359615 511134 359624
rect 510618 359136 510674 359145
rect 510618 359071 510674 359080
rect 509974 357640 510030 357649
rect 509974 357575 510030 357584
rect 509884 300756 509936 300762
rect 509884 300698 509936 300704
rect 509988 300082 510016 357575
rect 510066 356416 510122 356425
rect 510066 356351 510122 356360
rect 510080 349858 510108 356351
rect 510068 349852 510120 349858
rect 510068 349794 510120 349800
rect 510250 330304 510306 330313
rect 510250 330239 510306 330248
rect 510068 326460 510120 326466
rect 510068 326402 510120 326408
rect 510080 314226 510108 326402
rect 510158 325000 510214 325009
rect 510158 324935 510214 324944
rect 510172 318209 510200 324935
rect 510264 320210 510292 330239
rect 510342 328128 510398 328137
rect 510342 328063 510398 328072
rect 510252 320204 510304 320210
rect 510252 320146 510304 320152
rect 510158 318200 510214 318209
rect 510158 318135 510214 318144
rect 510068 314220 510120 314226
rect 510068 314162 510120 314168
rect 509976 300076 510028 300082
rect 509976 300018 510028 300024
rect 510356 300014 510384 328063
rect 510436 323604 510488 323610
rect 510436 323546 510488 323552
rect 510448 319938 510476 323546
rect 510528 322244 510580 322250
rect 510528 322186 510580 322192
rect 510436 319932 510488 319938
rect 510436 319874 510488 319880
rect 510540 319870 510568 322186
rect 510528 319864 510580 319870
rect 510528 319806 510580 319812
rect 510632 300694 510660 359071
rect 510894 355872 510950 355881
rect 510894 355807 510950 355816
rect 510710 353152 510766 353161
rect 510710 353087 510766 353096
rect 510620 300688 510672 300694
rect 510620 300630 510672 300636
rect 510344 300008 510396 300014
rect 510344 299950 510396 299956
rect 509792 295180 509844 295186
rect 509792 295122 509844 295128
rect 510724 295118 510752 353087
rect 510908 345014 510936 355807
rect 510816 344986 510936 345014
rect 510816 300830 510844 344986
rect 510894 344448 510950 344457
rect 510894 344383 510950 344392
rect 510908 303414 510936 344383
rect 510986 342816 511042 342825
rect 510986 342751 511042 342760
rect 511000 303482 511028 342751
rect 511092 320278 511120 359615
rect 511170 348800 511226 348809
rect 511170 348735 511226 348744
rect 511184 321842 511212 348735
rect 511172 321836 511224 321842
rect 511172 321778 511224 321784
rect 511276 321162 511304 404330
rect 513392 387122 513420 600086
rect 515404 599616 515456 599622
rect 515404 599558 515456 599564
rect 513380 387116 513432 387122
rect 513380 387058 513432 387064
rect 512092 386572 512144 386578
rect 512092 386514 512144 386520
rect 512000 386436 512052 386442
rect 512000 386378 512052 386384
rect 512012 374921 512040 386378
rect 512104 377641 512132 386514
rect 512276 386504 512328 386510
rect 512276 386446 512328 386452
rect 512184 385416 512236 385422
rect 512184 385358 512236 385364
rect 512090 377632 512146 377641
rect 512090 377567 512146 377576
rect 512196 376553 512224 385358
rect 512288 378185 512316 386446
rect 513286 384704 513342 384713
rect 513286 384639 513342 384648
rect 512458 384160 512514 384169
rect 512458 384095 512514 384104
rect 512472 383722 512500 384095
rect 513300 383790 513328 384639
rect 513288 383784 513340 383790
rect 513288 383726 513340 383732
rect 512460 383716 512512 383722
rect 512460 383658 512512 383664
rect 512642 383616 512698 383625
rect 512642 383551 512698 383560
rect 512656 383042 512684 383551
rect 513010 383072 513066 383081
rect 512644 383036 512696 383042
rect 513010 383007 513066 383016
rect 512644 382978 512696 382984
rect 513024 382974 513052 383007
rect 513012 382968 513064 382974
rect 513012 382910 513064 382916
rect 512458 382528 512514 382537
rect 512458 382463 512460 382472
rect 512512 382463 512514 382472
rect 512460 382434 512512 382440
rect 513102 381984 513158 381993
rect 513102 381919 513158 381928
rect 512550 379808 512606 379817
rect 512550 379743 512552 379752
rect 512604 379743 512606 379752
rect 512552 379714 512604 379720
rect 512918 379264 512974 379273
rect 512918 379199 512974 379208
rect 512458 378720 512514 378729
rect 512458 378655 512514 378664
rect 512472 378282 512500 378655
rect 512460 378276 512512 378282
rect 512460 378218 512512 378224
rect 512932 378214 512960 379199
rect 512920 378208 512972 378214
rect 512274 378176 512330 378185
rect 512920 378150 512972 378156
rect 512274 378111 512330 378120
rect 512642 377088 512698 377097
rect 512642 377023 512698 377032
rect 512656 376786 512684 377023
rect 512644 376780 512696 376786
rect 512644 376722 512696 376728
rect 512182 376544 512238 376553
rect 512182 376479 512238 376488
rect 513116 376038 513144 381919
rect 513286 381440 513342 381449
rect 513286 381375 513342 381384
rect 513300 380934 513328 381375
rect 513288 380928 513340 380934
rect 513194 380896 513250 380905
rect 513288 380870 513340 380876
rect 513194 380831 513250 380840
rect 513208 377466 513236 380831
rect 513286 380352 513342 380361
rect 513286 380287 513342 380296
rect 513300 379574 513328 380287
rect 513288 379568 513340 379574
rect 513288 379510 513340 379516
rect 513196 377460 513248 377466
rect 513196 377402 513248 377408
rect 513104 376032 513156 376038
rect 512642 376000 512698 376009
rect 513104 375974 513156 375980
rect 512642 375935 512698 375944
rect 512656 375426 512684 375935
rect 512828 375488 512880 375494
rect 512826 375456 512828 375465
rect 512880 375456 512882 375465
rect 512644 375420 512696 375426
rect 512826 375391 512882 375400
rect 512644 375362 512696 375368
rect 511998 374912 512054 374921
rect 511998 374847 512054 374856
rect 513286 374368 513342 374377
rect 513286 374303 513342 374312
rect 513300 374066 513328 374303
rect 513288 374060 513340 374066
rect 513288 374002 513340 374008
rect 512642 373824 512698 373833
rect 512642 373759 512644 373768
rect 512696 373759 512698 373768
rect 512644 373730 512696 373736
rect 512458 373280 512514 373289
rect 512458 373215 512514 373224
rect 512472 372774 512500 373215
rect 512460 372768 512512 372774
rect 512090 372736 512146 372745
rect 512460 372710 512512 372716
rect 512090 372671 512092 372680
rect 512144 372671 512146 372680
rect 514760 372700 514812 372706
rect 512092 372642 512144 372648
rect 514760 372642 514812 372648
rect 512826 372192 512882 372201
rect 512826 372127 512882 372136
rect 512182 371648 512238 371657
rect 512182 371583 512238 371592
rect 512090 368384 512146 368393
rect 512090 368319 512146 368328
rect 511998 367840 512054 367849
rect 511998 367775 512054 367784
rect 512012 367402 512040 367775
rect 512000 367396 512052 367402
rect 512000 367338 512052 367344
rect 511998 366208 512054 366217
rect 511998 366143 512000 366152
rect 512052 366143 512054 366152
rect 512000 366114 512052 366120
rect 512104 366058 512132 368319
rect 512012 366030 512132 366058
rect 511356 352096 511408 352102
rect 511356 352038 511408 352044
rect 511368 321230 511396 352038
rect 511908 324964 511960 324970
rect 511908 324906 511960 324912
rect 511356 321224 511408 321230
rect 511356 321166 511408 321172
rect 511264 321156 511316 321162
rect 511264 321098 511316 321104
rect 511080 320272 511132 320278
rect 511080 320214 511132 320220
rect 511920 320006 511948 324906
rect 511908 320000 511960 320006
rect 511908 319942 511960 319948
rect 510988 303476 511040 303482
rect 510988 303418 511040 303424
rect 510896 303408 510948 303414
rect 510896 303350 510948 303356
rect 510804 300824 510856 300830
rect 510804 300766 510856 300772
rect 512012 300286 512040 366030
rect 512196 364334 512224 371583
rect 512840 371278 512868 372127
rect 512828 371272 512880 371278
rect 512828 371214 512880 371220
rect 512642 371104 512698 371113
rect 512642 371039 512698 371048
rect 512656 369986 512684 371039
rect 513286 370016 513342 370025
rect 512644 369980 512696 369986
rect 513286 369951 513342 369960
rect 512644 369922 512696 369928
rect 513300 369918 513328 369951
rect 513288 369912 513340 369918
rect 513288 369854 513340 369860
rect 513286 369472 513342 369481
rect 513286 369407 513342 369416
rect 512826 368928 512882 368937
rect 512826 368863 512882 368872
rect 512840 368558 512868 368863
rect 513300 368626 513328 369407
rect 513288 368620 513340 368626
rect 513288 368562 513340 368568
rect 512828 368552 512880 368558
rect 512828 368494 512880 368500
rect 514116 367396 514168 367402
rect 514116 367338 514168 367344
rect 513286 367296 513342 367305
rect 513286 367231 513288 367240
rect 513340 367231 513342 367240
rect 513288 367202 513340 367208
rect 513286 366752 513342 366761
rect 513286 366687 513342 366696
rect 513300 365770 513328 366687
rect 513288 365764 513340 365770
rect 513288 365706 513340 365712
rect 513286 365664 513342 365673
rect 513342 365622 513420 365650
rect 513286 365599 513342 365608
rect 512642 365120 512698 365129
rect 512642 365055 512698 365064
rect 512656 364410 512684 365055
rect 513286 364576 513342 364585
rect 513286 364511 513288 364520
rect 513340 364511 513342 364520
rect 513288 364482 513340 364488
rect 512644 364404 512696 364410
rect 512644 364346 512696 364352
rect 512104 364306 512224 364334
rect 513392 364334 513420 365622
rect 513392 364306 513604 364334
rect 512104 305697 512132 364306
rect 512182 364032 512238 364041
rect 512182 363967 512238 363976
rect 512196 363322 512224 363967
rect 513286 363488 513342 363497
rect 513286 363423 513342 363432
rect 512184 363316 512236 363322
rect 512184 363258 512236 363264
rect 513300 362982 513328 363423
rect 513288 362976 513340 362982
rect 513010 362944 513066 362953
rect 513288 362918 513340 362924
rect 513010 362879 513066 362888
rect 512182 362400 512238 362409
rect 512182 362335 512184 362344
rect 512236 362335 512238 362344
rect 512184 362306 512236 362312
rect 512366 361856 512422 361865
rect 512366 361791 512422 361800
rect 512274 358592 512330 358601
rect 512274 358527 512330 358536
rect 512182 358048 512238 358057
rect 512182 357983 512238 357992
rect 512196 357746 512224 357983
rect 512184 357740 512236 357746
rect 512184 357682 512236 357688
rect 512184 357604 512236 357610
rect 512184 357546 512236 357552
rect 512090 305688 512146 305697
rect 512090 305623 512146 305632
rect 512000 300280 512052 300286
rect 512000 300222 512052 300228
rect 512196 297838 512224 357546
rect 512288 301578 512316 358527
rect 512380 357610 512408 361791
rect 513024 361690 513052 362879
rect 513012 361684 513064 361690
rect 513012 361626 513064 361632
rect 513010 361312 513066 361321
rect 513010 361247 513066 361256
rect 513024 360330 513052 361247
rect 513012 360324 513064 360330
rect 513012 360266 513064 360272
rect 513288 360256 513340 360262
rect 513286 360224 513288 360233
rect 513340 360224 513342 360233
rect 513286 360159 513342 360168
rect 512368 357604 512420 357610
rect 512368 357546 512420 357552
rect 513286 356960 513342 356969
rect 513286 356895 513342 356904
rect 513300 356114 513328 356895
rect 513288 356108 513340 356114
rect 513288 356050 513340 356056
rect 512366 355328 512422 355337
rect 512366 355263 512422 355272
rect 512276 301572 512328 301578
rect 512276 301514 512328 301520
rect 512380 301510 512408 355263
rect 513286 354784 513342 354793
rect 513286 354719 513288 354728
rect 513340 354719 513342 354728
rect 513288 354690 513340 354696
rect 512458 354240 512514 354249
rect 512458 354175 512514 354184
rect 512472 353666 512500 354175
rect 513194 353696 513250 353705
rect 512460 353660 512512 353666
rect 513194 353631 513250 353640
rect 512460 353602 512512 353608
rect 513208 353530 513236 353631
rect 513196 353524 513248 353530
rect 513196 353466 513248 353472
rect 512458 352608 512514 352617
rect 512458 352543 512460 352552
rect 512512 352543 512514 352552
rect 512460 352514 512512 352520
rect 513286 352064 513342 352073
rect 513286 351999 513288 352008
rect 513340 351999 513342 352008
rect 513288 351970 513340 351976
rect 513286 351520 513342 351529
rect 513286 351455 513342 351464
rect 512458 350976 512514 350985
rect 513300 350946 513328 351455
rect 512458 350911 512514 350920
rect 513288 350940 513340 350946
rect 512472 350810 512500 350911
rect 513288 350882 513340 350888
rect 512460 350804 512512 350810
rect 512460 350746 512512 350752
rect 512458 350432 512514 350441
rect 512458 350367 512514 350376
rect 512472 349586 512500 350367
rect 513286 349888 513342 349897
rect 513286 349823 513342 349832
rect 513300 349722 513328 349823
rect 513288 349716 513340 349722
rect 513288 349658 513340 349664
rect 512460 349580 512512 349586
rect 512460 349522 512512 349528
rect 512458 349344 512514 349353
rect 512458 349279 512514 349288
rect 512472 349178 512500 349279
rect 512460 349172 512512 349178
rect 512460 349114 512512 349120
rect 513010 348256 513066 348265
rect 513010 348191 513066 348200
rect 513024 347954 513052 348191
rect 513012 347948 513064 347954
rect 513012 347890 513064 347896
rect 512458 347712 512514 347721
rect 512458 347647 512460 347656
rect 512512 347647 512514 347656
rect 512460 347618 512512 347624
rect 512826 347168 512882 347177
rect 512826 347103 512882 347112
rect 512840 346458 512868 347103
rect 513286 346624 513342 346633
rect 513286 346559 513288 346568
rect 513340 346559 513342 346568
rect 513288 346530 513340 346536
rect 512828 346452 512880 346458
rect 512828 346394 512880 346400
rect 512458 346080 512514 346089
rect 512458 346015 512514 346024
rect 512472 345642 512500 346015
rect 512460 345636 512512 345642
rect 512460 345578 512512 345584
rect 512458 345536 512514 345545
rect 512458 345471 512514 345480
rect 512472 302938 512500 345471
rect 513010 344992 513066 345001
rect 513010 344927 513066 344936
rect 513024 343738 513052 344927
rect 513288 344412 513340 344418
rect 513288 344354 513340 344360
rect 513300 343913 513328 344354
rect 513286 343904 513342 343913
rect 513286 343839 513342 343848
rect 513012 343732 513064 343738
rect 513012 343674 513064 343680
rect 513010 343360 513066 343369
rect 513010 343295 513066 343304
rect 513024 343194 513052 343295
rect 513012 343188 513064 343194
rect 513012 343130 513064 343136
rect 512550 342272 512606 342281
rect 512550 342207 512606 342216
rect 512564 302977 512592 342207
rect 513286 341728 513342 341737
rect 513286 341663 513342 341672
rect 513300 341290 513328 341663
rect 513288 341284 513340 341290
rect 513288 341226 513340 341232
rect 513286 341184 513342 341193
rect 513286 341119 513288 341128
rect 513340 341119 513342 341128
rect 513288 341090 513340 341096
rect 513286 340640 513342 340649
rect 513342 340598 513420 340626
rect 513286 340575 513342 340584
rect 513102 340096 513158 340105
rect 513102 340031 513158 340040
rect 513116 339658 513144 340031
rect 513104 339652 513156 339658
rect 513104 339594 513156 339600
rect 513288 339584 513340 339590
rect 513286 339552 513288 339561
rect 513340 339552 513342 339561
rect 513286 339487 513342 339496
rect 512642 339008 512698 339017
rect 512642 338943 512698 338952
rect 512656 304298 512684 338943
rect 513012 338700 513064 338706
rect 513012 338642 513064 338648
rect 513024 338473 513052 338642
rect 513010 338464 513066 338473
rect 513010 338399 513066 338408
rect 512734 337920 512790 337929
rect 512734 337855 512790 337864
rect 512748 337074 512776 337855
rect 512826 337376 512882 337385
rect 512826 337311 512882 337320
rect 512736 337068 512788 337074
rect 512736 337010 512788 337016
rect 512840 337006 512868 337311
rect 513288 337204 513340 337210
rect 513288 337146 513340 337152
rect 512828 337000 512880 337006
rect 512828 336942 512880 336948
rect 513300 336841 513328 337146
rect 513286 336832 513342 336841
rect 513286 336767 513342 336776
rect 512734 336288 512790 336297
rect 512734 336223 512790 336232
rect 512748 335986 512776 336223
rect 512736 335980 512788 335986
rect 512736 335922 512788 335928
rect 513010 335200 513066 335209
rect 513010 335135 513066 335144
rect 513024 334762 513052 335135
rect 513012 334756 513064 334762
rect 513012 334698 513064 334704
rect 512734 334656 512790 334665
rect 512734 334591 512790 334600
rect 513288 334620 513340 334626
rect 512748 304366 512776 334591
rect 513288 334562 513340 334568
rect 513300 334121 513328 334562
rect 513286 334112 513342 334121
rect 513286 334047 513342 334056
rect 512826 332480 512882 332489
rect 512826 332415 512882 332424
rect 512840 331634 512868 332415
rect 512828 331628 512880 331634
rect 512828 331570 512880 331576
rect 512826 329760 512882 329769
rect 512826 329695 512882 329704
rect 512840 329186 512868 329695
rect 512828 329180 512880 329186
rect 512828 329122 512880 329128
rect 512826 327040 512882 327049
rect 512826 326975 512882 326984
rect 512736 304360 512788 304366
rect 512736 304302 512788 304308
rect 512644 304292 512696 304298
rect 512644 304234 512696 304240
rect 512550 302968 512606 302977
rect 512460 302932 512512 302938
rect 512550 302903 512606 302912
rect 512460 302874 512512 302880
rect 512840 302841 512868 326975
rect 513392 318170 513420 340598
rect 513470 333568 513526 333577
rect 513470 333503 513526 333512
rect 513484 321774 513512 333503
rect 513472 321768 513524 321774
rect 513472 321710 513524 321716
rect 513380 318164 513432 318170
rect 513380 318106 513432 318112
rect 512826 302832 512882 302841
rect 512826 302767 512882 302776
rect 512368 301504 512420 301510
rect 512368 301446 512420 301452
rect 513576 300422 513604 364306
rect 513656 362364 513708 362370
rect 513656 362306 513708 362312
rect 513668 300558 513696 362306
rect 514024 357740 514076 357746
rect 514024 357682 514076 357688
rect 513748 353660 513800 353666
rect 513748 353602 513800 353608
rect 513760 303210 513788 353602
rect 513840 349172 513892 349178
rect 513840 349114 513892 349120
rect 513748 303204 513800 303210
rect 513748 303146 513800 303152
rect 513852 303142 513880 349114
rect 513932 347676 513984 347682
rect 513932 347618 513984 347624
rect 513944 303346 513972 347618
rect 514036 320346 514064 357682
rect 514024 320340 514076 320346
rect 514024 320282 514076 320288
rect 513932 303340 513984 303346
rect 513932 303282 513984 303288
rect 513840 303136 513892 303142
rect 513840 303078 513892 303084
rect 513656 300552 513708 300558
rect 513656 300494 513708 300500
rect 513564 300416 513616 300422
rect 513564 300358 513616 300364
rect 512184 297832 512236 297838
rect 512184 297774 512236 297780
rect 510712 295112 510764 295118
rect 510712 295054 510764 295060
rect 507768 294500 507820 294506
rect 507768 294442 507820 294448
rect 507492 292528 507544 292534
rect 507492 292470 507544 292476
rect 514128 292262 514156 367338
rect 514208 366172 514260 366178
rect 514208 366114 514260 366120
rect 514220 295254 514248 366114
rect 514208 295248 514260 295254
rect 514208 295190 514260 295196
rect 514772 292398 514800 372642
rect 514852 363316 514904 363322
rect 514852 363258 514904 363264
rect 514864 300490 514892 363258
rect 515036 352572 515088 352578
rect 515036 352514 515088 352520
rect 514944 349580 514996 349586
rect 514944 349522 514996 349528
rect 514852 300484 514904 300490
rect 514852 300426 514904 300432
rect 514760 292392 514812 292398
rect 514760 292334 514812 292340
rect 514116 292256 514168 292262
rect 514116 292198 514168 292204
rect 507400 291780 507452 291786
rect 507400 291722 507452 291728
rect 514956 289474 514984 349522
rect 515048 303074 515076 352514
rect 515128 350804 515180 350810
rect 515128 350746 515180 350752
rect 515036 303068 515088 303074
rect 515036 303010 515088 303016
rect 515140 303006 515168 350746
rect 515220 345636 515272 345642
rect 515220 345578 515272 345584
rect 515232 303278 515260 345578
rect 515312 337068 515364 337074
rect 515312 337010 515364 337016
rect 515220 303272 515272 303278
rect 515220 303214 515272 303220
rect 515128 303000 515180 303006
rect 515128 302942 515180 302948
rect 515324 297770 515352 337010
rect 515416 319530 515444 599558
rect 519544 590708 519596 590714
rect 519544 590650 519596 590656
rect 518164 536852 518216 536858
rect 518164 536794 518216 536800
rect 515496 484424 515548 484430
rect 515496 484366 515548 484372
rect 515508 319598 515536 484366
rect 515588 382492 515640 382498
rect 515588 382434 515640 382440
rect 515600 358494 515628 382434
rect 515680 379772 515732 379778
rect 515680 379714 515732 379720
rect 515692 359854 515720 379714
rect 516416 376780 516468 376786
rect 516416 376722 516468 376728
rect 516232 375488 516284 375494
rect 516232 375430 516284 375436
rect 515680 359848 515732 359854
rect 515680 359790 515732 359796
rect 515588 358488 515640 358494
rect 515588 358430 515640 358436
rect 516140 337000 516192 337006
rect 516140 336942 516192 336948
rect 515588 335980 515640 335986
rect 515588 335922 515640 335928
rect 515496 319592 515548 319598
rect 515496 319534 515548 319540
rect 515404 319524 515456 319530
rect 515404 319466 515456 319472
rect 515312 297764 515364 297770
rect 515312 297706 515364 297712
rect 515600 297566 515628 335922
rect 516152 318102 516180 336942
rect 516140 318096 516192 318102
rect 516140 318038 516192 318044
rect 515588 297560 515640 297566
rect 515588 297502 515640 297508
rect 516244 297430 516272 375430
rect 516324 373788 516376 373794
rect 516324 373730 516376 373736
rect 516336 300218 516364 373730
rect 516428 305658 516456 376722
rect 517520 371272 517572 371278
rect 517520 371214 517572 371220
rect 516968 369980 517020 369986
rect 516968 369922 517020 369928
rect 516508 368552 516560 368558
rect 516508 368494 516560 368500
rect 516416 305652 516468 305658
rect 516416 305594 516468 305600
rect 516520 300354 516548 368494
rect 516692 347948 516744 347954
rect 516692 347890 516744 347896
rect 516600 346452 516652 346458
rect 516600 346394 516652 346400
rect 516508 300348 516560 300354
rect 516508 300290 516560 300296
rect 516324 300212 516376 300218
rect 516324 300154 516376 300160
rect 516232 297424 516284 297430
rect 516232 297366 516284 297372
rect 516612 289610 516640 346394
rect 516704 294642 516732 347890
rect 516784 339652 516836 339658
rect 516784 339594 516836 339600
rect 516692 294636 516744 294642
rect 516692 294578 516744 294584
rect 516796 292058 516824 339594
rect 516876 329180 516928 329186
rect 516876 329122 516928 329128
rect 516888 297634 516916 329122
rect 516876 297628 516928 297634
rect 516876 297570 516928 297576
rect 516980 292330 517008 369922
rect 517532 300150 517560 371214
rect 517888 367260 517940 367266
rect 517888 367202 517940 367208
rect 517612 361684 517664 361690
rect 517612 361626 517664 361632
rect 517520 300144 517572 300150
rect 517520 300086 517572 300092
rect 517624 295050 517652 361626
rect 517704 360324 517756 360330
rect 517704 360266 517756 360272
rect 517612 295044 517664 295050
rect 517612 294986 517664 294992
rect 517716 294982 517744 360266
rect 517796 353524 517848 353530
rect 517796 353466 517848 353472
rect 517704 294976 517756 294982
rect 517704 294918 517756 294924
rect 516968 292324 517020 292330
rect 516968 292266 517020 292272
rect 516784 292052 516836 292058
rect 516784 291994 516836 292000
rect 517808 289746 517836 353466
rect 517900 305833 517928 367202
rect 517980 354748 518032 354754
rect 517980 354690 518032 354696
rect 517886 305824 517942 305833
rect 517886 305759 517942 305768
rect 517992 294846 518020 354690
rect 518072 346588 518124 346594
rect 518072 346530 518124 346536
rect 518084 297974 518112 346530
rect 518176 319666 518204 536794
rect 518256 382968 518308 382974
rect 518256 382910 518308 382916
rect 518268 358698 518296 382910
rect 518900 360256 518952 360262
rect 518900 360198 518952 360204
rect 518256 358692 518308 358698
rect 518256 358634 518308 358640
rect 518256 343732 518308 343738
rect 518256 343674 518308 343680
rect 518164 319660 518216 319666
rect 518164 319602 518216 319608
rect 518072 297968 518124 297974
rect 518072 297910 518124 297916
rect 518268 297906 518296 343674
rect 518348 343188 518400 343194
rect 518348 343130 518400 343136
rect 518256 297900 518308 297906
rect 518256 297842 518308 297848
rect 518360 297702 518388 343130
rect 518348 297696 518400 297702
rect 518348 297638 518400 297644
rect 517980 294840 518032 294846
rect 517980 294782 518032 294788
rect 517796 289740 517848 289746
rect 517796 289682 517848 289688
rect 516600 289604 516652 289610
rect 516600 289546 516652 289552
rect 518912 289542 518940 360198
rect 518992 350940 519044 350946
rect 518992 350882 519044 350888
rect 519004 294710 519032 350882
rect 519176 349716 519228 349722
rect 519176 349658 519228 349664
rect 519084 344412 519136 344418
rect 519084 344354 519136 344360
rect 518992 294704 519044 294710
rect 518992 294646 519044 294652
rect 518900 289536 518952 289542
rect 518900 289478 518952 289484
rect 514944 289468 514996 289474
rect 514944 289410 514996 289416
rect 519096 289406 519124 344354
rect 519188 294778 519216 349658
rect 519360 341148 519412 341154
rect 519360 341090 519412 341096
rect 519268 338700 519320 338706
rect 519268 338642 519320 338648
rect 519176 294772 519228 294778
rect 519176 294714 519228 294720
rect 519280 291990 519308 338642
rect 519372 298042 519400 341090
rect 519452 334756 519504 334762
rect 519452 334698 519504 334704
rect 519360 298036 519412 298042
rect 519360 297978 519412 297984
rect 519268 291984 519320 291990
rect 519268 291926 519320 291932
rect 519464 291854 519492 334698
rect 519556 319802 519584 590650
rect 520292 520946 520320 600086
rect 520280 520940 520332 520946
rect 520280 520882 520332 520888
rect 519634 502344 519690 502353
rect 519634 502279 519690 502288
rect 519544 319796 519596 319802
rect 519544 319738 519596 319744
rect 519648 319734 519676 502279
rect 525812 464370 525840 600086
rect 547878 516760 547934 516769
rect 547878 516695 547934 516704
rect 545120 514072 545172 514078
rect 545120 514014 545172 514020
rect 535460 512644 535512 512650
rect 535460 512586 535512 512592
rect 532700 508564 532752 508570
rect 532700 508506 532752 508512
rect 529940 505776 529992 505782
rect 529940 505718 529992 505724
rect 529952 480254 529980 505718
rect 532712 480254 532740 508506
rect 535472 480254 535500 512586
rect 538220 509924 538272 509930
rect 538220 509866 538272 509872
rect 538232 480254 538260 509866
rect 529952 480226 530256 480254
rect 532712 480226 533200 480254
rect 535472 480226 536144 480254
rect 538232 480226 539088 480254
rect 525800 464364 525852 464370
rect 525800 464306 525852 464312
rect 521750 462904 521806 462913
rect 521750 462839 521806 462848
rect 521764 460972 521792 462839
rect 527640 462460 527692 462466
rect 527640 462402 527692 462408
rect 524696 461100 524748 461106
rect 524696 461042 524748 461048
rect 524708 460972 524736 461042
rect 527652 460972 527680 462402
rect 530228 460986 530256 480226
rect 533172 460986 533200 480226
rect 536116 460986 536144 480226
rect 539060 460986 539088 480226
rect 542360 462392 542412 462398
rect 542360 462334 542412 462340
rect 530228 460958 530610 460986
rect 533172 460958 533554 460986
rect 536116 460958 536498 460986
rect 539060 460958 539442 460986
rect 542372 460972 542400 462334
rect 545132 460986 545160 514014
rect 547892 460986 547920 516695
rect 553860 461032 553912 461038
rect 545132 460958 545330 460986
rect 547892 460958 548274 460986
rect 550928 460970 551218 460986
rect 553912 460980 554162 460986
rect 553860 460974 554162 460980
rect 550916 460964 551218 460970
rect 550968 460958 551218 460964
rect 553872 460958 554162 460974
rect 550916 460906 550968 460912
rect 557538 442912 557594 442921
rect 557538 442847 557594 442856
rect 521212 421598 521240 425068
rect 522304 423496 522356 423502
rect 522304 423438 522356 423444
rect 521200 421592 521252 421598
rect 521200 421534 521252 421540
rect 522316 388686 522344 423438
rect 522500 423434 522528 425068
rect 523788 423570 523816 425068
rect 524708 425054 525090 425082
rect 523776 423564 523828 423570
rect 523776 423506 523828 423512
rect 522488 423428 522540 423434
rect 522488 423370 522540 423376
rect 523684 423428 523736 423434
rect 523684 423370 523736 423376
rect 523696 388754 523724 423370
rect 524708 412634 524736 425054
rect 526364 423366 526392 425068
rect 526352 423360 526404 423366
rect 526352 423302 526404 423308
rect 526444 423360 526496 423366
rect 526444 423302 526496 423308
rect 524432 412606 524736 412634
rect 523684 388748 523736 388754
rect 523684 388690 523736 388696
rect 522304 388680 522356 388686
rect 522304 388622 522356 388628
rect 524432 388618 524460 412606
rect 526456 388822 526484 423302
rect 527652 416090 527680 425068
rect 528940 423298 528968 425068
rect 530228 423638 530256 425068
rect 529204 423632 529256 423638
rect 529204 423574 529256 423580
rect 530216 423632 530268 423638
rect 530216 423574 530268 423580
rect 530584 423632 530636 423638
rect 530584 423574 530636 423580
rect 528928 423292 528980 423298
rect 528928 423234 528980 423240
rect 527640 416084 527692 416090
rect 527640 416026 527692 416032
rect 526444 388816 526496 388822
rect 526444 388758 526496 388764
rect 524420 388612 524472 388618
rect 524420 388554 524472 388560
rect 529216 388482 529244 423574
rect 530596 388550 530624 423574
rect 531516 423230 531544 425068
rect 532804 423638 532832 425068
rect 532792 423632 532844 423638
rect 532792 423574 532844 423580
rect 531504 423224 531556 423230
rect 531504 423166 531556 423172
rect 533436 421592 533488 421598
rect 533436 421534 533488 421540
rect 530584 388544 530636 388550
rect 530584 388486 530636 388492
rect 529204 388476 529256 388482
rect 529204 388418 529256 388424
rect 519728 383036 519780 383042
rect 519728 382978 519780 382984
rect 519740 358630 519768 382978
rect 522304 378276 522356 378282
rect 522304 378218 522356 378224
rect 520280 375420 520332 375426
rect 520280 375362 520332 375368
rect 519728 358624 519780 358630
rect 519728 358566 519780 358572
rect 519728 339584 519780 339590
rect 519728 339526 519780 339532
rect 519636 319728 519688 319734
rect 519636 319670 519688 319676
rect 519740 297498 519768 339526
rect 519728 297492 519780 297498
rect 519728 297434 519780 297440
rect 520292 292466 520320 375362
rect 520372 374060 520424 374066
rect 520372 374002 520424 374008
rect 520280 292460 520332 292466
rect 520280 292402 520332 292408
rect 520384 292194 520412 374002
rect 521660 369912 521712 369918
rect 521660 369854 521712 369860
rect 520464 368620 520516 368626
rect 520464 368562 520516 368568
rect 520372 292188 520424 292194
rect 520372 292130 520424 292136
rect 520476 292126 520504 368562
rect 520556 364540 520608 364546
rect 520556 364482 520608 364488
rect 520568 294914 520596 364482
rect 520648 341284 520700 341290
rect 520648 341226 520700 341232
rect 520556 294908 520608 294914
rect 520556 294850 520608 294856
rect 520464 292120 520516 292126
rect 520464 292062 520516 292068
rect 519452 291848 519504 291854
rect 519452 291790 519504 291796
rect 519084 289400 519136 289406
rect 519084 289342 519136 289348
rect 520660 289134 520688 341226
rect 520740 337204 520792 337210
rect 520740 337146 520792 337152
rect 520752 291922 520780 337146
rect 520924 334620 520976 334626
rect 520924 334562 520976 334568
rect 520832 331628 520884 331634
rect 520832 331570 520884 331576
rect 520844 304434 520872 331570
rect 520936 307086 520964 334562
rect 520924 307080 520976 307086
rect 520924 307022 520976 307028
rect 520832 304428 520884 304434
rect 520832 304370 520884 304376
rect 520740 291916 520792 291922
rect 520740 291858 520792 291864
rect 520648 289128 520700 289134
rect 520648 289070 520700 289076
rect 507308 288992 507360 288998
rect 507308 288934 507360 288940
rect 521672 286414 521700 369854
rect 521752 364404 521804 364410
rect 521752 364346 521804 364352
rect 521764 289202 521792 364346
rect 522316 359786 522344 378218
rect 523040 372768 523092 372774
rect 523040 372710 523092 372716
rect 522304 359780 522356 359786
rect 522304 359722 522356 359728
rect 521844 356108 521896 356114
rect 521844 356050 521896 356056
rect 521856 289678 521884 356050
rect 521844 289672 521896 289678
rect 521844 289614 521896 289620
rect 521752 289196 521804 289202
rect 521752 289138 521804 289144
rect 523052 286482 523080 372710
rect 523132 365764 523184 365770
rect 523132 365706 523184 365712
rect 523040 286476 523092 286482
rect 523040 286418 523092 286424
rect 521660 286408 521712 286414
rect 521660 286350 521712 286356
rect 523144 286346 523172 365706
rect 523224 362976 523276 362982
rect 523224 362918 523276 362924
rect 523236 289270 523264 362918
rect 523316 352028 523368 352034
rect 523316 351970 523368 351976
rect 523328 289338 523356 351970
rect 533448 320074 533476 421534
rect 534092 392630 534120 425068
rect 535012 425054 535394 425082
rect 536300 425054 536682 425082
rect 537588 425054 537970 425082
rect 538876 425054 539258 425082
rect 540164 425054 540546 425082
rect 535012 412634 535040 425054
rect 536300 412634 536328 425054
rect 537588 412634 537616 425054
rect 538876 412634 538904 425054
rect 540164 412634 540192 425054
rect 541820 420238 541848 425068
rect 542740 425054 543122 425082
rect 544028 425054 544410 425082
rect 541808 420232 541860 420238
rect 541808 420174 541860 420180
rect 542740 412634 542768 425054
rect 544028 412634 544056 425054
rect 545684 423162 545712 425068
rect 546604 425054 546986 425082
rect 545672 423156 545724 423162
rect 545672 423098 545724 423104
rect 546604 412634 546632 425054
rect 548260 423094 548288 425068
rect 549548 423502 549576 425068
rect 549536 423496 549588 423502
rect 549536 423438 549588 423444
rect 548248 423088 548300 423094
rect 548248 423030 548300 423036
rect 550836 423026 550864 425068
rect 552124 423434 552152 425068
rect 552112 423428 552164 423434
rect 552112 423370 552164 423376
rect 550824 423020 550876 423026
rect 550824 422962 550876 422968
rect 553412 422958 553440 425068
rect 554700 423366 554728 425068
rect 557552 424386 557580 442847
rect 557540 424380 557592 424386
rect 557540 424322 557592 424328
rect 554688 423360 554740 423366
rect 554688 423302 554740 423308
rect 553400 422952 553452 422958
rect 553400 422894 553452 422900
rect 534184 412606 535040 412634
rect 535472 412606 536328 412634
rect 536852 412606 537616 412634
rect 538232 412606 538904 412634
rect 539612 412606 540192 412634
rect 542372 412606 542768 412634
rect 543752 412606 544056 412634
rect 546512 412606 546632 412634
rect 534184 393990 534212 412606
rect 534172 393984 534224 393990
rect 534172 393926 534224 393932
rect 534080 392624 534132 392630
rect 534080 392566 534132 392572
rect 535472 389910 535500 412606
rect 536852 395350 536880 412606
rect 538232 396778 538260 412606
rect 539612 398138 539640 412606
rect 539600 398132 539652 398138
rect 539600 398074 539652 398080
rect 538220 396772 538272 396778
rect 538220 396714 538272 396720
rect 536840 395344 536892 395350
rect 536840 395286 536892 395292
rect 542372 391338 542400 412606
rect 543752 399498 543780 412606
rect 546512 400926 546540 412606
rect 546500 400920 546552 400926
rect 546500 400862 546552 400868
rect 543740 399492 543792 399498
rect 543740 399434 543792 399440
rect 542360 391332 542412 391338
rect 542360 391274 542412 391280
rect 535460 389904 535512 389910
rect 535460 389846 535512 389852
rect 553952 386640 554004 386646
rect 553952 386582 554004 386588
rect 534724 383784 534776 383790
rect 534724 383726 534776 383732
rect 534736 360126 534764 383726
rect 548524 383716 548576 383722
rect 548524 383658 548576 383664
rect 547144 380928 547196 380934
rect 547144 380870 547196 380876
rect 544384 376032 544436 376038
rect 544384 375974 544436 375980
rect 534724 360120 534776 360126
rect 534724 360062 534776 360068
rect 544396 358562 544424 375974
rect 547156 359922 547184 380870
rect 547236 378208 547288 378214
rect 547236 378150 547288 378156
rect 547248 360194 547276 378150
rect 547236 360188 547288 360194
rect 547236 360130 547288 360136
rect 548536 359990 548564 383658
rect 549904 379568 549956 379574
rect 549904 379510 549956 379516
rect 548616 377460 548668 377466
rect 548616 377402 548668 377408
rect 548524 359984 548576 359990
rect 548524 359926 548576 359932
rect 547144 359916 547196 359922
rect 547144 359858 547196 359864
rect 548628 358766 548656 377402
rect 549916 360058 549944 379510
rect 553964 377890 553992 386582
rect 563428 385484 563480 385490
rect 563428 385426 563480 385432
rect 553964 377862 554438 377890
rect 563440 377876 563468 385426
rect 552032 360194 552322 360210
rect 552020 360188 552322 360194
rect 552072 360182 552322 360188
rect 552020 360130 552072 360136
rect 566740 360120 566792 360126
rect 549904 360052 549956 360058
rect 549904 359994 549956 360000
rect 550836 359786 550864 360060
rect 553780 359854 553808 360060
rect 554976 360058 555266 360074
rect 554964 360052 555266 360058
rect 555016 360046 555266 360052
rect 554964 359994 555016 360000
rect 553768 359848 553820 359854
rect 553768 359790 553820 359796
rect 550824 359780 550876 359786
rect 550824 359722 550876 359728
rect 556724 358766 556752 360060
rect 558196 359922 558224 360060
rect 558184 359916 558236 359922
rect 558184 359858 558236 359864
rect 548616 358760 548668 358766
rect 548616 358702 548668 358708
rect 556712 358760 556764 358766
rect 556712 358702 556764 358708
rect 559668 358562 559696 360060
rect 544384 358556 544436 358562
rect 544384 358498 544436 358504
rect 559656 358556 559708 358562
rect 559656 358498 559708 358504
rect 561140 358494 561168 360060
rect 562612 358698 562640 360060
rect 562600 358692 562652 358698
rect 562600 358634 562652 358640
rect 564084 358630 564112 360060
rect 565280 360046 565570 360074
rect 566792 360068 567042 360074
rect 566740 360062 567042 360068
rect 566752 360046 567042 360062
rect 565280 359990 565308 360046
rect 565268 359984 565320 359990
rect 565268 359926 565320 359932
rect 564072 358624 564124 358630
rect 564072 358566 564124 358572
rect 561128 358488 561180 358494
rect 561128 358430 561180 358436
rect 533436 320068 533488 320074
rect 533436 320010 533488 320016
rect 543740 319456 543792 319462
rect 543740 319398 543792 319404
rect 533344 319388 533396 319394
rect 533344 319330 533396 319336
rect 529940 316940 529992 316946
rect 529940 316882 529992 316888
rect 523316 289332 523368 289338
rect 523316 289274 523368 289280
rect 523224 289264 523276 289270
rect 523224 289206 523276 289212
rect 523132 286340 523184 286346
rect 523132 286282 523184 286288
rect 505284 280832 505336 280838
rect 505284 280774 505336 280780
rect 504732 268388 504784 268394
rect 504732 268330 504784 268336
rect 529952 209273 529980 316882
rect 530032 304496 530084 304502
rect 530032 304438 530084 304444
rect 530044 226250 530072 304438
rect 531320 286612 531372 286618
rect 531320 286554 531372 286560
rect 531228 268524 531280 268530
rect 531228 268466 531280 268472
rect 531240 267458 531268 268466
rect 531332 267734 531360 286554
rect 531332 267706 531544 267734
rect 531240 267430 531360 267458
rect 531332 261089 531360 267430
rect 531318 261080 531374 261089
rect 531318 261015 531374 261024
rect 531516 258074 531544 267706
rect 531332 258046 531544 258074
rect 531332 243681 531360 258046
rect 531318 243672 531374 243681
rect 531318 243607 531374 243616
rect 530122 226264 530178 226273
rect 530044 226222 530122 226250
rect 530122 226199 530178 226208
rect 529938 209264 529994 209273
rect 529938 209199 529994 209208
rect 462412 201136 462464 201142
rect 462412 201078 462464 201084
rect 460756 200728 460808 200734
rect 460756 200670 460808 200676
rect 462320 200728 462372 200734
rect 462320 200670 462372 200676
rect 460676 200246 461072 200274
rect 460940 200184 460992 200190
rect 460940 200126 460992 200132
rect 459560 161492 459612 161498
rect 459560 161434 459612 161440
rect 460204 161492 460256 161498
rect 460204 161434 460256 161440
rect 459284 146260 459336 146266
rect 459284 146202 459336 146208
rect 460216 143546 460244 161434
rect 460204 143540 460256 143546
rect 460204 143482 460256 143488
rect 460848 143540 460900 143546
rect 460848 143482 460900 143488
rect 460860 142254 460888 143482
rect 460848 142248 460900 142254
rect 460848 142190 460900 142196
rect 459192 122052 459244 122058
rect 459192 121994 459244 122000
rect 457732 113146 458128 113174
rect 454684 107024 454736 107030
rect 454684 106966 454736 106972
rect 457732 104938 457760 113146
rect 389528 104910 389864 104938
rect 395692 104910 396028 104938
rect 401856 104910 402192 104938
rect 408020 104910 408448 104938
rect 414184 104910 414520 104938
rect 420348 104910 420684 104938
rect 426512 104910 426848 104938
rect 432676 104910 433012 104938
rect 438840 104910 439176 104938
rect 445004 104910 445340 104938
rect 451168 104910 451228 104938
rect 457332 104910 457760 104938
rect 386236 95192 386288 95198
rect 386236 95134 386288 95140
rect 460860 67697 460888 142190
rect 460294 67688 460350 67697
rect 460294 67623 460350 67632
rect 460846 67688 460902 67697
rect 460846 67623 460902 67632
rect 386144 62076 386196 62082
rect 386144 62018 386196 62024
rect 386144 51128 386196 51134
rect 386144 51070 386196 51076
rect 386052 34468 386104 34474
rect 386052 34410 386104 34416
rect 386156 31754 386184 51070
rect 460308 45554 460336 67623
rect 460216 45526 460336 45554
rect 460216 31754 460244 45526
rect 386144 31748 386196 31754
rect 386144 31690 386196 31696
rect 460204 31748 460256 31754
rect 460204 31690 460256 31696
rect 385960 31476 386012 31482
rect 385960 31418 386012 31424
rect 460952 28286 460980 200126
rect 461044 28422 461072 200246
rect 461584 199436 461636 199442
rect 461584 199378 461636 199384
rect 461596 41410 461624 199378
rect 461584 41404 461636 41410
rect 461584 41346 461636 41352
rect 462332 28490 462360 200670
rect 462320 28484 462372 28490
rect 462320 28426 462372 28432
rect 461032 28416 461084 28422
rect 461032 28358 461084 28364
rect 462424 28354 462452 201078
rect 528560 182844 528612 182850
rect 528560 182786 528612 182792
rect 524420 171828 524472 171834
rect 524420 171770 524472 171776
rect 485780 162308 485832 162314
rect 485780 162250 485832 162256
rect 481916 142248 481968 142254
rect 481916 142190 481968 142196
rect 481928 139890 481956 142190
rect 485792 139890 485820 162250
rect 489920 162172 489972 162178
rect 489920 162114 489972 162120
rect 489932 139890 489960 162114
rect 521660 160744 521712 160750
rect 521660 160686 521712 160692
rect 496820 160540 496872 160546
rect 496820 160482 496872 160488
rect 494060 160404 494112 160410
rect 494060 160346 494112 160352
rect 494072 139890 494100 160346
rect 496832 151814 496860 160482
rect 500960 160472 501012 160478
rect 500960 160414 501012 160420
rect 500972 151814 501000 160414
rect 509240 160336 509292 160342
rect 509240 160278 509292 160284
rect 505100 160268 505152 160274
rect 505100 160210 505152 160216
rect 505112 151814 505140 160210
rect 509252 151814 509280 160278
rect 513380 160200 513432 160206
rect 513380 160142 513432 160148
rect 513392 151814 513420 160142
rect 517520 160132 517572 160138
rect 517520 160074 517572 160080
rect 496832 151786 497688 151814
rect 500972 151786 501644 151814
rect 505112 151786 505600 151814
rect 509252 151786 509556 151814
rect 513392 151786 513512 151814
rect 497660 139890 497688 151786
rect 501616 139890 501644 151786
rect 505572 139890 505600 151786
rect 509528 139890 509556 151786
rect 513484 139890 513512 151786
rect 517532 139890 517560 160074
rect 521672 139890 521700 160686
rect 524432 151814 524460 171770
rect 528572 151814 528600 182786
rect 524432 151786 525380 151814
rect 528572 151786 529336 151814
rect 525352 139890 525380 151786
rect 529308 139890 529336 151786
rect 533356 140078 533384 319330
rect 539600 318300 539652 318306
rect 539600 318242 539652 318248
rect 533436 313948 533488 313954
rect 533436 313890 533488 313896
rect 533448 167006 533476 313890
rect 538864 311296 538916 311302
rect 538864 311238 538916 311244
rect 537484 309800 537536 309806
rect 537484 309742 537536 309748
rect 536840 284980 536892 284986
rect 536840 284922 536892 284928
rect 533436 167000 533488 167006
rect 533436 166942 533488 166948
rect 536852 151814 536880 284922
rect 537496 153202 537524 309742
rect 537484 153196 537536 153202
rect 537484 153138 537536 153144
rect 536852 151786 537248 151814
rect 533988 142180 534040 142186
rect 533988 142122 534040 142128
rect 533344 140072 533396 140078
rect 533344 140014 533396 140020
rect 534000 139890 534028 142122
rect 481928 139862 482264 139890
rect 485792 139862 486220 139890
rect 489932 139862 490176 139890
rect 494072 139862 494132 139890
rect 497660 139862 498088 139890
rect 501616 139862 502044 139890
rect 505572 139862 506000 139890
rect 509528 139862 509956 139890
rect 513484 139862 513912 139890
rect 517532 139862 517868 139890
rect 521672 139862 521824 139890
rect 525352 139862 525780 139890
rect 529308 139862 529736 139890
rect 533692 139862 534028 139890
rect 537220 139890 537248 151786
rect 537220 139862 537648 139890
rect 538876 137850 538904 311238
rect 538956 287768 539008 287774
rect 538956 287710 539008 287716
rect 538968 138009 538996 287710
rect 538954 138000 539010 138009
rect 538954 137935 539010 137944
rect 539414 137864 539470 137873
rect 538876 137822 538996 137850
rect 538968 136610 538996 137822
rect 539414 137799 539470 137808
rect 538956 136604 539008 136610
rect 538956 136546 539008 136552
rect 539428 129713 539456 137799
rect 539508 136604 539560 136610
rect 539508 136546 539560 136552
rect 539520 135969 539548 136546
rect 539506 135960 539562 135969
rect 539506 135895 539562 135904
rect 539414 129704 539470 129713
rect 539414 129639 539470 129648
rect 539612 95169 539640 318242
rect 540980 318232 541032 318238
rect 540980 318174 541032 318180
rect 539876 315376 539928 315382
rect 539876 315318 539928 315324
rect 539692 312588 539744 312594
rect 539692 312530 539744 312536
rect 539704 97209 539732 312530
rect 539784 308508 539836 308514
rect 539784 308450 539836 308456
rect 539796 99249 539824 308450
rect 539888 117337 539916 315318
rect 540244 283688 540296 283694
rect 540244 283630 540296 283636
rect 540152 280900 540204 280906
rect 540152 280842 540204 280848
rect 540060 274032 540112 274038
rect 540060 273974 540112 273980
rect 539968 272604 540020 272610
rect 539968 272546 540020 272552
rect 539874 117328 539930 117337
rect 539874 117263 539930 117272
rect 539980 108769 540008 272546
rect 540072 112849 540100 273974
rect 540164 127265 540192 280842
rect 540256 131345 540284 283630
rect 540336 275392 540388 275398
rect 540336 275334 540388 275340
rect 540242 131336 540298 131345
rect 540242 131271 540298 131280
rect 540150 127256 540206 127265
rect 540150 127191 540206 127200
rect 540348 125225 540376 275334
rect 540428 142180 540480 142186
rect 540428 142122 540480 142128
rect 540334 125216 540390 125225
rect 540334 125151 540390 125160
rect 540058 112840 540114 112849
rect 540058 112775 540114 112784
rect 539966 108760 540022 108769
rect 539966 108695 540022 108704
rect 539782 99240 539838 99249
rect 539782 99175 539838 99184
rect 539690 97200 539746 97209
rect 539690 97135 539746 97144
rect 539598 95160 539654 95169
rect 539598 95095 539654 95104
rect 536840 41404 536892 41410
rect 536840 41346 536892 41352
rect 536852 41041 536880 41346
rect 536838 41032 536894 41041
rect 536838 40967 536894 40976
rect 540440 34241 540468 142122
rect 540992 82385 541020 318174
rect 541072 317076 541124 317082
rect 541072 317018 541124 317024
rect 541084 110945 541112 317018
rect 543096 317008 543148 317014
rect 543096 316950 543148 316956
rect 542728 314084 542780 314090
rect 542728 314026 542780 314032
rect 542636 312656 542688 312662
rect 542636 312598 542688 312604
rect 542452 309868 542504 309874
rect 542452 309810 542504 309816
rect 541440 278044 541492 278050
rect 541440 277986 541492 277992
rect 541348 276684 541400 276690
rect 541348 276626 541400 276632
rect 541256 275324 541308 275330
rect 541256 275266 541308 275272
rect 541164 273964 541216 273970
rect 541164 273906 541216 273912
rect 541070 110936 541126 110945
rect 541070 110871 541126 110880
rect 541176 102785 541204 273906
rect 541268 104825 541296 275266
rect 541360 106865 541388 276626
rect 541452 115025 541480 277986
rect 541438 115016 541494 115025
rect 541438 114951 541494 114960
rect 541346 106856 541402 106865
rect 541346 106791 541402 106800
rect 541254 104816 541310 104825
rect 541254 104751 541310 104760
rect 541162 102776 541218 102785
rect 541162 102711 541218 102720
rect 542464 90545 542492 309810
rect 542544 140072 542596 140078
rect 542544 140014 542596 140020
rect 542556 100745 542584 140014
rect 542648 121145 542676 312598
rect 542740 123185 542768 314026
rect 543004 272536 543056 272542
rect 543004 272478 543056 272484
rect 542820 271244 542872 271250
rect 542820 271186 542872 271192
rect 542726 123176 542782 123185
rect 542726 123111 542782 123120
rect 542634 121136 542690 121145
rect 542634 121071 542690 121080
rect 542542 100736 542598 100745
rect 542542 100671 542598 100680
rect 542450 90536 542506 90545
rect 542450 90471 542506 90480
rect 542832 84425 542860 271186
rect 542912 268456 542964 268462
rect 542912 268398 542964 268404
rect 542924 86465 542952 268398
rect 543016 92585 543044 272478
rect 543108 119105 543136 316950
rect 543188 316872 543240 316878
rect 543188 316814 543240 316820
rect 543094 119096 543150 119105
rect 543094 119031 543150 119040
rect 543002 92576 543058 92585
rect 543002 92511 543058 92520
rect 543200 88505 543228 316814
rect 543186 88496 543242 88505
rect 543186 88431 543242 88440
rect 542910 86456 542966 86465
rect 542910 86391 542966 86400
rect 542818 84416 542874 84425
rect 542818 84351 542874 84360
rect 540978 82376 541034 82385
rect 540978 82311 541034 82320
rect 543752 51134 543780 319398
rect 569236 318714 569264 616830
rect 569316 430636 569368 430642
rect 569316 430578 569368 430584
rect 569328 321298 569356 430578
rect 569408 364404 569460 364410
rect 569408 364346 569460 364352
rect 569420 321366 569448 364346
rect 570616 321502 570644 670686
rect 570604 321496 570656 321502
rect 570604 321438 570656 321444
rect 569408 321360 569460 321366
rect 569408 321302 569460 321308
rect 569316 321292 569368 321298
rect 569316 321234 569368 321240
rect 571996 320142 572024 696934
rect 580170 683904 580226 683913
rect 580170 683839 580226 683848
rect 580184 683194 580212 683839
rect 573364 683188 573416 683194
rect 573364 683130 573416 683136
rect 580172 683188 580224 683194
rect 580172 683130 580224 683136
rect 573376 321434 573404 683130
rect 580172 670744 580224 670750
rect 580170 670712 580172 670721
rect 580224 670712 580226 670721
rect 580170 670647 580226 670656
rect 580262 644056 580318 644065
rect 580262 643991 580318 644000
rect 580170 617536 580226 617545
rect 580170 617471 580226 617480
rect 580184 616894 580212 617471
rect 580172 616888 580224 616894
rect 580172 616830 580224 616836
rect 580276 599622 580304 643991
rect 580354 630864 580410 630873
rect 580354 630799 580410 630808
rect 580264 599616 580316 599622
rect 580264 599558 580316 599564
rect 580170 591016 580226 591025
rect 580170 590951 580226 590960
rect 580184 590714 580212 590951
rect 580172 590708 580224 590714
rect 580172 590650 580224 590656
rect 580170 577688 580226 577697
rect 580170 577623 580226 577632
rect 580184 576910 580212 577623
rect 574744 576904 574796 576910
rect 574744 576846 574796 576852
rect 580172 576904 580224 576910
rect 580172 576846 580224 576852
rect 574756 321978 574784 576846
rect 580262 564360 580318 564369
rect 580262 564295 580318 564304
rect 580170 537840 580226 537849
rect 580170 537775 580226 537784
rect 580184 536858 580212 537775
rect 580172 536852 580224 536858
rect 580172 536794 580224 536800
rect 580170 484664 580226 484673
rect 580170 484599 580226 484608
rect 580184 484430 580212 484599
rect 580172 484424 580224 484430
rect 580172 484366 580224 484372
rect 580170 458144 580226 458153
rect 580170 458079 580226 458088
rect 580184 456822 580212 458079
rect 576124 456816 576176 456822
rect 576124 456758 576176 456764
rect 580172 456816 580224 456822
rect 580172 456758 580224 456764
rect 574744 321972 574796 321978
rect 574744 321914 574796 321920
rect 573364 321428 573416 321434
rect 573364 321370 573416 321376
rect 571984 320136 572036 320142
rect 571984 320078 572036 320084
rect 576136 318782 576164 456758
rect 580170 431624 580226 431633
rect 580170 431559 580226 431568
rect 580184 430642 580212 431559
rect 580172 430636 580224 430642
rect 580172 430578 580224 430584
rect 580170 404968 580226 404977
rect 580170 404903 580226 404912
rect 580184 404394 580212 404903
rect 580172 404388 580224 404394
rect 580172 404330 580224 404336
rect 580170 365120 580226 365129
rect 580170 365055 580226 365064
rect 580184 364410 580212 365055
rect 580172 364404 580224 364410
rect 580172 364346 580224 364352
rect 580172 352096 580224 352102
rect 580172 352038 580224 352044
rect 580184 351937 580212 352038
rect 580170 351928 580226 351937
rect 580170 351863 580226 351872
rect 580170 325272 580226 325281
rect 580170 325207 580226 325216
rect 580184 321910 580212 325207
rect 580172 321904 580224 321910
rect 580172 321846 580224 321852
rect 580276 321570 580304 564295
rect 580368 421598 580396 630799
rect 580446 524512 580502 524521
rect 580446 524447 580502 524456
rect 580356 421592 580408 421598
rect 580356 421534 580408 421540
rect 580354 418296 580410 418305
rect 580354 418231 580410 418240
rect 580368 323610 580396 418231
rect 580356 323604 580408 323610
rect 580356 323546 580408 323552
rect 580460 322250 580488 524447
rect 580538 511320 580594 511329
rect 580538 511255 580594 511264
rect 580448 322244 580500 322250
rect 580448 322186 580500 322192
rect 580264 321564 580316 321570
rect 580264 321506 580316 321512
rect 580552 320890 580580 511255
rect 580630 471472 580686 471481
rect 580630 471407 580686 471416
rect 580644 324970 580672 471407
rect 580722 378448 580778 378457
rect 580722 378383 580778 378392
rect 580632 324964 580684 324970
rect 580632 324906 580684 324912
rect 580736 320958 580764 378383
rect 580724 320952 580776 320958
rect 580724 320894 580776 320900
rect 580540 320884 580592 320890
rect 580540 320826 580592 320832
rect 576124 318776 576176 318782
rect 576124 318718 576176 318724
rect 569224 318708 569276 318714
rect 569224 318650 569276 318656
rect 580172 313268 580224 313274
rect 580172 313210 580224 313216
rect 580184 312089 580212 313210
rect 580170 312080 580226 312089
rect 580170 312015 580226 312024
rect 544384 311160 544436 311166
rect 544384 311102 544436 311108
rect 544396 73166 544424 311102
rect 548524 308440 548576 308446
rect 548524 308382 548576 308388
rect 547144 302864 547196 302870
rect 547144 302806 547196 302812
rect 547156 193186 547184 302806
rect 547144 193180 547196 193186
rect 547144 193122 547196 193128
rect 544384 73160 544436 73166
rect 544384 73102 544436 73108
rect 548536 60722 548564 308382
rect 576124 307148 576176 307154
rect 576124 307090 576176 307096
rect 562324 305924 562376 305930
rect 562324 305866 562376 305872
rect 559564 301708 559616 301714
rect 559564 301650 559616 301656
rect 551284 299940 551336 299946
rect 551284 299882 551336 299888
rect 551296 179382 551324 299882
rect 558184 293276 558236 293282
rect 558184 293218 558236 293224
rect 555424 269884 555476 269890
rect 555424 269826 555476 269832
rect 551284 179376 551336 179382
rect 551284 179318 551336 179324
rect 555436 139398 555464 269826
rect 558196 233238 558224 293218
rect 558184 233232 558236 233238
rect 558184 233174 558236 233180
rect 555424 139392 555476 139398
rect 555424 139334 555476 139340
rect 559576 100706 559604 301650
rect 559564 100700 559616 100706
rect 559564 100642 559616 100648
rect 548524 60716 548576 60722
rect 548524 60658 548576 60664
rect 540612 51128 540664 51134
rect 540612 51070 540664 51076
rect 543740 51128 543792 51134
rect 543740 51070 543792 51076
rect 540624 48929 540652 51070
rect 540610 48920 540666 48929
rect 540610 48855 540666 48864
rect 540426 34232 540482 34241
rect 540426 34167 540482 34176
rect 562336 33114 562364 305866
rect 566464 298104 566516 298110
rect 566464 298046 566516 298052
rect 562324 33108 562376 33114
rect 562324 33050 562376 33056
rect 462412 28348 462464 28354
rect 462412 28290 462464 28296
rect 460940 28280 460992 28286
rect 460940 28222 460992 28228
rect 566476 6866 566504 298046
rect 573364 295996 573416 296002
rect 573364 295938 573416 295944
rect 570604 294432 570656 294438
rect 570604 294374 570656 294380
rect 569224 290488 569276 290494
rect 569224 290430 569276 290436
rect 569236 113150 569264 290430
rect 569224 113144 569276 113150
rect 569224 113086 569276 113092
rect 570616 86970 570644 294374
rect 572076 291712 572128 291718
rect 572076 291654 572128 291660
rect 571984 286544 572036 286550
rect 571984 286486 572036 286492
rect 570604 86964 570656 86970
rect 570604 86906 570656 86912
rect 571996 20670 572024 286486
rect 572088 245614 572116 291654
rect 572076 245608 572128 245614
rect 572076 245550 572128 245556
rect 573376 46918 573404 295938
rect 574744 288924 574796 288930
rect 574744 288866 574796 288872
rect 574756 126954 574784 288866
rect 576136 206990 576164 307090
rect 580172 299464 580224 299470
rect 580172 299406 580224 299412
rect 580184 298761 580212 299406
rect 580170 298752 580226 298761
rect 580170 298687 580226 298696
rect 580264 283620 580316 283626
rect 580264 283562 580316 283568
rect 580276 272241 580304 283562
rect 580262 272232 580318 272241
rect 580262 272167 580318 272176
rect 580356 271176 580408 271182
rect 580356 271118 580408 271124
rect 580264 269816 580316 269822
rect 580264 269758 580316 269764
rect 580172 245608 580224 245614
rect 580170 245576 580172 245585
rect 580224 245576 580226 245585
rect 580170 245511 580226 245520
rect 580172 233232 580224 233238
rect 580172 233174 580224 233180
rect 580184 232393 580212 233174
rect 580170 232384 580226 232393
rect 580170 232319 580226 232328
rect 580276 219065 580304 269758
rect 580368 258913 580396 271118
rect 580354 258904 580410 258913
rect 580354 258839 580410 258848
rect 580262 219056 580318 219065
rect 580262 218991 580318 219000
rect 576124 206984 576176 206990
rect 576124 206926 576176 206932
rect 579804 206984 579856 206990
rect 579804 206926 579856 206932
rect 579816 205737 579844 206926
rect 579802 205728 579858 205737
rect 579802 205663 579858 205672
rect 580172 193180 580224 193186
rect 580172 193122 580224 193128
rect 580184 192545 580212 193122
rect 580170 192536 580226 192545
rect 580170 192471 580226 192480
rect 580172 179376 580224 179382
rect 580172 179318 580224 179324
rect 580184 179217 580212 179318
rect 580170 179208 580226 179217
rect 580170 179143 580226 179152
rect 580172 167000 580224 167006
rect 580172 166942 580224 166948
rect 580184 165889 580212 166942
rect 580170 165880 580226 165889
rect 580170 165815 580226 165824
rect 580172 153196 580224 153202
rect 580172 153138 580224 153144
rect 580184 152697 580212 153138
rect 580170 152688 580226 152697
rect 580170 152623 580226 152632
rect 580172 139392 580224 139398
rect 580170 139360 580172 139369
rect 580224 139360 580226 139369
rect 580170 139295 580226 139304
rect 574744 126948 574796 126954
rect 574744 126890 574796 126896
rect 580172 126948 580224 126954
rect 580172 126890 580224 126896
rect 580184 126041 580212 126890
rect 580170 126032 580226 126041
rect 580170 125967 580226 125976
rect 579804 113144 579856 113150
rect 579804 113086 579856 113092
rect 579816 112849 579844 113086
rect 579802 112840 579858 112849
rect 579802 112775 579858 112784
rect 580172 100700 580224 100706
rect 580172 100642 580224 100648
rect 580184 99521 580212 100642
rect 580170 99512 580226 99521
rect 580170 99447 580226 99456
rect 580172 86964 580224 86970
rect 580172 86906 580224 86912
rect 580184 86193 580212 86906
rect 580170 86184 580226 86193
rect 580170 86119 580226 86128
rect 580172 73160 580224 73166
rect 580172 73102 580224 73108
rect 580184 73001 580212 73102
rect 580170 72992 580226 73001
rect 580170 72927 580226 72936
rect 580172 60716 580224 60722
rect 580172 60658 580224 60664
rect 580184 59673 580212 60658
rect 580170 59664 580226 59673
rect 580170 59599 580226 59608
rect 573364 46912 573416 46918
rect 573364 46854 573416 46860
rect 580172 46912 580224 46918
rect 580172 46854 580224 46860
rect 580184 46345 580212 46854
rect 580170 46336 580226 46345
rect 580170 46271 580226 46280
rect 580170 33144 580226 33153
rect 580170 33079 580172 33088
rect 580224 33079 580226 33088
rect 580172 33050 580224 33056
rect 571984 20664 572036 20670
rect 571984 20606 572036 20612
rect 579988 20664 580040 20670
rect 579988 20606 580040 20612
rect 580000 19825 580028 20606
rect 579986 19816 580042 19825
rect 579986 19751 580042 19760
rect 566464 6860 566516 6866
rect 566464 6802 566516 6808
rect 580172 6860 580224 6866
rect 580172 6802 580224 6808
rect 580184 6633 580212 6802
rect 580170 6624 580226 6633
rect 580170 6559 580226 6568
rect 385868 3528 385920 3534
rect 385868 3470 385920 3476
rect 381726 3431 381782 3440
rect 385776 3460 385828 3466
rect 385776 3402 385828 3408
rect 360844 3198 360896 3204
rect 365074 3224 365130 3233
rect 365074 3159 365130 3168
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9926 -960 10038 480
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14710 -960 14822 480
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 18206 -960 18318 480
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22990 -960 23102 480
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26486 -960 26598 480
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 31270 -960 31382 480
rect 32374 -960 32486 480
rect 33570 -960 33682 480
rect 34766 -960 34878 480
rect 35962 -960 36074 480
rect 37158 -960 37270 480
rect 38354 -960 38466 480
rect 39550 -960 39662 480
rect 40654 -960 40766 480
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45438 -960 45550 480
rect 46634 -960 46746 480
rect 47830 -960 47942 480
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53718 -960 53830 480
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 57214 -960 57326 480
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61998 -960 62110 480
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67886 -960 67998 480
rect 69082 -960 69194 480
rect 70278 -960 70390 480
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 76166 -960 76278 480
rect 77362 -960 77474 480
rect 78558 -960 78670 480
rect 79662 -960 79774 480
rect 80858 -960 80970 480
rect 82054 -960 82166 480
rect 83250 -960 83362 480
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 86838 -960 86950 480
rect 87942 -960 88054 480
rect 89138 -960 89250 480
rect 90334 -960 90446 480
rect 91530 -960 91642 480
rect 92726 -960 92838 480
rect 93922 -960 94034 480
rect 95118 -960 95230 480
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98614 -960 98726 480
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104502 -960 104614 480
rect 105698 -960 105810 480
rect 106894 -960 107006 480
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112782 -960 112894 480
rect 113978 -960 114090 480
rect 115174 -960 115286 480
rect 116370 -960 116482 480
rect 117566 -960 117678 480
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 123454 -960 123566 480
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 148294 -960 148406 480
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 174238 -960 174350 480
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 179022 -960 179134 480
rect 180218 -960 180330 480
rect 181414 -960 181526 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 199078 -960 199190 480
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220422 -960 220534 480
rect 221526 -960 221638 480
rect 222722 -960 222834 480
rect 223918 -960 224030 480
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236982 -960 237094 480
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248758 -960 248870 480
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273598 -960 273710 480
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 279486 -960 279598 480
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293654 -960 293766 480
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 304326 -960 304438 480
rect 305522 -960 305634 480
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318494 -960 318606 480
rect 319690 -960 319802 480
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 354006 -960 354118 480
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370566 -960 370678 480
rect 371670 -960 371782 480
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 378846 -960 378958 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 387126 -960 387238 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396510 -960 396622 480
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409574 -960 409686 480
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 413070 -960 413182 480
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417854 -960 417966 480
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 421350 -960 421462 480
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 427238 -960 427350 480
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435518 -960 435630 480
rect 436714 -960 436826 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 446190 -960 446302 480
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 460358 -960 460470 480
rect 461554 -960 461666 480
rect 462750 -960 462862 480
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 471030 -960 471142 480
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474526 -960 474638 480
rect 475722 -960 475834 480
rect 476918 -960 477030 480
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482806 -960 482918 480
rect 484002 -960 484114 480
rect 485198 -960 485310 480
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 491086 -960 491198 480
rect 492282 -960 492394 480
rect 493478 -960 493590 480
rect 494674 -960 494786 480
rect 495870 -960 495982 480
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499366 -960 499478 480
rect 500562 -960 500674 480
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 504150 -960 504262 480
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507646 -960 507758 480
rect 508842 -960 508954 480
rect 510038 -960 510150 480
rect 511234 -960 511346 480
rect 512430 -960 512542 480
rect 513534 -960 513646 480
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 518318 -960 518430 480
rect 519514 -960 519626 480
rect 520710 -960 520822 480
rect 521814 -960 521926 480
rect 523010 -960 523122 480
rect 524206 -960 524318 480
rect 525402 -960 525514 480
rect 526598 -960 526710 480
rect 527794 -960 527906 480
rect 528990 -960 529102 480
rect 530094 -960 530206 480
rect 531290 -960 531402 480
rect 532486 -960 532598 480
rect 533682 -960 533794 480
rect 534878 -960 534990 480
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538374 -960 538486 480
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 543158 -960 543270 480
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546654 -960 546766 480
rect 547850 -960 547962 480
rect 549046 -960 549158 480
rect 550242 -960 550354 480
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 557326 -960 557438 480
rect 558522 -960 558634 480
rect 559718 -960 559830 480
rect 560822 -960 560934 480
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564410 -960 564522 480
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 40498 700304 40554 700360
rect 24306 686432 24362 686488
rect 202786 700440 202842 700496
rect 300122 689288 300178 689344
rect 3238 684256 3294 684312
rect 3146 658180 3148 658200
rect 3148 658180 3200 658200
rect 3200 658180 3202 658200
rect 3146 658144 3202 658180
rect 3238 579944 3294 580000
rect 3330 566888 3386 566944
rect 3698 632032 3754 632088
rect 3606 475632 3662 475688
rect 3514 462576 3570 462632
rect 3422 449520 3478 449576
rect 4066 553832 4122 553888
rect 3974 527856 4030 527912
rect 3882 514800 3938 514856
rect 361762 678988 361764 679008
rect 361764 678988 361816 679008
rect 361816 678988 361818 679008
rect 361762 678952 361818 678988
rect 361762 667956 361818 667992
rect 361762 667936 361764 667956
rect 361764 667936 361816 667956
rect 361816 667936 361818 667956
rect 361762 656940 361818 656976
rect 361762 656920 361764 656940
rect 361764 656920 361816 656940
rect 361816 656920 361818 656940
rect 361762 645924 361818 645960
rect 361762 645904 361764 645924
rect 361764 645904 361816 645924
rect 361816 645904 361818 645924
rect 361578 634888 361634 634944
rect 361578 623872 361634 623928
rect 361578 612856 361634 612912
rect 361762 601840 361818 601896
rect 361762 590824 361818 590880
rect 361762 579808 361818 579864
rect 361578 568812 361634 568848
rect 361578 568792 361580 568812
rect 361580 568792 361632 568812
rect 361632 568792 361634 568812
rect 361670 557776 361726 557832
rect 361762 546760 361818 546816
rect 361578 535744 361634 535800
rect 361578 524748 361634 524784
rect 361578 524728 361580 524748
rect 361580 524728 361632 524748
rect 361632 524728 361634 524748
rect 3790 501744 3846 501800
rect 3698 423544 3754 423600
rect 361762 513712 361818 513768
rect 361762 502696 361818 502752
rect 361762 491680 361818 491736
rect 361762 480664 361818 480720
rect 361762 469648 361818 469704
rect 361762 458632 361818 458688
rect 362222 447616 362278 447672
rect 361762 436600 361818 436656
rect 362314 425584 362370 425640
rect 361578 414568 361634 414624
rect 3974 410488 4030 410544
rect 361578 403552 361634 403608
rect 3790 397432 3846 397488
rect 3514 358400 3570 358456
rect 3422 345344 3478 345400
rect 3606 306176 3662 306232
rect 3422 267144 3478 267200
rect 3330 162832 3386 162888
rect 3238 149776 3294 149832
rect 3054 98640 3110 98696
rect 3514 254088 3570 254144
rect 3422 45464 3478 45520
rect 3698 293120 3754 293176
rect 361578 392536 361634 392592
rect 361578 381520 361634 381576
rect 3882 371320 3938 371376
rect 3790 241032 3846 241088
rect 3698 84632 3754 84688
rect 3606 71576 3662 71632
rect 3606 58520 3662 58576
rect 361578 370504 361634 370560
rect 362222 359488 362278 359544
rect 361762 348472 361818 348528
rect 361762 337456 361818 337512
rect 362222 326440 362278 326496
rect 3974 319232 4030 319288
rect 361762 315424 361818 315480
rect 3882 214920 3938 214976
rect 3974 201864 4030 201920
rect 4066 188808 4122 188864
rect 360842 305632 360898 305688
rect 20902 73616 20958 73672
rect 11702 48864 11758 48920
rect 19246 49544 19302 49600
rect 21454 73616 21510 73672
rect 359554 46416 359610 46472
rect 2870 32408 2926 32464
rect 3422 19352 3478 19408
rect 3422 6432 3478 6488
rect 2870 3576 2926 3632
rect 1674 3440 1730 3496
rect 570 3304 626 3360
rect 8758 3984 8814 4040
rect 9954 3712 10010 3768
rect 13542 3848 13598 3904
rect 17038 3168 17094 3224
rect 361762 304408 361818 304464
rect 362222 302776 362278 302832
rect 361762 293392 361818 293448
rect 361762 282376 361818 282432
rect 361762 271360 361818 271416
rect 361762 260344 361818 260400
rect 361762 249328 361818 249384
rect 361762 238312 361818 238368
rect 361762 227296 361818 227352
rect 361670 216316 361672 216336
rect 361672 216316 361724 216336
rect 361724 216316 361726 216336
rect 361670 216280 361726 216316
rect 361762 205264 361818 205320
rect 361762 194248 361818 194304
rect 361762 183232 361818 183288
rect 361762 172216 361818 172272
rect 361762 161200 361818 161256
rect 361762 150184 361818 150240
rect 361762 139168 361818 139224
rect 361302 46552 361358 46608
rect 361762 128152 361818 128208
rect 361762 117136 361818 117192
rect 361762 106120 361818 106176
rect 361762 95140 361764 95160
rect 361764 95140 361816 95160
rect 361816 95140 361818 95160
rect 361762 95104 361818 95140
rect 361762 84124 361764 84144
rect 361764 84124 361816 84144
rect 361816 84124 361818 84144
rect 361762 84088 361818 84124
rect 361762 73108 361764 73128
rect 361764 73108 361816 73128
rect 361816 73108 361818 73128
rect 361762 73072 361818 73108
rect 361762 62076 361818 62112
rect 361762 62056 361764 62076
rect 361764 62056 361816 62076
rect 361816 62056 361818 62076
rect 361762 51076 361764 51096
rect 361764 51076 361816 51096
rect 361816 51076 361818 51096
rect 361762 51040 361818 51076
rect 362222 3984 362278 4040
rect 363694 302912 363750 302968
rect 363786 297336 363842 297392
rect 367834 305768 367890 305824
rect 365166 297608 365222 297664
rect 368202 297472 368258 297528
rect 374734 286320 374790 286376
rect 374642 3848 374698 3904
rect 381542 306040 381598 306096
rect 381450 303048 381506 303104
rect 374826 3712 374882 3768
rect 381726 305904 381782 305960
rect 381542 3576 381598 3632
rect 384302 46688 384358 46744
rect 384486 46824 384542 46880
rect 384854 291760 384910 291816
rect 381726 3440 381782 3496
rect 429842 700576 429898 700632
rect 420090 682760 420146 682816
rect 427818 337048 427874 337104
rect 428094 334464 428150 334520
rect 420458 334328 420514 334384
rect 424138 334328 424194 334384
rect 421838 162696 421894 162752
rect 425886 162696 425942 162752
rect 428646 162696 428702 162752
rect 432786 332832 432842 332888
rect 432694 329160 432750 329216
rect 432602 325488 432658 325544
rect 432786 321816 432842 321872
rect 432694 318144 432750 318200
rect 432602 314472 432658 314528
rect 432050 310800 432106 310856
rect 432694 307128 432750 307184
rect 439962 322632 440018 322688
rect 442446 320048 442502 320104
rect 442722 321136 442778 321192
rect 444194 421912 444250 421968
rect 444838 322768 444894 322824
rect 446862 683304 446918 683360
rect 447046 683168 447102 683224
rect 447138 383832 447194 383888
rect 447138 383152 447194 383208
rect 447230 382472 447286 382528
rect 447138 381792 447194 381848
rect 447230 381112 447286 381168
rect 447138 380432 447194 380488
rect 447230 379752 447286 379808
rect 447138 379072 447194 379128
rect 447230 378392 447286 378448
rect 447138 377712 447194 377768
rect 447230 377032 447286 377088
rect 447138 376352 447194 376408
rect 447230 375672 447286 375728
rect 447138 374992 447194 375048
rect 447230 374312 447286 374368
rect 447138 373632 447194 373688
rect 447230 372952 447286 373008
rect 447138 372272 447194 372328
rect 447230 371592 447286 371648
rect 447138 370912 447194 370968
rect 447230 370232 447286 370288
rect 447138 369552 447194 369608
rect 447230 368872 447286 368928
rect 447230 368192 447286 368248
rect 447138 367512 447194 367568
rect 447138 366832 447194 366888
rect 447230 366152 447286 366208
rect 447230 365472 447286 365528
rect 447138 364792 447194 364848
rect 447230 364112 447286 364168
rect 447138 363432 447194 363488
rect 447138 362752 447194 362808
rect 447230 362072 447286 362128
rect 447230 361392 447286 361448
rect 447138 360712 447194 360768
rect 447138 360032 447194 360088
rect 447230 359352 447286 359408
rect 447414 355952 447470 356008
rect 447690 354592 447746 354648
rect 447598 353912 447654 353968
rect 447874 353232 447930 353288
rect 447138 351908 447140 351928
rect 447140 351908 447192 351928
rect 447192 351908 447194 351928
rect 447138 351872 447194 351908
rect 447138 350548 447140 350568
rect 447140 350548 447192 350568
rect 447192 350548 447194 350568
rect 447138 350512 447194 350548
rect 447598 349832 447654 349888
rect 447138 347112 447194 347168
rect 447230 341672 447286 341728
rect 447138 341012 447194 341048
rect 447138 340992 447140 341012
rect 447140 340992 447192 341012
rect 447192 340992 447194 341012
rect 447230 340312 447286 340368
rect 447138 339632 447194 339688
rect 447230 338952 447286 339008
rect 447138 338272 447194 338328
rect 447138 337592 447194 337648
rect 447230 336912 447286 336968
rect 447138 336232 447194 336288
rect 447138 335552 447194 335608
rect 447230 334872 447286 334928
rect 447138 334192 447194 334248
rect 447230 333512 447286 333568
rect 447138 332832 447194 332888
rect 447138 330132 447194 330168
rect 447138 330112 447140 330132
rect 447140 330112 447192 330132
rect 447192 330112 447194 330132
rect 447138 329432 447194 329488
rect 447046 322496 447102 322552
rect 447782 330792 447838 330848
rect 448242 355272 448298 355328
rect 448150 352552 448206 352608
rect 448242 351192 448298 351248
rect 448150 332152 448206 332208
rect 448058 330112 448114 330168
rect 447966 329432 448022 329488
rect 448334 348472 448390 348528
rect 448334 344392 448390 344448
rect 449070 386960 449126 387016
rect 448978 358672 449034 358728
rect 449070 357312 449126 357368
rect 448426 343032 448482 343088
rect 448334 331472 448390 331528
rect 448426 330792 448482 330848
rect 543462 700304 543518 700360
rect 527178 699760 527234 699816
rect 559654 699760 559710 699816
rect 580170 697176 580226 697232
rect 460202 668072 460258 668128
rect 458086 659912 458142 659968
rect 457810 657464 457866 657520
rect 457718 652840 457774 652896
rect 457626 650120 457682 650176
rect 457534 645904 457590 645960
rect 457442 643184 457498 643240
rect 457350 623872 457406 623928
rect 457258 621016 457314 621072
rect 450450 516840 450506 516896
rect 450450 514664 450506 514720
rect 457994 635432 458050 635488
rect 457902 618296 457958 618352
rect 459374 647672 459430 647728
rect 459282 640328 459338 640384
rect 459190 637880 459246 637936
rect 459098 633392 459154 633448
rect 459006 630672 459062 630728
rect 458822 615984 458878 616040
rect 458730 611360 458786 611416
rect 458638 608640 458694 608696
rect 458914 614080 458970 614136
rect 459190 599528 459246 599584
rect 459098 598168 459154 598224
rect 459006 595584 459062 595640
rect 459466 628088 459522 628144
rect 459374 591232 459430 591288
rect 459282 589872 459338 589928
rect 460110 625776 460166 625832
rect 460018 606328 460074 606384
rect 459926 603608 459982 603664
rect 459834 601840 459890 601896
rect 450542 512352 450598 512408
rect 450358 510176 450414 510232
rect 449990 507592 450046 507648
rect 449806 503444 449862 503500
rect 449346 347792 449402 347848
rect 449346 343712 449402 343768
rect 449530 357992 449586 358048
rect 449622 356632 449678 356688
rect 449714 346432 449770 346488
rect 449806 345752 449862 345808
rect 449806 345072 449862 345128
rect 449438 342352 449494 342408
rect 450082 505416 450138 505472
rect 450174 503240 450230 503296
rect 450266 338000 450322 338056
rect 450266 337048 450322 337104
rect 449990 333920 450046 333976
rect 449898 328500 449954 328536
rect 449898 328480 449900 328500
rect 449900 328480 449952 328500
rect 449952 328480 449954 328500
rect 449898 327800 449954 327856
rect 449990 326168 450046 326224
rect 450266 327528 450322 327584
rect 450634 505416 450690 505472
rect 450542 338000 450598 338056
rect 461766 597624 461822 597680
rect 463054 501064 463110 501120
rect 464342 388320 464398 388376
rect 467102 518064 467158 518120
rect 482742 517520 482798 517576
rect 494058 515480 494114 515536
rect 492126 512420 492182 512476
rect 494150 508816 494206 508872
rect 500958 516840 501014 516896
rect 502246 516840 502302 516896
rect 507122 516704 507178 516760
rect 494242 505688 494298 505744
rect 495070 505724 495072 505744
rect 495072 505724 495124 505744
rect 495124 505724 495126 505744
rect 495070 505688 495126 505724
rect 494702 501200 494758 501256
rect 473726 462848 473782 462904
rect 489182 496848 489238 496904
rect 472162 389000 472218 389056
rect 474370 389000 474426 389056
rect 475106 389000 475162 389056
rect 477314 389000 477370 389056
rect 479522 389000 479578 389056
rect 472898 388864 472954 388920
rect 509698 370096 509754 370152
rect 450450 334328 450506 334384
rect 450450 326848 450506 326904
rect 509882 360304 509938 360360
rect 450450 325488 450506 325544
rect 450358 324400 450414 324456
rect 450082 324128 450138 324184
rect 450634 323720 450690 323776
rect 509698 322904 509754 322960
rect 471058 322632 471114 322688
rect 482374 322632 482430 322688
rect 471886 322496 471942 322552
rect 459190 322360 459246 322416
rect 451738 158208 451794 158264
rect 451738 156848 451794 156904
rect 451830 145968 451886 146024
rect 451554 144608 451610 144664
rect 451554 139204 451556 139224
rect 451556 139204 451608 139224
rect 451608 139204 451610 139224
rect 451554 139168 451610 139204
rect 451554 136484 451556 136504
rect 451556 136484 451608 136504
rect 451608 136484 451610 136504
rect 451554 136448 451610 136484
rect 452014 148688 452070 148744
rect 452014 135124 452016 135144
rect 452016 135124 452068 135144
rect 452068 135124 452070 135144
rect 452014 135088 452070 135124
rect 452198 155488 452254 155544
rect 452474 154128 452530 154184
rect 452474 152768 452530 152824
rect 452566 151444 452568 151464
rect 452568 151444 452620 151464
rect 452620 151444 452622 151464
rect 452566 151408 452622 151444
rect 452382 150048 452438 150104
rect 452566 147364 452568 147384
rect 452568 147364 452620 147384
rect 452620 147364 452622 147384
rect 452566 147328 452622 147364
rect 452566 143248 452622 143304
rect 452566 141924 452568 141944
rect 452568 141924 452620 141944
rect 452620 141924 452622 141944
rect 452566 141888 452622 141924
rect 452566 140528 452622 140584
rect 452566 137844 452568 137864
rect 452568 137844 452620 137864
rect 452620 137844 452622 137864
rect 452566 137808 452622 137844
rect 452290 133728 452346 133784
rect 451922 128288 451978 128344
rect 451738 125568 451794 125624
rect 452290 132404 452292 132424
rect 452292 132404 452344 132424
rect 452344 132404 452346 132424
rect 452290 132368 452346 132404
rect 452566 131044 452568 131064
rect 452568 131044 452620 131064
rect 452620 131044 452622 131064
rect 452566 131008 452622 131044
rect 452106 129684 452108 129704
rect 452108 129684 452160 129704
rect 452160 129684 452162 129704
rect 452106 129648 452162 129684
rect 452566 126948 452622 126984
rect 452566 126928 452568 126948
rect 452568 126928 452620 126948
rect 452620 126928 452622 126948
rect 452014 124208 452070 124264
rect 451738 122848 451794 122904
rect 451922 121488 451978 121544
rect 456062 318008 456118 318064
rect 458638 320592 458694 320648
rect 460570 321408 460626 321464
rect 460846 321272 460902 321328
rect 459742 319776 459798 319832
rect 460570 318280 460626 318336
rect 456798 262656 456854 262712
rect 456798 248784 456854 248840
rect 457994 234912 458050 234968
rect 457810 221040 457866 221096
rect 459466 318144 459522 318200
rect 459558 207168 459614 207224
rect 469126 321272 469182 321328
rect 471334 319912 471390 319968
rect 480994 321000 481050 321056
rect 481822 321136 481878 321192
rect 481546 320048 481602 320104
rect 501142 315288 501198 315344
rect 501694 313928 501750 313984
rect 507122 321816 507178 321872
rect 507306 321544 507362 321600
rect 509698 320728 509754 320784
rect 507582 320184 507638 320240
rect 511078 359624 511134 359680
rect 510618 359080 510674 359136
rect 509974 357584 510030 357640
rect 510066 356360 510122 356416
rect 510250 330248 510306 330304
rect 510158 324944 510214 325000
rect 510342 328072 510398 328128
rect 510158 318144 510214 318200
rect 510894 355816 510950 355872
rect 510710 353096 510766 353152
rect 510894 344392 510950 344448
rect 510986 342760 511042 342816
rect 511170 348744 511226 348800
rect 512090 377576 512146 377632
rect 513286 384648 513342 384704
rect 512458 384104 512514 384160
rect 512642 383560 512698 383616
rect 513010 383016 513066 383072
rect 512458 382492 512514 382528
rect 512458 382472 512460 382492
rect 512460 382472 512512 382492
rect 512512 382472 512514 382492
rect 513102 381928 513158 381984
rect 512550 379772 512606 379808
rect 512550 379752 512552 379772
rect 512552 379752 512604 379772
rect 512604 379752 512606 379772
rect 512918 379208 512974 379264
rect 512458 378664 512514 378720
rect 512274 378120 512330 378176
rect 512642 377032 512698 377088
rect 512182 376488 512238 376544
rect 513286 381384 513342 381440
rect 513194 380840 513250 380896
rect 513286 380296 513342 380352
rect 512642 375944 512698 376000
rect 512826 375436 512828 375456
rect 512828 375436 512880 375456
rect 512880 375436 512882 375456
rect 512826 375400 512882 375436
rect 511998 374856 512054 374912
rect 513286 374312 513342 374368
rect 512642 373788 512698 373824
rect 512642 373768 512644 373788
rect 512644 373768 512696 373788
rect 512696 373768 512698 373788
rect 512458 373224 512514 373280
rect 512090 372700 512146 372736
rect 512090 372680 512092 372700
rect 512092 372680 512144 372700
rect 512144 372680 512146 372700
rect 512826 372136 512882 372192
rect 512182 371592 512238 371648
rect 512090 368328 512146 368384
rect 511998 367784 512054 367840
rect 511998 366172 512054 366208
rect 511998 366152 512000 366172
rect 512000 366152 512052 366172
rect 512052 366152 512054 366172
rect 512642 371048 512698 371104
rect 513286 369960 513342 370016
rect 513286 369416 513342 369472
rect 512826 368872 512882 368928
rect 513286 367260 513342 367296
rect 513286 367240 513288 367260
rect 513288 367240 513340 367260
rect 513340 367240 513342 367260
rect 513286 366696 513342 366752
rect 513286 365608 513342 365664
rect 512642 365064 512698 365120
rect 513286 364540 513342 364576
rect 513286 364520 513288 364540
rect 513288 364520 513340 364540
rect 513340 364520 513342 364540
rect 512182 363976 512238 364032
rect 513286 363432 513342 363488
rect 513010 362888 513066 362944
rect 512182 362364 512238 362400
rect 512182 362344 512184 362364
rect 512184 362344 512236 362364
rect 512236 362344 512238 362364
rect 512366 361800 512422 361856
rect 512274 358536 512330 358592
rect 512182 357992 512238 358048
rect 512090 305632 512146 305688
rect 513010 361256 513066 361312
rect 513286 360204 513288 360224
rect 513288 360204 513340 360224
rect 513340 360204 513342 360224
rect 513286 360168 513342 360204
rect 513286 356904 513342 356960
rect 512366 355272 512422 355328
rect 513286 354748 513342 354784
rect 513286 354728 513288 354748
rect 513288 354728 513340 354748
rect 513340 354728 513342 354748
rect 512458 354184 512514 354240
rect 513194 353640 513250 353696
rect 512458 352572 512514 352608
rect 512458 352552 512460 352572
rect 512460 352552 512512 352572
rect 512512 352552 512514 352572
rect 513286 352028 513342 352064
rect 513286 352008 513288 352028
rect 513288 352008 513340 352028
rect 513340 352008 513342 352028
rect 513286 351464 513342 351520
rect 512458 350920 512514 350976
rect 512458 350376 512514 350432
rect 513286 349832 513342 349888
rect 512458 349288 512514 349344
rect 513010 348200 513066 348256
rect 512458 347676 512514 347712
rect 512458 347656 512460 347676
rect 512460 347656 512512 347676
rect 512512 347656 512514 347676
rect 512826 347112 512882 347168
rect 513286 346588 513342 346624
rect 513286 346568 513288 346588
rect 513288 346568 513340 346588
rect 513340 346568 513342 346588
rect 512458 346024 512514 346080
rect 512458 345480 512514 345536
rect 513010 344936 513066 344992
rect 513286 343848 513342 343904
rect 513010 343304 513066 343360
rect 512550 342216 512606 342272
rect 513286 341672 513342 341728
rect 513286 341148 513342 341184
rect 513286 341128 513288 341148
rect 513288 341128 513340 341148
rect 513340 341128 513342 341148
rect 513286 340584 513342 340640
rect 513102 340040 513158 340096
rect 513286 339532 513288 339552
rect 513288 339532 513340 339552
rect 513340 339532 513342 339552
rect 513286 339496 513342 339532
rect 512642 338952 512698 339008
rect 513010 338408 513066 338464
rect 512734 337864 512790 337920
rect 512826 337320 512882 337376
rect 513286 336776 513342 336832
rect 512734 336232 512790 336288
rect 513010 335144 513066 335200
rect 512734 334600 512790 334656
rect 513286 334056 513342 334112
rect 512826 332424 512882 332480
rect 512826 329704 512882 329760
rect 512826 326984 512882 327040
rect 512550 302912 512606 302968
rect 513470 333512 513526 333568
rect 512826 302776 512882 302832
rect 517886 305768 517942 305824
rect 519634 502288 519690 502344
rect 547878 516704 547934 516760
rect 521750 462848 521806 462904
rect 557538 442856 557594 442912
rect 531318 261024 531374 261080
rect 531318 243616 531374 243672
rect 530122 226208 530178 226264
rect 529938 209208 529994 209264
rect 460294 67632 460350 67688
rect 460846 67632 460902 67688
rect 538954 137944 539010 138000
rect 539414 137808 539470 137864
rect 539506 135904 539562 135960
rect 539414 129648 539470 129704
rect 539874 117272 539930 117328
rect 540242 131280 540298 131336
rect 540150 127200 540206 127256
rect 540334 125160 540390 125216
rect 540058 112784 540114 112840
rect 539966 108704 540022 108760
rect 539782 99184 539838 99240
rect 539690 97144 539746 97200
rect 539598 95104 539654 95160
rect 536838 40976 536894 41032
rect 541070 110880 541126 110936
rect 541438 114960 541494 115016
rect 541346 106800 541402 106856
rect 541254 104760 541310 104816
rect 541162 102720 541218 102776
rect 542726 123120 542782 123176
rect 542634 121080 542690 121136
rect 542542 100680 542598 100736
rect 542450 90480 542506 90536
rect 543094 119040 543150 119096
rect 543002 92520 543058 92576
rect 543186 88440 543242 88496
rect 542910 86400 542966 86456
rect 542818 84360 542874 84416
rect 540978 82320 541034 82376
rect 580170 683848 580226 683904
rect 580170 670692 580172 670712
rect 580172 670692 580224 670712
rect 580224 670692 580226 670712
rect 580170 670656 580226 670692
rect 580262 644000 580318 644056
rect 580170 617480 580226 617536
rect 580354 630808 580410 630864
rect 580170 590960 580226 591016
rect 580170 577632 580226 577688
rect 580262 564304 580318 564360
rect 580170 537784 580226 537840
rect 580170 484608 580226 484664
rect 580170 458088 580226 458144
rect 580170 431568 580226 431624
rect 580170 404912 580226 404968
rect 580170 365064 580226 365120
rect 580170 351872 580226 351928
rect 580170 325216 580226 325272
rect 580446 524456 580502 524512
rect 580354 418240 580410 418296
rect 580538 511264 580594 511320
rect 580630 471416 580686 471472
rect 580722 378392 580778 378448
rect 580170 312024 580226 312080
rect 540610 48864 540666 48920
rect 540426 34176 540482 34232
rect 580170 298696 580226 298752
rect 580262 272176 580318 272232
rect 580170 245556 580172 245576
rect 580172 245556 580224 245576
rect 580224 245556 580226 245576
rect 580170 245520 580226 245556
rect 580170 232328 580226 232384
rect 580354 258848 580410 258904
rect 580262 219000 580318 219056
rect 579802 205672 579858 205728
rect 580170 192480 580226 192536
rect 580170 179152 580226 179208
rect 580170 165824 580226 165880
rect 580170 152632 580226 152688
rect 580170 139340 580172 139360
rect 580172 139340 580224 139360
rect 580224 139340 580226 139360
rect 580170 139304 580226 139340
rect 580170 125976 580226 126032
rect 579802 112784 579858 112840
rect 580170 99456 580226 99512
rect 580170 86128 580226 86184
rect 580170 72936 580226 72992
rect 580170 59608 580226 59664
rect 580170 46280 580226 46336
rect 580170 33108 580226 33144
rect 580170 33088 580172 33108
rect 580172 33088 580224 33108
rect 580224 33088 580226 33108
rect 579986 19760 580042 19816
rect 580170 6568 580226 6624
rect 365074 3168 365130 3224
<< metal3 >>
rect 429837 700634 429903 700637
rect 447910 700634 447916 700636
rect 429837 700632 447916 700634
rect 429837 700576 429842 700632
rect 429898 700576 447916 700632
rect 429837 700574 447916 700576
rect 429837 700571 429903 700574
rect 447910 700572 447916 700574
rect 447980 700572 447986 700636
rect 202781 700498 202847 700501
rect 449566 700498 449572 700500
rect 202781 700496 449572 700498
rect 202781 700440 202786 700496
rect 202842 700440 449572 700496
rect 202781 700438 449572 700440
rect 202781 700435 202847 700438
rect 449566 700436 449572 700438
rect 449636 700436 449642 700500
rect 40493 700362 40559 700365
rect 447726 700362 447732 700364
rect 40493 700360 447732 700362
rect 40493 700304 40498 700360
rect 40554 700304 447732 700360
rect 40493 700302 447732 700304
rect 40493 700299 40559 700302
rect 447726 700300 447732 700302
rect 447796 700300 447802 700364
rect 530526 700300 530532 700364
rect 530596 700362 530602 700364
rect 543457 700362 543523 700365
rect 530596 700360 543523 700362
rect 530596 700304 543462 700360
rect 543518 700304 543523 700360
rect 530596 700302 543523 700304
rect 530596 700300 530602 700302
rect 543457 700299 543523 700302
rect 527173 699820 527239 699821
rect 527173 699818 527220 699820
rect 527128 699816 527220 699818
rect 527128 699760 527178 699816
rect 527128 699758 527220 699760
rect 527173 699756 527220 699758
rect 527284 699756 527290 699820
rect 558126 699756 558132 699820
rect 558196 699818 558202 699820
rect 559649 699818 559715 699821
rect 558196 699816 559715 699818
rect 558196 699760 559654 699816
rect 559710 699760 559715 699816
rect 558196 699758 559715 699760
rect 558196 699756 558202 699758
rect 527173 699755 527239 699756
rect 559649 699755 559715 699758
rect -960 697220 480 697460
rect 580165 697234 580231 697237
rect 583520 697234 584960 697324
rect 580165 697232 584960 697234
rect 580165 697176 580170 697232
rect 580226 697176 584960 697232
rect 580165 697174 584960 697176
rect 580165 697171 580231 697174
rect 583520 697084 584960 697174
rect 300117 689346 300183 689349
rect 444230 689346 444236 689348
rect 300117 689344 444236 689346
rect 300117 689288 300122 689344
rect 300178 689288 444236 689344
rect 300117 689286 444236 689288
rect 300117 689283 300183 689286
rect 444230 689284 444236 689286
rect 444300 689284 444306 689348
rect 24301 686490 24367 686493
rect 446254 686490 446260 686492
rect 24301 686488 446260 686490
rect 24301 686432 24306 686488
rect 24362 686432 446260 686488
rect 24301 686430 446260 686432
rect 24301 686427 24367 686430
rect 446254 686428 446260 686430
rect 446324 686428 446330 686492
rect -960 684314 480 684404
rect 3233 684314 3299 684317
rect -960 684312 3299 684314
rect -960 684256 3238 684312
rect 3294 684256 3299 684312
rect -960 684254 3299 684256
rect -960 684164 480 684254
rect 3233 684251 3299 684254
rect 580165 683906 580231 683909
rect 583520 683906 584960 683996
rect 580165 683904 584960 683906
rect 580165 683848 580170 683904
rect 580226 683848 584960 683904
rect 580165 683846 584960 683848
rect 580165 683843 580231 683846
rect 583520 683756 584960 683846
rect 3734 683300 3740 683364
rect 3804 683362 3810 683364
rect 446857 683362 446923 683365
rect 3804 683360 446923 683362
rect 3804 683304 446862 683360
rect 446918 683304 446923 683360
rect 3804 683302 446923 683304
rect 3804 683300 3810 683302
rect 446857 683299 446923 683302
rect 3550 683164 3556 683228
rect 3620 683226 3626 683228
rect 447041 683226 447107 683229
rect 3620 683224 447107 683226
rect 3620 683168 447046 683224
rect 447102 683168 447107 683224
rect 3620 683166 447107 683168
rect 3620 683164 3626 683166
rect 447041 683163 447107 683166
rect 3366 682756 3372 682820
rect 3436 682818 3442 682820
rect 420085 682818 420151 682821
rect 3436 682816 420151 682818
rect 3436 682760 420090 682816
rect 420146 682760 420151 682816
rect 3436 682758 420151 682760
rect 3436 682756 3442 682758
rect 420085 682755 420151 682758
rect 361757 679010 361823 679013
rect 359812 679008 361823 679010
rect 359812 678952 361762 679008
rect 361818 678952 361823 679008
rect 359812 678950 361823 678952
rect 361757 678947 361823 678950
rect -960 671258 480 671348
rect 3734 671258 3740 671260
rect -960 671198 3740 671258
rect -960 671108 480 671198
rect 3734 671196 3740 671198
rect 3804 671196 3810 671260
rect 580165 670714 580231 670717
rect 583520 670714 584960 670804
rect 580165 670712 584960 670714
rect 580165 670656 580170 670712
rect 580226 670656 584960 670712
rect 580165 670654 584960 670656
rect 580165 670651 580231 670654
rect 583520 670564 584960 670654
rect 460197 668130 460263 668133
rect 460197 668128 460306 668130
rect 460197 668072 460202 668128
rect 460258 668072 460306 668128
rect 460197 668067 460306 668072
rect 361757 667994 361823 667997
rect 359812 667992 361823 667994
rect 359812 667936 361762 667992
rect 361818 667936 361823 667992
rect 460246 667964 460306 668067
rect 359812 667934 361823 667936
rect 361757 667931 361823 667934
rect 457846 665212 457852 665276
rect 457916 665274 457922 665276
rect 460062 665274 460122 665448
rect 457916 665214 460122 665274
rect 457916 665212 457922 665214
rect 458030 662492 458036 662556
rect 458100 662554 458106 662556
rect 460062 662554 460122 663000
rect 458100 662494 460122 662554
rect 458100 662492 458106 662494
rect 458081 659970 458147 659973
rect 460062 659970 460122 660552
rect 458081 659968 460122 659970
rect 458081 659912 458086 659968
rect 458142 659912 460122 659968
rect 458081 659910 460122 659912
rect 458081 659907 458147 659910
rect -960 658202 480 658292
rect 3141 658202 3207 658205
rect -960 658200 3207 658202
rect -960 658144 3146 658200
rect 3202 658144 3207 658200
rect -960 658142 3207 658144
rect -960 658052 480 658142
rect 3141 658139 3207 658142
rect 457805 657522 457871 657525
rect 460062 657522 460122 658104
rect 457805 657520 460122 657522
rect 457805 657464 457810 657520
rect 457866 657464 460122 657520
rect 457805 657462 460122 657464
rect 457805 657459 457871 657462
rect 583520 657236 584960 657476
rect 361757 656978 361823 656981
rect 359812 656976 361823 656978
rect 359812 656920 361762 656976
rect 361818 656920 361823 656976
rect 359812 656918 361823 656920
rect 361757 656915 361823 656918
rect 459502 655624 459508 655688
rect 459572 655686 459578 655688
rect 459572 655626 460092 655686
rect 459572 655624 459578 655626
rect 457713 652898 457779 652901
rect 460062 652898 460122 653208
rect 457713 652896 460122 652898
rect 457713 652840 457718 652896
rect 457774 652840 460122 652896
rect 457713 652838 460122 652840
rect 457713 652835 457779 652838
rect 457621 650178 457687 650181
rect 460062 650178 460122 650760
rect 457621 650176 460122 650178
rect 457621 650120 457626 650176
rect 457682 650120 460122 650176
rect 457621 650118 460122 650120
rect 457621 650115 457687 650118
rect 459369 647730 459435 647733
rect 460062 647730 460122 648312
rect 459369 647728 460122 647730
rect 459369 647672 459374 647728
rect 459430 647672 460122 647728
rect 459369 647670 460122 647672
rect 459369 647667 459435 647670
rect 361757 645962 361823 645965
rect 359812 645960 361823 645962
rect 359812 645904 361762 645960
rect 361818 645904 361823 645960
rect 359812 645902 361823 645904
rect 361757 645899 361823 645902
rect 457529 645962 457595 645965
rect 457529 645960 460092 645962
rect 457529 645904 457534 645960
rect 457590 645904 460092 645960
rect 457529 645902 460092 645904
rect 457529 645899 457595 645902
rect -960 644996 480 645236
rect 580257 644058 580323 644061
rect 583520 644058 584960 644148
rect 580257 644056 584960 644058
rect 580257 644000 580262 644056
rect 580318 644000 584960 644056
rect 580257 643998 584960 644000
rect 580257 643995 580323 643998
rect 583520 643908 584960 643998
rect 457437 643242 457503 643245
rect 460062 643242 460122 643416
rect 457437 643240 460122 643242
rect 457437 643184 457442 643240
rect 457498 643184 460122 643240
rect 457437 643182 460122 643184
rect 457437 643179 457503 643182
rect 459277 640386 459343 640389
rect 460062 640386 460122 640968
rect 459277 640384 460122 640386
rect 459277 640328 459282 640384
rect 459338 640328 460122 640384
rect 459277 640326 460122 640328
rect 459277 640323 459343 640326
rect 459185 637938 459251 637941
rect 460062 637938 460122 638520
rect 459185 637936 460122 637938
rect 459185 637880 459190 637936
rect 459246 637880 460122 637936
rect 459185 637878 460122 637880
rect 459185 637875 459251 637878
rect 457989 635490 458055 635493
rect 460062 635490 460122 636072
rect 457989 635488 460122 635490
rect 457989 635432 457994 635488
rect 458050 635432 460122 635488
rect 457989 635430 460122 635432
rect 457989 635427 458055 635430
rect 361573 634946 361639 634949
rect 359812 634944 361639 634946
rect 359812 634888 361578 634944
rect 361634 634888 361639 634944
rect 359812 634886 361639 634888
rect 361573 634883 361639 634886
rect 459093 633450 459159 633453
rect 460062 633450 460122 633624
rect 459093 633448 460122 633450
rect 459093 633392 459098 633448
rect 459154 633392 460122 633448
rect 459093 633390 460122 633392
rect 459093 633387 459159 633390
rect -960 632090 480 632180
rect 3693 632090 3759 632093
rect -960 632088 3759 632090
rect -960 632032 3698 632088
rect 3754 632032 3759 632088
rect -960 632030 3759 632032
rect -960 631940 480 632030
rect 3693 632027 3759 632030
rect 459001 630730 459067 630733
rect 460062 630730 460122 631176
rect 580349 630866 580415 630869
rect 583520 630866 584960 630956
rect 580349 630864 584960 630866
rect 580349 630808 580354 630864
rect 580410 630808 584960 630864
rect 580349 630806 584960 630808
rect 580349 630803 580415 630806
rect 459001 630728 460122 630730
rect 459001 630672 459006 630728
rect 459062 630672 460122 630728
rect 583520 630716 584960 630806
rect 459001 630670 460122 630672
rect 459001 630667 459067 630670
rect 459461 628146 459527 628149
rect 460062 628146 460122 628728
rect 459461 628144 460122 628146
rect 459461 628088 459466 628144
rect 459522 628088 460122 628144
rect 459461 628086 460122 628088
rect 459461 628083 459527 628086
rect 460062 625837 460122 626280
rect 460062 625832 460171 625837
rect 460062 625776 460110 625832
rect 460166 625776 460171 625832
rect 460062 625774 460171 625776
rect 460105 625771 460171 625774
rect 361573 623930 361639 623933
rect 359812 623928 361639 623930
rect 359812 623872 361578 623928
rect 361634 623872 361639 623928
rect 359812 623870 361639 623872
rect 361573 623867 361639 623870
rect 457345 623930 457411 623933
rect 457345 623928 460092 623930
rect 457345 623872 457350 623928
rect 457406 623872 460092 623928
rect 457345 623870 460092 623872
rect 457345 623867 457411 623870
rect 457253 621074 457319 621077
rect 460062 621074 460122 621384
rect 457253 621072 460122 621074
rect 457253 621016 457258 621072
rect 457314 621016 460122 621072
rect 457253 621014 460122 621016
rect 457253 621011 457319 621014
rect -960 619170 480 619260
rect 3550 619170 3556 619172
rect -960 619110 3556 619170
rect -960 619020 480 619110
rect 3550 619108 3556 619110
rect 3620 619108 3626 619172
rect 457897 618354 457963 618357
rect 460062 618354 460122 618936
rect 457897 618352 460122 618354
rect 457897 618296 457902 618352
rect 457958 618296 460122 618352
rect 457897 618294 460122 618296
rect 457897 618291 457963 618294
rect 580165 617538 580231 617541
rect 583520 617538 584960 617628
rect 580165 617536 584960 617538
rect 580165 617480 580170 617536
rect 580226 617480 584960 617536
rect 580165 617478 584960 617480
rect 580165 617475 580231 617478
rect 583520 617388 584960 617478
rect 458817 616042 458883 616045
rect 460062 616042 460122 616488
rect 458817 616040 460122 616042
rect 458817 615984 458822 616040
rect 458878 615984 460122 616040
rect 458817 615982 460122 615984
rect 458817 615979 458883 615982
rect 458909 614138 458975 614141
rect 458909 614136 460092 614138
rect 458909 614080 458914 614136
rect 458970 614080 460092 614136
rect 458909 614078 460092 614080
rect 458909 614075 458975 614078
rect 361573 612914 361639 612917
rect 359812 612912 361639 612914
rect 359812 612856 361578 612912
rect 361634 612856 361639 612912
rect 359812 612854 361639 612856
rect 361573 612851 361639 612854
rect 458725 611418 458791 611421
rect 460062 611418 460122 611592
rect 458725 611416 460122 611418
rect 458725 611360 458730 611416
rect 458786 611360 460122 611416
rect 458725 611358 460122 611360
rect 458725 611355 458791 611358
rect 458633 608698 458699 608701
rect 460062 608698 460122 609144
rect 458633 608696 460122 608698
rect 458633 608640 458638 608696
rect 458694 608640 460122 608696
rect 458633 608638 460122 608640
rect 458633 608635 458699 608638
rect 460062 606389 460122 606696
rect 460013 606384 460122 606389
rect 460013 606328 460018 606384
rect 460074 606328 460122 606384
rect 460013 606326 460122 606328
rect 460013 606323 460079 606326
rect -960 606114 480 606204
rect 3366 606114 3372 606116
rect -960 606054 3372 606114
rect -960 605964 480 606054
rect 3366 606052 3372 606054
rect 3436 606052 3442 606116
rect 459921 603666 459987 603669
rect 460062 603666 460122 604248
rect 583520 604060 584960 604300
rect 459921 603664 460122 603666
rect 459921 603608 459926 603664
rect 459982 603608 460122 603664
rect 459921 603606 460122 603608
rect 459921 603603 459987 603606
rect 361757 601898 361823 601901
rect 359812 601896 361823 601898
rect 359812 601840 361762 601896
rect 361818 601840 361823 601896
rect 359812 601838 361823 601840
rect 361757 601835 361823 601838
rect 459829 601898 459895 601901
rect 459829 601896 460092 601898
rect 459829 601840 459834 601896
rect 459890 601840 460092 601896
rect 459829 601838 460092 601840
rect 459829 601835 459895 601838
rect 459185 599586 459251 599589
rect 474406 599586 474412 599588
rect 459185 599584 474412 599586
rect 459185 599528 459190 599584
rect 459246 599528 474412 599584
rect 459185 599526 474412 599528
rect 459185 599523 459251 599526
rect 474406 599524 474412 599526
rect 474476 599524 474482 599588
rect 459093 598226 459159 598229
rect 472014 598226 472020 598228
rect 459093 598224 472020 598226
rect 459093 598168 459098 598224
rect 459154 598168 472020 598224
rect 459093 598166 472020 598168
rect 459093 598163 459159 598166
rect 472014 598164 472020 598166
rect 472084 598164 472090 598228
rect 457846 597620 457852 597684
rect 457916 597682 457922 597684
rect 461761 597682 461827 597685
rect 457916 597680 461827 597682
rect 457916 597624 461766 597680
rect 461822 597624 461827 597680
rect 457916 597622 461827 597624
rect 457916 597620 457922 597622
rect 461761 597619 461827 597622
rect 459001 595642 459067 595645
rect 472198 595642 472204 595644
rect 459001 595640 472204 595642
rect 459001 595584 459006 595640
rect 459062 595584 472204 595640
rect 459001 595582 472204 595584
rect 459001 595579 459067 595582
rect 472198 595580 472204 595582
rect 472268 595580 472274 595644
rect 459502 595444 459508 595508
rect 459572 595506 459578 595508
rect 478822 595506 478828 595508
rect 459572 595446 478828 595506
rect 459572 595444 459578 595446
rect 478822 595444 478828 595446
rect 478892 595444 478898 595508
rect -960 592908 480 593148
rect 459369 591290 459435 591293
rect 476430 591290 476436 591292
rect 459369 591288 476436 591290
rect 459369 591232 459374 591288
rect 459430 591232 476436 591288
rect 459369 591230 476436 591232
rect 459369 591227 459435 591230
rect 476430 591228 476436 591230
rect 476500 591228 476506 591292
rect 580165 591018 580231 591021
rect 583520 591018 584960 591108
rect 580165 591016 584960 591018
rect 580165 590960 580170 591016
rect 580226 590960 584960 591016
rect 580165 590958 584960 590960
rect 580165 590955 580231 590958
rect 361757 590882 361823 590885
rect 359812 590880 361823 590882
rect 359812 590824 361762 590880
rect 361818 590824 361823 590880
rect 583520 590868 584960 590958
rect 359812 590822 361823 590824
rect 361757 590819 361823 590822
rect 459277 589930 459343 589933
rect 474774 589930 474780 589932
rect 459277 589928 474780 589930
rect 459277 589872 459282 589928
rect 459338 589872 474780 589928
rect 459277 589870 474780 589872
rect 459277 589867 459343 589870
rect 474774 589868 474780 589870
rect 474844 589868 474850 589932
rect -960 580002 480 580092
rect 3233 580002 3299 580005
rect -960 580000 3299 580002
rect -960 579944 3238 580000
rect 3294 579944 3299 580000
rect -960 579942 3299 579944
rect -960 579852 480 579942
rect 3233 579939 3299 579942
rect 361757 579866 361823 579869
rect 359812 579864 361823 579866
rect 359812 579808 361762 579864
rect 361818 579808 361823 579864
rect 359812 579806 361823 579808
rect 361757 579803 361823 579806
rect 580165 577690 580231 577693
rect 583520 577690 584960 577780
rect 580165 577688 584960 577690
rect 580165 577632 580170 577688
rect 580226 577632 584960 577688
rect 580165 577630 584960 577632
rect 580165 577627 580231 577630
rect 583520 577540 584960 577630
rect 361573 568850 361639 568853
rect 359812 568848 361639 568850
rect 359812 568792 361578 568848
rect 361634 568792 361639 568848
rect 359812 568790 361639 568792
rect 361573 568787 361639 568790
rect -960 566946 480 567036
rect 3325 566946 3391 566949
rect -960 566944 3391 566946
rect -960 566888 3330 566944
rect 3386 566888 3391 566944
rect -960 566886 3391 566888
rect -960 566796 480 566886
rect 3325 566883 3391 566886
rect 580257 564362 580323 564365
rect 583520 564362 584960 564452
rect 580257 564360 584960 564362
rect 580257 564304 580262 564360
rect 580318 564304 584960 564360
rect 580257 564302 584960 564304
rect 580257 564299 580323 564302
rect 583520 564212 584960 564302
rect 361665 557834 361731 557837
rect 359812 557832 361731 557834
rect 359812 557776 361670 557832
rect 361726 557776 361731 557832
rect 359812 557774 361731 557776
rect 361665 557771 361731 557774
rect -960 553890 480 553980
rect 4061 553890 4127 553893
rect -960 553888 4127 553890
rect -960 553832 4066 553888
rect 4122 553832 4127 553888
rect -960 553830 4127 553832
rect -960 553740 480 553830
rect 4061 553827 4127 553830
rect 583520 551020 584960 551260
rect 361757 546818 361823 546821
rect 359812 546816 361823 546818
rect 359812 546760 361762 546816
rect 361818 546760 361823 546816
rect 359812 546758 361823 546760
rect 361757 546755 361823 546758
rect -960 540684 480 540924
rect 580165 537842 580231 537845
rect 583520 537842 584960 537932
rect 580165 537840 584960 537842
rect 580165 537784 580170 537840
rect 580226 537784 584960 537840
rect 580165 537782 584960 537784
rect 580165 537779 580231 537782
rect 583520 537692 584960 537782
rect 361573 535802 361639 535805
rect 359812 535800 361639 535802
rect 359812 535744 361578 535800
rect 361634 535744 361639 535800
rect 359812 535742 361639 535744
rect 361573 535739 361639 535742
rect -960 527914 480 528004
rect 3969 527914 4035 527917
rect -960 527912 4035 527914
rect -960 527856 3974 527912
rect 4030 527856 4035 527912
rect -960 527854 4035 527856
rect -960 527764 480 527854
rect 3969 527851 4035 527854
rect 361573 524786 361639 524789
rect 359812 524784 361639 524786
rect 359812 524728 361578 524784
rect 361634 524728 361639 524784
rect 359812 524726 361639 524728
rect 361573 524723 361639 524726
rect 580441 524514 580507 524517
rect 583520 524514 584960 524604
rect 580441 524512 584960 524514
rect 580441 524456 580446 524512
rect 580502 524456 584960 524512
rect 580441 524454 584960 524456
rect 580441 524451 580507 524454
rect 583520 524364 584960 524454
rect 458030 518060 458036 518124
rect 458100 518122 458106 518124
rect 467097 518122 467163 518125
rect 458100 518120 467163 518122
rect 458100 518064 467102 518120
rect 467158 518064 467163 518120
rect 458100 518062 467163 518064
rect 458100 518060 458106 518062
rect 467097 518059 467163 518062
rect 482737 517580 482803 517581
rect 482686 517516 482692 517580
rect 482756 517578 482803 517580
rect 482756 517576 482848 517578
rect 482798 517520 482848 517576
rect 482756 517518 482848 517520
rect 482756 517516 482803 517518
rect 482737 517515 482803 517516
rect 450445 516898 450511 516901
rect 500953 516898 501019 516901
rect 502241 516898 502307 516901
rect 450445 516896 502307 516898
rect 450445 516840 450450 516896
rect 450506 516840 500958 516896
rect 501014 516840 502246 516896
rect 502302 516840 502307 516896
rect 450445 516838 502307 516840
rect 450445 516835 450511 516838
rect 500953 516835 501019 516838
rect 502241 516835 502307 516838
rect 451038 516762 451044 516764
rect 450678 516702 451044 516762
rect 450678 516528 450738 516702
rect 451038 516700 451044 516702
rect 451108 516762 451114 516764
rect 507117 516762 507183 516765
rect 547873 516762 547939 516765
rect 451108 516760 547939 516762
rect 451108 516704 507122 516760
rect 507178 516704 547878 516760
rect 547934 516704 547939 516760
rect 451108 516702 547939 516704
rect 451108 516700 451114 516702
rect 507117 516699 507183 516702
rect 547873 516699 547939 516702
rect 491894 515538 491954 515984
rect 494053 515538 494119 515541
rect 491894 515536 494119 515538
rect 491894 515480 494058 515536
rect 494114 515480 494119 515536
rect 491894 515478 494119 515480
rect 494053 515475 494119 515478
rect -960 514858 480 514948
rect 3877 514858 3943 514861
rect -960 514856 3943 514858
rect -960 514800 3882 514856
rect 3938 514800 3943 514856
rect -960 514798 3943 514800
rect -960 514708 480 514798
rect 3877 514795 3943 514798
rect 450445 514722 450511 514725
rect 450445 514720 450554 514722
rect 450445 514664 450450 514720
rect 450506 514664 450554 514720
rect 450445 514659 450554 514664
rect 450494 514384 450554 514659
rect 450486 514320 450492 514384
rect 450556 514320 450562 514384
rect 361757 513770 361823 513773
rect 359812 513768 361823 513770
rect 359812 513712 361762 513768
rect 361818 513712 361823 513768
rect 359812 513710 361823 513712
rect 361757 513707 361823 513710
rect 492121 512478 492187 512481
rect 491924 512476 492187 512478
rect 491924 512420 492126 512476
rect 492182 512420 492187 512476
rect 491924 512418 492187 512420
rect 492121 512415 492187 512418
rect 450537 512410 450603 512413
rect 450494 512408 450603 512410
rect 450494 512352 450542 512408
rect 450598 512352 450603 512408
rect 450494 512347 450603 512352
rect 450494 512176 450554 512347
rect 580533 511322 580599 511325
rect 583520 511322 584960 511412
rect 580533 511320 584960 511322
rect 580533 511264 580538 511320
rect 580594 511264 584960 511320
rect 580533 511262 584960 511264
rect 580533 511259 580599 511262
rect 583520 511172 584960 511262
rect 450353 510234 450419 510237
rect 450310 510232 450419 510234
rect 450310 510176 450358 510232
rect 450414 510176 450419 510232
rect 450310 510171 450419 510176
rect 450310 510000 450370 510171
rect 491894 508874 491954 508912
rect 494145 508874 494211 508877
rect 491894 508872 494211 508874
rect 491894 508816 494150 508872
rect 494206 508816 494211 508872
rect 491894 508814 494211 508816
rect 494145 508811 494211 508814
rect 449985 507650 450051 507653
rect 450126 507650 450186 507824
rect 449985 507648 450186 507650
rect 449985 507592 449990 507648
rect 450046 507592 450186 507648
rect 449985 507590 450186 507592
rect 449985 507587 450051 507590
rect 494237 505746 494303 505749
rect 495065 505746 495131 505749
rect 491894 505744 495131 505746
rect 491894 505688 494242 505744
rect 494298 505688 495070 505744
rect 495126 505688 495131 505744
rect 491894 505686 495131 505688
rect 450126 505477 450186 505648
rect 450077 505474 450186 505477
rect 450629 505474 450695 505477
rect 450077 505472 450695 505474
rect 450077 505416 450082 505472
rect 450138 505416 450634 505472
rect 450690 505416 450695 505472
rect 450077 505414 450695 505416
rect 450077 505411 450143 505414
rect 450629 505411 450695 505414
rect 491894 505376 491954 505686
rect 494237 505683 494303 505686
rect 495065 505683 495131 505686
rect 449801 503502 449867 503505
rect 449801 503500 450156 503502
rect 449801 503444 449806 503500
rect 449862 503472 450156 503500
rect 449862 503444 450186 503472
rect 449801 503442 450186 503444
rect 449801 503439 449867 503442
rect 450126 503301 450186 503442
rect 450126 503296 450235 503301
rect 450126 503240 450174 503296
rect 450230 503240 450235 503296
rect 450126 503238 450235 503240
rect 450169 503235 450235 503238
rect 361757 502754 361823 502757
rect 359812 502752 361823 502754
rect 359812 502696 361762 502752
rect 361818 502696 361823 502752
rect 359812 502694 361823 502696
rect 361757 502691 361823 502694
rect 519629 502346 519695 502349
rect 527214 502346 527220 502348
rect 519629 502344 527220 502346
rect 519629 502288 519634 502344
rect 519690 502288 527220 502344
rect 519629 502286 527220 502288
rect 519629 502283 519695 502286
rect 527214 502284 527220 502286
rect 527284 502284 527290 502348
rect -960 501802 480 501892
rect 3785 501802 3851 501805
rect -960 501800 3851 501802
rect -960 501744 3790 501800
rect 3846 501744 3851 501800
rect -960 501742 3851 501744
rect -960 501652 480 501742
rect 3785 501739 3851 501742
rect 491894 501666 491954 501840
rect 470550 501606 491954 501666
rect 450678 501122 450738 501296
rect 463049 501122 463115 501125
rect 470550 501122 470610 501606
rect 491894 501258 491954 501606
rect 494697 501258 494763 501261
rect 491894 501256 494763 501258
rect 491894 501200 494702 501256
rect 494758 501200 494763 501256
rect 491894 501198 494763 501200
rect 494697 501195 494763 501198
rect 450678 501120 470610 501122
rect 450678 501064 463054 501120
rect 463110 501064 470610 501120
rect 450678 501062 470610 501064
rect 463049 501059 463115 501062
rect 583520 497844 584960 498084
rect 489177 496906 489243 496909
rect 489310 496906 489316 496908
rect 489177 496904 489316 496906
rect 489177 496848 489182 496904
rect 489238 496848 489316 496904
rect 489177 496846 489316 496848
rect 489177 496843 489243 496846
rect 489310 496844 489316 496846
rect 489380 496844 489386 496908
rect 361757 491738 361823 491741
rect 359812 491736 361823 491738
rect 359812 491680 361762 491736
rect 361818 491680 361823 491736
rect 359812 491678 361823 491680
rect 361757 491675 361823 491678
rect -960 488596 480 488836
rect 580165 484666 580231 484669
rect 583520 484666 584960 484756
rect 580165 484664 584960 484666
rect 580165 484608 580170 484664
rect 580226 484608 584960 484664
rect 580165 484606 584960 484608
rect 580165 484603 580231 484606
rect 583520 484516 584960 484606
rect 361757 480722 361823 480725
rect 359812 480720 361823 480722
rect 359812 480664 361762 480720
rect 361818 480664 361823 480720
rect 359812 480662 361823 480664
rect 361757 480659 361823 480662
rect -960 475690 480 475780
rect 3601 475690 3667 475693
rect -960 475688 3667 475690
rect -960 475632 3606 475688
rect 3662 475632 3667 475688
rect -960 475630 3667 475632
rect -960 475540 480 475630
rect 3601 475627 3667 475630
rect 580625 471474 580691 471477
rect 583520 471474 584960 471564
rect 580625 471472 584960 471474
rect 580625 471416 580630 471472
rect 580686 471416 584960 471472
rect 580625 471414 584960 471416
rect 580625 471411 580691 471414
rect 583520 471324 584960 471414
rect 361757 469706 361823 469709
rect 359812 469704 361823 469706
rect 359812 469648 361762 469704
rect 361818 469648 361823 469704
rect 359812 469646 361823 469648
rect 361757 469643 361823 469646
rect 473721 462906 473787 462909
rect 482686 462906 482692 462908
rect 473721 462904 482692 462906
rect 473721 462848 473726 462904
rect 473782 462848 482692 462904
rect 473721 462846 482692 462848
rect 473721 462843 473787 462846
rect 482686 462844 482692 462846
rect 482756 462906 482762 462908
rect 521745 462906 521811 462909
rect 482756 462904 521811 462906
rect 482756 462848 521750 462904
rect 521806 462848 521811 462904
rect 482756 462846 521811 462848
rect 482756 462844 482762 462846
rect 521745 462843 521811 462846
rect -960 462634 480 462724
rect 3509 462634 3575 462637
rect -960 462632 3575 462634
rect -960 462576 3514 462632
rect 3570 462576 3575 462632
rect -960 462574 3575 462576
rect -960 462484 480 462574
rect 3509 462571 3575 462574
rect 361757 458690 361823 458693
rect 359812 458688 361823 458690
rect 359812 458632 361762 458688
rect 361818 458632 361823 458688
rect 359812 458630 361823 458632
rect 361757 458627 361823 458630
rect 580165 458146 580231 458149
rect 583520 458146 584960 458236
rect 580165 458144 584960 458146
rect 580165 458088 580170 458144
rect 580226 458088 584960 458144
rect 580165 458086 584960 458088
rect 580165 458083 580231 458086
rect 583520 457996 584960 458086
rect -960 449578 480 449668
rect 3417 449578 3483 449581
rect -960 449576 3483 449578
rect -960 449520 3422 449576
rect 3478 449520 3483 449576
rect -960 449518 3483 449520
rect -960 449428 480 449518
rect 3417 449515 3483 449518
rect 362217 447674 362283 447677
rect 359812 447672 362283 447674
rect 359812 447616 362222 447672
rect 362278 447616 362283 447672
rect 359812 447614 362283 447616
rect 362217 447611 362283 447614
rect 583520 444668 584960 444908
rect 557533 442914 557599 442917
rect 555956 442912 557599 442914
rect 555956 442856 557538 442912
rect 557594 442856 557599 442912
rect 555956 442854 557599 442856
rect 557533 442851 557599 442854
rect -960 436508 480 436748
rect 361757 436658 361823 436661
rect 359812 436656 361823 436658
rect 359812 436600 361762 436656
rect 361818 436600 361823 436656
rect 359812 436598 361823 436600
rect 361757 436595 361823 436598
rect 580165 431626 580231 431629
rect 583520 431626 584960 431716
rect 580165 431624 584960 431626
rect 580165 431568 580170 431624
rect 580226 431568 584960 431624
rect 580165 431566 584960 431568
rect 580165 431563 580231 431566
rect 583520 431476 584960 431566
rect 362309 425642 362375 425645
rect 359812 425640 362375 425642
rect 359812 425584 362314 425640
rect 362370 425584 362375 425640
rect 359812 425582 362375 425584
rect 362309 425579 362375 425582
rect -960 423602 480 423692
rect 3693 423602 3759 423605
rect -960 423600 3759 423602
rect -960 423544 3698 423600
rect 3754 423544 3759 423600
rect -960 423542 3759 423544
rect -960 423452 480 423542
rect 3693 423539 3759 423542
rect 444046 421908 444052 421972
rect 444116 421970 444122 421972
rect 444189 421970 444255 421973
rect 444116 421968 444255 421970
rect 444116 421912 444194 421968
rect 444250 421912 444255 421968
rect 444116 421910 444255 421912
rect 444116 421908 444122 421910
rect 444189 421907 444255 421910
rect 580349 418298 580415 418301
rect 583520 418298 584960 418388
rect 580349 418296 584960 418298
rect 580349 418240 580354 418296
rect 580410 418240 584960 418296
rect 580349 418238 584960 418240
rect 580349 418235 580415 418238
rect 583520 418148 584960 418238
rect 361573 414626 361639 414629
rect 359812 414624 361639 414626
rect 359812 414568 361578 414624
rect 361634 414568 361639 414624
rect 359812 414566 361639 414568
rect 361573 414563 361639 414566
rect -960 410546 480 410636
rect 3969 410546 4035 410549
rect -960 410544 4035 410546
rect -960 410488 3974 410544
rect 4030 410488 4035 410544
rect -960 410486 4035 410488
rect -960 410396 480 410486
rect 3969 410483 4035 410486
rect 580165 404970 580231 404973
rect 583520 404970 584960 405060
rect 580165 404968 584960 404970
rect 580165 404912 580170 404968
rect 580226 404912 584960 404968
rect 580165 404910 584960 404912
rect 580165 404907 580231 404910
rect 583520 404820 584960 404910
rect 361573 403610 361639 403613
rect 359812 403608 361639 403610
rect 359812 403552 361578 403608
rect 361634 403552 361639 403608
rect 359812 403550 361639 403552
rect 361573 403547 361639 403550
rect -960 397490 480 397580
rect 3785 397490 3851 397493
rect -960 397488 3851 397490
rect -960 397432 3790 397488
rect 3846 397432 3851 397488
rect -960 397430 3851 397432
rect -960 397340 480 397430
rect 3785 397427 3851 397430
rect 361573 392594 361639 392597
rect 359812 392592 361639 392594
rect 359812 392536 361578 392592
rect 361634 392536 361639 392592
rect 359812 392534 361639 392536
rect 361573 392531 361639 392534
rect 583520 391628 584960 391868
rect 472157 389060 472223 389061
rect 474365 389060 474431 389061
rect 472157 389058 472204 389060
rect 472112 389056 472204 389058
rect 472112 389000 472162 389056
rect 472112 388998 472204 389000
rect 472157 388996 472204 388998
rect 472268 388996 472274 389060
rect 474365 389058 474412 389060
rect 474320 389056 474412 389058
rect 474320 389000 474370 389056
rect 474320 388998 474412 389000
rect 474365 388996 474412 388998
rect 474476 388996 474482 389060
rect 474774 388996 474780 389060
rect 474844 389058 474850 389060
rect 475101 389058 475167 389061
rect 474844 389056 475167 389058
rect 474844 389000 475106 389056
rect 475162 389000 475167 389056
rect 474844 388998 475167 389000
rect 474844 388996 474850 388998
rect 472157 388995 472223 388996
rect 474365 388995 474431 388996
rect 475101 388995 475167 388998
rect 476430 388996 476436 389060
rect 476500 389058 476506 389060
rect 477309 389058 477375 389061
rect 476500 389056 477375 389058
rect 476500 389000 477314 389056
rect 477370 389000 477375 389056
rect 476500 388998 477375 389000
rect 476500 388996 476506 388998
rect 477309 388995 477375 388998
rect 478822 388996 478828 389060
rect 478892 389058 478898 389060
rect 479517 389058 479583 389061
rect 478892 389056 479583 389058
rect 478892 389000 479522 389056
rect 479578 389000 479583 389056
rect 478892 388998 479583 389000
rect 478892 388996 478898 388998
rect 479517 388995 479583 388998
rect 472014 388860 472020 388924
rect 472084 388922 472090 388924
rect 472893 388922 472959 388925
rect 472084 388920 472959 388922
rect 472084 388864 472898 388920
rect 472954 388864 472959 388920
rect 472084 388862 472959 388864
rect 472084 388860 472090 388862
rect 472893 388859 472959 388862
rect 448278 388316 448284 388380
rect 448348 388378 448354 388380
rect 464337 388378 464403 388381
rect 448348 388376 464403 388378
rect 448348 388320 464342 388376
rect 464398 388320 464403 388376
rect 448348 388318 464403 388320
rect 448348 388316 448354 388318
rect 464337 388315 464403 388318
rect 449065 387018 449131 387021
rect 489310 387018 489316 387020
rect 449065 387016 489316 387018
rect 449065 386960 449070 387016
rect 449126 386960 489316 387016
rect 449065 386958 489316 386960
rect 449065 386955 449131 386958
rect 489310 386956 489316 386958
rect 489380 386956 489386 387020
rect 513281 384706 513347 384709
rect 509956 384704 513347 384706
rect 509956 384648 513286 384704
rect 513342 384648 513347 384704
rect 509956 384646 513347 384648
rect 513281 384643 513347 384646
rect -960 384284 480 384524
rect 512453 384162 512519 384165
rect 509956 384160 512519 384162
rect 509956 384104 512458 384160
rect 512514 384104 512519 384160
rect 509956 384102 512519 384104
rect 512453 384099 512519 384102
rect 447133 383890 447199 383893
rect 447133 383888 450156 383890
rect 447133 383832 447138 383888
rect 447194 383832 450156 383888
rect 447133 383830 450156 383832
rect 447133 383827 447199 383830
rect 512637 383618 512703 383621
rect 509956 383616 512703 383618
rect 509956 383560 512642 383616
rect 512698 383560 512703 383616
rect 509956 383558 512703 383560
rect 512637 383555 512703 383558
rect 447133 383210 447199 383213
rect 447133 383208 450156 383210
rect 447133 383152 447138 383208
rect 447194 383152 450156 383208
rect 447133 383150 450156 383152
rect 447133 383147 447199 383150
rect 513005 383074 513071 383077
rect 509956 383072 513071 383074
rect 509956 383016 513010 383072
rect 513066 383016 513071 383072
rect 509956 383014 513071 383016
rect 513005 383011 513071 383014
rect 447225 382530 447291 382533
rect 512453 382530 512519 382533
rect 447225 382528 450156 382530
rect 447225 382472 447230 382528
rect 447286 382472 450156 382528
rect 447225 382470 450156 382472
rect 509956 382528 512519 382530
rect 509956 382472 512458 382528
rect 512514 382472 512519 382528
rect 509956 382470 512519 382472
rect 447225 382467 447291 382470
rect 512453 382467 512519 382470
rect 513097 381986 513163 381989
rect 509956 381984 513163 381986
rect 509956 381928 513102 381984
rect 513158 381928 513163 381984
rect 509956 381926 513163 381928
rect 513097 381923 513163 381926
rect 447133 381850 447199 381853
rect 447133 381848 450156 381850
rect 447133 381792 447138 381848
rect 447194 381792 450156 381848
rect 447133 381790 450156 381792
rect 447133 381787 447199 381790
rect 361573 381578 361639 381581
rect 359812 381576 361639 381578
rect 359812 381520 361578 381576
rect 361634 381520 361639 381576
rect 359812 381518 361639 381520
rect 361573 381515 361639 381518
rect 513281 381442 513347 381445
rect 509956 381440 513347 381442
rect 509956 381384 513286 381440
rect 513342 381384 513347 381440
rect 509956 381382 513347 381384
rect 513281 381379 513347 381382
rect 447225 381170 447291 381173
rect 447225 381168 450156 381170
rect 447225 381112 447230 381168
rect 447286 381112 450156 381168
rect 447225 381110 450156 381112
rect 447225 381107 447291 381110
rect 513189 380898 513255 380901
rect 509956 380896 513255 380898
rect 509956 380840 513194 380896
rect 513250 380840 513255 380896
rect 509956 380838 513255 380840
rect 513189 380835 513255 380838
rect 447133 380490 447199 380493
rect 447133 380488 450156 380490
rect 447133 380432 447138 380488
rect 447194 380432 450156 380488
rect 447133 380430 450156 380432
rect 447133 380427 447199 380430
rect 513281 380354 513347 380357
rect 509956 380352 513347 380354
rect 509956 380296 513286 380352
rect 513342 380296 513347 380352
rect 509956 380294 513347 380296
rect 513281 380291 513347 380294
rect 447225 379810 447291 379813
rect 512545 379810 512611 379813
rect 447225 379808 450156 379810
rect 447225 379752 447230 379808
rect 447286 379752 450156 379808
rect 447225 379750 450156 379752
rect 509956 379808 512611 379810
rect 509956 379752 512550 379808
rect 512606 379752 512611 379808
rect 509956 379750 512611 379752
rect 447225 379747 447291 379750
rect 512545 379747 512611 379750
rect 512913 379266 512979 379269
rect 509956 379264 512979 379266
rect 509956 379208 512918 379264
rect 512974 379208 512979 379264
rect 509956 379206 512979 379208
rect 512913 379203 512979 379206
rect 447133 379130 447199 379133
rect 447133 379128 450156 379130
rect 447133 379072 447138 379128
rect 447194 379072 450156 379128
rect 447133 379070 450156 379072
rect 447133 379067 447199 379070
rect 512453 378722 512519 378725
rect 509956 378720 512519 378722
rect 509956 378664 512458 378720
rect 512514 378664 512519 378720
rect 509956 378662 512519 378664
rect 512453 378659 512519 378662
rect 447225 378450 447291 378453
rect 580717 378450 580783 378453
rect 583520 378450 584960 378540
rect 447225 378448 450156 378450
rect 447225 378392 447230 378448
rect 447286 378392 450156 378448
rect 447225 378390 450156 378392
rect 580717 378448 584960 378450
rect 580717 378392 580722 378448
rect 580778 378392 584960 378448
rect 580717 378390 584960 378392
rect 447225 378387 447291 378390
rect 580717 378387 580783 378390
rect 583520 378300 584960 378390
rect 512269 378178 512335 378181
rect 509956 378176 512335 378178
rect 509956 378120 512274 378176
rect 512330 378120 512335 378176
rect 509956 378118 512335 378120
rect 512269 378115 512335 378118
rect 447133 377770 447199 377773
rect 447133 377768 450156 377770
rect 447133 377712 447138 377768
rect 447194 377712 450156 377768
rect 447133 377710 450156 377712
rect 447133 377707 447199 377710
rect 512085 377634 512151 377637
rect 509956 377632 512151 377634
rect 509956 377576 512090 377632
rect 512146 377576 512151 377632
rect 509956 377574 512151 377576
rect 512085 377571 512151 377574
rect 447225 377090 447291 377093
rect 512637 377090 512703 377093
rect 447225 377088 450156 377090
rect 447225 377032 447230 377088
rect 447286 377032 450156 377088
rect 447225 377030 450156 377032
rect 509956 377088 512703 377090
rect 509956 377032 512642 377088
rect 512698 377032 512703 377088
rect 509956 377030 512703 377032
rect 447225 377027 447291 377030
rect 512637 377027 512703 377030
rect 512177 376546 512243 376549
rect 509956 376544 512243 376546
rect 509956 376488 512182 376544
rect 512238 376488 512243 376544
rect 509956 376486 512243 376488
rect 512177 376483 512243 376486
rect 447133 376410 447199 376413
rect 447133 376408 450156 376410
rect 447133 376352 447138 376408
rect 447194 376352 450156 376408
rect 447133 376350 450156 376352
rect 447133 376347 447199 376350
rect 512637 376002 512703 376005
rect 509956 376000 512703 376002
rect 509956 375944 512642 376000
rect 512698 375944 512703 376000
rect 509956 375942 512703 375944
rect 512637 375939 512703 375942
rect 447225 375730 447291 375733
rect 447225 375728 450156 375730
rect 447225 375672 447230 375728
rect 447286 375672 450156 375728
rect 447225 375670 450156 375672
rect 447225 375667 447291 375670
rect 512821 375458 512887 375461
rect 509956 375456 512887 375458
rect 509956 375400 512826 375456
rect 512882 375400 512887 375456
rect 509956 375398 512887 375400
rect 512821 375395 512887 375398
rect 447133 375050 447199 375053
rect 447133 375048 450156 375050
rect 447133 374992 447138 375048
rect 447194 374992 450156 375048
rect 447133 374990 450156 374992
rect 447133 374987 447199 374990
rect 511993 374914 512059 374917
rect 509956 374912 512059 374914
rect 509956 374856 511998 374912
rect 512054 374856 512059 374912
rect 509956 374854 512059 374856
rect 511993 374851 512059 374854
rect 447225 374370 447291 374373
rect 513281 374370 513347 374373
rect 447225 374368 450156 374370
rect 447225 374312 447230 374368
rect 447286 374312 450156 374368
rect 447225 374310 450156 374312
rect 509956 374368 513347 374370
rect 509956 374312 513286 374368
rect 513342 374312 513347 374368
rect 509956 374310 513347 374312
rect 447225 374307 447291 374310
rect 513281 374307 513347 374310
rect 512637 373826 512703 373829
rect 509956 373824 512703 373826
rect 509956 373768 512642 373824
rect 512698 373768 512703 373824
rect 509956 373766 512703 373768
rect 512637 373763 512703 373766
rect 447133 373690 447199 373693
rect 447133 373688 450156 373690
rect 447133 373632 447138 373688
rect 447194 373632 450156 373688
rect 447133 373630 450156 373632
rect 447133 373627 447199 373630
rect 512453 373282 512519 373285
rect 509956 373280 512519 373282
rect 509956 373224 512458 373280
rect 512514 373224 512519 373280
rect 509956 373222 512519 373224
rect 512453 373219 512519 373222
rect 447225 373010 447291 373013
rect 447225 373008 450156 373010
rect 447225 372952 447230 373008
rect 447286 372952 450156 373008
rect 447225 372950 450156 372952
rect 447225 372947 447291 372950
rect 512085 372738 512151 372741
rect 509956 372736 512151 372738
rect 509956 372680 512090 372736
rect 512146 372680 512151 372736
rect 509956 372678 512151 372680
rect 512085 372675 512151 372678
rect 447133 372330 447199 372333
rect 447133 372328 450156 372330
rect 447133 372272 447138 372328
rect 447194 372272 450156 372328
rect 447133 372270 450156 372272
rect 447133 372267 447199 372270
rect 512821 372194 512887 372197
rect 509956 372192 512887 372194
rect 509956 372136 512826 372192
rect 512882 372136 512887 372192
rect 509956 372134 512887 372136
rect 512821 372131 512887 372134
rect 447225 371650 447291 371653
rect 512177 371650 512243 371653
rect 447225 371648 450156 371650
rect 447225 371592 447230 371648
rect 447286 371592 450156 371648
rect 447225 371590 450156 371592
rect 509956 371648 512243 371650
rect 509956 371592 512182 371648
rect 512238 371592 512243 371648
rect 509956 371590 512243 371592
rect 447225 371587 447291 371590
rect 512177 371587 512243 371590
rect -960 371378 480 371468
rect 3877 371378 3943 371381
rect -960 371376 3943 371378
rect -960 371320 3882 371376
rect 3938 371320 3943 371376
rect -960 371318 3943 371320
rect -960 371228 480 371318
rect 3877 371315 3943 371318
rect 512637 371106 512703 371109
rect 509956 371104 512703 371106
rect 509956 371048 512642 371104
rect 512698 371048 512703 371104
rect 509956 371046 512703 371048
rect 512637 371043 512703 371046
rect 447133 370970 447199 370973
rect 447133 370968 450156 370970
rect 447133 370912 447138 370968
rect 447194 370912 450156 370968
rect 447133 370910 450156 370912
rect 447133 370907 447199 370910
rect 361573 370562 361639 370565
rect 359812 370560 361639 370562
rect 359812 370504 361578 370560
rect 361634 370504 361639 370560
rect 359812 370502 361639 370504
rect 361573 370499 361639 370502
rect 447225 370290 447291 370293
rect 447225 370288 450156 370290
rect 447225 370232 447230 370288
rect 447286 370232 450156 370288
rect 447225 370230 450156 370232
rect 447225 370227 447291 370230
rect 509742 370157 509802 370532
rect 509693 370152 509802 370157
rect 509693 370096 509698 370152
rect 509754 370096 509802 370152
rect 509693 370094 509802 370096
rect 509693 370091 509759 370094
rect 513281 370018 513347 370021
rect 509956 370016 513347 370018
rect 509956 369960 513286 370016
rect 513342 369960 513347 370016
rect 509956 369958 513347 369960
rect 513281 369955 513347 369958
rect 447133 369610 447199 369613
rect 447133 369608 450156 369610
rect 447133 369552 447138 369608
rect 447194 369552 450156 369608
rect 447133 369550 450156 369552
rect 447133 369547 447199 369550
rect 513281 369474 513347 369477
rect 509956 369472 513347 369474
rect 509956 369416 513286 369472
rect 513342 369416 513347 369472
rect 509956 369414 513347 369416
rect 513281 369411 513347 369414
rect 447225 368930 447291 368933
rect 512821 368930 512887 368933
rect 447225 368928 450156 368930
rect 447225 368872 447230 368928
rect 447286 368872 450156 368928
rect 447225 368870 450156 368872
rect 509956 368928 512887 368930
rect 509956 368872 512826 368928
rect 512882 368872 512887 368928
rect 509956 368870 512887 368872
rect 447225 368867 447291 368870
rect 512821 368867 512887 368870
rect 512085 368386 512151 368389
rect 509956 368384 512151 368386
rect 509956 368328 512090 368384
rect 512146 368328 512151 368384
rect 509956 368326 512151 368328
rect 512085 368323 512151 368326
rect 447225 368250 447291 368253
rect 447225 368248 450156 368250
rect 447225 368192 447230 368248
rect 447286 368192 450156 368248
rect 447225 368190 450156 368192
rect 447225 368187 447291 368190
rect 511993 367842 512059 367845
rect 509956 367840 512059 367842
rect 509956 367784 511998 367840
rect 512054 367784 512059 367840
rect 509956 367782 512059 367784
rect 511993 367779 512059 367782
rect 447133 367570 447199 367573
rect 447133 367568 450156 367570
rect 447133 367512 447138 367568
rect 447194 367512 450156 367568
rect 447133 367510 450156 367512
rect 447133 367507 447199 367510
rect 513281 367298 513347 367301
rect 509956 367296 513347 367298
rect 509956 367240 513286 367296
rect 513342 367240 513347 367296
rect 509956 367238 513347 367240
rect 513281 367235 513347 367238
rect 447133 366890 447199 366893
rect 447133 366888 450156 366890
rect 447133 366832 447138 366888
rect 447194 366832 450156 366888
rect 447133 366830 450156 366832
rect 447133 366827 447199 366830
rect 513281 366754 513347 366757
rect 509956 366752 513347 366754
rect 509956 366696 513286 366752
rect 513342 366696 513347 366752
rect 509956 366694 513347 366696
rect 513281 366691 513347 366694
rect 447225 366210 447291 366213
rect 511993 366210 512059 366213
rect 447225 366208 450156 366210
rect 447225 366152 447230 366208
rect 447286 366152 450156 366208
rect 447225 366150 450156 366152
rect 509956 366208 512059 366210
rect 509956 366152 511998 366208
rect 512054 366152 512059 366208
rect 509956 366150 512059 366152
rect 447225 366147 447291 366150
rect 511993 366147 512059 366150
rect 513281 365666 513347 365669
rect 509956 365664 513347 365666
rect 509956 365608 513286 365664
rect 513342 365608 513347 365664
rect 509956 365606 513347 365608
rect 513281 365603 513347 365606
rect 447225 365530 447291 365533
rect 447225 365528 450156 365530
rect 447225 365472 447230 365528
rect 447286 365472 450156 365528
rect 447225 365470 450156 365472
rect 447225 365467 447291 365470
rect 512637 365122 512703 365125
rect 509956 365120 512703 365122
rect 509956 365064 512642 365120
rect 512698 365064 512703 365120
rect 509956 365062 512703 365064
rect 512637 365059 512703 365062
rect 580165 365122 580231 365125
rect 583520 365122 584960 365212
rect 580165 365120 584960 365122
rect 580165 365064 580170 365120
rect 580226 365064 584960 365120
rect 580165 365062 584960 365064
rect 580165 365059 580231 365062
rect 583520 364972 584960 365062
rect 447133 364850 447199 364853
rect 447133 364848 450156 364850
rect 447133 364792 447138 364848
rect 447194 364792 450156 364848
rect 447133 364790 450156 364792
rect 447133 364787 447199 364790
rect 513281 364578 513347 364581
rect 509956 364576 513347 364578
rect 509956 364520 513286 364576
rect 513342 364520 513347 364576
rect 509956 364518 513347 364520
rect 513281 364515 513347 364518
rect 447225 364170 447291 364173
rect 447225 364168 450156 364170
rect 447225 364112 447230 364168
rect 447286 364112 450156 364168
rect 447225 364110 450156 364112
rect 447225 364107 447291 364110
rect 512177 364034 512243 364037
rect 509956 364032 512243 364034
rect 509956 363976 512182 364032
rect 512238 363976 512243 364032
rect 509956 363974 512243 363976
rect 512177 363971 512243 363974
rect 447133 363490 447199 363493
rect 513281 363490 513347 363493
rect 447133 363488 450156 363490
rect 447133 363432 447138 363488
rect 447194 363432 450156 363488
rect 447133 363430 450156 363432
rect 509956 363488 513347 363490
rect 509956 363432 513286 363488
rect 513342 363432 513347 363488
rect 509956 363430 513347 363432
rect 447133 363427 447199 363430
rect 513281 363427 513347 363430
rect 513005 362946 513071 362949
rect 509956 362944 513071 362946
rect 509956 362888 513010 362944
rect 513066 362888 513071 362944
rect 509956 362886 513071 362888
rect 513005 362883 513071 362886
rect 447133 362810 447199 362813
rect 447133 362808 450156 362810
rect 447133 362752 447138 362808
rect 447194 362752 450156 362808
rect 447133 362750 450156 362752
rect 447133 362747 447199 362750
rect 512177 362402 512243 362405
rect 509956 362400 512243 362402
rect 509956 362344 512182 362400
rect 512238 362344 512243 362400
rect 509956 362342 512243 362344
rect 512177 362339 512243 362342
rect 447225 362130 447291 362133
rect 447225 362128 450156 362130
rect 447225 362072 447230 362128
rect 447286 362072 450156 362128
rect 447225 362070 450156 362072
rect 447225 362067 447291 362070
rect 512361 361858 512427 361861
rect 509956 361856 512427 361858
rect 509956 361800 512366 361856
rect 512422 361800 512427 361856
rect 509956 361798 512427 361800
rect 512361 361795 512427 361798
rect 447225 361450 447291 361453
rect 447225 361448 450156 361450
rect 447225 361392 447230 361448
rect 447286 361392 450156 361448
rect 447225 361390 450156 361392
rect 447225 361387 447291 361390
rect 513005 361314 513071 361317
rect 509956 361312 513071 361314
rect 509956 361256 513010 361312
rect 513066 361256 513071 361312
rect 509956 361254 513071 361256
rect 513005 361251 513071 361254
rect 447133 360770 447199 360773
rect 447133 360768 450156 360770
rect 447133 360712 447138 360768
rect 447194 360712 450156 360768
rect 447133 360710 450156 360712
rect 447133 360707 447199 360710
rect 509926 360365 509986 360740
rect 509877 360360 509986 360365
rect 509877 360304 509882 360360
rect 509938 360304 509986 360360
rect 509877 360302 509986 360304
rect 509877 360299 509943 360302
rect 513281 360226 513347 360229
rect 509956 360224 513347 360226
rect 509956 360168 513286 360224
rect 513342 360168 513347 360224
rect 509956 360166 513347 360168
rect 513281 360163 513347 360166
rect 447133 360090 447199 360093
rect 447133 360088 450156 360090
rect 447133 360032 447138 360088
rect 447194 360032 450156 360088
rect 447133 360030 450156 360032
rect 447133 360027 447199 360030
rect 511073 359682 511139 359685
rect 509956 359680 511139 359682
rect 509956 359624 511078 359680
rect 511134 359624 511139 359680
rect 509956 359622 511139 359624
rect 511073 359619 511139 359622
rect 362217 359546 362283 359549
rect 359812 359544 362283 359546
rect 359812 359488 362222 359544
rect 362278 359488 362283 359544
rect 359812 359486 362283 359488
rect 362217 359483 362283 359486
rect 447225 359410 447291 359413
rect 447225 359408 450156 359410
rect 447225 359352 447230 359408
rect 447286 359352 450156 359408
rect 447225 359350 450156 359352
rect 447225 359347 447291 359350
rect 510613 359138 510679 359141
rect 509956 359136 510679 359138
rect 509956 359080 510618 359136
rect 510674 359080 510679 359136
rect 509956 359078 510679 359080
rect 510613 359075 510679 359078
rect 448973 358730 449039 358733
rect 448973 358728 450156 358730
rect 448973 358672 448978 358728
rect 449034 358672 450156 358728
rect 448973 358670 450156 358672
rect 448973 358667 449039 358670
rect 512269 358594 512335 358597
rect 509956 358592 512335 358594
rect -960 358458 480 358548
rect 509956 358536 512274 358592
rect 512330 358536 512335 358592
rect 509956 358534 512335 358536
rect 512269 358531 512335 358534
rect 3509 358458 3575 358461
rect -960 358456 3575 358458
rect -960 358400 3514 358456
rect 3570 358400 3575 358456
rect -960 358398 3575 358400
rect -960 358308 480 358398
rect 3509 358395 3575 358398
rect 449525 358050 449591 358053
rect 512177 358050 512243 358053
rect 449525 358048 450156 358050
rect 449525 357992 449530 358048
rect 449586 357992 450156 358048
rect 449525 357990 450156 357992
rect 509956 358048 512243 358050
rect 509956 357992 512182 358048
rect 512238 357992 512243 358048
rect 509956 357990 512243 357992
rect 449525 357987 449591 357990
rect 512177 357987 512243 357990
rect 509969 357642 510035 357645
rect 509926 357640 510035 357642
rect 509926 357584 509974 357640
rect 510030 357584 510035 357640
rect 509926 357579 510035 357584
rect 509926 357476 509986 357579
rect 449065 357370 449131 357373
rect 449065 357368 450156 357370
rect 449065 357312 449070 357368
rect 449126 357312 450156 357368
rect 449065 357310 450156 357312
rect 449065 357307 449131 357310
rect 513281 356962 513347 356965
rect 509956 356960 513347 356962
rect 509956 356904 513286 356960
rect 513342 356904 513347 356960
rect 509956 356902 513347 356904
rect 513281 356899 513347 356902
rect 449617 356690 449683 356693
rect 449617 356688 450156 356690
rect 449617 356632 449622 356688
rect 449678 356632 450156 356688
rect 449617 356630 450156 356632
rect 449617 356627 449683 356630
rect 510061 356418 510127 356421
rect 509956 356416 510127 356418
rect 509956 356360 510066 356416
rect 510122 356360 510127 356416
rect 509956 356358 510127 356360
rect 510061 356355 510127 356358
rect 447409 356010 447475 356013
rect 447409 356008 450156 356010
rect 447409 355952 447414 356008
rect 447470 355952 450156 356008
rect 447409 355950 450156 355952
rect 447409 355947 447475 355950
rect 510889 355874 510955 355877
rect 509956 355872 510955 355874
rect 509956 355816 510894 355872
rect 510950 355816 510955 355872
rect 509956 355814 510955 355816
rect 510889 355811 510955 355814
rect 448237 355330 448303 355333
rect 512361 355330 512427 355333
rect 448237 355328 450156 355330
rect 448237 355272 448242 355328
rect 448298 355272 450156 355328
rect 448237 355270 450156 355272
rect 509956 355328 512427 355330
rect 509956 355272 512366 355328
rect 512422 355272 512427 355328
rect 509956 355270 512427 355272
rect 448237 355267 448303 355270
rect 512361 355267 512427 355270
rect 513281 354786 513347 354789
rect 509956 354784 513347 354786
rect 509956 354728 513286 354784
rect 513342 354728 513347 354784
rect 509956 354726 513347 354728
rect 513281 354723 513347 354726
rect 447685 354650 447751 354653
rect 447685 354648 450156 354650
rect 447685 354592 447690 354648
rect 447746 354592 450156 354648
rect 447685 354590 450156 354592
rect 447685 354587 447751 354590
rect 512453 354242 512519 354245
rect 509956 354240 512519 354242
rect 509956 354184 512458 354240
rect 512514 354184 512519 354240
rect 509956 354182 512519 354184
rect 512453 354179 512519 354182
rect 447593 353970 447659 353973
rect 447593 353968 450156 353970
rect 447593 353912 447598 353968
rect 447654 353912 450156 353968
rect 447593 353910 450156 353912
rect 447593 353907 447659 353910
rect 513189 353698 513255 353701
rect 509956 353696 513255 353698
rect 509956 353640 513194 353696
rect 513250 353640 513255 353696
rect 509956 353638 513255 353640
rect 513189 353635 513255 353638
rect 447869 353290 447935 353293
rect 447869 353288 450156 353290
rect 447869 353232 447874 353288
rect 447930 353232 450156 353288
rect 447869 353230 450156 353232
rect 447869 353227 447935 353230
rect 510705 353154 510771 353157
rect 509956 353152 510771 353154
rect 509956 353096 510710 353152
rect 510766 353096 510771 353152
rect 509956 353094 510771 353096
rect 510705 353091 510771 353094
rect 448145 352610 448211 352613
rect 512453 352610 512519 352613
rect 448145 352608 450156 352610
rect 448145 352552 448150 352608
rect 448206 352552 450156 352608
rect 448145 352550 450156 352552
rect 509956 352608 512519 352610
rect 509956 352552 512458 352608
rect 512514 352552 512519 352608
rect 509956 352550 512519 352552
rect 448145 352547 448211 352550
rect 512453 352547 512519 352550
rect 513281 352066 513347 352069
rect 509956 352064 513347 352066
rect 509956 352008 513286 352064
rect 513342 352008 513347 352064
rect 509956 352006 513347 352008
rect 513281 352003 513347 352006
rect 447133 351930 447199 351933
rect 580165 351930 580231 351933
rect 583520 351930 584960 352020
rect 447133 351928 450156 351930
rect 447133 351872 447138 351928
rect 447194 351872 450156 351928
rect 447133 351870 450156 351872
rect 580165 351928 584960 351930
rect 580165 351872 580170 351928
rect 580226 351872 584960 351928
rect 580165 351870 584960 351872
rect 447133 351867 447199 351870
rect 580165 351867 580231 351870
rect 583520 351780 584960 351870
rect 513281 351522 513347 351525
rect 509956 351520 513347 351522
rect 509956 351464 513286 351520
rect 513342 351464 513347 351520
rect 509956 351462 513347 351464
rect 513281 351459 513347 351462
rect 448237 351250 448303 351253
rect 448237 351248 450156 351250
rect 448237 351192 448242 351248
rect 448298 351192 450156 351248
rect 448237 351190 450156 351192
rect 448237 351187 448303 351190
rect 512453 350978 512519 350981
rect 509956 350976 512519 350978
rect 509956 350920 512458 350976
rect 512514 350920 512519 350976
rect 509956 350918 512519 350920
rect 512453 350915 512519 350918
rect 447133 350570 447199 350573
rect 447133 350568 450156 350570
rect 447133 350512 447138 350568
rect 447194 350512 450156 350568
rect 447133 350510 450156 350512
rect 447133 350507 447199 350510
rect 512453 350434 512519 350437
rect 509956 350432 512519 350434
rect 509956 350376 512458 350432
rect 512514 350376 512519 350432
rect 509956 350374 512519 350376
rect 512453 350371 512519 350374
rect 447593 349890 447659 349893
rect 513281 349890 513347 349893
rect 447593 349888 450156 349890
rect 447593 349832 447598 349888
rect 447654 349832 450156 349888
rect 447593 349830 450156 349832
rect 509956 349888 513347 349890
rect 509956 349832 513286 349888
rect 513342 349832 513347 349888
rect 509956 349830 513347 349832
rect 447593 349827 447659 349830
rect 513281 349827 513347 349830
rect 512453 349346 512519 349349
rect 509956 349344 512519 349346
rect 509956 349288 512458 349344
rect 512514 349288 512519 349344
rect 509956 349286 512519 349288
rect 512453 349283 512519 349286
rect 448278 349148 448284 349212
rect 448348 349210 448354 349212
rect 448348 349150 450156 349210
rect 448348 349148 448354 349150
rect 511165 348802 511231 348805
rect 509956 348800 511231 348802
rect 509956 348744 511170 348800
rect 511226 348744 511231 348800
rect 509956 348742 511231 348744
rect 511165 348739 511231 348742
rect 361757 348530 361823 348533
rect 359812 348528 361823 348530
rect 359812 348472 361762 348528
rect 361818 348472 361823 348528
rect 359812 348470 361823 348472
rect 361757 348467 361823 348470
rect 448329 348530 448395 348533
rect 448329 348528 450156 348530
rect 448329 348472 448334 348528
rect 448390 348472 450156 348528
rect 448329 348470 450156 348472
rect 448329 348467 448395 348470
rect 513005 348258 513071 348261
rect 509956 348256 513071 348258
rect 509956 348200 513010 348256
rect 513066 348200 513071 348256
rect 509956 348198 513071 348200
rect 513005 348195 513071 348198
rect 449341 347850 449407 347853
rect 449341 347848 450156 347850
rect 449341 347792 449346 347848
rect 449402 347792 450156 347848
rect 449341 347790 450156 347792
rect 449341 347787 449407 347790
rect 512453 347714 512519 347717
rect 509956 347712 512519 347714
rect 509956 347656 512458 347712
rect 512514 347656 512519 347712
rect 509956 347654 512519 347656
rect 512453 347651 512519 347654
rect 447133 347170 447199 347173
rect 512821 347170 512887 347173
rect 447133 347168 450156 347170
rect 447133 347112 447138 347168
rect 447194 347112 450156 347168
rect 447133 347110 450156 347112
rect 509956 347168 512887 347170
rect 509956 347112 512826 347168
rect 512882 347112 512887 347168
rect 509956 347110 512887 347112
rect 447133 347107 447199 347110
rect 512821 347107 512887 347110
rect 513281 346626 513347 346629
rect 509956 346624 513347 346626
rect 509956 346568 513286 346624
rect 513342 346568 513347 346624
rect 509956 346566 513347 346568
rect 513281 346563 513347 346566
rect 449709 346490 449775 346493
rect 449709 346488 450156 346490
rect 449709 346432 449714 346488
rect 449770 346432 450156 346488
rect 449709 346430 450156 346432
rect 449709 346427 449775 346430
rect 512453 346082 512519 346085
rect 509956 346080 512519 346082
rect 509956 346024 512458 346080
rect 512514 346024 512519 346080
rect 509956 346022 512519 346024
rect 512453 346019 512519 346022
rect 449801 345810 449867 345813
rect 449801 345808 450156 345810
rect 449801 345752 449806 345808
rect 449862 345752 450156 345808
rect 449801 345750 450156 345752
rect 449801 345747 449867 345750
rect 512453 345538 512519 345541
rect 509956 345536 512519 345538
rect -960 345402 480 345492
rect 509956 345480 512458 345536
rect 512514 345480 512519 345536
rect 509956 345478 512519 345480
rect 512453 345475 512519 345478
rect 3417 345402 3483 345405
rect -960 345400 3483 345402
rect -960 345344 3422 345400
rect 3478 345344 3483 345400
rect -960 345342 3483 345344
rect -960 345252 480 345342
rect 3417 345339 3483 345342
rect 449801 345130 449867 345133
rect 449801 345128 450156 345130
rect 449801 345072 449806 345128
rect 449862 345072 450156 345128
rect 449801 345070 450156 345072
rect 449801 345067 449867 345070
rect 513005 344994 513071 344997
rect 509956 344992 513071 344994
rect 509956 344936 513010 344992
rect 513066 344936 513071 344992
rect 509956 344934 513071 344936
rect 513005 344931 513071 344934
rect 448329 344450 448395 344453
rect 510889 344450 510955 344453
rect 448329 344448 450156 344450
rect 448329 344392 448334 344448
rect 448390 344392 450156 344448
rect 448329 344390 450156 344392
rect 509956 344448 510955 344450
rect 509956 344392 510894 344448
rect 510950 344392 510955 344448
rect 509956 344390 510955 344392
rect 448329 344387 448395 344390
rect 510889 344387 510955 344390
rect 513281 343906 513347 343909
rect 509956 343904 513347 343906
rect 509956 343848 513286 343904
rect 513342 343848 513347 343904
rect 509956 343846 513347 343848
rect 513281 343843 513347 343846
rect 449341 343770 449407 343773
rect 449341 343768 450156 343770
rect 449341 343712 449346 343768
rect 449402 343712 450156 343768
rect 449341 343710 450156 343712
rect 449341 343707 449407 343710
rect 513005 343362 513071 343365
rect 509956 343360 513071 343362
rect 509956 343304 513010 343360
rect 513066 343304 513071 343360
rect 509956 343302 513071 343304
rect 513005 343299 513071 343302
rect 448421 343090 448487 343093
rect 448421 343088 450156 343090
rect 448421 343032 448426 343088
rect 448482 343032 450156 343088
rect 448421 343030 450156 343032
rect 448421 343027 448487 343030
rect 510981 342818 511047 342821
rect 509956 342816 511047 342818
rect 509956 342760 510986 342816
rect 511042 342760 511047 342816
rect 509956 342758 511047 342760
rect 510981 342755 511047 342758
rect 449433 342410 449499 342413
rect 449433 342408 450156 342410
rect 449433 342352 449438 342408
rect 449494 342352 450156 342408
rect 449433 342350 450156 342352
rect 449433 342347 449499 342350
rect 512545 342274 512611 342277
rect 509956 342272 512611 342274
rect 509956 342216 512550 342272
rect 512606 342216 512611 342272
rect 509956 342214 512611 342216
rect 512545 342211 512611 342214
rect 447225 341730 447291 341733
rect 513281 341730 513347 341733
rect 447225 341728 450156 341730
rect 447225 341672 447230 341728
rect 447286 341672 450156 341728
rect 447225 341670 450156 341672
rect 509956 341728 513347 341730
rect 509956 341672 513286 341728
rect 513342 341672 513347 341728
rect 509956 341670 513347 341672
rect 447225 341667 447291 341670
rect 513281 341667 513347 341670
rect 513281 341186 513347 341189
rect 509956 341184 513347 341186
rect 509956 341128 513286 341184
rect 513342 341128 513347 341184
rect 509956 341126 513347 341128
rect 513281 341123 513347 341126
rect 447133 341050 447199 341053
rect 447133 341048 450156 341050
rect 447133 340992 447138 341048
rect 447194 340992 450156 341048
rect 447133 340990 450156 340992
rect 447133 340987 447199 340990
rect 513281 340642 513347 340645
rect 509956 340640 513347 340642
rect 509956 340584 513286 340640
rect 513342 340584 513347 340640
rect 509956 340582 513347 340584
rect 513281 340579 513347 340582
rect 447225 340370 447291 340373
rect 447225 340368 450156 340370
rect 447225 340312 447230 340368
rect 447286 340312 450156 340368
rect 447225 340310 450156 340312
rect 447225 340307 447291 340310
rect 513097 340098 513163 340101
rect 509956 340096 513163 340098
rect 509956 340040 513102 340096
rect 513158 340040 513163 340096
rect 509956 340038 513163 340040
rect 513097 340035 513163 340038
rect 447133 339690 447199 339693
rect 447133 339688 450156 339690
rect 447133 339632 447138 339688
rect 447194 339632 450156 339688
rect 447133 339630 450156 339632
rect 447133 339627 447199 339630
rect 513281 339554 513347 339557
rect 509956 339552 513347 339554
rect 509956 339496 513286 339552
rect 513342 339496 513347 339552
rect 509956 339494 513347 339496
rect 513281 339491 513347 339494
rect 447225 339010 447291 339013
rect 512637 339010 512703 339013
rect 447225 339008 450156 339010
rect 447225 338952 447230 339008
rect 447286 338952 450156 339008
rect 447225 338950 450156 338952
rect 509956 339008 512703 339010
rect 509956 338952 512642 339008
rect 512698 338952 512703 339008
rect 509956 338950 512703 338952
rect 447225 338947 447291 338950
rect 512637 338947 512703 338950
rect 513005 338466 513071 338469
rect 509956 338464 513071 338466
rect 509956 338408 513010 338464
rect 513066 338408 513071 338464
rect 583520 338452 584960 338692
rect 509956 338406 513071 338408
rect 513005 338403 513071 338406
rect 447133 338330 447199 338333
rect 447133 338328 450156 338330
rect 447133 338272 447138 338328
rect 447194 338272 450156 338328
rect 447133 338270 450156 338272
rect 447133 338267 447199 338270
rect 450261 338058 450327 338061
rect 450537 338058 450603 338061
rect 450261 338056 450603 338058
rect 450261 338000 450266 338056
rect 450322 338000 450542 338056
rect 450598 338000 450603 338056
rect 450261 337998 450603 338000
rect 450261 337995 450327 337998
rect 450537 337995 450603 337998
rect 512729 337922 512795 337925
rect 509956 337920 512795 337922
rect 509956 337864 512734 337920
rect 512790 337864 512795 337920
rect 509956 337862 512795 337864
rect 512729 337859 512795 337862
rect 447133 337650 447199 337653
rect 447133 337648 450156 337650
rect 447133 337592 447138 337648
rect 447194 337592 450156 337648
rect 447133 337590 450156 337592
rect 447133 337587 447199 337590
rect 361757 337514 361823 337517
rect 359812 337512 361823 337514
rect 359812 337456 361762 337512
rect 361818 337456 361823 337512
rect 359812 337454 361823 337456
rect 361757 337451 361823 337454
rect 512821 337378 512887 337381
rect 509956 337376 512887 337378
rect 509956 337320 512826 337376
rect 512882 337320 512887 337376
rect 509956 337318 512887 337320
rect 512821 337315 512887 337318
rect 427813 337106 427879 337109
rect 450261 337106 450327 337109
rect 427813 337104 450327 337106
rect 427813 337048 427818 337104
rect 427874 337048 450266 337104
rect 450322 337048 450327 337104
rect 427813 337046 450327 337048
rect 427813 337043 427879 337046
rect 450261 337043 450327 337046
rect 447225 336970 447291 336973
rect 447225 336968 450156 336970
rect 447225 336912 447230 336968
rect 447286 336912 450156 336968
rect 447225 336910 450156 336912
rect 447225 336907 447291 336910
rect 513281 336834 513347 336837
rect 509956 336832 513347 336834
rect 509956 336776 513286 336832
rect 513342 336776 513347 336832
rect 509956 336774 513347 336776
rect 513281 336771 513347 336774
rect 447133 336290 447199 336293
rect 512729 336290 512795 336293
rect 447133 336288 450156 336290
rect 447133 336232 447138 336288
rect 447194 336232 450156 336288
rect 447133 336230 450156 336232
rect 509956 336288 512795 336290
rect 509956 336232 512734 336288
rect 512790 336232 512795 336288
rect 509956 336230 512795 336232
rect 447133 336227 447199 336230
rect 512729 336227 512795 336230
rect 511206 335746 511212 335748
rect 509956 335686 511212 335746
rect 511206 335684 511212 335686
rect 511276 335684 511282 335748
rect 447133 335610 447199 335613
rect 447133 335608 450156 335610
rect 447133 335552 447138 335608
rect 447194 335552 450156 335608
rect 447133 335550 450156 335552
rect 447133 335547 447199 335550
rect 513005 335202 513071 335205
rect 509956 335200 513071 335202
rect 509956 335144 513010 335200
rect 513066 335144 513071 335200
rect 509956 335142 513071 335144
rect 513005 335139 513071 335142
rect 447225 334930 447291 334933
rect 447225 334928 450156 334930
rect 447225 334872 447230 334928
rect 447286 334872 450156 334928
rect 447225 334870 450156 334872
rect 447225 334867 447291 334870
rect 512729 334658 512795 334661
rect 509956 334656 512795 334658
rect 509956 334600 512734 334656
rect 512790 334600 512795 334656
rect 509956 334598 512795 334600
rect 512729 334595 512795 334598
rect 428089 334522 428155 334525
rect 428406 334522 428412 334524
rect 428089 334520 428412 334522
rect 428089 334464 428094 334520
rect 428150 334464 428412 334520
rect 428089 334462 428412 334464
rect 428089 334459 428155 334462
rect 428406 334460 428412 334462
rect 428476 334460 428482 334524
rect 420453 334386 420519 334389
rect 424133 334386 424199 334389
rect 425830 334386 425836 334388
rect 420453 334384 421482 334386
rect 420453 334328 420458 334384
rect 420514 334328 421482 334384
rect 420453 334326 421482 334328
rect 420453 334323 420519 334326
rect 421422 334116 421482 334326
rect 424133 334384 425836 334386
rect 424133 334328 424138 334384
rect 424194 334328 425836 334384
rect 424133 334326 425836 334328
rect 424133 334323 424199 334326
rect 425830 334324 425836 334326
rect 425900 334386 425906 334388
rect 450445 334386 450511 334389
rect 425900 334384 450511 334386
rect 425900 334328 450450 334384
rect 450506 334328 450511 334384
rect 425900 334326 450511 334328
rect 425900 334324 425906 334326
rect 450445 334323 450511 334326
rect 447133 334250 447199 334253
rect 447133 334248 450156 334250
rect 447133 334192 447138 334248
rect 447194 334192 450156 334248
rect 447133 334190 450156 334192
rect 447133 334187 447199 334190
rect 421414 334052 421420 334116
rect 421484 334114 421490 334116
rect 513281 334114 513347 334117
rect 421484 334054 448530 334114
rect 509956 334112 513347 334114
rect 509956 334056 513286 334112
rect 513342 334056 513347 334112
rect 509956 334054 513347 334056
rect 421484 334052 421490 334054
rect 448470 333978 448530 334054
rect 513281 334051 513347 334054
rect 449985 333978 450051 333981
rect 448470 333976 450051 333978
rect 448470 333920 449990 333976
rect 450046 333920 450051 333976
rect 448470 333918 450051 333920
rect 449985 333915 450051 333918
rect 447225 333570 447291 333573
rect 513465 333570 513531 333573
rect 447225 333568 450156 333570
rect 447225 333512 447230 333568
rect 447286 333512 450156 333568
rect 447225 333510 450156 333512
rect 509956 333568 513531 333570
rect 509956 333512 513470 333568
rect 513526 333512 513531 333568
rect 509956 333510 513531 333512
rect 447225 333507 447291 333510
rect 513465 333507 513531 333510
rect 510654 333026 510660 333028
rect 509956 332966 510660 333026
rect 510654 332964 510660 332966
rect 510724 332964 510730 333028
rect 432781 332890 432847 332893
rect 429916 332888 432847 332890
rect 429916 332832 432786 332888
rect 432842 332832 432847 332888
rect 429916 332830 432847 332832
rect 432781 332827 432847 332830
rect 447133 332890 447199 332893
rect 447133 332888 450156 332890
rect 447133 332832 447138 332888
rect 447194 332832 450156 332888
rect 447133 332830 450156 332832
rect 447133 332827 447199 332830
rect 512821 332482 512887 332485
rect 509956 332480 512887 332482
rect -960 332196 480 332436
rect 509956 332424 512826 332480
rect 512882 332424 512887 332480
rect 509956 332422 512887 332424
rect 512821 332419 512887 332422
rect 448145 332210 448211 332213
rect 448145 332208 450156 332210
rect 448145 332152 448150 332208
rect 448206 332152 450156 332208
rect 448145 332150 450156 332152
rect 448145 332147 448211 332150
rect 514702 331938 514708 331940
rect 509956 331878 514708 331938
rect 514702 331876 514708 331878
rect 514772 331876 514778 331940
rect 448329 331530 448395 331533
rect 448329 331528 450156 331530
rect 448329 331472 448334 331528
rect 448390 331472 450156 331528
rect 448329 331470 450156 331472
rect 448329 331467 448395 331470
rect 514886 331394 514892 331396
rect 509956 331334 514892 331394
rect 514886 331332 514892 331334
rect 514956 331332 514962 331396
rect 447777 330850 447843 330853
rect 448421 330850 448487 330853
rect 517830 330850 517836 330852
rect 447777 330848 450156 330850
rect 447777 330792 447782 330848
rect 447838 330792 448426 330848
rect 448482 330792 450156 330848
rect 447777 330790 450156 330792
rect 509956 330790 517836 330850
rect 447777 330787 447843 330790
rect 448421 330787 448487 330790
rect 517830 330788 517836 330790
rect 517900 330788 517906 330852
rect 510245 330306 510311 330309
rect 509956 330304 510311 330306
rect 509956 330248 510250 330304
rect 510306 330248 510311 330304
rect 509956 330246 510311 330248
rect 510245 330243 510311 330246
rect 447133 330170 447199 330173
rect 448053 330170 448119 330173
rect 447133 330168 450156 330170
rect 447133 330112 447138 330168
rect 447194 330112 448058 330168
rect 448114 330112 450156 330168
rect 447133 330110 450156 330112
rect 447133 330107 447199 330110
rect 448053 330107 448119 330110
rect 512821 329762 512887 329765
rect 509956 329760 512887 329762
rect 509956 329704 512826 329760
rect 512882 329704 512887 329760
rect 509956 329702 512887 329704
rect 512821 329699 512887 329702
rect 447133 329490 447199 329493
rect 447961 329490 448027 329493
rect 447133 329488 450156 329490
rect 447133 329432 447138 329488
rect 447194 329432 447966 329488
rect 448022 329432 450156 329488
rect 447133 329430 450156 329432
rect 447133 329427 447199 329430
rect 447961 329427 448027 329430
rect 432689 329218 432755 329221
rect 515070 329218 515076 329220
rect 429916 329216 432755 329218
rect 429916 329160 432694 329216
rect 432750 329160 432755 329216
rect 429916 329158 432755 329160
rect 509956 329158 515076 329218
rect 432689 329155 432755 329158
rect 515070 329156 515076 329158
rect 515140 329156 515146 329220
rect 450126 328674 450186 328780
rect 450670 328748 450676 328812
rect 450740 328748 450746 328812
rect 450678 328674 450738 328748
rect 514334 328674 514340 328676
rect 450126 328614 450738 328674
rect 509956 328614 514340 328674
rect 449893 328538 449959 328541
rect 450126 328538 450186 328614
rect 514334 328612 514340 328614
rect 514404 328612 514410 328676
rect 449893 328536 450186 328538
rect 449893 328480 449898 328536
rect 449954 328480 450186 328536
rect 449893 328478 450186 328480
rect 449893 328475 449959 328478
rect 450486 328402 450492 328404
rect 450126 328342 450492 328402
rect 449893 327858 449959 327861
rect 450126 327858 450186 328342
rect 450486 328340 450492 328342
rect 450556 328340 450562 328404
rect 510337 328130 510403 328133
rect 509956 328128 510403 328130
rect 509956 328072 510342 328128
rect 510398 328072 510403 328128
rect 509956 328070 510403 328072
rect 510337 328067 510403 328070
rect 449893 327856 450186 327858
rect 449893 327800 449898 327856
rect 449954 327800 450186 327856
rect 449893 327798 450186 327800
rect 449893 327795 449959 327798
rect 450261 327586 450327 327589
rect 510470 327586 510476 327588
rect 450261 327584 450370 327586
rect 450261 327528 450266 327584
rect 450322 327528 450370 327584
rect 450261 327523 450370 327528
rect 509956 327526 510476 327586
rect 510470 327524 510476 327526
rect 510540 327524 510546 327588
rect 450310 327420 450370 327523
rect 512821 327042 512887 327045
rect 509956 327040 512887 327042
rect 509956 326984 512826 327040
rect 512882 326984 512887 327040
rect 509956 326982 512887 326984
rect 512821 326979 512887 326982
rect 450445 326906 450511 326909
rect 450445 326904 450554 326906
rect 450445 326848 450450 326904
rect 450506 326848 450554 326904
rect 450445 326843 450554 326848
rect 450494 326740 450554 326843
rect 362217 326498 362283 326501
rect 510838 326498 510844 326500
rect 359812 326496 362283 326498
rect 359812 326440 362222 326496
rect 362278 326440 362283 326496
rect 359812 326438 362283 326440
rect 509956 326438 510844 326498
rect 362217 326435 362283 326438
rect 510838 326436 510844 326438
rect 510908 326436 510914 326500
rect 449985 326226 450051 326229
rect 449985 326224 450186 326226
rect 449985 326168 449990 326224
rect 450046 326168 450186 326224
rect 449985 326166 450186 326168
rect 449985 326163 450051 326166
rect 450126 326060 450186 326166
rect 509926 325818 509986 325924
rect 518934 325818 518940 325820
rect 509926 325758 518940 325818
rect 518934 325756 518940 325758
rect 519004 325756 519010 325820
rect 432597 325546 432663 325549
rect 429916 325544 432663 325546
rect 429916 325488 432602 325544
rect 432658 325488 432663 325544
rect 429916 325486 432663 325488
rect 432597 325483 432663 325486
rect 450445 325546 450511 325549
rect 450445 325544 450554 325546
rect 450445 325488 450450 325544
rect 450506 325488 450554 325544
rect 450445 325483 450554 325488
rect 450494 325380 450554 325483
rect 509926 325002 509986 325380
rect 580165 325274 580231 325277
rect 583520 325274 584960 325364
rect 580165 325272 584960 325274
rect 580165 325216 580170 325272
rect 580226 325216 584960 325272
rect 580165 325214 584960 325216
rect 580165 325211 580231 325214
rect 583520 325124 584960 325214
rect 510153 325002 510219 325005
rect 509926 325000 510219 325002
rect 509926 324944 510158 325000
rect 510214 324944 510219 325000
rect 509926 324942 510219 324944
rect 510153 324939 510219 324942
rect 514150 324866 514156 324868
rect 509956 324806 514156 324866
rect 514150 324804 514156 324806
rect 514220 324804 514226 324868
rect 450310 324461 450370 324700
rect 450310 324456 450419 324461
rect 450310 324400 450358 324456
rect 450414 324400 450419 324456
rect 450310 324398 450419 324400
rect 450353 324395 450419 324398
rect 510286 324322 510292 324324
rect 509956 324262 510292 324322
rect 510286 324260 510292 324262
rect 510356 324260 510362 324324
rect 450077 324186 450143 324189
rect 450077 324184 450738 324186
rect 450077 324128 450082 324184
rect 450138 324128 450738 324184
rect 450077 324126 450738 324128
rect 450077 324123 450143 324126
rect 450678 323781 450738 324126
rect 450629 323776 450738 323781
rect 511022 323778 511028 323780
rect 450629 323720 450634 323776
rect 450690 323720 450738 323776
rect 450629 323718 450738 323720
rect 509956 323718 511028 323778
rect 450629 323715 450695 323718
rect 511022 323716 511028 323718
rect 511092 323716 511098 323780
rect 509742 322965 509802 323204
rect 509693 322960 509802 322965
rect 509693 322904 509698 322960
rect 509754 322904 509802 322960
rect 509693 322902 509802 322904
rect 509693 322899 509759 322902
rect 444833 322826 444899 322829
rect 444833 322824 480270 322826
rect 444833 322768 444838 322824
rect 444894 322768 480270 322824
rect 444833 322766 480270 322768
rect 444833 322763 444899 322766
rect 439957 322690 440023 322693
rect 471053 322690 471119 322693
rect 439957 322688 471119 322690
rect 439957 322632 439962 322688
rect 440018 322632 471058 322688
rect 471114 322632 471119 322688
rect 439957 322630 471119 322632
rect 480210 322690 480270 322766
rect 482369 322690 482435 322693
rect 480210 322688 482435 322690
rect 480210 322632 482374 322688
rect 482430 322632 482435 322688
rect 480210 322630 482435 322632
rect 439957 322627 440023 322630
rect 471053 322627 471119 322630
rect 482369 322627 482435 322630
rect 447041 322554 447107 322557
rect 471881 322554 471947 322557
rect 447041 322552 471947 322554
rect 447041 322496 447046 322552
rect 447102 322496 471886 322552
rect 471942 322496 471947 322552
rect 447041 322494 471947 322496
rect 447041 322491 447107 322494
rect 471881 322491 471947 322494
rect 447910 322356 447916 322420
rect 447980 322418 447986 322420
rect 459185 322418 459251 322421
rect 447980 322416 459251 322418
rect 447980 322360 459190 322416
rect 459246 322360 459251 322416
rect 447980 322358 459251 322360
rect 447980 322356 447986 322358
rect 459185 322355 459251 322358
rect 432781 321874 432847 321877
rect 429916 321872 432847 321874
rect 429916 321816 432786 321872
rect 432842 321816 432847 321872
rect 429916 321814 432847 321816
rect 432781 321811 432847 321814
rect 507117 321874 507183 321877
rect 510470 321874 510476 321876
rect 507117 321872 510476 321874
rect 507117 321816 507122 321872
rect 507178 321816 510476 321872
rect 507117 321814 510476 321816
rect 507117 321811 507183 321814
rect 510470 321812 510476 321814
rect 510540 321812 510546 321876
rect 515070 321738 515076 321740
rect 514710 321678 515076 321738
rect 507301 321602 507367 321605
rect 514710 321602 514770 321678
rect 515070 321676 515076 321678
rect 515140 321676 515146 321740
rect 507301 321600 514770 321602
rect 507301 321544 507306 321600
rect 507362 321544 514770 321600
rect 507301 321542 514770 321544
rect 507301 321539 507367 321542
rect 444046 321404 444052 321468
rect 444116 321466 444122 321468
rect 460565 321466 460631 321469
rect 444116 321464 460631 321466
rect 444116 321408 460570 321464
rect 460626 321408 460631 321464
rect 444116 321406 460631 321408
rect 444116 321404 444122 321406
rect 460565 321403 460631 321406
rect 447726 321268 447732 321332
rect 447796 321330 447802 321332
rect 460841 321330 460907 321333
rect 447796 321328 460907 321330
rect 447796 321272 460846 321328
rect 460902 321272 460907 321328
rect 447796 321270 460907 321272
rect 447796 321268 447802 321270
rect 460841 321267 460907 321270
rect 469121 321330 469187 321333
rect 530526 321330 530532 321332
rect 469121 321328 530532 321330
rect 469121 321272 469126 321328
rect 469182 321272 530532 321328
rect 469121 321270 530532 321272
rect 469121 321267 469187 321270
rect 530526 321268 530532 321270
rect 530596 321268 530602 321332
rect 442717 321194 442783 321197
rect 481817 321194 481883 321197
rect 442717 321192 481883 321194
rect 442717 321136 442722 321192
rect 442778 321136 481822 321192
rect 481878 321136 481883 321192
rect 442717 321134 481883 321136
rect 442717 321131 442783 321134
rect 481817 321131 481883 321134
rect 449566 320996 449572 321060
rect 449636 321058 449642 321060
rect 480989 321058 481055 321061
rect 449636 321056 481055 321058
rect 449636 321000 480994 321056
rect 481050 321000 481055 321056
rect 449636 320998 481055 321000
rect 449636 320996 449642 320998
rect 480989 320995 481055 320998
rect 460790 320724 460796 320788
rect 460860 320786 460866 320788
rect 509693 320786 509759 320789
rect 460860 320784 509759 320786
rect 460860 320728 509698 320784
rect 509754 320728 509759 320784
rect 460860 320726 509759 320728
rect 460860 320724 460866 320726
rect 509693 320723 509759 320726
rect 458633 320650 458699 320653
rect 558126 320650 558132 320652
rect 458633 320648 558132 320650
rect 458633 320592 458638 320648
rect 458694 320592 558132 320648
rect 458633 320590 558132 320592
rect 458633 320587 458699 320590
rect 558126 320588 558132 320590
rect 558196 320588 558202 320652
rect 507577 320242 507643 320245
rect 514334 320242 514340 320244
rect 507577 320240 514340 320242
rect 507577 320184 507582 320240
rect 507638 320184 514340 320240
rect 507577 320182 514340 320184
rect 507577 320179 507643 320182
rect 514334 320180 514340 320182
rect 514404 320180 514410 320244
rect 442441 320106 442507 320109
rect 481541 320106 481607 320109
rect 442441 320104 481607 320106
rect 442441 320048 442446 320104
rect 442502 320048 481546 320104
rect 481602 320048 481607 320104
rect 442441 320046 481607 320048
rect 442441 320043 442507 320046
rect 481541 320043 481607 320046
rect 446254 319908 446260 319972
rect 446324 319970 446330 319972
rect 471329 319970 471395 319973
rect 446324 319968 471395 319970
rect 446324 319912 471334 319968
rect 471390 319912 471395 319968
rect 446324 319910 471395 319912
rect 446324 319908 446330 319910
rect 471329 319907 471395 319910
rect 444230 319772 444236 319836
rect 444300 319834 444306 319836
rect 459737 319834 459803 319837
rect 444300 319832 459803 319834
rect 444300 319776 459742 319832
rect 459798 319776 459803 319832
rect 444300 319774 459803 319776
rect 444300 319772 444306 319774
rect 459737 319771 459803 319774
rect -960 319290 480 319380
rect 3969 319290 4035 319293
rect -960 319288 4035 319290
rect -960 319232 3974 319288
rect 4030 319232 4035 319288
rect -960 319230 4035 319232
rect -960 319140 480 319230
rect 3969 319227 4035 319230
rect 460565 318338 460631 318341
rect 511206 318338 511212 318340
rect 460565 318336 511212 318338
rect 460565 318280 460570 318336
rect 460626 318280 511212 318336
rect 460565 318278 511212 318280
rect 460565 318275 460631 318278
rect 511206 318276 511212 318278
rect 511276 318276 511282 318340
rect 432689 318202 432755 318205
rect 429916 318200 432755 318202
rect 429916 318144 432694 318200
rect 432750 318144 432755 318200
rect 429916 318142 432755 318144
rect 432689 318139 432755 318142
rect 459461 318202 459527 318205
rect 510153 318202 510219 318205
rect 459461 318200 510219 318202
rect 459461 318144 459466 318200
rect 459522 318144 510158 318200
rect 510214 318144 510219 318200
rect 459461 318142 510219 318144
rect 459461 318139 459527 318142
rect 510153 318139 510219 318142
rect 456057 318066 456123 318069
rect 518934 318066 518940 318068
rect 456057 318064 518940 318066
rect 456057 318008 456062 318064
rect 456118 318008 518940 318064
rect 456057 318006 518940 318008
rect 456057 318003 456123 318006
rect 518934 318004 518940 318006
rect 519004 318004 519010 318068
rect 509182 316644 509188 316708
rect 509252 316706 509258 316708
rect 510286 316706 510292 316708
rect 509252 316646 510292 316706
rect 509252 316644 509258 316646
rect 510286 316644 510292 316646
rect 510356 316644 510362 316708
rect 361757 315482 361823 315485
rect 359812 315480 361823 315482
rect 359812 315424 361762 315480
rect 361818 315424 361823 315480
rect 359812 315422 361823 315424
rect 361757 315419 361823 315422
rect 501137 315346 501203 315349
rect 538438 315346 538444 315348
rect 501137 315344 538444 315346
rect 501137 315288 501142 315344
rect 501198 315288 538444 315344
rect 501137 315286 538444 315288
rect 501137 315283 501203 315286
rect 538438 315284 538444 315286
rect 538508 315284 538514 315348
rect 432597 314530 432663 314533
rect 429916 314528 432663 314530
rect 429916 314472 432602 314528
rect 432658 314472 432663 314528
rect 429916 314470 432663 314472
rect 432597 314467 432663 314470
rect 501689 313986 501755 313989
rect 538254 313986 538260 313988
rect 501689 313984 538260 313986
rect 501689 313928 501694 313984
rect 501750 313928 538260 313984
rect 501689 313926 538260 313928
rect 501689 313923 501755 313926
rect 538254 313924 538260 313926
rect 538324 313924 538330 313988
rect 580165 312082 580231 312085
rect 583520 312082 584960 312172
rect 580165 312080 584960 312082
rect 580165 312024 580170 312080
rect 580226 312024 584960 312080
rect 580165 312022 584960 312024
rect 580165 312019 580231 312022
rect 583520 311932 584960 312022
rect 432045 310858 432111 310861
rect 429916 310856 432111 310858
rect 429916 310800 432050 310856
rect 432106 310800 432111 310856
rect 429916 310798 432111 310800
rect 432045 310795 432111 310798
rect 432689 307186 432755 307189
rect 429916 307184 432755 307186
rect 429916 307128 432694 307184
rect 432750 307128 432755 307184
rect 429916 307126 432755 307128
rect 432689 307123 432755 307126
rect -960 306234 480 306324
rect 3601 306234 3667 306237
rect -960 306232 3667 306234
rect -960 306176 3606 306232
rect 3662 306176 3667 306232
rect -960 306174 3667 306176
rect -960 306084 480 306174
rect 3601 306171 3667 306174
rect 381537 306098 381603 306101
rect 508998 306098 509004 306100
rect 381537 306096 509004 306098
rect 381537 306040 381542 306096
rect 381598 306040 509004 306096
rect 381537 306038 509004 306040
rect 381537 306035 381603 306038
rect 508998 306036 509004 306038
rect 509068 306036 509074 306100
rect 381721 305962 381787 305965
rect 511022 305962 511028 305964
rect 381721 305960 511028 305962
rect 381721 305904 381726 305960
rect 381782 305904 511028 305960
rect 381721 305902 511028 305904
rect 381721 305899 381787 305902
rect 511022 305900 511028 305902
rect 511092 305900 511098 305964
rect 367829 305826 367895 305829
rect 517881 305826 517947 305829
rect 367829 305824 517947 305826
rect 367829 305768 367834 305824
rect 367890 305768 517886 305824
rect 517942 305768 517947 305824
rect 367829 305766 517947 305768
rect 367829 305763 367895 305766
rect 517881 305763 517947 305766
rect 360837 305690 360903 305693
rect 512085 305690 512151 305693
rect 360837 305688 512151 305690
rect 360837 305632 360842 305688
rect 360898 305632 512090 305688
rect 512146 305632 512151 305688
rect 360837 305630 512151 305632
rect 360837 305627 360903 305630
rect 512085 305627 512151 305630
rect 361757 304466 361823 304469
rect 359812 304464 361823 304466
rect 359812 304408 361762 304464
rect 361818 304408 361823 304464
rect 359812 304406 361823 304408
rect 361757 304403 361823 304406
rect 381445 303106 381511 303109
rect 510838 303106 510844 303108
rect 381445 303104 510844 303106
rect 381445 303048 381450 303104
rect 381506 303048 510844 303104
rect 381445 303046 510844 303048
rect 381445 303043 381511 303046
rect 510838 303044 510844 303046
rect 510908 303044 510914 303108
rect 363689 302970 363755 302973
rect 512545 302970 512611 302973
rect 363689 302968 512611 302970
rect 363689 302912 363694 302968
rect 363750 302912 512550 302968
rect 512606 302912 512611 302968
rect 363689 302910 512611 302912
rect 363689 302907 363755 302910
rect 512545 302907 512611 302910
rect 362217 302834 362283 302837
rect 512821 302834 512887 302837
rect 362217 302832 512887 302834
rect 362217 302776 362222 302832
rect 362278 302776 512826 302832
rect 512882 302776 512887 302832
rect 362217 302774 512887 302776
rect 362217 302771 362283 302774
rect 512821 302771 512887 302774
rect 580165 298754 580231 298757
rect 583520 298754 584960 298844
rect 580165 298752 584960 298754
rect 580165 298696 580170 298752
rect 580226 298696 584960 298752
rect 580165 298694 584960 298696
rect 580165 298691 580231 298694
rect 583520 298604 584960 298694
rect 365161 297666 365227 297669
rect 510654 297666 510660 297668
rect 365161 297664 510660 297666
rect 365161 297608 365166 297664
rect 365222 297608 510660 297664
rect 365161 297606 510660 297608
rect 365161 297603 365227 297606
rect 510654 297604 510660 297606
rect 510724 297604 510730 297668
rect 368197 297530 368263 297533
rect 514150 297530 514156 297532
rect 368197 297528 514156 297530
rect 368197 297472 368202 297528
rect 368258 297472 514156 297528
rect 368197 297470 514156 297472
rect 368197 297467 368263 297470
rect 514150 297468 514156 297470
rect 514220 297468 514226 297532
rect 363781 297394 363847 297397
rect 514886 297394 514892 297396
rect 363781 297392 514892 297394
rect 363781 297336 363786 297392
rect 363842 297336 514892 297392
rect 363781 297334 514892 297336
rect 363781 297331 363847 297334
rect 514886 297332 514892 297334
rect 514956 297332 514962 297396
rect 361757 293450 361823 293453
rect 359812 293448 361823 293450
rect 359812 293392 361762 293448
rect 361818 293392 361823 293448
rect 359812 293390 361823 293392
rect 361757 293387 361823 293390
rect -960 293178 480 293268
rect 3693 293178 3759 293181
rect -960 293176 3759 293178
rect -960 293120 3698 293176
rect 3754 293120 3759 293176
rect -960 293118 3759 293120
rect -960 293028 480 293118
rect 3693 293115 3759 293118
rect 384849 291818 384915 291821
rect 514702 291818 514708 291820
rect 384849 291816 514708 291818
rect 384849 291760 384854 291816
rect 384910 291760 514708 291816
rect 384849 291758 514708 291760
rect 384849 291755 384915 291758
rect 514702 291756 514708 291758
rect 514772 291756 514778 291820
rect 374729 286378 374795 286381
rect 517830 286378 517836 286380
rect 374729 286376 517836 286378
rect 374729 286320 374734 286376
rect 374790 286320 517836 286376
rect 374729 286318 517836 286320
rect 374729 286315 374795 286318
rect 517830 286316 517836 286318
rect 517900 286316 517906 286380
rect 583520 285276 584960 285516
rect 361757 282434 361823 282437
rect 359812 282432 361823 282434
rect 359812 282376 361762 282432
rect 361818 282376 361823 282432
rect 359812 282374 361823 282376
rect 361757 282371 361823 282374
rect -960 279972 480 280212
rect 580257 272234 580323 272237
rect 583520 272234 584960 272324
rect 580257 272232 584960 272234
rect 580257 272176 580262 272232
rect 580318 272176 584960 272232
rect 580257 272174 584960 272176
rect 580257 272171 580323 272174
rect 583520 272084 584960 272174
rect 361757 271418 361823 271421
rect 359812 271416 361823 271418
rect 359812 271360 361762 271416
rect 361818 271360 361823 271416
rect 359812 271358 361823 271360
rect 361757 271355 361823 271358
rect -960 267202 480 267292
rect 3417 267202 3483 267205
rect -960 267200 3483 267202
rect -960 267144 3422 267200
rect 3478 267144 3483 267200
rect -960 267142 3483 267144
rect -960 267052 480 267142
rect 3417 267139 3483 267142
rect 456793 262714 456859 262717
rect 456793 262712 460092 262714
rect 456793 262656 456798 262712
rect 456854 262656 460092 262712
rect 456793 262654 460092 262656
rect 456793 262651 456859 262654
rect 531313 261082 531379 261085
rect 529828 261080 531379 261082
rect 529828 261024 531318 261080
rect 531374 261024 531379 261080
rect 529828 261022 531379 261024
rect 531313 261019 531379 261022
rect 361757 260402 361823 260405
rect 359812 260400 361823 260402
rect 359812 260344 361762 260400
rect 361818 260344 361823 260400
rect 359812 260342 361823 260344
rect 361757 260339 361823 260342
rect 580349 258906 580415 258909
rect 583520 258906 584960 258996
rect 580349 258904 584960 258906
rect 580349 258848 580354 258904
rect 580410 258848 584960 258904
rect 580349 258846 584960 258848
rect 580349 258843 580415 258846
rect 583520 258756 584960 258846
rect -960 254146 480 254236
rect 3509 254146 3575 254149
rect -960 254144 3575 254146
rect -960 254088 3514 254144
rect 3570 254088 3575 254144
rect -960 254086 3575 254088
rect -960 253996 480 254086
rect 3509 254083 3575 254086
rect 361757 249386 361823 249389
rect 359812 249384 361823 249386
rect 359812 249328 361762 249384
rect 361818 249328 361823 249384
rect 359812 249326 361823 249328
rect 361757 249323 361823 249326
rect 456793 248842 456859 248845
rect 456793 248840 460092 248842
rect 456793 248784 456798 248840
rect 456854 248784 460092 248840
rect 456793 248782 460092 248784
rect 456793 248779 456859 248782
rect 580165 245578 580231 245581
rect 583520 245578 584960 245668
rect 580165 245576 584960 245578
rect 580165 245520 580170 245576
rect 580226 245520 584960 245576
rect 580165 245518 584960 245520
rect 580165 245515 580231 245518
rect 583520 245428 584960 245518
rect 531313 243674 531379 243677
rect 529828 243672 531379 243674
rect 529828 243616 531318 243672
rect 531374 243616 531379 243672
rect 529828 243614 531379 243616
rect 531313 243611 531379 243614
rect -960 241090 480 241180
rect 3785 241090 3851 241093
rect -960 241088 3851 241090
rect -960 241032 3790 241088
rect 3846 241032 3851 241088
rect -960 241030 3851 241032
rect -960 240940 480 241030
rect 3785 241027 3851 241030
rect 361757 238370 361823 238373
rect 359812 238368 361823 238370
rect 359812 238312 361762 238368
rect 361818 238312 361823 238368
rect 359812 238310 361823 238312
rect 361757 238307 361823 238310
rect 457989 234970 458055 234973
rect 457989 234968 460092 234970
rect 457989 234912 457994 234968
rect 458050 234912 460092 234968
rect 457989 234910 460092 234912
rect 457989 234907 458055 234910
rect 580165 232386 580231 232389
rect 583520 232386 584960 232476
rect 580165 232384 584960 232386
rect 580165 232328 580170 232384
rect 580226 232328 584960 232384
rect 580165 232326 584960 232328
rect 580165 232323 580231 232326
rect 583520 232236 584960 232326
rect -960 227884 480 228124
rect 361757 227354 361823 227357
rect 359812 227352 361823 227354
rect 359812 227296 361762 227352
rect 361818 227296 361823 227352
rect 359812 227294 361823 227296
rect 361757 227291 361823 227294
rect 530117 226266 530183 226269
rect 529828 226264 530183 226266
rect 529828 226208 530122 226264
rect 530178 226208 530183 226264
rect 529828 226206 530183 226208
rect 530117 226203 530183 226206
rect 457805 221098 457871 221101
rect 457805 221096 460092 221098
rect 457805 221040 457810 221096
rect 457866 221040 460092 221096
rect 457805 221038 460092 221040
rect 457805 221035 457871 221038
rect 580257 219058 580323 219061
rect 583520 219058 584960 219148
rect 580257 219056 584960 219058
rect 580257 219000 580262 219056
rect 580318 219000 584960 219056
rect 580257 218998 584960 219000
rect 580257 218995 580323 218998
rect 583520 218908 584960 218998
rect 361665 216338 361731 216341
rect 359812 216336 361731 216338
rect 359812 216280 361670 216336
rect 361726 216280 361731 216336
rect 359812 216278 361731 216280
rect 361665 216275 361731 216278
rect -960 214978 480 215068
rect 3877 214978 3943 214981
rect -960 214976 3943 214978
rect -960 214920 3882 214976
rect 3938 214920 3943 214976
rect -960 214918 3943 214920
rect -960 214828 480 214918
rect 3877 214915 3943 214918
rect 529933 209266 529999 209269
rect 529798 209264 529999 209266
rect 529798 209208 529938 209264
rect 529994 209208 529999 209264
rect 529798 209206 529999 209208
rect 529798 208828 529858 209206
rect 529933 209203 529999 209206
rect 459553 207226 459619 207229
rect 459553 207224 460092 207226
rect 459553 207168 459558 207224
rect 459614 207168 460092 207224
rect 459553 207166 460092 207168
rect 459553 207163 459619 207166
rect 579797 205730 579863 205733
rect 583520 205730 584960 205820
rect 579797 205728 584960 205730
rect 579797 205672 579802 205728
rect 579858 205672 584960 205728
rect 579797 205670 584960 205672
rect 579797 205667 579863 205670
rect 583520 205580 584960 205670
rect 361757 205322 361823 205325
rect 359812 205320 361823 205322
rect 359812 205264 361762 205320
rect 361818 205264 361823 205320
rect 359812 205262 361823 205264
rect 361757 205259 361823 205262
rect -960 201922 480 202012
rect 3969 201922 4035 201925
rect -960 201920 4035 201922
rect -960 201864 3974 201920
rect 4030 201864 4035 201920
rect -960 201862 4035 201864
rect -960 201772 480 201862
rect 3969 201859 4035 201862
rect 361757 194306 361823 194309
rect 359812 194304 361823 194306
rect 359812 194248 361762 194304
rect 361818 194248 361823 194304
rect 359812 194246 361823 194248
rect 361757 194243 361823 194246
rect 580165 192538 580231 192541
rect 583520 192538 584960 192628
rect 580165 192536 584960 192538
rect 580165 192480 580170 192536
rect 580226 192480 584960 192536
rect 580165 192478 584960 192480
rect 580165 192475 580231 192478
rect 583520 192388 584960 192478
rect -960 188866 480 188956
rect 4061 188866 4127 188869
rect -960 188864 4127 188866
rect -960 188808 4066 188864
rect 4122 188808 4127 188864
rect -960 188806 4127 188808
rect -960 188716 480 188806
rect 4061 188803 4127 188806
rect 361757 183290 361823 183293
rect 359812 183288 361823 183290
rect 359812 183232 361762 183288
rect 361818 183232 361823 183288
rect 359812 183230 361823 183232
rect 361757 183227 361823 183230
rect 580165 179210 580231 179213
rect 583520 179210 584960 179300
rect 580165 179208 584960 179210
rect 580165 179152 580170 179208
rect 580226 179152 584960 179208
rect 580165 179150 584960 179152
rect 580165 179147 580231 179150
rect 583520 179060 584960 179150
rect -960 175796 480 176036
rect 361757 172274 361823 172277
rect 359812 172272 361823 172274
rect 359812 172216 361762 172272
rect 361818 172216 361823 172272
rect 359812 172214 361823 172216
rect 361757 172211 361823 172214
rect 580165 165882 580231 165885
rect 583520 165882 584960 165972
rect 580165 165880 584960 165882
rect 580165 165824 580170 165880
rect 580226 165824 584960 165880
rect 580165 165822 584960 165824
rect 580165 165819 580231 165822
rect 583520 165732 584960 165822
rect -960 162890 480 162980
rect 3325 162890 3391 162893
rect -960 162888 3391 162890
rect -960 162832 3330 162888
rect 3386 162832 3391 162888
rect -960 162830 3391 162832
rect -960 162740 480 162830
rect 3325 162827 3391 162830
rect 421414 162692 421420 162756
rect 421484 162754 421490 162756
rect 421833 162754 421899 162757
rect 425881 162756 425947 162757
rect 425830 162754 425836 162756
rect 421484 162752 421899 162754
rect 421484 162696 421838 162752
rect 421894 162696 421899 162752
rect 421484 162694 421899 162696
rect 425790 162694 425836 162754
rect 425900 162752 425947 162756
rect 425942 162696 425947 162752
rect 421484 162692 421490 162694
rect 421833 162691 421899 162694
rect 425830 162692 425836 162694
rect 425900 162692 425947 162696
rect 428406 162692 428412 162756
rect 428476 162754 428482 162756
rect 428641 162754 428707 162757
rect 428476 162752 428707 162754
rect 428476 162696 428646 162752
rect 428702 162696 428707 162752
rect 428476 162694 428707 162696
rect 428476 162692 428482 162694
rect 425881 162691 425947 162692
rect 428641 162691 428707 162694
rect 361757 161258 361823 161261
rect 359812 161256 361823 161258
rect 359812 161200 361762 161256
rect 361818 161200 361823 161256
rect 359812 161198 361823 161200
rect 361757 161195 361823 161198
rect 451733 158266 451799 158269
rect 449788 158264 451799 158266
rect 449788 158208 451738 158264
rect 451794 158208 451799 158264
rect 449788 158206 451799 158208
rect 451733 158203 451799 158206
rect 451733 156906 451799 156909
rect 449788 156904 451799 156906
rect 449788 156848 451738 156904
rect 451794 156848 451799 156904
rect 449788 156846 451799 156848
rect 451733 156843 451799 156846
rect 452193 155546 452259 155549
rect 449788 155544 452259 155546
rect 449788 155488 452198 155544
rect 452254 155488 452259 155544
rect 449788 155486 452259 155488
rect 452193 155483 452259 155486
rect 452469 154186 452535 154189
rect 449788 154184 452535 154186
rect 449788 154128 452474 154184
rect 452530 154128 452535 154184
rect 449788 154126 452535 154128
rect 452469 154123 452535 154126
rect 452469 152826 452535 152829
rect 449788 152824 452535 152826
rect 449788 152768 452474 152824
rect 452530 152768 452535 152824
rect 449788 152766 452535 152768
rect 452469 152763 452535 152766
rect 580165 152690 580231 152693
rect 583520 152690 584960 152780
rect 580165 152688 584960 152690
rect 580165 152632 580170 152688
rect 580226 152632 584960 152688
rect 580165 152630 584960 152632
rect 580165 152627 580231 152630
rect 583520 152540 584960 152630
rect 452561 151466 452627 151469
rect 449788 151464 452627 151466
rect 449788 151408 452566 151464
rect 452622 151408 452627 151464
rect 449788 151406 452627 151408
rect 452561 151403 452627 151406
rect 361757 150242 361823 150245
rect 359812 150240 361823 150242
rect 359812 150184 361762 150240
rect 361818 150184 361823 150240
rect 359812 150182 361823 150184
rect 361757 150179 361823 150182
rect 452377 150106 452443 150109
rect 449788 150104 452443 150106
rect 449788 150048 452382 150104
rect 452438 150048 452443 150104
rect 449788 150046 452443 150048
rect 452377 150043 452443 150046
rect -960 149834 480 149924
rect 3233 149834 3299 149837
rect -960 149832 3299 149834
rect -960 149776 3238 149832
rect 3294 149776 3299 149832
rect -960 149774 3299 149776
rect -960 149684 480 149774
rect 3233 149771 3299 149774
rect 452009 148746 452075 148749
rect 449788 148744 452075 148746
rect 449788 148688 452014 148744
rect 452070 148688 452075 148744
rect 449788 148686 452075 148688
rect 452009 148683 452075 148686
rect 452561 147386 452627 147389
rect 449788 147384 452627 147386
rect 449788 147328 452566 147384
rect 452622 147328 452627 147384
rect 449788 147326 452627 147328
rect 452561 147323 452627 147326
rect 451825 146026 451891 146029
rect 449788 146024 451891 146026
rect 449788 145968 451830 146024
rect 451886 145968 451891 146024
rect 449788 145966 451891 145968
rect 451825 145963 451891 145966
rect 451549 144666 451615 144669
rect 449788 144664 451615 144666
rect 449788 144608 451554 144664
rect 451610 144608 451615 144664
rect 449788 144606 451615 144608
rect 451549 144603 451615 144606
rect 452561 143306 452627 143309
rect 449788 143304 452627 143306
rect 449788 143248 452566 143304
rect 452622 143248 452627 143304
rect 449788 143246 452627 143248
rect 452561 143243 452627 143246
rect 452561 141946 452627 141949
rect 449788 141944 452627 141946
rect 449788 141888 452566 141944
rect 452622 141888 452627 141944
rect 449788 141886 452627 141888
rect 452561 141883 452627 141886
rect 452561 140586 452627 140589
rect 449788 140584 452627 140586
rect 449788 140528 452566 140584
rect 452622 140528 452627 140584
rect 449788 140526 452627 140528
rect 452561 140523 452627 140526
rect 580165 139362 580231 139365
rect 583520 139362 584960 139452
rect 580165 139360 584960 139362
rect 580165 139304 580170 139360
rect 580226 139304 584960 139360
rect 580165 139302 584960 139304
rect 580165 139299 580231 139302
rect 361757 139226 361823 139229
rect 451549 139226 451615 139229
rect 359812 139224 361823 139226
rect 359812 139168 361762 139224
rect 361818 139168 361823 139224
rect 359812 139166 361823 139168
rect 449788 139224 451615 139226
rect 449788 139168 451554 139224
rect 451610 139168 451615 139224
rect 583520 139212 584960 139302
rect 449788 139166 451615 139168
rect 361757 139163 361823 139166
rect 451549 139163 451615 139166
rect 538949 138002 539015 138005
rect 538949 138000 539610 138002
rect 538949 137944 538954 138000
rect 539010 137944 539610 138000
rect 538949 137942 539610 137944
rect 538949 137939 539015 137942
rect 452561 137866 452627 137869
rect 449788 137864 452627 137866
rect 449788 137808 452566 137864
rect 452622 137808 452627 137864
rect 449788 137806 452627 137808
rect 452561 137803 452627 137806
rect 538438 137804 538444 137868
rect 538508 137866 538514 137868
rect 539409 137866 539475 137869
rect 538508 137864 539475 137866
rect 538508 137808 539414 137864
rect 539470 137808 539475 137864
rect 538508 137806 539475 137808
rect 538508 137804 538514 137806
rect 539409 137803 539475 137806
rect 539550 137428 539610 137942
rect -960 136778 480 136868
rect 2814 136778 2820 136780
rect -960 136718 2820 136778
rect -960 136628 480 136718
rect 2814 136716 2820 136718
rect 2884 136716 2890 136780
rect 451549 136506 451615 136509
rect 449788 136504 451615 136506
rect 449788 136448 451554 136504
rect 451610 136448 451615 136504
rect 449788 136446 451615 136448
rect 451549 136443 451615 136446
rect 539501 135962 539567 135965
rect 539501 135960 539610 135962
rect 539501 135904 539506 135960
rect 539562 135904 539610 135960
rect 539501 135899 539610 135904
rect 539550 135388 539610 135899
rect 452009 135146 452075 135149
rect 449788 135144 452075 135146
rect 449788 135088 452014 135144
rect 452070 135088 452075 135144
rect 449788 135086 452075 135088
rect 452009 135083 452075 135086
rect 452285 133786 452351 133789
rect 449788 133784 452351 133786
rect 449788 133728 452290 133784
rect 452346 133728 452351 133784
rect 449788 133726 452351 133728
rect 452285 133723 452351 133726
rect 539358 133316 539364 133380
rect 539428 133316 539434 133380
rect 452285 132426 452351 132429
rect 449788 132424 452351 132426
rect 449788 132368 452290 132424
rect 452346 132368 452351 132424
rect 449788 132366 452351 132368
rect 452285 132363 452351 132366
rect 540237 131338 540303 131341
rect 539948 131336 540303 131338
rect 539948 131280 540242 131336
rect 540298 131280 540303 131336
rect 539948 131278 540303 131280
rect 540237 131275 540303 131278
rect 452561 131066 452627 131069
rect 449788 131064 452627 131066
rect 449788 131008 452566 131064
rect 452622 131008 452627 131064
rect 449788 131006 452627 131008
rect 452561 131003 452627 131006
rect 452101 129706 452167 129709
rect 449788 129704 452167 129706
rect 449788 129648 452106 129704
rect 452162 129648 452167 129704
rect 449788 129646 452167 129648
rect 452101 129643 452167 129646
rect 539409 129706 539475 129709
rect 539409 129704 539610 129706
rect 539409 129648 539414 129704
rect 539470 129648 539610 129704
rect 539409 129646 539610 129648
rect 539409 129643 539475 129646
rect 539550 129268 539610 129646
rect 451917 128346 451983 128349
rect 449788 128344 451983 128346
rect 449788 128288 451922 128344
rect 451978 128288 451983 128344
rect 449788 128286 451983 128288
rect 451917 128283 451983 128286
rect 361757 128210 361823 128213
rect 359812 128208 361823 128210
rect 359812 128152 361762 128208
rect 361818 128152 361823 128208
rect 359812 128150 361823 128152
rect 361757 128147 361823 128150
rect 540145 127258 540211 127261
rect 539948 127256 540211 127258
rect 539948 127200 540150 127256
rect 540206 127200 540211 127256
rect 539948 127198 540211 127200
rect 540145 127195 540211 127198
rect 452561 126986 452627 126989
rect 449788 126984 452627 126986
rect 449788 126928 452566 126984
rect 452622 126928 452627 126984
rect 449788 126926 452627 126928
rect 452561 126923 452627 126926
rect 580165 126034 580231 126037
rect 583520 126034 584960 126124
rect 580165 126032 584960 126034
rect 580165 125976 580170 126032
rect 580226 125976 584960 126032
rect 580165 125974 584960 125976
rect 580165 125971 580231 125974
rect 583520 125884 584960 125974
rect 451733 125626 451799 125629
rect 449788 125624 451799 125626
rect 449788 125568 451738 125624
rect 451794 125568 451799 125624
rect 449788 125566 451799 125568
rect 451733 125563 451799 125566
rect 540329 125218 540395 125221
rect 539948 125216 540395 125218
rect 539948 125160 540334 125216
rect 540390 125160 540395 125216
rect 539948 125158 540395 125160
rect 540329 125155 540395 125158
rect 452009 124266 452075 124269
rect 449788 124264 452075 124266
rect 449788 124208 452014 124264
rect 452070 124208 452075 124264
rect 449788 124206 452075 124208
rect 452009 124203 452075 124206
rect -960 123572 480 123812
rect 542721 123178 542787 123181
rect 539948 123176 542787 123178
rect 539948 123120 542726 123176
rect 542782 123120 542787 123176
rect 539948 123118 542787 123120
rect 542721 123115 542787 123118
rect 451733 122906 451799 122909
rect 449788 122904 451799 122906
rect 449788 122848 451738 122904
rect 451794 122848 451799 122904
rect 449788 122846 451799 122848
rect 451733 122843 451799 122846
rect 451917 121546 451983 121549
rect 449788 121544 451983 121546
rect 449788 121488 451922 121544
rect 451978 121488 451983 121544
rect 449788 121486 451983 121488
rect 451917 121483 451983 121486
rect 542629 121138 542695 121141
rect 539948 121136 542695 121138
rect 539948 121080 542634 121136
rect 542690 121080 542695 121136
rect 539948 121078 542695 121080
rect 542629 121075 542695 121078
rect 543089 119098 543155 119101
rect 539948 119096 543155 119098
rect 539948 119040 543094 119096
rect 543150 119040 543155 119096
rect 539948 119038 543155 119040
rect 543089 119035 543155 119038
rect 539869 117330 539935 117333
rect 539869 117328 539978 117330
rect 539869 117272 539874 117328
rect 539930 117272 539978 117328
rect 539869 117267 539978 117272
rect 361757 117194 361823 117197
rect 359812 117192 361823 117194
rect 359812 117136 361762 117192
rect 361818 117136 361823 117192
rect 359812 117134 361823 117136
rect 361757 117131 361823 117134
rect 539918 117028 539978 117267
rect 541433 115018 541499 115021
rect 539948 115016 541499 115018
rect 539948 114960 541438 115016
rect 541494 114960 541499 115016
rect 539948 114958 541499 114960
rect 541433 114955 541499 114958
rect 539918 112842 539978 112948
rect 540053 112842 540119 112845
rect 539918 112840 540119 112842
rect 539918 112784 540058 112840
rect 540114 112784 540119 112840
rect 539918 112782 540119 112784
rect 540053 112779 540119 112782
rect 579797 112842 579863 112845
rect 583520 112842 584960 112932
rect 579797 112840 584960 112842
rect 579797 112784 579802 112840
rect 579858 112784 584960 112840
rect 579797 112782 584960 112784
rect 579797 112779 579863 112782
rect 583520 112692 584960 112782
rect 541065 110938 541131 110941
rect 539948 110936 541131 110938
rect 539948 110880 541070 110936
rect 541126 110880 541131 110936
rect 539948 110878 541131 110880
rect 541065 110875 541131 110878
rect -960 110666 480 110756
rect 3366 110666 3372 110668
rect -960 110606 3372 110666
rect -960 110516 480 110606
rect 3366 110604 3372 110606
rect 3436 110604 3442 110668
rect 539918 108765 539978 108868
rect 539918 108760 540027 108765
rect 539918 108704 539966 108760
rect 540022 108704 540027 108760
rect 539918 108702 540027 108704
rect 539961 108699 540027 108702
rect 541341 106858 541407 106861
rect 539948 106856 541407 106858
rect 539948 106800 541346 106856
rect 541402 106800 541407 106856
rect 539948 106798 541407 106800
rect 541341 106795 541407 106798
rect 361757 106178 361823 106181
rect 359812 106176 361823 106178
rect 359812 106120 361762 106176
rect 361818 106120 361823 106176
rect 359812 106118 361823 106120
rect 361757 106115 361823 106118
rect 541249 104818 541315 104821
rect 539948 104816 541315 104818
rect 539948 104760 541254 104816
rect 541310 104760 541315 104816
rect 539948 104758 541315 104760
rect 541249 104755 541315 104758
rect 541157 102778 541223 102781
rect 539948 102776 541223 102778
rect 539948 102720 541162 102776
rect 541218 102720 541223 102776
rect 539948 102718 541223 102720
rect 541157 102715 541223 102718
rect 542537 100738 542603 100741
rect 539948 100736 542603 100738
rect 539948 100680 542542 100736
rect 542598 100680 542603 100736
rect 539948 100678 542603 100680
rect 542537 100675 542603 100678
rect 580165 99514 580231 99517
rect 583520 99514 584960 99604
rect 580165 99512 584960 99514
rect 580165 99456 580170 99512
rect 580226 99456 584960 99512
rect 580165 99454 584960 99456
rect 580165 99451 580231 99454
rect 583520 99364 584960 99454
rect 539777 99242 539843 99245
rect 539734 99240 539843 99242
rect 539734 99184 539782 99240
rect 539838 99184 539843 99240
rect 539734 99179 539843 99184
rect 2814 98636 2820 98700
rect 2884 98698 2890 98700
rect 3049 98698 3115 98701
rect 2884 98696 3115 98698
rect 2884 98640 3054 98696
rect 3110 98640 3115 98696
rect 539734 98668 539794 99179
rect 2884 98638 3115 98640
rect 2884 98636 2890 98638
rect 3049 98635 3115 98638
rect -960 97610 480 97700
rect 3550 97610 3556 97612
rect -960 97550 3556 97610
rect -960 97460 480 97550
rect 3550 97548 3556 97550
rect 3620 97548 3626 97612
rect 539685 97202 539751 97205
rect 539685 97200 539794 97202
rect 539685 97144 539690 97200
rect 539746 97144 539794 97200
rect 539685 97139 539794 97144
rect 539734 96628 539794 97139
rect 361757 95162 361823 95165
rect 539593 95162 539659 95165
rect 359812 95160 361823 95162
rect 359812 95104 361762 95160
rect 361818 95104 361823 95160
rect 359812 95102 361823 95104
rect 361757 95099 361823 95102
rect 539550 95160 539659 95162
rect 539550 95104 539598 95160
rect 539654 95104 539659 95160
rect 539550 95099 539659 95104
rect 539550 94588 539610 95099
rect 542997 92578 543063 92581
rect 539948 92576 543063 92578
rect 539948 92520 543002 92576
rect 543058 92520 543063 92576
rect 539948 92518 543063 92520
rect 542997 92515 543063 92518
rect 542445 90538 542511 90541
rect 539948 90536 542511 90538
rect 539948 90480 542450 90536
rect 542506 90480 542511 90536
rect 539948 90478 542511 90480
rect 542445 90475 542511 90478
rect 543181 88498 543247 88501
rect 539948 88496 543247 88498
rect 539948 88440 543186 88496
rect 543242 88440 543247 88496
rect 539948 88438 543247 88440
rect 543181 88435 543247 88438
rect 542905 86458 542971 86461
rect 539948 86456 542971 86458
rect 539948 86400 542910 86456
rect 542966 86400 542971 86456
rect 539948 86398 542971 86400
rect 542905 86395 542971 86398
rect 580165 86186 580231 86189
rect 583520 86186 584960 86276
rect 580165 86184 584960 86186
rect 580165 86128 580170 86184
rect 580226 86128 584960 86184
rect 580165 86126 584960 86128
rect 580165 86123 580231 86126
rect 583520 86036 584960 86126
rect -960 84690 480 84780
rect 3693 84690 3759 84693
rect -960 84688 3759 84690
rect -960 84632 3698 84688
rect 3754 84632 3759 84688
rect -960 84630 3759 84632
rect -960 84540 480 84630
rect 3693 84627 3759 84630
rect 542813 84418 542879 84421
rect 539948 84416 542879 84418
rect 539948 84360 542818 84416
rect 542874 84360 542879 84416
rect 539948 84358 542879 84360
rect 542813 84355 542879 84358
rect 361757 84146 361823 84149
rect 359812 84144 361823 84146
rect 359812 84088 361762 84144
rect 361818 84088 361823 84144
rect 359812 84086 361823 84088
rect 361757 84083 361823 84086
rect 540973 82378 541039 82381
rect 539948 82376 541039 82378
rect 539948 82320 540978 82376
rect 541034 82320 541039 82376
rect 539948 82318 541039 82320
rect 540973 82315 541039 82318
rect 20897 73674 20963 73677
rect 21449 73674 21515 73677
rect 20897 73672 21515 73674
rect 20897 73616 20902 73672
rect 20958 73616 21454 73672
rect 21510 73616 21515 73672
rect 20897 73614 21515 73616
rect 20897 73611 20963 73614
rect 21449 73611 21515 73614
rect 361757 73130 361823 73133
rect 359812 73128 361823 73130
rect 359812 73072 361762 73128
rect 361818 73072 361823 73128
rect 359812 73070 361823 73072
rect 361757 73067 361823 73070
rect 580165 72994 580231 72997
rect 583520 72994 584960 73084
rect 580165 72992 584960 72994
rect 580165 72936 580170 72992
rect 580226 72936 584960 72992
rect 580165 72934 584960 72936
rect 580165 72931 580231 72934
rect 583520 72844 584960 72934
rect -960 71634 480 71724
rect 3601 71634 3667 71637
rect -960 71632 3667 71634
rect -960 71576 3606 71632
rect 3662 71576 3667 71632
rect -960 71574 3667 71576
rect -960 71484 480 71574
rect 3601 71571 3667 71574
rect 460289 67690 460355 67693
rect 460841 67690 460907 67693
rect 460289 67688 460907 67690
rect 460289 67632 460294 67688
rect 460350 67632 460846 67688
rect 460902 67632 460907 67688
rect 460289 67630 460907 67632
rect 460289 67627 460355 67630
rect 460798 67627 460907 67630
rect 460798 67524 460858 67627
rect 361757 62114 361823 62117
rect 359812 62112 361823 62114
rect 359812 62056 361762 62112
rect 361818 62056 361823 62112
rect 359812 62054 361823 62056
rect 361757 62051 361823 62054
rect 580165 59666 580231 59669
rect 583520 59666 584960 59756
rect 580165 59664 584960 59666
rect 580165 59608 580170 59664
rect 580226 59608 584960 59664
rect 580165 59606 584960 59608
rect 580165 59603 580231 59606
rect 583520 59516 584960 59606
rect -960 58578 480 58668
rect 3601 58578 3667 58581
rect -960 58576 3667 58578
rect -960 58520 3606 58576
rect 3662 58520 3667 58576
rect -960 58518 3667 58520
rect -960 58428 480 58518
rect 3601 58515 3667 58518
rect 361757 51098 361823 51101
rect 359812 51096 361823 51098
rect 359812 51040 361762 51096
rect 361818 51040 361823 51096
rect 359812 51038 361823 51040
rect 361757 51035 361823 51038
rect 19241 49602 19307 49605
rect 22134 49602 22140 49604
rect 19241 49600 22140 49602
rect 19241 49544 19246 49600
rect 19302 49544 22140 49600
rect 19241 49542 22140 49544
rect 19241 49539 19307 49542
rect 22134 49540 22140 49542
rect 22204 49540 22210 49604
rect 11697 48922 11763 48925
rect 22318 48922 22324 48924
rect 11697 48920 22324 48922
rect 11697 48864 11702 48920
rect 11758 48864 22324 48920
rect 11697 48862 22324 48864
rect 11697 48859 11763 48862
rect 22318 48860 22324 48862
rect 22388 48860 22394 48924
rect 540605 48922 540671 48925
rect 540605 48920 540714 48922
rect 540605 48864 540610 48920
rect 540666 48864 540714 48920
rect 540605 48859 540714 48864
rect 540654 48348 540714 48859
rect 3550 46820 3556 46884
rect 3620 46882 3626 46884
rect 384481 46882 384547 46885
rect 3620 46880 384547 46882
rect 3620 46824 384486 46880
rect 384542 46824 384547 46880
rect 3620 46822 384547 46824
rect 3620 46820 3626 46822
rect 384481 46819 384547 46822
rect 3366 46684 3372 46748
rect 3436 46746 3442 46748
rect 384297 46746 384363 46749
rect 3436 46744 384363 46746
rect 3436 46688 384302 46744
rect 384358 46688 384363 46744
rect 3436 46686 384363 46688
rect 3436 46684 3442 46686
rect 384297 46683 384363 46686
rect 22134 46548 22140 46612
rect 22204 46610 22210 46612
rect 361297 46610 361363 46613
rect 22204 46608 361363 46610
rect 22204 46552 361302 46608
rect 361358 46552 361363 46608
rect 22204 46550 361363 46552
rect 22204 46548 22210 46550
rect 361297 46547 361363 46550
rect 22318 46412 22324 46476
rect 22388 46474 22394 46476
rect 359549 46474 359615 46477
rect 22388 46472 359615 46474
rect 22388 46416 359554 46472
rect 359610 46416 359615 46472
rect 22388 46414 359615 46416
rect 22388 46412 22394 46414
rect 359549 46411 359615 46414
rect 580165 46338 580231 46341
rect 583520 46338 584960 46428
rect 580165 46336 584960 46338
rect 580165 46280 580170 46336
rect 580226 46280 584960 46336
rect 580165 46278 584960 46280
rect 580165 46275 580231 46278
rect 583520 46188 584960 46278
rect -960 45522 480 45612
rect 3417 45522 3483 45525
rect -960 45520 3483 45522
rect -960 45464 3422 45520
rect 3478 45464 3483 45520
rect -960 45462 3483 45464
rect -960 45372 480 45462
rect 3417 45459 3483 45462
rect 536833 41034 536899 41037
rect 536833 41032 540132 41034
rect 536833 40976 536838 41032
rect 536894 40976 540132 41032
rect 536833 40974 540132 40976
rect 536833 40971 536899 40974
rect 540421 34234 540487 34237
rect 540421 34232 540530 34234
rect 540421 34176 540426 34232
rect 540482 34176 540530 34232
rect 540421 34171 540530 34176
rect 540470 33660 540530 34171
rect 580165 33146 580231 33149
rect 583520 33146 584960 33236
rect 580165 33144 584960 33146
rect 580165 33088 580170 33144
rect 580226 33088 584960 33144
rect 580165 33086 584960 33088
rect 580165 33083 580231 33086
rect 583520 32996 584960 33086
rect -960 32466 480 32556
rect 2865 32466 2931 32469
rect -960 32464 2931 32466
rect -960 32408 2870 32464
rect 2926 32408 2931 32464
rect -960 32406 2931 32408
rect -960 32316 480 32406
rect 2865 32403 2931 32406
rect 579981 19818 580047 19821
rect 583520 19818 584960 19908
rect 579981 19816 584960 19818
rect 579981 19760 579986 19816
rect 580042 19760 584960 19816
rect 579981 19758 584960 19760
rect 579981 19755 580047 19758
rect 583520 19668 584960 19758
rect -960 19410 480 19500
rect 3417 19410 3483 19413
rect -960 19408 3483 19410
rect -960 19352 3422 19408
rect 3478 19352 3483 19408
rect -960 19350 3483 19352
rect -960 19260 480 19350
rect 3417 19347 3483 19350
rect 580165 6626 580231 6629
rect 583520 6626 584960 6716
rect 580165 6624 584960 6626
rect -960 6490 480 6580
rect 580165 6568 580170 6624
rect 580226 6568 584960 6624
rect 580165 6566 584960 6568
rect 580165 6563 580231 6566
rect 3417 6490 3483 6493
rect -960 6488 3483 6490
rect -960 6432 3422 6488
rect 3478 6432 3483 6488
rect 583520 6476 584960 6566
rect -960 6430 3483 6432
rect -960 6340 480 6430
rect 3417 6427 3483 6430
rect 8753 4042 8819 4045
rect 362217 4042 362283 4045
rect 8753 4040 362283 4042
rect 8753 3984 8758 4040
rect 8814 3984 362222 4040
rect 362278 3984 362283 4040
rect 8753 3982 362283 3984
rect 8753 3979 8819 3982
rect 362217 3979 362283 3982
rect 13537 3906 13603 3909
rect 374637 3906 374703 3909
rect 13537 3904 374703 3906
rect 13537 3848 13542 3904
rect 13598 3848 374642 3904
rect 374698 3848 374703 3904
rect 13537 3846 374703 3848
rect 13537 3843 13603 3846
rect 374637 3843 374703 3846
rect 9949 3770 10015 3773
rect 374821 3770 374887 3773
rect 9949 3768 374887 3770
rect 9949 3712 9954 3768
rect 10010 3712 374826 3768
rect 374882 3712 374887 3768
rect 9949 3710 374887 3712
rect 9949 3707 10015 3710
rect 374821 3707 374887 3710
rect 2865 3634 2931 3637
rect 381537 3634 381603 3637
rect 2865 3632 381603 3634
rect 2865 3576 2870 3632
rect 2926 3576 381542 3632
rect 381598 3576 381603 3632
rect 2865 3574 381603 3576
rect 2865 3571 2931 3574
rect 381537 3571 381603 3574
rect 1669 3498 1735 3501
rect 381721 3498 381787 3501
rect 1669 3496 381787 3498
rect 1669 3440 1674 3496
rect 1730 3440 381726 3496
rect 381782 3440 381787 3496
rect 1669 3438 381787 3440
rect 1669 3435 1735 3438
rect 381721 3435 381787 3438
rect 565 3362 631 3365
rect 460790 3362 460796 3364
rect 565 3360 460796 3362
rect 565 3304 570 3360
rect 626 3304 460796 3360
rect 565 3302 460796 3304
rect 565 3299 631 3302
rect 460790 3300 460796 3302
rect 460860 3300 460866 3364
rect 17033 3226 17099 3229
rect 365069 3226 365135 3229
rect 17033 3224 365135 3226
rect 17033 3168 17038 3224
rect 17094 3168 365074 3224
rect 365130 3168 365135 3224
rect 17033 3166 365135 3168
rect 17033 3163 17099 3166
rect 365069 3163 365135 3166
<< via3 >>
rect 447916 700572 447980 700636
rect 449572 700436 449636 700500
rect 447732 700300 447796 700364
rect 530532 700300 530596 700364
rect 527220 699816 527284 699820
rect 527220 699760 527234 699816
rect 527234 699760 527284 699816
rect 527220 699756 527284 699760
rect 558132 699756 558196 699820
rect 444236 689284 444300 689348
rect 446260 686428 446324 686492
rect 3740 683300 3804 683364
rect 3556 683164 3620 683228
rect 3372 682756 3436 682820
rect 3740 671196 3804 671260
rect 457852 665212 457916 665276
rect 458036 662492 458100 662556
rect 459508 655624 459572 655688
rect 3556 619108 3620 619172
rect 3372 606052 3436 606116
rect 474412 599524 474476 599588
rect 472020 598164 472084 598228
rect 457852 597620 457916 597684
rect 472204 595580 472268 595644
rect 459508 595444 459572 595508
rect 478828 595444 478892 595508
rect 476436 591228 476500 591292
rect 474780 589868 474844 589932
rect 458036 518060 458100 518124
rect 482692 517576 482756 517580
rect 482692 517520 482742 517576
rect 482742 517520 482756 517576
rect 482692 517516 482756 517520
rect 451044 516700 451108 516764
rect 450492 514320 450556 514384
rect 527220 502284 527284 502348
rect 489316 496844 489380 496908
rect 482692 462844 482756 462908
rect 444052 421908 444116 421972
rect 472204 389056 472268 389060
rect 472204 389000 472218 389056
rect 472218 389000 472268 389056
rect 472204 388996 472268 389000
rect 474412 389056 474476 389060
rect 474412 389000 474426 389056
rect 474426 389000 474476 389056
rect 474412 388996 474476 389000
rect 474780 388996 474844 389060
rect 476436 388996 476500 389060
rect 478828 388996 478892 389060
rect 472020 388860 472084 388924
rect 448284 388316 448348 388380
rect 489316 386956 489380 387020
rect 448284 349148 448348 349212
rect 511212 335684 511276 335748
rect 428412 334460 428476 334524
rect 425836 334324 425900 334388
rect 421420 334052 421484 334116
rect 510660 332964 510724 333028
rect 514708 331876 514772 331940
rect 514892 331332 514956 331396
rect 517836 330788 517900 330852
rect 515076 329156 515140 329220
rect 450676 328748 450740 328812
rect 514340 328612 514404 328676
rect 450492 328340 450556 328404
rect 510476 327524 510540 327588
rect 510844 326436 510908 326500
rect 518940 325756 519004 325820
rect 514156 324804 514220 324868
rect 510292 324260 510356 324324
rect 511028 323716 511092 323780
rect 447916 322356 447980 322420
rect 510476 321812 510540 321876
rect 515076 321676 515140 321740
rect 444052 321404 444116 321468
rect 447732 321268 447796 321332
rect 530532 321268 530596 321332
rect 449572 320996 449636 321060
rect 460796 320724 460860 320788
rect 558132 320588 558196 320652
rect 514340 320180 514404 320244
rect 446260 319908 446324 319972
rect 444236 319772 444300 319836
rect 511212 318276 511276 318340
rect 518940 318004 519004 318068
rect 509188 316644 509252 316708
rect 510292 316644 510356 316708
rect 538444 315284 538508 315348
rect 538260 313924 538324 313988
rect 509004 306036 509068 306100
rect 511028 305900 511092 305964
rect 510844 303044 510908 303108
rect 510660 297604 510724 297668
rect 514156 297468 514220 297532
rect 514892 297332 514956 297396
rect 514708 291756 514772 291820
rect 517836 286316 517900 286380
rect 421420 162692 421484 162756
rect 425836 162752 425900 162756
rect 425836 162696 425886 162752
rect 425886 162696 425900 162752
rect 425836 162692 425900 162696
rect 428412 162692 428476 162756
rect 538444 137804 538508 137868
rect 2820 136716 2884 136780
rect 539364 133316 539428 133380
rect 3372 110604 3436 110668
rect 2820 98636 2884 98700
rect 3556 97548 3620 97612
rect 22140 49540 22204 49604
rect 22324 48860 22388 48924
rect 3556 46820 3620 46884
rect 3372 46684 3436 46748
rect 22140 46548 22204 46612
rect 22324 46412 22388 46476
rect 460796 3300 460860 3364
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 677494 -8106 711002
rect -8726 677258 -8694 677494
rect -8458 677258 -8374 677494
rect -8138 677258 -8106 677494
rect -8726 677174 -8106 677258
rect -8726 676938 -8694 677174
rect -8458 676938 -8374 677174
rect -8138 676938 -8106 677174
rect -8726 641494 -8106 676938
rect -8726 641258 -8694 641494
rect -8458 641258 -8374 641494
rect -8138 641258 -8106 641494
rect -8726 641174 -8106 641258
rect -8726 640938 -8694 641174
rect -8458 640938 -8374 641174
rect -8138 640938 -8106 641174
rect -8726 605494 -8106 640938
rect -8726 605258 -8694 605494
rect -8458 605258 -8374 605494
rect -8138 605258 -8106 605494
rect -8726 605174 -8106 605258
rect -8726 604938 -8694 605174
rect -8458 604938 -8374 605174
rect -8138 604938 -8106 605174
rect -8726 569494 -8106 604938
rect -8726 569258 -8694 569494
rect -8458 569258 -8374 569494
rect -8138 569258 -8106 569494
rect -8726 569174 -8106 569258
rect -8726 568938 -8694 569174
rect -8458 568938 -8374 569174
rect -8138 568938 -8106 569174
rect -8726 533494 -8106 568938
rect -8726 533258 -8694 533494
rect -8458 533258 -8374 533494
rect -8138 533258 -8106 533494
rect -8726 533174 -8106 533258
rect -8726 532938 -8694 533174
rect -8458 532938 -8374 533174
rect -8138 532938 -8106 533174
rect -8726 497494 -8106 532938
rect -8726 497258 -8694 497494
rect -8458 497258 -8374 497494
rect -8138 497258 -8106 497494
rect -8726 497174 -8106 497258
rect -8726 496938 -8694 497174
rect -8458 496938 -8374 497174
rect -8138 496938 -8106 497174
rect -8726 461494 -8106 496938
rect -8726 461258 -8694 461494
rect -8458 461258 -8374 461494
rect -8138 461258 -8106 461494
rect -8726 461174 -8106 461258
rect -8726 460938 -8694 461174
rect -8458 460938 -8374 461174
rect -8138 460938 -8106 461174
rect -8726 425494 -8106 460938
rect -8726 425258 -8694 425494
rect -8458 425258 -8374 425494
rect -8138 425258 -8106 425494
rect -8726 425174 -8106 425258
rect -8726 424938 -8694 425174
rect -8458 424938 -8374 425174
rect -8138 424938 -8106 425174
rect -8726 389494 -8106 424938
rect -8726 389258 -8694 389494
rect -8458 389258 -8374 389494
rect -8138 389258 -8106 389494
rect -8726 389174 -8106 389258
rect -8726 388938 -8694 389174
rect -8458 388938 -8374 389174
rect -8138 388938 -8106 389174
rect -8726 353494 -8106 388938
rect -8726 353258 -8694 353494
rect -8458 353258 -8374 353494
rect -8138 353258 -8106 353494
rect -8726 353174 -8106 353258
rect -8726 352938 -8694 353174
rect -8458 352938 -8374 353174
rect -8138 352938 -8106 353174
rect -8726 317494 -8106 352938
rect -8726 317258 -8694 317494
rect -8458 317258 -8374 317494
rect -8138 317258 -8106 317494
rect -8726 317174 -8106 317258
rect -8726 316938 -8694 317174
rect -8458 316938 -8374 317174
rect -8138 316938 -8106 317174
rect -8726 281494 -8106 316938
rect -8726 281258 -8694 281494
rect -8458 281258 -8374 281494
rect -8138 281258 -8106 281494
rect -8726 281174 -8106 281258
rect -8726 280938 -8694 281174
rect -8458 280938 -8374 281174
rect -8138 280938 -8106 281174
rect -8726 245494 -8106 280938
rect -8726 245258 -8694 245494
rect -8458 245258 -8374 245494
rect -8138 245258 -8106 245494
rect -8726 245174 -8106 245258
rect -8726 244938 -8694 245174
rect -8458 244938 -8374 245174
rect -8138 244938 -8106 245174
rect -8726 209494 -8106 244938
rect -8726 209258 -8694 209494
rect -8458 209258 -8374 209494
rect -8138 209258 -8106 209494
rect -8726 209174 -8106 209258
rect -8726 208938 -8694 209174
rect -8458 208938 -8374 209174
rect -8138 208938 -8106 209174
rect -8726 173494 -8106 208938
rect -8726 173258 -8694 173494
rect -8458 173258 -8374 173494
rect -8138 173258 -8106 173494
rect -8726 173174 -8106 173258
rect -8726 172938 -8694 173174
rect -8458 172938 -8374 173174
rect -8138 172938 -8106 173174
rect -8726 137494 -8106 172938
rect -8726 137258 -8694 137494
rect -8458 137258 -8374 137494
rect -8138 137258 -8106 137494
rect -8726 137174 -8106 137258
rect -8726 136938 -8694 137174
rect -8458 136938 -8374 137174
rect -8138 136938 -8106 137174
rect -8726 101494 -8106 136938
rect -8726 101258 -8694 101494
rect -8458 101258 -8374 101494
rect -8138 101258 -8106 101494
rect -8726 101174 -8106 101258
rect -8726 100938 -8694 101174
rect -8458 100938 -8374 101174
rect -8138 100938 -8106 101174
rect -8726 65494 -8106 100938
rect -8726 65258 -8694 65494
rect -8458 65258 -8374 65494
rect -8138 65258 -8106 65494
rect -8726 65174 -8106 65258
rect -8726 64938 -8694 65174
rect -8458 64938 -8374 65174
rect -8138 64938 -8106 65174
rect -8726 29494 -8106 64938
rect -8726 29258 -8694 29494
rect -8458 29258 -8374 29494
rect -8138 29258 -8106 29494
rect -8726 29174 -8106 29258
rect -8726 28938 -8694 29174
rect -8458 28938 -8374 29174
rect -8138 28938 -8106 29174
rect -8726 -7066 -8106 28938
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 673774 -7146 710042
rect -7766 673538 -7734 673774
rect -7498 673538 -7414 673774
rect -7178 673538 -7146 673774
rect -7766 673454 -7146 673538
rect -7766 673218 -7734 673454
rect -7498 673218 -7414 673454
rect -7178 673218 -7146 673454
rect -7766 637774 -7146 673218
rect -7766 637538 -7734 637774
rect -7498 637538 -7414 637774
rect -7178 637538 -7146 637774
rect -7766 637454 -7146 637538
rect -7766 637218 -7734 637454
rect -7498 637218 -7414 637454
rect -7178 637218 -7146 637454
rect -7766 601774 -7146 637218
rect -7766 601538 -7734 601774
rect -7498 601538 -7414 601774
rect -7178 601538 -7146 601774
rect -7766 601454 -7146 601538
rect -7766 601218 -7734 601454
rect -7498 601218 -7414 601454
rect -7178 601218 -7146 601454
rect -7766 565774 -7146 601218
rect -7766 565538 -7734 565774
rect -7498 565538 -7414 565774
rect -7178 565538 -7146 565774
rect -7766 565454 -7146 565538
rect -7766 565218 -7734 565454
rect -7498 565218 -7414 565454
rect -7178 565218 -7146 565454
rect -7766 529774 -7146 565218
rect -7766 529538 -7734 529774
rect -7498 529538 -7414 529774
rect -7178 529538 -7146 529774
rect -7766 529454 -7146 529538
rect -7766 529218 -7734 529454
rect -7498 529218 -7414 529454
rect -7178 529218 -7146 529454
rect -7766 493774 -7146 529218
rect -7766 493538 -7734 493774
rect -7498 493538 -7414 493774
rect -7178 493538 -7146 493774
rect -7766 493454 -7146 493538
rect -7766 493218 -7734 493454
rect -7498 493218 -7414 493454
rect -7178 493218 -7146 493454
rect -7766 457774 -7146 493218
rect -7766 457538 -7734 457774
rect -7498 457538 -7414 457774
rect -7178 457538 -7146 457774
rect -7766 457454 -7146 457538
rect -7766 457218 -7734 457454
rect -7498 457218 -7414 457454
rect -7178 457218 -7146 457454
rect -7766 421774 -7146 457218
rect -7766 421538 -7734 421774
rect -7498 421538 -7414 421774
rect -7178 421538 -7146 421774
rect -7766 421454 -7146 421538
rect -7766 421218 -7734 421454
rect -7498 421218 -7414 421454
rect -7178 421218 -7146 421454
rect -7766 385774 -7146 421218
rect -7766 385538 -7734 385774
rect -7498 385538 -7414 385774
rect -7178 385538 -7146 385774
rect -7766 385454 -7146 385538
rect -7766 385218 -7734 385454
rect -7498 385218 -7414 385454
rect -7178 385218 -7146 385454
rect -7766 349774 -7146 385218
rect -7766 349538 -7734 349774
rect -7498 349538 -7414 349774
rect -7178 349538 -7146 349774
rect -7766 349454 -7146 349538
rect -7766 349218 -7734 349454
rect -7498 349218 -7414 349454
rect -7178 349218 -7146 349454
rect -7766 313774 -7146 349218
rect -7766 313538 -7734 313774
rect -7498 313538 -7414 313774
rect -7178 313538 -7146 313774
rect -7766 313454 -7146 313538
rect -7766 313218 -7734 313454
rect -7498 313218 -7414 313454
rect -7178 313218 -7146 313454
rect -7766 277774 -7146 313218
rect -7766 277538 -7734 277774
rect -7498 277538 -7414 277774
rect -7178 277538 -7146 277774
rect -7766 277454 -7146 277538
rect -7766 277218 -7734 277454
rect -7498 277218 -7414 277454
rect -7178 277218 -7146 277454
rect -7766 241774 -7146 277218
rect -7766 241538 -7734 241774
rect -7498 241538 -7414 241774
rect -7178 241538 -7146 241774
rect -7766 241454 -7146 241538
rect -7766 241218 -7734 241454
rect -7498 241218 -7414 241454
rect -7178 241218 -7146 241454
rect -7766 205774 -7146 241218
rect -7766 205538 -7734 205774
rect -7498 205538 -7414 205774
rect -7178 205538 -7146 205774
rect -7766 205454 -7146 205538
rect -7766 205218 -7734 205454
rect -7498 205218 -7414 205454
rect -7178 205218 -7146 205454
rect -7766 169774 -7146 205218
rect -7766 169538 -7734 169774
rect -7498 169538 -7414 169774
rect -7178 169538 -7146 169774
rect -7766 169454 -7146 169538
rect -7766 169218 -7734 169454
rect -7498 169218 -7414 169454
rect -7178 169218 -7146 169454
rect -7766 133774 -7146 169218
rect -7766 133538 -7734 133774
rect -7498 133538 -7414 133774
rect -7178 133538 -7146 133774
rect -7766 133454 -7146 133538
rect -7766 133218 -7734 133454
rect -7498 133218 -7414 133454
rect -7178 133218 -7146 133454
rect -7766 97774 -7146 133218
rect -7766 97538 -7734 97774
rect -7498 97538 -7414 97774
rect -7178 97538 -7146 97774
rect -7766 97454 -7146 97538
rect -7766 97218 -7734 97454
rect -7498 97218 -7414 97454
rect -7178 97218 -7146 97454
rect -7766 61774 -7146 97218
rect -7766 61538 -7734 61774
rect -7498 61538 -7414 61774
rect -7178 61538 -7146 61774
rect -7766 61454 -7146 61538
rect -7766 61218 -7734 61454
rect -7498 61218 -7414 61454
rect -7178 61218 -7146 61454
rect -7766 25774 -7146 61218
rect -7766 25538 -7734 25774
rect -7498 25538 -7414 25774
rect -7178 25538 -7146 25774
rect -7766 25454 -7146 25538
rect -7766 25218 -7734 25454
rect -7498 25218 -7414 25454
rect -7178 25218 -7146 25454
rect -7766 -6106 -7146 25218
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 670054 -6186 709082
rect -6806 669818 -6774 670054
rect -6538 669818 -6454 670054
rect -6218 669818 -6186 670054
rect -6806 669734 -6186 669818
rect -6806 669498 -6774 669734
rect -6538 669498 -6454 669734
rect -6218 669498 -6186 669734
rect -6806 634054 -6186 669498
rect -6806 633818 -6774 634054
rect -6538 633818 -6454 634054
rect -6218 633818 -6186 634054
rect -6806 633734 -6186 633818
rect -6806 633498 -6774 633734
rect -6538 633498 -6454 633734
rect -6218 633498 -6186 633734
rect -6806 598054 -6186 633498
rect -6806 597818 -6774 598054
rect -6538 597818 -6454 598054
rect -6218 597818 -6186 598054
rect -6806 597734 -6186 597818
rect -6806 597498 -6774 597734
rect -6538 597498 -6454 597734
rect -6218 597498 -6186 597734
rect -6806 562054 -6186 597498
rect -6806 561818 -6774 562054
rect -6538 561818 -6454 562054
rect -6218 561818 -6186 562054
rect -6806 561734 -6186 561818
rect -6806 561498 -6774 561734
rect -6538 561498 -6454 561734
rect -6218 561498 -6186 561734
rect -6806 526054 -6186 561498
rect -6806 525818 -6774 526054
rect -6538 525818 -6454 526054
rect -6218 525818 -6186 526054
rect -6806 525734 -6186 525818
rect -6806 525498 -6774 525734
rect -6538 525498 -6454 525734
rect -6218 525498 -6186 525734
rect -6806 490054 -6186 525498
rect -6806 489818 -6774 490054
rect -6538 489818 -6454 490054
rect -6218 489818 -6186 490054
rect -6806 489734 -6186 489818
rect -6806 489498 -6774 489734
rect -6538 489498 -6454 489734
rect -6218 489498 -6186 489734
rect -6806 454054 -6186 489498
rect -6806 453818 -6774 454054
rect -6538 453818 -6454 454054
rect -6218 453818 -6186 454054
rect -6806 453734 -6186 453818
rect -6806 453498 -6774 453734
rect -6538 453498 -6454 453734
rect -6218 453498 -6186 453734
rect -6806 418054 -6186 453498
rect -6806 417818 -6774 418054
rect -6538 417818 -6454 418054
rect -6218 417818 -6186 418054
rect -6806 417734 -6186 417818
rect -6806 417498 -6774 417734
rect -6538 417498 -6454 417734
rect -6218 417498 -6186 417734
rect -6806 382054 -6186 417498
rect -6806 381818 -6774 382054
rect -6538 381818 -6454 382054
rect -6218 381818 -6186 382054
rect -6806 381734 -6186 381818
rect -6806 381498 -6774 381734
rect -6538 381498 -6454 381734
rect -6218 381498 -6186 381734
rect -6806 346054 -6186 381498
rect -6806 345818 -6774 346054
rect -6538 345818 -6454 346054
rect -6218 345818 -6186 346054
rect -6806 345734 -6186 345818
rect -6806 345498 -6774 345734
rect -6538 345498 -6454 345734
rect -6218 345498 -6186 345734
rect -6806 310054 -6186 345498
rect -6806 309818 -6774 310054
rect -6538 309818 -6454 310054
rect -6218 309818 -6186 310054
rect -6806 309734 -6186 309818
rect -6806 309498 -6774 309734
rect -6538 309498 -6454 309734
rect -6218 309498 -6186 309734
rect -6806 274054 -6186 309498
rect -6806 273818 -6774 274054
rect -6538 273818 -6454 274054
rect -6218 273818 -6186 274054
rect -6806 273734 -6186 273818
rect -6806 273498 -6774 273734
rect -6538 273498 -6454 273734
rect -6218 273498 -6186 273734
rect -6806 238054 -6186 273498
rect -6806 237818 -6774 238054
rect -6538 237818 -6454 238054
rect -6218 237818 -6186 238054
rect -6806 237734 -6186 237818
rect -6806 237498 -6774 237734
rect -6538 237498 -6454 237734
rect -6218 237498 -6186 237734
rect -6806 202054 -6186 237498
rect -6806 201818 -6774 202054
rect -6538 201818 -6454 202054
rect -6218 201818 -6186 202054
rect -6806 201734 -6186 201818
rect -6806 201498 -6774 201734
rect -6538 201498 -6454 201734
rect -6218 201498 -6186 201734
rect -6806 166054 -6186 201498
rect -6806 165818 -6774 166054
rect -6538 165818 -6454 166054
rect -6218 165818 -6186 166054
rect -6806 165734 -6186 165818
rect -6806 165498 -6774 165734
rect -6538 165498 -6454 165734
rect -6218 165498 -6186 165734
rect -6806 130054 -6186 165498
rect -6806 129818 -6774 130054
rect -6538 129818 -6454 130054
rect -6218 129818 -6186 130054
rect -6806 129734 -6186 129818
rect -6806 129498 -6774 129734
rect -6538 129498 -6454 129734
rect -6218 129498 -6186 129734
rect -6806 94054 -6186 129498
rect -6806 93818 -6774 94054
rect -6538 93818 -6454 94054
rect -6218 93818 -6186 94054
rect -6806 93734 -6186 93818
rect -6806 93498 -6774 93734
rect -6538 93498 -6454 93734
rect -6218 93498 -6186 93734
rect -6806 58054 -6186 93498
rect -6806 57818 -6774 58054
rect -6538 57818 -6454 58054
rect -6218 57818 -6186 58054
rect -6806 57734 -6186 57818
rect -6806 57498 -6774 57734
rect -6538 57498 -6454 57734
rect -6218 57498 -6186 57734
rect -6806 22054 -6186 57498
rect -6806 21818 -6774 22054
rect -6538 21818 -6454 22054
rect -6218 21818 -6186 22054
rect -6806 21734 -6186 21818
rect -6806 21498 -6774 21734
rect -6538 21498 -6454 21734
rect -6218 21498 -6186 21734
rect -6806 -5146 -6186 21498
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 666334 -5226 708122
rect -5846 666098 -5814 666334
rect -5578 666098 -5494 666334
rect -5258 666098 -5226 666334
rect -5846 666014 -5226 666098
rect -5846 665778 -5814 666014
rect -5578 665778 -5494 666014
rect -5258 665778 -5226 666014
rect -5846 630334 -5226 665778
rect -5846 630098 -5814 630334
rect -5578 630098 -5494 630334
rect -5258 630098 -5226 630334
rect -5846 630014 -5226 630098
rect -5846 629778 -5814 630014
rect -5578 629778 -5494 630014
rect -5258 629778 -5226 630014
rect -5846 594334 -5226 629778
rect -5846 594098 -5814 594334
rect -5578 594098 -5494 594334
rect -5258 594098 -5226 594334
rect -5846 594014 -5226 594098
rect -5846 593778 -5814 594014
rect -5578 593778 -5494 594014
rect -5258 593778 -5226 594014
rect -5846 558334 -5226 593778
rect -5846 558098 -5814 558334
rect -5578 558098 -5494 558334
rect -5258 558098 -5226 558334
rect -5846 558014 -5226 558098
rect -5846 557778 -5814 558014
rect -5578 557778 -5494 558014
rect -5258 557778 -5226 558014
rect -5846 522334 -5226 557778
rect -5846 522098 -5814 522334
rect -5578 522098 -5494 522334
rect -5258 522098 -5226 522334
rect -5846 522014 -5226 522098
rect -5846 521778 -5814 522014
rect -5578 521778 -5494 522014
rect -5258 521778 -5226 522014
rect -5846 486334 -5226 521778
rect -5846 486098 -5814 486334
rect -5578 486098 -5494 486334
rect -5258 486098 -5226 486334
rect -5846 486014 -5226 486098
rect -5846 485778 -5814 486014
rect -5578 485778 -5494 486014
rect -5258 485778 -5226 486014
rect -5846 450334 -5226 485778
rect -5846 450098 -5814 450334
rect -5578 450098 -5494 450334
rect -5258 450098 -5226 450334
rect -5846 450014 -5226 450098
rect -5846 449778 -5814 450014
rect -5578 449778 -5494 450014
rect -5258 449778 -5226 450014
rect -5846 414334 -5226 449778
rect -5846 414098 -5814 414334
rect -5578 414098 -5494 414334
rect -5258 414098 -5226 414334
rect -5846 414014 -5226 414098
rect -5846 413778 -5814 414014
rect -5578 413778 -5494 414014
rect -5258 413778 -5226 414014
rect -5846 378334 -5226 413778
rect -5846 378098 -5814 378334
rect -5578 378098 -5494 378334
rect -5258 378098 -5226 378334
rect -5846 378014 -5226 378098
rect -5846 377778 -5814 378014
rect -5578 377778 -5494 378014
rect -5258 377778 -5226 378014
rect -5846 342334 -5226 377778
rect -5846 342098 -5814 342334
rect -5578 342098 -5494 342334
rect -5258 342098 -5226 342334
rect -5846 342014 -5226 342098
rect -5846 341778 -5814 342014
rect -5578 341778 -5494 342014
rect -5258 341778 -5226 342014
rect -5846 306334 -5226 341778
rect -5846 306098 -5814 306334
rect -5578 306098 -5494 306334
rect -5258 306098 -5226 306334
rect -5846 306014 -5226 306098
rect -5846 305778 -5814 306014
rect -5578 305778 -5494 306014
rect -5258 305778 -5226 306014
rect -5846 270334 -5226 305778
rect -5846 270098 -5814 270334
rect -5578 270098 -5494 270334
rect -5258 270098 -5226 270334
rect -5846 270014 -5226 270098
rect -5846 269778 -5814 270014
rect -5578 269778 -5494 270014
rect -5258 269778 -5226 270014
rect -5846 234334 -5226 269778
rect -5846 234098 -5814 234334
rect -5578 234098 -5494 234334
rect -5258 234098 -5226 234334
rect -5846 234014 -5226 234098
rect -5846 233778 -5814 234014
rect -5578 233778 -5494 234014
rect -5258 233778 -5226 234014
rect -5846 198334 -5226 233778
rect -5846 198098 -5814 198334
rect -5578 198098 -5494 198334
rect -5258 198098 -5226 198334
rect -5846 198014 -5226 198098
rect -5846 197778 -5814 198014
rect -5578 197778 -5494 198014
rect -5258 197778 -5226 198014
rect -5846 162334 -5226 197778
rect -5846 162098 -5814 162334
rect -5578 162098 -5494 162334
rect -5258 162098 -5226 162334
rect -5846 162014 -5226 162098
rect -5846 161778 -5814 162014
rect -5578 161778 -5494 162014
rect -5258 161778 -5226 162014
rect -5846 126334 -5226 161778
rect -5846 126098 -5814 126334
rect -5578 126098 -5494 126334
rect -5258 126098 -5226 126334
rect -5846 126014 -5226 126098
rect -5846 125778 -5814 126014
rect -5578 125778 -5494 126014
rect -5258 125778 -5226 126014
rect -5846 90334 -5226 125778
rect -5846 90098 -5814 90334
rect -5578 90098 -5494 90334
rect -5258 90098 -5226 90334
rect -5846 90014 -5226 90098
rect -5846 89778 -5814 90014
rect -5578 89778 -5494 90014
rect -5258 89778 -5226 90014
rect -5846 54334 -5226 89778
rect -5846 54098 -5814 54334
rect -5578 54098 -5494 54334
rect -5258 54098 -5226 54334
rect -5846 54014 -5226 54098
rect -5846 53778 -5814 54014
rect -5578 53778 -5494 54014
rect -5258 53778 -5226 54014
rect -5846 18334 -5226 53778
rect -5846 18098 -5814 18334
rect -5578 18098 -5494 18334
rect -5258 18098 -5226 18334
rect -5846 18014 -5226 18098
rect -5846 17778 -5814 18014
rect -5578 17778 -5494 18014
rect -5258 17778 -5226 18014
rect -5846 -4186 -5226 17778
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 698614 -4266 707162
rect -4886 698378 -4854 698614
rect -4618 698378 -4534 698614
rect -4298 698378 -4266 698614
rect -4886 698294 -4266 698378
rect -4886 698058 -4854 698294
rect -4618 698058 -4534 698294
rect -4298 698058 -4266 698294
rect -4886 662614 -4266 698058
rect -4886 662378 -4854 662614
rect -4618 662378 -4534 662614
rect -4298 662378 -4266 662614
rect -4886 662294 -4266 662378
rect -4886 662058 -4854 662294
rect -4618 662058 -4534 662294
rect -4298 662058 -4266 662294
rect -4886 626614 -4266 662058
rect -4886 626378 -4854 626614
rect -4618 626378 -4534 626614
rect -4298 626378 -4266 626614
rect -4886 626294 -4266 626378
rect -4886 626058 -4854 626294
rect -4618 626058 -4534 626294
rect -4298 626058 -4266 626294
rect -4886 590614 -4266 626058
rect -4886 590378 -4854 590614
rect -4618 590378 -4534 590614
rect -4298 590378 -4266 590614
rect -4886 590294 -4266 590378
rect -4886 590058 -4854 590294
rect -4618 590058 -4534 590294
rect -4298 590058 -4266 590294
rect -4886 554614 -4266 590058
rect -4886 554378 -4854 554614
rect -4618 554378 -4534 554614
rect -4298 554378 -4266 554614
rect -4886 554294 -4266 554378
rect -4886 554058 -4854 554294
rect -4618 554058 -4534 554294
rect -4298 554058 -4266 554294
rect -4886 518614 -4266 554058
rect -4886 518378 -4854 518614
rect -4618 518378 -4534 518614
rect -4298 518378 -4266 518614
rect -4886 518294 -4266 518378
rect -4886 518058 -4854 518294
rect -4618 518058 -4534 518294
rect -4298 518058 -4266 518294
rect -4886 482614 -4266 518058
rect -4886 482378 -4854 482614
rect -4618 482378 -4534 482614
rect -4298 482378 -4266 482614
rect -4886 482294 -4266 482378
rect -4886 482058 -4854 482294
rect -4618 482058 -4534 482294
rect -4298 482058 -4266 482294
rect -4886 446614 -4266 482058
rect -4886 446378 -4854 446614
rect -4618 446378 -4534 446614
rect -4298 446378 -4266 446614
rect -4886 446294 -4266 446378
rect -4886 446058 -4854 446294
rect -4618 446058 -4534 446294
rect -4298 446058 -4266 446294
rect -4886 410614 -4266 446058
rect -4886 410378 -4854 410614
rect -4618 410378 -4534 410614
rect -4298 410378 -4266 410614
rect -4886 410294 -4266 410378
rect -4886 410058 -4854 410294
rect -4618 410058 -4534 410294
rect -4298 410058 -4266 410294
rect -4886 374614 -4266 410058
rect -4886 374378 -4854 374614
rect -4618 374378 -4534 374614
rect -4298 374378 -4266 374614
rect -4886 374294 -4266 374378
rect -4886 374058 -4854 374294
rect -4618 374058 -4534 374294
rect -4298 374058 -4266 374294
rect -4886 338614 -4266 374058
rect -4886 338378 -4854 338614
rect -4618 338378 -4534 338614
rect -4298 338378 -4266 338614
rect -4886 338294 -4266 338378
rect -4886 338058 -4854 338294
rect -4618 338058 -4534 338294
rect -4298 338058 -4266 338294
rect -4886 302614 -4266 338058
rect -4886 302378 -4854 302614
rect -4618 302378 -4534 302614
rect -4298 302378 -4266 302614
rect -4886 302294 -4266 302378
rect -4886 302058 -4854 302294
rect -4618 302058 -4534 302294
rect -4298 302058 -4266 302294
rect -4886 266614 -4266 302058
rect -4886 266378 -4854 266614
rect -4618 266378 -4534 266614
rect -4298 266378 -4266 266614
rect -4886 266294 -4266 266378
rect -4886 266058 -4854 266294
rect -4618 266058 -4534 266294
rect -4298 266058 -4266 266294
rect -4886 230614 -4266 266058
rect -4886 230378 -4854 230614
rect -4618 230378 -4534 230614
rect -4298 230378 -4266 230614
rect -4886 230294 -4266 230378
rect -4886 230058 -4854 230294
rect -4618 230058 -4534 230294
rect -4298 230058 -4266 230294
rect -4886 194614 -4266 230058
rect -4886 194378 -4854 194614
rect -4618 194378 -4534 194614
rect -4298 194378 -4266 194614
rect -4886 194294 -4266 194378
rect -4886 194058 -4854 194294
rect -4618 194058 -4534 194294
rect -4298 194058 -4266 194294
rect -4886 158614 -4266 194058
rect -4886 158378 -4854 158614
rect -4618 158378 -4534 158614
rect -4298 158378 -4266 158614
rect -4886 158294 -4266 158378
rect -4886 158058 -4854 158294
rect -4618 158058 -4534 158294
rect -4298 158058 -4266 158294
rect -4886 122614 -4266 158058
rect -4886 122378 -4854 122614
rect -4618 122378 -4534 122614
rect -4298 122378 -4266 122614
rect -4886 122294 -4266 122378
rect -4886 122058 -4854 122294
rect -4618 122058 -4534 122294
rect -4298 122058 -4266 122294
rect -4886 86614 -4266 122058
rect -4886 86378 -4854 86614
rect -4618 86378 -4534 86614
rect -4298 86378 -4266 86614
rect -4886 86294 -4266 86378
rect -4886 86058 -4854 86294
rect -4618 86058 -4534 86294
rect -4298 86058 -4266 86294
rect -4886 50614 -4266 86058
rect -4886 50378 -4854 50614
rect -4618 50378 -4534 50614
rect -4298 50378 -4266 50614
rect -4886 50294 -4266 50378
rect -4886 50058 -4854 50294
rect -4618 50058 -4534 50294
rect -4298 50058 -4266 50294
rect -4886 14614 -4266 50058
rect -4886 14378 -4854 14614
rect -4618 14378 -4534 14614
rect -4298 14378 -4266 14614
rect -4886 14294 -4266 14378
rect -4886 14058 -4854 14294
rect -4618 14058 -4534 14294
rect -4298 14058 -4266 14294
rect -4886 -3226 -4266 14058
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 694894 -3306 706202
rect -3926 694658 -3894 694894
rect -3658 694658 -3574 694894
rect -3338 694658 -3306 694894
rect -3926 694574 -3306 694658
rect -3926 694338 -3894 694574
rect -3658 694338 -3574 694574
rect -3338 694338 -3306 694574
rect -3926 658894 -3306 694338
rect -3926 658658 -3894 658894
rect -3658 658658 -3574 658894
rect -3338 658658 -3306 658894
rect -3926 658574 -3306 658658
rect -3926 658338 -3894 658574
rect -3658 658338 -3574 658574
rect -3338 658338 -3306 658574
rect -3926 622894 -3306 658338
rect -3926 622658 -3894 622894
rect -3658 622658 -3574 622894
rect -3338 622658 -3306 622894
rect -3926 622574 -3306 622658
rect -3926 622338 -3894 622574
rect -3658 622338 -3574 622574
rect -3338 622338 -3306 622574
rect -3926 586894 -3306 622338
rect -3926 586658 -3894 586894
rect -3658 586658 -3574 586894
rect -3338 586658 -3306 586894
rect -3926 586574 -3306 586658
rect -3926 586338 -3894 586574
rect -3658 586338 -3574 586574
rect -3338 586338 -3306 586574
rect -3926 550894 -3306 586338
rect -3926 550658 -3894 550894
rect -3658 550658 -3574 550894
rect -3338 550658 -3306 550894
rect -3926 550574 -3306 550658
rect -3926 550338 -3894 550574
rect -3658 550338 -3574 550574
rect -3338 550338 -3306 550574
rect -3926 514894 -3306 550338
rect -3926 514658 -3894 514894
rect -3658 514658 -3574 514894
rect -3338 514658 -3306 514894
rect -3926 514574 -3306 514658
rect -3926 514338 -3894 514574
rect -3658 514338 -3574 514574
rect -3338 514338 -3306 514574
rect -3926 478894 -3306 514338
rect -3926 478658 -3894 478894
rect -3658 478658 -3574 478894
rect -3338 478658 -3306 478894
rect -3926 478574 -3306 478658
rect -3926 478338 -3894 478574
rect -3658 478338 -3574 478574
rect -3338 478338 -3306 478574
rect -3926 442894 -3306 478338
rect -3926 442658 -3894 442894
rect -3658 442658 -3574 442894
rect -3338 442658 -3306 442894
rect -3926 442574 -3306 442658
rect -3926 442338 -3894 442574
rect -3658 442338 -3574 442574
rect -3338 442338 -3306 442574
rect -3926 406894 -3306 442338
rect -3926 406658 -3894 406894
rect -3658 406658 -3574 406894
rect -3338 406658 -3306 406894
rect -3926 406574 -3306 406658
rect -3926 406338 -3894 406574
rect -3658 406338 -3574 406574
rect -3338 406338 -3306 406574
rect -3926 370894 -3306 406338
rect -3926 370658 -3894 370894
rect -3658 370658 -3574 370894
rect -3338 370658 -3306 370894
rect -3926 370574 -3306 370658
rect -3926 370338 -3894 370574
rect -3658 370338 -3574 370574
rect -3338 370338 -3306 370574
rect -3926 334894 -3306 370338
rect -3926 334658 -3894 334894
rect -3658 334658 -3574 334894
rect -3338 334658 -3306 334894
rect -3926 334574 -3306 334658
rect -3926 334338 -3894 334574
rect -3658 334338 -3574 334574
rect -3338 334338 -3306 334574
rect -3926 298894 -3306 334338
rect -3926 298658 -3894 298894
rect -3658 298658 -3574 298894
rect -3338 298658 -3306 298894
rect -3926 298574 -3306 298658
rect -3926 298338 -3894 298574
rect -3658 298338 -3574 298574
rect -3338 298338 -3306 298574
rect -3926 262894 -3306 298338
rect -3926 262658 -3894 262894
rect -3658 262658 -3574 262894
rect -3338 262658 -3306 262894
rect -3926 262574 -3306 262658
rect -3926 262338 -3894 262574
rect -3658 262338 -3574 262574
rect -3338 262338 -3306 262574
rect -3926 226894 -3306 262338
rect -3926 226658 -3894 226894
rect -3658 226658 -3574 226894
rect -3338 226658 -3306 226894
rect -3926 226574 -3306 226658
rect -3926 226338 -3894 226574
rect -3658 226338 -3574 226574
rect -3338 226338 -3306 226574
rect -3926 190894 -3306 226338
rect -3926 190658 -3894 190894
rect -3658 190658 -3574 190894
rect -3338 190658 -3306 190894
rect -3926 190574 -3306 190658
rect -3926 190338 -3894 190574
rect -3658 190338 -3574 190574
rect -3338 190338 -3306 190574
rect -3926 154894 -3306 190338
rect -3926 154658 -3894 154894
rect -3658 154658 -3574 154894
rect -3338 154658 -3306 154894
rect -3926 154574 -3306 154658
rect -3926 154338 -3894 154574
rect -3658 154338 -3574 154574
rect -3338 154338 -3306 154574
rect -3926 118894 -3306 154338
rect -3926 118658 -3894 118894
rect -3658 118658 -3574 118894
rect -3338 118658 -3306 118894
rect -3926 118574 -3306 118658
rect -3926 118338 -3894 118574
rect -3658 118338 -3574 118574
rect -3338 118338 -3306 118574
rect -3926 82894 -3306 118338
rect -3926 82658 -3894 82894
rect -3658 82658 -3574 82894
rect -3338 82658 -3306 82894
rect -3926 82574 -3306 82658
rect -3926 82338 -3894 82574
rect -3658 82338 -3574 82574
rect -3338 82338 -3306 82574
rect -3926 46894 -3306 82338
rect -3926 46658 -3894 46894
rect -3658 46658 -3574 46894
rect -3338 46658 -3306 46894
rect -3926 46574 -3306 46658
rect -3926 46338 -3894 46574
rect -3658 46338 -3574 46574
rect -3338 46338 -3306 46574
rect -3926 10894 -3306 46338
rect -3926 10658 -3894 10894
rect -3658 10658 -3574 10894
rect -3338 10658 -3306 10894
rect -3926 10574 -3306 10658
rect -3926 10338 -3894 10574
rect -3658 10338 -3574 10574
rect -3338 10338 -3306 10574
rect -3926 -2266 -3306 10338
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 691174 -2346 705242
rect -2966 690938 -2934 691174
rect -2698 690938 -2614 691174
rect -2378 690938 -2346 691174
rect -2966 690854 -2346 690938
rect -2966 690618 -2934 690854
rect -2698 690618 -2614 690854
rect -2378 690618 -2346 690854
rect -2966 655174 -2346 690618
rect -2966 654938 -2934 655174
rect -2698 654938 -2614 655174
rect -2378 654938 -2346 655174
rect -2966 654854 -2346 654938
rect -2966 654618 -2934 654854
rect -2698 654618 -2614 654854
rect -2378 654618 -2346 654854
rect -2966 619174 -2346 654618
rect -2966 618938 -2934 619174
rect -2698 618938 -2614 619174
rect -2378 618938 -2346 619174
rect -2966 618854 -2346 618938
rect -2966 618618 -2934 618854
rect -2698 618618 -2614 618854
rect -2378 618618 -2346 618854
rect -2966 583174 -2346 618618
rect -2966 582938 -2934 583174
rect -2698 582938 -2614 583174
rect -2378 582938 -2346 583174
rect -2966 582854 -2346 582938
rect -2966 582618 -2934 582854
rect -2698 582618 -2614 582854
rect -2378 582618 -2346 582854
rect -2966 547174 -2346 582618
rect -2966 546938 -2934 547174
rect -2698 546938 -2614 547174
rect -2378 546938 -2346 547174
rect -2966 546854 -2346 546938
rect -2966 546618 -2934 546854
rect -2698 546618 -2614 546854
rect -2378 546618 -2346 546854
rect -2966 511174 -2346 546618
rect -2966 510938 -2934 511174
rect -2698 510938 -2614 511174
rect -2378 510938 -2346 511174
rect -2966 510854 -2346 510938
rect -2966 510618 -2934 510854
rect -2698 510618 -2614 510854
rect -2378 510618 -2346 510854
rect -2966 475174 -2346 510618
rect -2966 474938 -2934 475174
rect -2698 474938 -2614 475174
rect -2378 474938 -2346 475174
rect -2966 474854 -2346 474938
rect -2966 474618 -2934 474854
rect -2698 474618 -2614 474854
rect -2378 474618 -2346 474854
rect -2966 439174 -2346 474618
rect -2966 438938 -2934 439174
rect -2698 438938 -2614 439174
rect -2378 438938 -2346 439174
rect -2966 438854 -2346 438938
rect -2966 438618 -2934 438854
rect -2698 438618 -2614 438854
rect -2378 438618 -2346 438854
rect -2966 403174 -2346 438618
rect -2966 402938 -2934 403174
rect -2698 402938 -2614 403174
rect -2378 402938 -2346 403174
rect -2966 402854 -2346 402938
rect -2966 402618 -2934 402854
rect -2698 402618 -2614 402854
rect -2378 402618 -2346 402854
rect -2966 367174 -2346 402618
rect -2966 366938 -2934 367174
rect -2698 366938 -2614 367174
rect -2378 366938 -2346 367174
rect -2966 366854 -2346 366938
rect -2966 366618 -2934 366854
rect -2698 366618 -2614 366854
rect -2378 366618 -2346 366854
rect -2966 331174 -2346 366618
rect -2966 330938 -2934 331174
rect -2698 330938 -2614 331174
rect -2378 330938 -2346 331174
rect -2966 330854 -2346 330938
rect -2966 330618 -2934 330854
rect -2698 330618 -2614 330854
rect -2378 330618 -2346 330854
rect -2966 295174 -2346 330618
rect -2966 294938 -2934 295174
rect -2698 294938 -2614 295174
rect -2378 294938 -2346 295174
rect -2966 294854 -2346 294938
rect -2966 294618 -2934 294854
rect -2698 294618 -2614 294854
rect -2378 294618 -2346 294854
rect -2966 259174 -2346 294618
rect -2966 258938 -2934 259174
rect -2698 258938 -2614 259174
rect -2378 258938 -2346 259174
rect -2966 258854 -2346 258938
rect -2966 258618 -2934 258854
rect -2698 258618 -2614 258854
rect -2378 258618 -2346 258854
rect -2966 223174 -2346 258618
rect -2966 222938 -2934 223174
rect -2698 222938 -2614 223174
rect -2378 222938 -2346 223174
rect -2966 222854 -2346 222938
rect -2966 222618 -2934 222854
rect -2698 222618 -2614 222854
rect -2378 222618 -2346 222854
rect -2966 187174 -2346 222618
rect -2966 186938 -2934 187174
rect -2698 186938 -2614 187174
rect -2378 186938 -2346 187174
rect -2966 186854 -2346 186938
rect -2966 186618 -2934 186854
rect -2698 186618 -2614 186854
rect -2378 186618 -2346 186854
rect -2966 151174 -2346 186618
rect -2966 150938 -2934 151174
rect -2698 150938 -2614 151174
rect -2378 150938 -2346 151174
rect -2966 150854 -2346 150938
rect -2966 150618 -2934 150854
rect -2698 150618 -2614 150854
rect -2378 150618 -2346 150854
rect -2966 115174 -2346 150618
rect -2966 114938 -2934 115174
rect -2698 114938 -2614 115174
rect -2378 114938 -2346 115174
rect -2966 114854 -2346 114938
rect -2966 114618 -2934 114854
rect -2698 114618 -2614 114854
rect -2378 114618 -2346 114854
rect -2966 79174 -2346 114618
rect -2966 78938 -2934 79174
rect -2698 78938 -2614 79174
rect -2378 78938 -2346 79174
rect -2966 78854 -2346 78938
rect -2966 78618 -2934 78854
rect -2698 78618 -2614 78854
rect -2378 78618 -2346 78854
rect -2966 43174 -2346 78618
rect -2966 42938 -2934 43174
rect -2698 42938 -2614 43174
rect -2378 42938 -2346 43174
rect -2966 42854 -2346 42938
rect -2966 42618 -2934 42854
rect -2698 42618 -2614 42854
rect -2378 42618 -2346 42854
rect -2966 7174 -2346 42618
rect -2966 6938 -2934 7174
rect -2698 6938 -2614 7174
rect -2378 6938 -2346 7174
rect -2966 6854 -2346 6938
rect -2966 6618 -2934 6854
rect -2698 6618 -2614 6854
rect -2378 6618 -2346 6854
rect -2966 -1306 -2346 6618
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 687454 -1386 704282
rect -2006 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 -1386 687454
rect -2006 687134 -1386 687218
rect -2006 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 -1386 687134
rect -2006 651454 -1386 686898
rect -2006 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 -1386 651454
rect -2006 651134 -1386 651218
rect -2006 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 -1386 651134
rect -2006 615454 -1386 650898
rect -2006 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 -1386 615454
rect -2006 615134 -1386 615218
rect -2006 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 -1386 615134
rect -2006 579454 -1386 614898
rect -2006 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 -1386 579454
rect -2006 579134 -1386 579218
rect -2006 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 -1386 579134
rect -2006 543454 -1386 578898
rect -2006 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 -1386 543454
rect -2006 543134 -1386 543218
rect -2006 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 -1386 543134
rect -2006 507454 -1386 542898
rect -2006 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 -1386 507454
rect -2006 507134 -1386 507218
rect -2006 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 -1386 507134
rect -2006 471454 -1386 506898
rect -2006 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 -1386 471454
rect -2006 471134 -1386 471218
rect -2006 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 -1386 471134
rect -2006 435454 -1386 470898
rect -2006 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 -1386 435454
rect -2006 435134 -1386 435218
rect -2006 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 -1386 435134
rect -2006 399454 -1386 434898
rect -2006 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 -1386 399454
rect -2006 399134 -1386 399218
rect -2006 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 -1386 399134
rect -2006 363454 -1386 398898
rect -2006 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 -1386 363454
rect -2006 363134 -1386 363218
rect -2006 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 -1386 363134
rect -2006 327454 -1386 362898
rect -2006 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 -1386 327454
rect -2006 327134 -1386 327218
rect -2006 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 -1386 327134
rect -2006 291454 -1386 326898
rect -2006 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 -1386 291454
rect -2006 291134 -1386 291218
rect -2006 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 -1386 291134
rect -2006 255454 -1386 290898
rect -2006 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 -1386 255454
rect -2006 255134 -1386 255218
rect -2006 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 -1386 255134
rect -2006 219454 -1386 254898
rect -2006 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 -1386 219454
rect -2006 219134 -1386 219218
rect -2006 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 -1386 219134
rect -2006 183454 -1386 218898
rect -2006 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 -1386 183454
rect -2006 183134 -1386 183218
rect -2006 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 -1386 183134
rect -2006 147454 -1386 182898
rect -2006 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 -1386 147454
rect -2006 147134 -1386 147218
rect -2006 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 -1386 147134
rect -2006 111454 -1386 146898
rect -2006 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 -1386 111454
rect -2006 111134 -1386 111218
rect -2006 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 -1386 111134
rect -2006 75454 -1386 110898
rect -2006 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 -1386 75454
rect -2006 75134 -1386 75218
rect -2006 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 -1386 75134
rect -2006 39454 -1386 74898
rect -2006 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 -1386 39454
rect -2006 39134 -1386 39218
rect -2006 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 -1386 39134
rect -2006 3454 -1386 38898
rect -2006 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 -1386 3454
rect -2006 3134 -1386 3218
rect -2006 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 -1386 3134
rect -2006 -346 -1386 2898
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect 1794 704838 2414 711590
rect 1794 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 2414 704838
rect 1794 704518 2414 704602
rect 1794 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 2414 704518
rect 1794 687454 2414 704282
rect 1794 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 2414 687454
rect 1794 687134 2414 687218
rect 1794 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 2414 687134
rect 1794 651454 2414 686898
rect 5514 705798 6134 711590
rect 5514 705562 5546 705798
rect 5782 705562 5866 705798
rect 6102 705562 6134 705798
rect 5514 705478 6134 705562
rect 5514 705242 5546 705478
rect 5782 705242 5866 705478
rect 6102 705242 6134 705478
rect 5514 691174 6134 705242
rect 5514 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 6134 691174
rect 5514 690854 6134 690938
rect 5514 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 6134 690854
rect 3739 683364 3805 683365
rect 3739 683300 3740 683364
rect 3804 683300 3805 683364
rect 3739 683299 3805 683300
rect 3555 683228 3621 683229
rect 3555 683164 3556 683228
rect 3620 683164 3621 683228
rect 3555 683163 3621 683164
rect 3371 682820 3437 682821
rect 3371 682756 3372 682820
rect 3436 682756 3437 682820
rect 3371 682755 3437 682756
rect 1794 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 2414 651454
rect 1794 651134 2414 651218
rect 1794 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 2414 651134
rect 1794 615454 2414 650898
rect 1794 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 2414 615454
rect 1794 615134 2414 615218
rect 1794 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 2414 615134
rect 1794 579454 2414 614898
rect 3374 606117 3434 682755
rect 3558 619173 3618 683163
rect 3742 671261 3802 683299
rect 3739 671260 3805 671261
rect 3739 671196 3740 671260
rect 3804 671196 3805 671260
rect 3739 671195 3805 671196
rect 5514 655174 6134 690618
rect 5514 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 6134 655174
rect 5514 654854 6134 654938
rect 5514 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 6134 654854
rect 5514 619174 6134 654618
rect 3555 619172 3621 619173
rect 3555 619108 3556 619172
rect 3620 619108 3621 619172
rect 3555 619107 3621 619108
rect 5514 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 6134 619174
rect 5514 618854 6134 618938
rect 5514 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 6134 618854
rect 3371 606116 3437 606117
rect 3371 606052 3372 606116
rect 3436 606052 3437 606116
rect 3371 606051 3437 606052
rect 1794 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 2414 579454
rect 1794 579134 2414 579218
rect 1794 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 2414 579134
rect 1794 543454 2414 578898
rect 1794 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 2414 543454
rect 1794 543134 2414 543218
rect 1794 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 2414 543134
rect 1794 507454 2414 542898
rect 1794 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 2414 507454
rect 1794 507134 2414 507218
rect 1794 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 2414 507134
rect 1794 471454 2414 506898
rect 1794 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 2414 471454
rect 1794 471134 2414 471218
rect 1794 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 2414 471134
rect 1794 435454 2414 470898
rect 1794 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 2414 435454
rect 1794 435134 2414 435218
rect 1794 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 2414 435134
rect 1794 399454 2414 434898
rect 1794 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 2414 399454
rect 1794 399134 2414 399218
rect 1794 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 2414 399134
rect 1794 363454 2414 398898
rect 1794 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 2414 363454
rect 1794 363134 2414 363218
rect 1794 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 2414 363134
rect 1794 327454 2414 362898
rect 1794 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 2414 327454
rect 1794 327134 2414 327218
rect 1794 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 2414 327134
rect 1794 291454 2414 326898
rect 1794 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 2414 291454
rect 1794 291134 2414 291218
rect 1794 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 2414 291134
rect 1794 255454 2414 290898
rect 1794 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 2414 255454
rect 1794 255134 2414 255218
rect 1794 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 2414 255134
rect 1794 219454 2414 254898
rect 1794 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 2414 219454
rect 1794 219134 2414 219218
rect 1794 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 2414 219134
rect 1794 183454 2414 218898
rect 1794 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 2414 183454
rect 1794 183134 2414 183218
rect 1794 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 2414 183134
rect 1794 147454 2414 182898
rect 1794 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 2414 147454
rect 1794 147134 2414 147218
rect 1794 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 2414 147134
rect 1794 111454 2414 146898
rect 5514 583174 6134 618618
rect 5514 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 6134 583174
rect 5514 582854 6134 582938
rect 5514 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 6134 582854
rect 5514 547174 6134 582618
rect 5514 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 6134 547174
rect 5514 546854 6134 546938
rect 5514 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 6134 546854
rect 5514 511174 6134 546618
rect 5514 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 6134 511174
rect 5514 510854 6134 510938
rect 5514 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 6134 510854
rect 5514 475174 6134 510618
rect 5514 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 6134 475174
rect 5514 474854 6134 474938
rect 5514 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 6134 474854
rect 5514 439174 6134 474618
rect 5514 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 6134 439174
rect 5514 438854 6134 438938
rect 5514 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 6134 438854
rect 5514 403174 6134 438618
rect 5514 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 6134 403174
rect 5514 402854 6134 402938
rect 5514 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 6134 402854
rect 5514 367174 6134 402618
rect 5514 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 6134 367174
rect 5514 366854 6134 366938
rect 5514 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 6134 366854
rect 5514 331174 6134 366618
rect 5514 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 6134 331174
rect 5514 330854 6134 330938
rect 5514 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 6134 330854
rect 5514 295174 6134 330618
rect 5514 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 6134 295174
rect 5514 294854 6134 294938
rect 5514 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 6134 294854
rect 5514 259174 6134 294618
rect 5514 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 6134 259174
rect 5514 258854 6134 258938
rect 5514 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 6134 258854
rect 5514 223174 6134 258618
rect 5514 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 6134 223174
rect 5514 222854 6134 222938
rect 5514 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 6134 222854
rect 5514 187174 6134 222618
rect 5514 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 6134 187174
rect 5514 186854 6134 186938
rect 5514 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 6134 186854
rect 5514 151174 6134 186618
rect 5514 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 6134 151174
rect 5514 150854 6134 150938
rect 5514 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 6134 150854
rect 2819 136780 2885 136781
rect 2819 136716 2820 136780
rect 2884 136716 2885 136780
rect 2819 136715 2885 136716
rect 1794 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 2414 111454
rect 1794 111134 2414 111218
rect 1794 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 2414 111134
rect 1794 75454 2414 110898
rect 2822 98701 2882 136715
rect 5514 115174 6134 150618
rect 5514 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 6134 115174
rect 5514 114854 6134 114938
rect 5514 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 6134 114854
rect 3371 110668 3437 110669
rect 3371 110604 3372 110668
rect 3436 110604 3437 110668
rect 3371 110603 3437 110604
rect 2819 98700 2885 98701
rect 2819 98636 2820 98700
rect 2884 98636 2885 98700
rect 2819 98635 2885 98636
rect 1794 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 2414 75454
rect 1794 75134 2414 75218
rect 1794 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 2414 75134
rect 1794 39454 2414 74898
rect 3374 46749 3434 110603
rect 3555 97612 3621 97613
rect 3555 97548 3556 97612
rect 3620 97548 3621 97612
rect 3555 97547 3621 97548
rect 3558 46885 3618 97547
rect 5514 79174 6134 114618
rect 5514 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 6134 79174
rect 5514 78854 6134 78938
rect 5514 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 6134 78854
rect 3555 46884 3621 46885
rect 3555 46820 3556 46884
rect 3620 46820 3621 46884
rect 3555 46819 3621 46820
rect 3371 46748 3437 46749
rect 3371 46684 3372 46748
rect 3436 46684 3437 46748
rect 3371 46683 3437 46684
rect 1794 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 2414 39454
rect 1794 39134 2414 39218
rect 1794 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 2414 39134
rect 1794 3454 2414 38898
rect 1794 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 2414 3454
rect 1794 3134 2414 3218
rect 1794 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 2414 3134
rect 1794 -346 2414 2898
rect 1794 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 2414 -346
rect 1794 -666 2414 -582
rect 1794 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 2414 -666
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 1794 -7654 2414 -902
rect 5514 43174 6134 78618
rect 5514 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 6134 43174
rect 5514 42854 6134 42938
rect 5514 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 6134 42854
rect 5514 7174 6134 42618
rect 5514 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 6134 7174
rect 5514 6854 6134 6938
rect 5514 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 6134 6854
rect 5514 -1306 6134 6618
rect 5514 -1542 5546 -1306
rect 5782 -1542 5866 -1306
rect 6102 -1542 6134 -1306
rect 5514 -1626 6134 -1542
rect 5514 -1862 5546 -1626
rect 5782 -1862 5866 -1626
rect 6102 -1862 6134 -1626
rect 5514 -7654 6134 -1862
rect 9234 706758 9854 711590
rect 9234 706522 9266 706758
rect 9502 706522 9586 706758
rect 9822 706522 9854 706758
rect 9234 706438 9854 706522
rect 9234 706202 9266 706438
rect 9502 706202 9586 706438
rect 9822 706202 9854 706438
rect 9234 694894 9854 706202
rect 9234 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 9854 694894
rect 9234 694574 9854 694658
rect 9234 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 9854 694574
rect 9234 658894 9854 694338
rect 9234 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 9854 658894
rect 9234 658574 9854 658658
rect 9234 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 9854 658574
rect 9234 622894 9854 658338
rect 9234 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 9854 622894
rect 9234 622574 9854 622658
rect 9234 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 9854 622574
rect 9234 586894 9854 622338
rect 9234 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 9854 586894
rect 9234 586574 9854 586658
rect 9234 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 9854 586574
rect 9234 550894 9854 586338
rect 9234 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 9854 550894
rect 9234 550574 9854 550658
rect 9234 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 9854 550574
rect 9234 514894 9854 550338
rect 9234 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 9854 514894
rect 9234 514574 9854 514658
rect 9234 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 9854 514574
rect 9234 478894 9854 514338
rect 9234 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 9854 478894
rect 9234 478574 9854 478658
rect 9234 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 9854 478574
rect 9234 442894 9854 478338
rect 9234 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 9854 442894
rect 9234 442574 9854 442658
rect 9234 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 9854 442574
rect 9234 406894 9854 442338
rect 9234 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 9854 406894
rect 9234 406574 9854 406658
rect 9234 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 9854 406574
rect 9234 370894 9854 406338
rect 9234 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 9854 370894
rect 9234 370574 9854 370658
rect 9234 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 9854 370574
rect 9234 334894 9854 370338
rect 9234 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 9854 334894
rect 9234 334574 9854 334658
rect 9234 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 9854 334574
rect 9234 298894 9854 334338
rect 9234 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 9854 298894
rect 9234 298574 9854 298658
rect 9234 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 9854 298574
rect 9234 262894 9854 298338
rect 9234 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 9854 262894
rect 9234 262574 9854 262658
rect 9234 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 9854 262574
rect 9234 226894 9854 262338
rect 9234 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 9854 226894
rect 9234 226574 9854 226658
rect 9234 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 9854 226574
rect 9234 190894 9854 226338
rect 9234 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 9854 190894
rect 9234 190574 9854 190658
rect 9234 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 9854 190574
rect 9234 154894 9854 190338
rect 9234 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 9854 154894
rect 9234 154574 9854 154658
rect 9234 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 9854 154574
rect 9234 118894 9854 154338
rect 9234 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 9854 118894
rect 9234 118574 9854 118658
rect 9234 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 9854 118574
rect 9234 82894 9854 118338
rect 9234 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 9854 82894
rect 9234 82574 9854 82658
rect 9234 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 9854 82574
rect 9234 46894 9854 82338
rect 9234 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 9854 46894
rect 9234 46574 9854 46658
rect 9234 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 9854 46574
rect 9234 10894 9854 46338
rect 9234 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 9854 10894
rect 9234 10574 9854 10658
rect 9234 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 9854 10574
rect 9234 -2266 9854 10338
rect 9234 -2502 9266 -2266
rect 9502 -2502 9586 -2266
rect 9822 -2502 9854 -2266
rect 9234 -2586 9854 -2502
rect 9234 -2822 9266 -2586
rect 9502 -2822 9586 -2586
rect 9822 -2822 9854 -2586
rect 9234 -7654 9854 -2822
rect 12954 707718 13574 711590
rect 12954 707482 12986 707718
rect 13222 707482 13306 707718
rect 13542 707482 13574 707718
rect 12954 707398 13574 707482
rect 12954 707162 12986 707398
rect 13222 707162 13306 707398
rect 13542 707162 13574 707398
rect 12954 698614 13574 707162
rect 12954 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 13574 698614
rect 12954 698294 13574 698378
rect 12954 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 13574 698294
rect 12954 662614 13574 698058
rect 12954 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 13574 662614
rect 12954 662294 13574 662378
rect 12954 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 13574 662294
rect 12954 626614 13574 662058
rect 12954 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 13574 626614
rect 12954 626294 13574 626378
rect 12954 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 13574 626294
rect 12954 590614 13574 626058
rect 12954 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 13574 590614
rect 12954 590294 13574 590378
rect 12954 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 13574 590294
rect 12954 554614 13574 590058
rect 12954 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 13574 554614
rect 12954 554294 13574 554378
rect 12954 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 13574 554294
rect 12954 518614 13574 554058
rect 12954 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 13574 518614
rect 12954 518294 13574 518378
rect 12954 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 13574 518294
rect 12954 482614 13574 518058
rect 12954 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 13574 482614
rect 12954 482294 13574 482378
rect 12954 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 13574 482294
rect 12954 446614 13574 482058
rect 12954 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 13574 446614
rect 12954 446294 13574 446378
rect 12954 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 13574 446294
rect 12954 410614 13574 446058
rect 12954 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 13574 410614
rect 12954 410294 13574 410378
rect 12954 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 13574 410294
rect 12954 374614 13574 410058
rect 12954 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 13574 374614
rect 12954 374294 13574 374378
rect 12954 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 13574 374294
rect 12954 338614 13574 374058
rect 12954 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 13574 338614
rect 12954 338294 13574 338378
rect 12954 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 13574 338294
rect 12954 302614 13574 338058
rect 12954 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 13574 302614
rect 12954 302294 13574 302378
rect 12954 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 13574 302294
rect 12954 266614 13574 302058
rect 12954 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 13574 266614
rect 12954 266294 13574 266378
rect 12954 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 13574 266294
rect 12954 230614 13574 266058
rect 12954 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 13574 230614
rect 12954 230294 13574 230378
rect 12954 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 13574 230294
rect 12954 194614 13574 230058
rect 12954 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 13574 194614
rect 12954 194294 13574 194378
rect 12954 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 13574 194294
rect 12954 158614 13574 194058
rect 12954 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 13574 158614
rect 12954 158294 13574 158378
rect 12954 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 13574 158294
rect 12954 122614 13574 158058
rect 12954 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 13574 122614
rect 12954 122294 13574 122378
rect 12954 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 13574 122294
rect 12954 86614 13574 122058
rect 12954 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 13574 86614
rect 12954 86294 13574 86378
rect 12954 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 13574 86294
rect 12954 50614 13574 86058
rect 12954 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 13574 50614
rect 12954 50294 13574 50378
rect 12954 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 13574 50294
rect 12954 14614 13574 50058
rect 12954 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 13574 14614
rect 12954 14294 13574 14378
rect 12954 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 13574 14294
rect 12954 -3226 13574 14058
rect 12954 -3462 12986 -3226
rect 13222 -3462 13306 -3226
rect 13542 -3462 13574 -3226
rect 12954 -3546 13574 -3462
rect 12954 -3782 12986 -3546
rect 13222 -3782 13306 -3546
rect 13542 -3782 13574 -3546
rect 12954 -7654 13574 -3782
rect 16674 708678 17294 711590
rect 16674 708442 16706 708678
rect 16942 708442 17026 708678
rect 17262 708442 17294 708678
rect 16674 708358 17294 708442
rect 16674 708122 16706 708358
rect 16942 708122 17026 708358
rect 17262 708122 17294 708358
rect 16674 666334 17294 708122
rect 16674 666098 16706 666334
rect 16942 666098 17026 666334
rect 17262 666098 17294 666334
rect 16674 666014 17294 666098
rect 16674 665778 16706 666014
rect 16942 665778 17026 666014
rect 17262 665778 17294 666014
rect 16674 630334 17294 665778
rect 16674 630098 16706 630334
rect 16942 630098 17026 630334
rect 17262 630098 17294 630334
rect 16674 630014 17294 630098
rect 16674 629778 16706 630014
rect 16942 629778 17026 630014
rect 17262 629778 17294 630014
rect 16674 594334 17294 629778
rect 16674 594098 16706 594334
rect 16942 594098 17026 594334
rect 17262 594098 17294 594334
rect 16674 594014 17294 594098
rect 16674 593778 16706 594014
rect 16942 593778 17026 594014
rect 17262 593778 17294 594014
rect 16674 558334 17294 593778
rect 16674 558098 16706 558334
rect 16942 558098 17026 558334
rect 17262 558098 17294 558334
rect 16674 558014 17294 558098
rect 16674 557778 16706 558014
rect 16942 557778 17026 558014
rect 17262 557778 17294 558014
rect 16674 522334 17294 557778
rect 16674 522098 16706 522334
rect 16942 522098 17026 522334
rect 17262 522098 17294 522334
rect 16674 522014 17294 522098
rect 16674 521778 16706 522014
rect 16942 521778 17026 522014
rect 17262 521778 17294 522014
rect 16674 486334 17294 521778
rect 16674 486098 16706 486334
rect 16942 486098 17026 486334
rect 17262 486098 17294 486334
rect 16674 486014 17294 486098
rect 16674 485778 16706 486014
rect 16942 485778 17026 486014
rect 17262 485778 17294 486014
rect 16674 450334 17294 485778
rect 16674 450098 16706 450334
rect 16942 450098 17026 450334
rect 17262 450098 17294 450334
rect 16674 450014 17294 450098
rect 16674 449778 16706 450014
rect 16942 449778 17026 450014
rect 17262 449778 17294 450014
rect 16674 414334 17294 449778
rect 16674 414098 16706 414334
rect 16942 414098 17026 414334
rect 17262 414098 17294 414334
rect 16674 414014 17294 414098
rect 16674 413778 16706 414014
rect 16942 413778 17026 414014
rect 17262 413778 17294 414014
rect 16674 378334 17294 413778
rect 16674 378098 16706 378334
rect 16942 378098 17026 378334
rect 17262 378098 17294 378334
rect 16674 378014 17294 378098
rect 16674 377778 16706 378014
rect 16942 377778 17026 378014
rect 17262 377778 17294 378014
rect 16674 342334 17294 377778
rect 16674 342098 16706 342334
rect 16942 342098 17026 342334
rect 17262 342098 17294 342334
rect 16674 342014 17294 342098
rect 16674 341778 16706 342014
rect 16942 341778 17026 342014
rect 17262 341778 17294 342014
rect 16674 306334 17294 341778
rect 16674 306098 16706 306334
rect 16942 306098 17026 306334
rect 17262 306098 17294 306334
rect 16674 306014 17294 306098
rect 16674 305778 16706 306014
rect 16942 305778 17026 306014
rect 17262 305778 17294 306014
rect 16674 270334 17294 305778
rect 16674 270098 16706 270334
rect 16942 270098 17026 270334
rect 17262 270098 17294 270334
rect 16674 270014 17294 270098
rect 16674 269778 16706 270014
rect 16942 269778 17026 270014
rect 17262 269778 17294 270014
rect 16674 234334 17294 269778
rect 16674 234098 16706 234334
rect 16942 234098 17026 234334
rect 17262 234098 17294 234334
rect 16674 234014 17294 234098
rect 16674 233778 16706 234014
rect 16942 233778 17026 234014
rect 17262 233778 17294 234014
rect 16674 198334 17294 233778
rect 16674 198098 16706 198334
rect 16942 198098 17026 198334
rect 17262 198098 17294 198334
rect 16674 198014 17294 198098
rect 16674 197778 16706 198014
rect 16942 197778 17026 198014
rect 17262 197778 17294 198014
rect 16674 162334 17294 197778
rect 16674 162098 16706 162334
rect 16942 162098 17026 162334
rect 17262 162098 17294 162334
rect 16674 162014 17294 162098
rect 16674 161778 16706 162014
rect 16942 161778 17026 162014
rect 17262 161778 17294 162014
rect 16674 126334 17294 161778
rect 16674 126098 16706 126334
rect 16942 126098 17026 126334
rect 17262 126098 17294 126334
rect 16674 126014 17294 126098
rect 16674 125778 16706 126014
rect 16942 125778 17026 126014
rect 17262 125778 17294 126014
rect 16674 90334 17294 125778
rect 16674 90098 16706 90334
rect 16942 90098 17026 90334
rect 17262 90098 17294 90334
rect 16674 90014 17294 90098
rect 16674 89778 16706 90014
rect 16942 89778 17026 90014
rect 17262 89778 17294 90014
rect 16674 54334 17294 89778
rect 16674 54098 16706 54334
rect 16942 54098 17026 54334
rect 17262 54098 17294 54334
rect 16674 54014 17294 54098
rect 16674 53778 16706 54014
rect 16942 53778 17026 54014
rect 17262 53778 17294 54014
rect 16674 18334 17294 53778
rect 16674 18098 16706 18334
rect 16942 18098 17026 18334
rect 17262 18098 17294 18334
rect 16674 18014 17294 18098
rect 16674 17778 16706 18014
rect 16942 17778 17026 18014
rect 17262 17778 17294 18014
rect 16674 -4186 17294 17778
rect 16674 -4422 16706 -4186
rect 16942 -4422 17026 -4186
rect 17262 -4422 17294 -4186
rect 16674 -4506 17294 -4422
rect 16674 -4742 16706 -4506
rect 16942 -4742 17026 -4506
rect 17262 -4742 17294 -4506
rect 16674 -7654 17294 -4742
rect 20394 709638 21014 711590
rect 20394 709402 20426 709638
rect 20662 709402 20746 709638
rect 20982 709402 21014 709638
rect 20394 709318 21014 709402
rect 20394 709082 20426 709318
rect 20662 709082 20746 709318
rect 20982 709082 21014 709318
rect 20394 670054 21014 709082
rect 20394 669818 20426 670054
rect 20662 669818 20746 670054
rect 20982 669818 21014 670054
rect 20394 669734 21014 669818
rect 20394 669498 20426 669734
rect 20662 669498 20746 669734
rect 20982 669498 21014 669734
rect 20394 634054 21014 669498
rect 27834 711558 28454 711590
rect 27834 711322 27866 711558
rect 28102 711322 28186 711558
rect 28422 711322 28454 711558
rect 27834 711238 28454 711322
rect 27834 711002 27866 711238
rect 28102 711002 28186 711238
rect 28422 711002 28454 711238
rect 27834 677494 28454 711002
rect 27834 677258 27866 677494
rect 28102 677258 28186 677494
rect 28422 677258 28454 677494
rect 27834 677174 28454 677258
rect 27834 676938 27866 677174
rect 28102 676938 28186 677174
rect 28422 676938 28454 677174
rect 24208 651454 24528 651486
rect 24208 651218 24250 651454
rect 24486 651218 24528 651454
rect 24208 651134 24528 651218
rect 24208 650898 24250 651134
rect 24486 650898 24528 651134
rect 24208 650866 24528 650898
rect 20394 633818 20426 634054
rect 20662 633818 20746 634054
rect 20982 633818 21014 634054
rect 20394 633734 21014 633818
rect 20394 633498 20426 633734
rect 20662 633498 20746 633734
rect 20982 633498 21014 633734
rect 20394 598054 21014 633498
rect 27834 641494 28454 676938
rect 37794 704838 38414 711590
rect 37794 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 38414 704838
rect 37794 704518 38414 704602
rect 37794 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 38414 704518
rect 37794 687454 38414 704282
rect 37794 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 38414 687454
rect 37794 687134 38414 687218
rect 37794 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 38414 687134
rect 37794 674393 38414 686898
rect 41514 705798 42134 711590
rect 41514 705562 41546 705798
rect 41782 705562 41866 705798
rect 42102 705562 42134 705798
rect 41514 705478 42134 705562
rect 41514 705242 41546 705478
rect 41782 705242 41866 705478
rect 42102 705242 42134 705478
rect 41514 691174 42134 705242
rect 41514 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 42134 691174
rect 41514 690854 42134 690938
rect 41514 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 42134 690854
rect 41514 674393 42134 690618
rect 45234 706758 45854 711590
rect 45234 706522 45266 706758
rect 45502 706522 45586 706758
rect 45822 706522 45854 706758
rect 45234 706438 45854 706522
rect 45234 706202 45266 706438
rect 45502 706202 45586 706438
rect 45822 706202 45854 706438
rect 45234 694894 45854 706202
rect 45234 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 45854 694894
rect 45234 694574 45854 694658
rect 45234 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 45854 694574
rect 45234 674393 45854 694338
rect 48954 707718 49574 711590
rect 48954 707482 48986 707718
rect 49222 707482 49306 707718
rect 49542 707482 49574 707718
rect 48954 707398 49574 707482
rect 48954 707162 48986 707398
rect 49222 707162 49306 707398
rect 49542 707162 49574 707398
rect 48954 698614 49574 707162
rect 48954 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 49574 698614
rect 48954 698294 49574 698378
rect 48954 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 49574 698294
rect 48954 674393 49574 698058
rect 63834 711558 64454 711590
rect 63834 711322 63866 711558
rect 64102 711322 64186 711558
rect 64422 711322 64454 711558
rect 63834 711238 64454 711322
rect 63834 711002 63866 711238
rect 64102 711002 64186 711238
rect 64422 711002 64454 711238
rect 63834 677494 64454 711002
rect 63834 677258 63866 677494
rect 64102 677258 64186 677494
rect 64422 677258 64454 677494
rect 63834 677174 64454 677258
rect 63834 676938 63866 677174
rect 64102 676938 64186 677174
rect 64422 676938 64454 677174
rect 63834 674393 64454 676938
rect 73794 704838 74414 711590
rect 73794 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 74414 704838
rect 73794 704518 74414 704602
rect 73794 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 74414 704518
rect 73794 687454 74414 704282
rect 73794 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 74414 687454
rect 73794 687134 74414 687218
rect 73794 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 74414 687134
rect 73794 674393 74414 686898
rect 77514 705798 78134 711590
rect 77514 705562 77546 705798
rect 77782 705562 77866 705798
rect 78102 705562 78134 705798
rect 77514 705478 78134 705562
rect 77514 705242 77546 705478
rect 77782 705242 77866 705478
rect 78102 705242 78134 705478
rect 77514 691174 78134 705242
rect 77514 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 78134 691174
rect 77514 690854 78134 690938
rect 77514 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 78134 690854
rect 77514 674393 78134 690618
rect 81234 706758 81854 711590
rect 81234 706522 81266 706758
rect 81502 706522 81586 706758
rect 81822 706522 81854 706758
rect 81234 706438 81854 706522
rect 81234 706202 81266 706438
rect 81502 706202 81586 706438
rect 81822 706202 81854 706438
rect 81234 694894 81854 706202
rect 81234 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 81854 694894
rect 81234 694574 81854 694658
rect 81234 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 81854 694574
rect 81234 674393 81854 694338
rect 84954 707718 85574 711590
rect 84954 707482 84986 707718
rect 85222 707482 85306 707718
rect 85542 707482 85574 707718
rect 84954 707398 85574 707482
rect 84954 707162 84986 707398
rect 85222 707162 85306 707398
rect 85542 707162 85574 707398
rect 84954 698614 85574 707162
rect 84954 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 85574 698614
rect 84954 698294 85574 698378
rect 84954 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 85574 698294
rect 84954 674393 85574 698058
rect 99834 711558 100454 711590
rect 99834 711322 99866 711558
rect 100102 711322 100186 711558
rect 100422 711322 100454 711558
rect 99834 711238 100454 711322
rect 99834 711002 99866 711238
rect 100102 711002 100186 711238
rect 100422 711002 100454 711238
rect 99834 677494 100454 711002
rect 99834 677258 99866 677494
rect 100102 677258 100186 677494
rect 100422 677258 100454 677494
rect 99834 677174 100454 677258
rect 99834 676938 99866 677174
rect 100102 676938 100186 677174
rect 100422 676938 100454 677174
rect 99834 674393 100454 676938
rect 109794 704838 110414 711590
rect 109794 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 110414 704838
rect 109794 704518 110414 704602
rect 109794 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 110414 704518
rect 109794 687454 110414 704282
rect 109794 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 110414 687454
rect 109794 687134 110414 687218
rect 109794 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 110414 687134
rect 109794 674393 110414 686898
rect 113514 705798 114134 711590
rect 113514 705562 113546 705798
rect 113782 705562 113866 705798
rect 114102 705562 114134 705798
rect 113514 705478 114134 705562
rect 113514 705242 113546 705478
rect 113782 705242 113866 705478
rect 114102 705242 114134 705478
rect 113514 691174 114134 705242
rect 113514 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 114134 691174
rect 113514 690854 114134 690938
rect 113514 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 114134 690854
rect 113514 674393 114134 690618
rect 117234 706758 117854 711590
rect 117234 706522 117266 706758
rect 117502 706522 117586 706758
rect 117822 706522 117854 706758
rect 117234 706438 117854 706522
rect 117234 706202 117266 706438
rect 117502 706202 117586 706438
rect 117822 706202 117854 706438
rect 117234 694894 117854 706202
rect 117234 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 117854 694894
rect 117234 694574 117854 694658
rect 117234 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 117854 694574
rect 117234 674393 117854 694338
rect 120954 707718 121574 711590
rect 120954 707482 120986 707718
rect 121222 707482 121306 707718
rect 121542 707482 121574 707718
rect 120954 707398 121574 707482
rect 120954 707162 120986 707398
rect 121222 707162 121306 707398
rect 121542 707162 121574 707398
rect 120954 698614 121574 707162
rect 120954 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 121574 698614
rect 120954 698294 121574 698378
rect 120954 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 121574 698294
rect 120954 674393 121574 698058
rect 135834 711558 136454 711590
rect 135834 711322 135866 711558
rect 136102 711322 136186 711558
rect 136422 711322 136454 711558
rect 135834 711238 136454 711322
rect 135834 711002 135866 711238
rect 136102 711002 136186 711238
rect 136422 711002 136454 711238
rect 135834 677494 136454 711002
rect 135834 677258 135866 677494
rect 136102 677258 136186 677494
rect 136422 677258 136454 677494
rect 135834 677174 136454 677258
rect 135834 676938 135866 677174
rect 136102 676938 136186 677174
rect 136422 676938 136454 677174
rect 135834 674393 136454 676938
rect 145794 704838 146414 711590
rect 145794 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 146414 704838
rect 145794 704518 146414 704602
rect 145794 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 146414 704518
rect 145794 687454 146414 704282
rect 145794 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 146414 687454
rect 145794 687134 146414 687218
rect 145794 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 146414 687134
rect 145794 674393 146414 686898
rect 149514 705798 150134 711590
rect 149514 705562 149546 705798
rect 149782 705562 149866 705798
rect 150102 705562 150134 705798
rect 149514 705478 150134 705562
rect 149514 705242 149546 705478
rect 149782 705242 149866 705478
rect 150102 705242 150134 705478
rect 149514 691174 150134 705242
rect 149514 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 150134 691174
rect 149514 690854 150134 690938
rect 149514 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 150134 690854
rect 149514 674393 150134 690618
rect 153234 706758 153854 711590
rect 153234 706522 153266 706758
rect 153502 706522 153586 706758
rect 153822 706522 153854 706758
rect 153234 706438 153854 706522
rect 153234 706202 153266 706438
rect 153502 706202 153586 706438
rect 153822 706202 153854 706438
rect 153234 694894 153854 706202
rect 153234 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 153854 694894
rect 153234 694574 153854 694658
rect 153234 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 153854 694574
rect 153234 674393 153854 694338
rect 156954 707718 157574 711590
rect 156954 707482 156986 707718
rect 157222 707482 157306 707718
rect 157542 707482 157574 707718
rect 156954 707398 157574 707482
rect 156954 707162 156986 707398
rect 157222 707162 157306 707398
rect 157542 707162 157574 707398
rect 156954 698614 157574 707162
rect 156954 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 157574 698614
rect 156954 698294 157574 698378
rect 156954 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 157574 698294
rect 156954 674393 157574 698058
rect 171834 711558 172454 711590
rect 171834 711322 171866 711558
rect 172102 711322 172186 711558
rect 172422 711322 172454 711558
rect 171834 711238 172454 711322
rect 171834 711002 171866 711238
rect 172102 711002 172186 711238
rect 172422 711002 172454 711238
rect 171834 677494 172454 711002
rect 171834 677258 171866 677494
rect 172102 677258 172186 677494
rect 172422 677258 172454 677494
rect 171834 677174 172454 677258
rect 171834 676938 171866 677174
rect 172102 676938 172186 677174
rect 172422 676938 172454 677174
rect 171834 674393 172454 676938
rect 181794 704838 182414 711590
rect 181794 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 182414 704838
rect 181794 704518 182414 704602
rect 181794 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 182414 704518
rect 181794 687454 182414 704282
rect 181794 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 182414 687454
rect 181794 687134 182414 687218
rect 181794 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 182414 687134
rect 181794 674393 182414 686898
rect 185514 705798 186134 711590
rect 185514 705562 185546 705798
rect 185782 705562 185866 705798
rect 186102 705562 186134 705798
rect 185514 705478 186134 705562
rect 185514 705242 185546 705478
rect 185782 705242 185866 705478
rect 186102 705242 186134 705478
rect 185514 691174 186134 705242
rect 185514 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 186134 691174
rect 185514 690854 186134 690938
rect 185514 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 186134 690854
rect 185514 674393 186134 690618
rect 189234 706758 189854 711590
rect 189234 706522 189266 706758
rect 189502 706522 189586 706758
rect 189822 706522 189854 706758
rect 189234 706438 189854 706522
rect 189234 706202 189266 706438
rect 189502 706202 189586 706438
rect 189822 706202 189854 706438
rect 189234 694894 189854 706202
rect 189234 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 189854 694894
rect 189234 694574 189854 694658
rect 189234 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 189854 694574
rect 189234 674393 189854 694338
rect 192954 707718 193574 711590
rect 192954 707482 192986 707718
rect 193222 707482 193306 707718
rect 193542 707482 193574 707718
rect 192954 707398 193574 707482
rect 192954 707162 192986 707398
rect 193222 707162 193306 707398
rect 193542 707162 193574 707398
rect 192954 698614 193574 707162
rect 192954 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 193574 698614
rect 192954 698294 193574 698378
rect 192954 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 193574 698294
rect 192954 684676 193574 698058
rect 207834 711558 208454 711590
rect 207834 711322 207866 711558
rect 208102 711322 208186 711558
rect 208422 711322 208454 711558
rect 207834 711238 208454 711322
rect 207834 711002 207866 711238
rect 208102 711002 208186 711238
rect 208422 711002 208454 711238
rect 207834 677494 208454 711002
rect 207834 677258 207866 677494
rect 208102 677258 208186 677494
rect 208422 677258 208454 677494
rect 207834 677174 208454 677258
rect 207834 676938 207866 677174
rect 208102 676938 208186 677174
rect 208422 676938 208454 677174
rect 207834 674393 208454 676938
rect 217794 704838 218414 711590
rect 217794 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 218414 704838
rect 217794 704518 218414 704602
rect 217794 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 218414 704518
rect 217794 687454 218414 704282
rect 217794 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 218414 687454
rect 217794 687134 218414 687218
rect 217794 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 218414 687134
rect 217794 674393 218414 686898
rect 221514 705798 222134 711590
rect 221514 705562 221546 705798
rect 221782 705562 221866 705798
rect 222102 705562 222134 705798
rect 221514 705478 222134 705562
rect 221514 705242 221546 705478
rect 221782 705242 221866 705478
rect 222102 705242 222134 705478
rect 221514 691174 222134 705242
rect 221514 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 222134 691174
rect 221514 690854 222134 690938
rect 221514 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 222134 690854
rect 221514 674393 222134 690618
rect 225234 706758 225854 711590
rect 225234 706522 225266 706758
rect 225502 706522 225586 706758
rect 225822 706522 225854 706758
rect 225234 706438 225854 706522
rect 225234 706202 225266 706438
rect 225502 706202 225586 706438
rect 225822 706202 225854 706438
rect 225234 694894 225854 706202
rect 225234 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 225854 694894
rect 225234 694574 225854 694658
rect 225234 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 225854 694574
rect 225234 674393 225854 694338
rect 228954 707718 229574 711590
rect 228954 707482 228986 707718
rect 229222 707482 229306 707718
rect 229542 707482 229574 707718
rect 228954 707398 229574 707482
rect 228954 707162 228986 707398
rect 229222 707162 229306 707398
rect 229542 707162 229574 707398
rect 228954 698614 229574 707162
rect 228954 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 229574 698614
rect 228954 698294 229574 698378
rect 228954 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 229574 698294
rect 228954 674393 229574 698058
rect 243834 711558 244454 711590
rect 243834 711322 243866 711558
rect 244102 711322 244186 711558
rect 244422 711322 244454 711558
rect 243834 711238 244454 711322
rect 243834 711002 243866 711238
rect 244102 711002 244186 711238
rect 244422 711002 244454 711238
rect 243834 677494 244454 711002
rect 243834 677258 243866 677494
rect 244102 677258 244186 677494
rect 244422 677258 244454 677494
rect 243834 677174 244454 677258
rect 243834 676938 243866 677174
rect 244102 676938 244186 677174
rect 244422 676938 244454 677174
rect 243834 674393 244454 676938
rect 253794 704838 254414 711590
rect 253794 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 254414 704838
rect 253794 704518 254414 704602
rect 253794 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 254414 704518
rect 253794 687454 254414 704282
rect 253794 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 254414 687454
rect 253794 687134 254414 687218
rect 253794 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 254414 687134
rect 253794 674393 254414 686898
rect 257514 705798 258134 711590
rect 257514 705562 257546 705798
rect 257782 705562 257866 705798
rect 258102 705562 258134 705798
rect 257514 705478 258134 705562
rect 257514 705242 257546 705478
rect 257782 705242 257866 705478
rect 258102 705242 258134 705478
rect 257514 691174 258134 705242
rect 257514 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 258134 691174
rect 257514 690854 258134 690938
rect 257514 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 258134 690854
rect 257514 674393 258134 690618
rect 261234 706758 261854 711590
rect 261234 706522 261266 706758
rect 261502 706522 261586 706758
rect 261822 706522 261854 706758
rect 261234 706438 261854 706522
rect 261234 706202 261266 706438
rect 261502 706202 261586 706438
rect 261822 706202 261854 706438
rect 261234 694894 261854 706202
rect 261234 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 261854 694894
rect 261234 694574 261854 694658
rect 261234 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 261854 694574
rect 261234 674393 261854 694338
rect 264954 707718 265574 711590
rect 264954 707482 264986 707718
rect 265222 707482 265306 707718
rect 265542 707482 265574 707718
rect 264954 707398 265574 707482
rect 264954 707162 264986 707398
rect 265222 707162 265306 707398
rect 265542 707162 265574 707398
rect 264954 698614 265574 707162
rect 264954 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 265574 698614
rect 264954 698294 265574 698378
rect 264954 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 265574 698294
rect 264954 674393 265574 698058
rect 279834 711558 280454 711590
rect 279834 711322 279866 711558
rect 280102 711322 280186 711558
rect 280422 711322 280454 711558
rect 279834 711238 280454 711322
rect 279834 711002 279866 711238
rect 280102 711002 280186 711238
rect 280422 711002 280454 711238
rect 279834 677494 280454 711002
rect 279834 677258 279866 677494
rect 280102 677258 280186 677494
rect 280422 677258 280454 677494
rect 279834 677174 280454 677258
rect 279834 676938 279866 677174
rect 280102 676938 280186 677174
rect 280422 676938 280454 677174
rect 279834 674393 280454 676938
rect 289794 704838 290414 711590
rect 289794 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 290414 704838
rect 289794 704518 290414 704602
rect 289794 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 290414 704518
rect 289794 687454 290414 704282
rect 289794 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 290414 687454
rect 289794 687134 290414 687218
rect 289794 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 290414 687134
rect 289794 674393 290414 686898
rect 293514 705798 294134 711590
rect 293514 705562 293546 705798
rect 293782 705562 293866 705798
rect 294102 705562 294134 705798
rect 293514 705478 294134 705562
rect 293514 705242 293546 705478
rect 293782 705242 293866 705478
rect 294102 705242 294134 705478
rect 293514 691174 294134 705242
rect 293514 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 294134 691174
rect 293514 690854 294134 690938
rect 293514 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 294134 690854
rect 293514 674393 294134 690618
rect 297234 706758 297854 711590
rect 297234 706522 297266 706758
rect 297502 706522 297586 706758
rect 297822 706522 297854 706758
rect 297234 706438 297854 706522
rect 297234 706202 297266 706438
rect 297502 706202 297586 706438
rect 297822 706202 297854 706438
rect 297234 694894 297854 706202
rect 297234 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 297854 694894
rect 297234 694574 297854 694658
rect 297234 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 297854 694574
rect 297234 674393 297854 694338
rect 300954 707718 301574 711590
rect 300954 707482 300986 707718
rect 301222 707482 301306 707718
rect 301542 707482 301574 707718
rect 300954 707398 301574 707482
rect 300954 707162 300986 707398
rect 301222 707162 301306 707398
rect 301542 707162 301574 707398
rect 300954 698614 301574 707162
rect 300954 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 301574 698614
rect 300954 698294 301574 698378
rect 300954 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 301574 698294
rect 300954 684676 301574 698058
rect 325794 704838 326414 711590
rect 325794 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 326414 704838
rect 325794 704518 326414 704602
rect 325794 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 326414 704518
rect 325794 687454 326414 704282
rect 325794 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 326414 687454
rect 325794 687134 326414 687218
rect 325794 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 326414 687134
rect 325794 674393 326414 686898
rect 329514 705798 330134 711590
rect 329514 705562 329546 705798
rect 329782 705562 329866 705798
rect 330102 705562 330134 705798
rect 329514 705478 330134 705562
rect 329514 705242 329546 705478
rect 329782 705242 329866 705478
rect 330102 705242 330134 705478
rect 329514 691174 330134 705242
rect 329514 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 330134 691174
rect 329514 690854 330134 690938
rect 329514 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 330134 690854
rect 329514 674393 330134 690618
rect 333234 706758 333854 711590
rect 333234 706522 333266 706758
rect 333502 706522 333586 706758
rect 333822 706522 333854 706758
rect 333234 706438 333854 706522
rect 333234 706202 333266 706438
rect 333502 706202 333586 706438
rect 333822 706202 333854 706438
rect 333234 694894 333854 706202
rect 333234 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 333854 694894
rect 333234 694574 333854 694658
rect 333234 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 333854 694574
rect 333234 674393 333854 694338
rect 336954 707718 337574 711590
rect 336954 707482 336986 707718
rect 337222 707482 337306 707718
rect 337542 707482 337574 707718
rect 336954 707398 337574 707482
rect 336954 707162 336986 707398
rect 337222 707162 337306 707398
rect 337542 707162 337574 707398
rect 336954 698614 337574 707162
rect 336954 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 337574 698614
rect 336954 698294 337574 698378
rect 336954 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 337574 698294
rect 336954 674393 337574 698058
rect 351834 711558 352454 711590
rect 351834 711322 351866 711558
rect 352102 711322 352186 711558
rect 352422 711322 352454 711558
rect 351834 711238 352454 711322
rect 351834 711002 351866 711238
rect 352102 711002 352186 711238
rect 352422 711002 352454 711238
rect 351834 677494 352454 711002
rect 351834 677258 351866 677494
rect 352102 677258 352186 677494
rect 352422 677258 352454 677494
rect 351834 677174 352454 677258
rect 351834 676938 351866 677174
rect 352102 676938 352186 677174
rect 352422 676938 352454 677174
rect 351834 674393 352454 676938
rect 361794 704838 362414 711590
rect 361794 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 362414 704838
rect 361794 704518 362414 704602
rect 361794 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 362414 704518
rect 361794 687454 362414 704282
rect 361794 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 362414 687454
rect 361794 687134 362414 687218
rect 361794 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 362414 687134
rect 39568 655174 39888 655206
rect 39568 654938 39610 655174
rect 39846 654938 39888 655174
rect 39568 654854 39888 654938
rect 39568 654618 39610 654854
rect 39846 654618 39888 654854
rect 39568 654586 39888 654618
rect 70288 655174 70608 655206
rect 70288 654938 70330 655174
rect 70566 654938 70608 655174
rect 70288 654854 70608 654938
rect 70288 654618 70330 654854
rect 70566 654618 70608 654854
rect 70288 654586 70608 654618
rect 101008 655174 101328 655206
rect 101008 654938 101050 655174
rect 101286 654938 101328 655174
rect 101008 654854 101328 654938
rect 101008 654618 101050 654854
rect 101286 654618 101328 654854
rect 101008 654586 101328 654618
rect 131728 655174 132048 655206
rect 131728 654938 131770 655174
rect 132006 654938 132048 655174
rect 131728 654854 132048 654938
rect 131728 654618 131770 654854
rect 132006 654618 132048 654854
rect 131728 654586 132048 654618
rect 162448 655174 162768 655206
rect 162448 654938 162490 655174
rect 162726 654938 162768 655174
rect 162448 654854 162768 654938
rect 162448 654618 162490 654854
rect 162726 654618 162768 654854
rect 162448 654586 162768 654618
rect 193168 655174 193488 655206
rect 193168 654938 193210 655174
rect 193446 654938 193488 655174
rect 193168 654854 193488 654938
rect 193168 654618 193210 654854
rect 193446 654618 193488 654854
rect 193168 654586 193488 654618
rect 223888 655174 224208 655206
rect 223888 654938 223930 655174
rect 224166 654938 224208 655174
rect 223888 654854 224208 654938
rect 223888 654618 223930 654854
rect 224166 654618 224208 654854
rect 223888 654586 224208 654618
rect 254608 655174 254928 655206
rect 254608 654938 254650 655174
rect 254886 654938 254928 655174
rect 254608 654854 254928 654938
rect 254608 654618 254650 654854
rect 254886 654618 254928 654854
rect 254608 654586 254928 654618
rect 285328 655174 285648 655206
rect 285328 654938 285370 655174
rect 285606 654938 285648 655174
rect 285328 654854 285648 654938
rect 285328 654618 285370 654854
rect 285606 654618 285648 654854
rect 285328 654586 285648 654618
rect 316048 655174 316368 655206
rect 316048 654938 316090 655174
rect 316326 654938 316368 655174
rect 316048 654854 316368 654938
rect 316048 654618 316090 654854
rect 316326 654618 316368 654854
rect 316048 654586 316368 654618
rect 346768 655174 347088 655206
rect 346768 654938 346810 655174
rect 347046 654938 347088 655174
rect 346768 654854 347088 654938
rect 346768 654618 346810 654854
rect 347046 654618 347088 654854
rect 346768 654586 347088 654618
rect 54928 651454 55248 651486
rect 54928 651218 54970 651454
rect 55206 651218 55248 651454
rect 54928 651134 55248 651218
rect 54928 650898 54970 651134
rect 55206 650898 55248 651134
rect 54928 650866 55248 650898
rect 85648 651454 85968 651486
rect 85648 651218 85690 651454
rect 85926 651218 85968 651454
rect 85648 651134 85968 651218
rect 85648 650898 85690 651134
rect 85926 650898 85968 651134
rect 85648 650866 85968 650898
rect 116368 651454 116688 651486
rect 116368 651218 116410 651454
rect 116646 651218 116688 651454
rect 116368 651134 116688 651218
rect 116368 650898 116410 651134
rect 116646 650898 116688 651134
rect 116368 650866 116688 650898
rect 147088 651454 147408 651486
rect 147088 651218 147130 651454
rect 147366 651218 147408 651454
rect 147088 651134 147408 651218
rect 147088 650898 147130 651134
rect 147366 650898 147408 651134
rect 147088 650866 147408 650898
rect 177808 651454 178128 651486
rect 177808 651218 177850 651454
rect 178086 651218 178128 651454
rect 177808 651134 178128 651218
rect 177808 650898 177850 651134
rect 178086 650898 178128 651134
rect 177808 650866 178128 650898
rect 208528 651454 208848 651486
rect 208528 651218 208570 651454
rect 208806 651218 208848 651454
rect 208528 651134 208848 651218
rect 208528 650898 208570 651134
rect 208806 650898 208848 651134
rect 208528 650866 208848 650898
rect 239248 651454 239568 651486
rect 239248 651218 239290 651454
rect 239526 651218 239568 651454
rect 239248 651134 239568 651218
rect 239248 650898 239290 651134
rect 239526 650898 239568 651134
rect 239248 650866 239568 650898
rect 269968 651454 270288 651486
rect 269968 651218 270010 651454
rect 270246 651218 270288 651454
rect 269968 651134 270288 651218
rect 269968 650898 270010 651134
rect 270246 650898 270288 651134
rect 269968 650866 270288 650898
rect 300688 651454 301008 651486
rect 300688 651218 300730 651454
rect 300966 651218 301008 651454
rect 300688 651134 301008 651218
rect 300688 650898 300730 651134
rect 300966 650898 301008 651134
rect 300688 650866 301008 650898
rect 331408 651454 331728 651486
rect 331408 651218 331450 651454
rect 331686 651218 331728 651454
rect 331408 651134 331728 651218
rect 331408 650898 331450 651134
rect 331686 650898 331728 651134
rect 331408 650866 331728 650898
rect 361794 651454 362414 686898
rect 361794 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 362414 651454
rect 361794 651134 362414 651218
rect 361794 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 362414 651134
rect 27834 641258 27866 641494
rect 28102 641258 28186 641494
rect 28422 641258 28454 641494
rect 27834 641174 28454 641258
rect 27834 640938 27866 641174
rect 28102 640938 28186 641174
rect 28422 640938 28454 641174
rect 24208 615454 24528 615486
rect 24208 615218 24250 615454
rect 24486 615218 24528 615454
rect 24208 615134 24528 615218
rect 24208 614898 24250 615134
rect 24486 614898 24528 615134
rect 24208 614866 24528 614898
rect 20394 597818 20426 598054
rect 20662 597818 20746 598054
rect 20982 597818 21014 598054
rect 20394 597734 21014 597818
rect 20394 597498 20426 597734
rect 20662 597498 20746 597734
rect 20982 597498 21014 597734
rect 20394 562054 21014 597498
rect 27834 605494 28454 640938
rect 39568 619174 39888 619206
rect 39568 618938 39610 619174
rect 39846 618938 39888 619174
rect 39568 618854 39888 618938
rect 39568 618618 39610 618854
rect 39846 618618 39888 618854
rect 39568 618586 39888 618618
rect 70288 619174 70608 619206
rect 70288 618938 70330 619174
rect 70566 618938 70608 619174
rect 70288 618854 70608 618938
rect 70288 618618 70330 618854
rect 70566 618618 70608 618854
rect 70288 618586 70608 618618
rect 101008 619174 101328 619206
rect 101008 618938 101050 619174
rect 101286 618938 101328 619174
rect 101008 618854 101328 618938
rect 101008 618618 101050 618854
rect 101286 618618 101328 618854
rect 101008 618586 101328 618618
rect 131728 619174 132048 619206
rect 131728 618938 131770 619174
rect 132006 618938 132048 619174
rect 131728 618854 132048 618938
rect 131728 618618 131770 618854
rect 132006 618618 132048 618854
rect 131728 618586 132048 618618
rect 162448 619174 162768 619206
rect 162448 618938 162490 619174
rect 162726 618938 162768 619174
rect 162448 618854 162768 618938
rect 162448 618618 162490 618854
rect 162726 618618 162768 618854
rect 162448 618586 162768 618618
rect 193168 619174 193488 619206
rect 193168 618938 193210 619174
rect 193446 618938 193488 619174
rect 193168 618854 193488 618938
rect 193168 618618 193210 618854
rect 193446 618618 193488 618854
rect 193168 618586 193488 618618
rect 223888 619174 224208 619206
rect 223888 618938 223930 619174
rect 224166 618938 224208 619174
rect 223888 618854 224208 618938
rect 223888 618618 223930 618854
rect 224166 618618 224208 618854
rect 223888 618586 224208 618618
rect 254608 619174 254928 619206
rect 254608 618938 254650 619174
rect 254886 618938 254928 619174
rect 254608 618854 254928 618938
rect 254608 618618 254650 618854
rect 254886 618618 254928 618854
rect 254608 618586 254928 618618
rect 285328 619174 285648 619206
rect 285328 618938 285370 619174
rect 285606 618938 285648 619174
rect 285328 618854 285648 618938
rect 285328 618618 285370 618854
rect 285606 618618 285648 618854
rect 285328 618586 285648 618618
rect 316048 619174 316368 619206
rect 316048 618938 316090 619174
rect 316326 618938 316368 619174
rect 316048 618854 316368 618938
rect 316048 618618 316090 618854
rect 316326 618618 316368 618854
rect 316048 618586 316368 618618
rect 346768 619174 347088 619206
rect 346768 618938 346810 619174
rect 347046 618938 347088 619174
rect 346768 618854 347088 618938
rect 346768 618618 346810 618854
rect 347046 618618 347088 618854
rect 346768 618586 347088 618618
rect 54928 615454 55248 615486
rect 54928 615218 54970 615454
rect 55206 615218 55248 615454
rect 54928 615134 55248 615218
rect 54928 614898 54970 615134
rect 55206 614898 55248 615134
rect 54928 614866 55248 614898
rect 85648 615454 85968 615486
rect 85648 615218 85690 615454
rect 85926 615218 85968 615454
rect 85648 615134 85968 615218
rect 85648 614898 85690 615134
rect 85926 614898 85968 615134
rect 85648 614866 85968 614898
rect 116368 615454 116688 615486
rect 116368 615218 116410 615454
rect 116646 615218 116688 615454
rect 116368 615134 116688 615218
rect 116368 614898 116410 615134
rect 116646 614898 116688 615134
rect 116368 614866 116688 614898
rect 147088 615454 147408 615486
rect 147088 615218 147130 615454
rect 147366 615218 147408 615454
rect 147088 615134 147408 615218
rect 147088 614898 147130 615134
rect 147366 614898 147408 615134
rect 147088 614866 147408 614898
rect 177808 615454 178128 615486
rect 177808 615218 177850 615454
rect 178086 615218 178128 615454
rect 177808 615134 178128 615218
rect 177808 614898 177850 615134
rect 178086 614898 178128 615134
rect 177808 614866 178128 614898
rect 208528 615454 208848 615486
rect 208528 615218 208570 615454
rect 208806 615218 208848 615454
rect 208528 615134 208848 615218
rect 208528 614898 208570 615134
rect 208806 614898 208848 615134
rect 208528 614866 208848 614898
rect 239248 615454 239568 615486
rect 239248 615218 239290 615454
rect 239526 615218 239568 615454
rect 239248 615134 239568 615218
rect 239248 614898 239290 615134
rect 239526 614898 239568 615134
rect 239248 614866 239568 614898
rect 269968 615454 270288 615486
rect 269968 615218 270010 615454
rect 270246 615218 270288 615454
rect 269968 615134 270288 615218
rect 269968 614898 270010 615134
rect 270246 614898 270288 615134
rect 269968 614866 270288 614898
rect 300688 615454 301008 615486
rect 300688 615218 300730 615454
rect 300966 615218 301008 615454
rect 300688 615134 301008 615218
rect 300688 614898 300730 615134
rect 300966 614898 301008 615134
rect 300688 614866 301008 614898
rect 331408 615454 331728 615486
rect 331408 615218 331450 615454
rect 331686 615218 331728 615454
rect 331408 615134 331728 615218
rect 331408 614898 331450 615134
rect 331686 614898 331728 615134
rect 331408 614866 331728 614898
rect 361794 615454 362414 650898
rect 361794 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 362414 615454
rect 361794 615134 362414 615218
rect 361794 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 362414 615134
rect 27834 605258 27866 605494
rect 28102 605258 28186 605494
rect 28422 605258 28454 605494
rect 27834 605174 28454 605258
rect 27834 604938 27866 605174
rect 28102 604938 28186 605174
rect 28422 604938 28454 605174
rect 24208 579454 24528 579486
rect 24208 579218 24250 579454
rect 24486 579218 24528 579454
rect 24208 579134 24528 579218
rect 24208 578898 24250 579134
rect 24486 578898 24528 579134
rect 24208 578866 24528 578898
rect 20394 561818 20426 562054
rect 20662 561818 20746 562054
rect 20982 561818 21014 562054
rect 20394 561734 21014 561818
rect 20394 561498 20426 561734
rect 20662 561498 20746 561734
rect 20982 561498 21014 561734
rect 20394 526054 21014 561498
rect 27834 569494 28454 604938
rect 39568 583174 39888 583206
rect 39568 582938 39610 583174
rect 39846 582938 39888 583174
rect 39568 582854 39888 582938
rect 39568 582618 39610 582854
rect 39846 582618 39888 582854
rect 39568 582586 39888 582618
rect 70288 583174 70608 583206
rect 70288 582938 70330 583174
rect 70566 582938 70608 583174
rect 70288 582854 70608 582938
rect 70288 582618 70330 582854
rect 70566 582618 70608 582854
rect 70288 582586 70608 582618
rect 101008 583174 101328 583206
rect 101008 582938 101050 583174
rect 101286 582938 101328 583174
rect 101008 582854 101328 582938
rect 101008 582618 101050 582854
rect 101286 582618 101328 582854
rect 101008 582586 101328 582618
rect 131728 583174 132048 583206
rect 131728 582938 131770 583174
rect 132006 582938 132048 583174
rect 131728 582854 132048 582938
rect 131728 582618 131770 582854
rect 132006 582618 132048 582854
rect 131728 582586 132048 582618
rect 162448 583174 162768 583206
rect 162448 582938 162490 583174
rect 162726 582938 162768 583174
rect 162448 582854 162768 582938
rect 162448 582618 162490 582854
rect 162726 582618 162768 582854
rect 162448 582586 162768 582618
rect 193168 583174 193488 583206
rect 193168 582938 193210 583174
rect 193446 582938 193488 583174
rect 193168 582854 193488 582938
rect 193168 582618 193210 582854
rect 193446 582618 193488 582854
rect 193168 582586 193488 582618
rect 223888 583174 224208 583206
rect 223888 582938 223930 583174
rect 224166 582938 224208 583174
rect 223888 582854 224208 582938
rect 223888 582618 223930 582854
rect 224166 582618 224208 582854
rect 223888 582586 224208 582618
rect 254608 583174 254928 583206
rect 254608 582938 254650 583174
rect 254886 582938 254928 583174
rect 254608 582854 254928 582938
rect 254608 582618 254650 582854
rect 254886 582618 254928 582854
rect 254608 582586 254928 582618
rect 285328 583174 285648 583206
rect 285328 582938 285370 583174
rect 285606 582938 285648 583174
rect 285328 582854 285648 582938
rect 285328 582618 285370 582854
rect 285606 582618 285648 582854
rect 285328 582586 285648 582618
rect 316048 583174 316368 583206
rect 316048 582938 316090 583174
rect 316326 582938 316368 583174
rect 316048 582854 316368 582938
rect 316048 582618 316090 582854
rect 316326 582618 316368 582854
rect 316048 582586 316368 582618
rect 346768 583174 347088 583206
rect 346768 582938 346810 583174
rect 347046 582938 347088 583174
rect 346768 582854 347088 582938
rect 346768 582618 346810 582854
rect 347046 582618 347088 582854
rect 346768 582586 347088 582618
rect 54928 579454 55248 579486
rect 54928 579218 54970 579454
rect 55206 579218 55248 579454
rect 54928 579134 55248 579218
rect 54928 578898 54970 579134
rect 55206 578898 55248 579134
rect 54928 578866 55248 578898
rect 85648 579454 85968 579486
rect 85648 579218 85690 579454
rect 85926 579218 85968 579454
rect 85648 579134 85968 579218
rect 85648 578898 85690 579134
rect 85926 578898 85968 579134
rect 85648 578866 85968 578898
rect 116368 579454 116688 579486
rect 116368 579218 116410 579454
rect 116646 579218 116688 579454
rect 116368 579134 116688 579218
rect 116368 578898 116410 579134
rect 116646 578898 116688 579134
rect 116368 578866 116688 578898
rect 147088 579454 147408 579486
rect 147088 579218 147130 579454
rect 147366 579218 147408 579454
rect 147088 579134 147408 579218
rect 147088 578898 147130 579134
rect 147366 578898 147408 579134
rect 147088 578866 147408 578898
rect 177808 579454 178128 579486
rect 177808 579218 177850 579454
rect 178086 579218 178128 579454
rect 177808 579134 178128 579218
rect 177808 578898 177850 579134
rect 178086 578898 178128 579134
rect 177808 578866 178128 578898
rect 208528 579454 208848 579486
rect 208528 579218 208570 579454
rect 208806 579218 208848 579454
rect 208528 579134 208848 579218
rect 208528 578898 208570 579134
rect 208806 578898 208848 579134
rect 208528 578866 208848 578898
rect 239248 579454 239568 579486
rect 239248 579218 239290 579454
rect 239526 579218 239568 579454
rect 239248 579134 239568 579218
rect 239248 578898 239290 579134
rect 239526 578898 239568 579134
rect 239248 578866 239568 578898
rect 269968 579454 270288 579486
rect 269968 579218 270010 579454
rect 270246 579218 270288 579454
rect 269968 579134 270288 579218
rect 269968 578898 270010 579134
rect 270246 578898 270288 579134
rect 269968 578866 270288 578898
rect 300688 579454 301008 579486
rect 300688 579218 300730 579454
rect 300966 579218 301008 579454
rect 300688 579134 301008 579218
rect 300688 578898 300730 579134
rect 300966 578898 301008 579134
rect 300688 578866 301008 578898
rect 331408 579454 331728 579486
rect 331408 579218 331450 579454
rect 331686 579218 331728 579454
rect 331408 579134 331728 579218
rect 331408 578898 331450 579134
rect 331686 578898 331728 579134
rect 331408 578866 331728 578898
rect 361794 579454 362414 614898
rect 361794 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 362414 579454
rect 361794 579134 362414 579218
rect 361794 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 362414 579134
rect 27834 569258 27866 569494
rect 28102 569258 28186 569494
rect 28422 569258 28454 569494
rect 27834 569174 28454 569258
rect 27834 568938 27866 569174
rect 28102 568938 28186 569174
rect 28422 568938 28454 569174
rect 24208 543454 24528 543486
rect 24208 543218 24250 543454
rect 24486 543218 24528 543454
rect 24208 543134 24528 543218
rect 24208 542898 24250 543134
rect 24486 542898 24528 543134
rect 24208 542866 24528 542898
rect 20394 525818 20426 526054
rect 20662 525818 20746 526054
rect 20982 525818 21014 526054
rect 20394 525734 21014 525818
rect 20394 525498 20426 525734
rect 20662 525498 20746 525734
rect 20982 525498 21014 525734
rect 20394 490054 21014 525498
rect 27834 533494 28454 568938
rect 39568 547174 39888 547206
rect 39568 546938 39610 547174
rect 39846 546938 39888 547174
rect 39568 546854 39888 546938
rect 39568 546618 39610 546854
rect 39846 546618 39888 546854
rect 39568 546586 39888 546618
rect 70288 547174 70608 547206
rect 70288 546938 70330 547174
rect 70566 546938 70608 547174
rect 70288 546854 70608 546938
rect 70288 546618 70330 546854
rect 70566 546618 70608 546854
rect 70288 546586 70608 546618
rect 101008 547174 101328 547206
rect 101008 546938 101050 547174
rect 101286 546938 101328 547174
rect 101008 546854 101328 546938
rect 101008 546618 101050 546854
rect 101286 546618 101328 546854
rect 101008 546586 101328 546618
rect 131728 547174 132048 547206
rect 131728 546938 131770 547174
rect 132006 546938 132048 547174
rect 131728 546854 132048 546938
rect 131728 546618 131770 546854
rect 132006 546618 132048 546854
rect 131728 546586 132048 546618
rect 162448 547174 162768 547206
rect 162448 546938 162490 547174
rect 162726 546938 162768 547174
rect 162448 546854 162768 546938
rect 162448 546618 162490 546854
rect 162726 546618 162768 546854
rect 162448 546586 162768 546618
rect 193168 547174 193488 547206
rect 193168 546938 193210 547174
rect 193446 546938 193488 547174
rect 193168 546854 193488 546938
rect 193168 546618 193210 546854
rect 193446 546618 193488 546854
rect 193168 546586 193488 546618
rect 223888 547174 224208 547206
rect 223888 546938 223930 547174
rect 224166 546938 224208 547174
rect 223888 546854 224208 546938
rect 223888 546618 223930 546854
rect 224166 546618 224208 546854
rect 223888 546586 224208 546618
rect 254608 547174 254928 547206
rect 254608 546938 254650 547174
rect 254886 546938 254928 547174
rect 254608 546854 254928 546938
rect 254608 546618 254650 546854
rect 254886 546618 254928 546854
rect 254608 546586 254928 546618
rect 285328 547174 285648 547206
rect 285328 546938 285370 547174
rect 285606 546938 285648 547174
rect 285328 546854 285648 546938
rect 285328 546618 285370 546854
rect 285606 546618 285648 546854
rect 285328 546586 285648 546618
rect 316048 547174 316368 547206
rect 316048 546938 316090 547174
rect 316326 546938 316368 547174
rect 316048 546854 316368 546938
rect 316048 546618 316090 546854
rect 316326 546618 316368 546854
rect 316048 546586 316368 546618
rect 346768 547174 347088 547206
rect 346768 546938 346810 547174
rect 347046 546938 347088 547174
rect 346768 546854 347088 546938
rect 346768 546618 346810 546854
rect 347046 546618 347088 546854
rect 346768 546586 347088 546618
rect 54928 543454 55248 543486
rect 54928 543218 54970 543454
rect 55206 543218 55248 543454
rect 54928 543134 55248 543218
rect 54928 542898 54970 543134
rect 55206 542898 55248 543134
rect 54928 542866 55248 542898
rect 85648 543454 85968 543486
rect 85648 543218 85690 543454
rect 85926 543218 85968 543454
rect 85648 543134 85968 543218
rect 85648 542898 85690 543134
rect 85926 542898 85968 543134
rect 85648 542866 85968 542898
rect 116368 543454 116688 543486
rect 116368 543218 116410 543454
rect 116646 543218 116688 543454
rect 116368 543134 116688 543218
rect 116368 542898 116410 543134
rect 116646 542898 116688 543134
rect 116368 542866 116688 542898
rect 147088 543454 147408 543486
rect 147088 543218 147130 543454
rect 147366 543218 147408 543454
rect 147088 543134 147408 543218
rect 147088 542898 147130 543134
rect 147366 542898 147408 543134
rect 147088 542866 147408 542898
rect 177808 543454 178128 543486
rect 177808 543218 177850 543454
rect 178086 543218 178128 543454
rect 177808 543134 178128 543218
rect 177808 542898 177850 543134
rect 178086 542898 178128 543134
rect 177808 542866 178128 542898
rect 208528 543454 208848 543486
rect 208528 543218 208570 543454
rect 208806 543218 208848 543454
rect 208528 543134 208848 543218
rect 208528 542898 208570 543134
rect 208806 542898 208848 543134
rect 208528 542866 208848 542898
rect 239248 543454 239568 543486
rect 239248 543218 239290 543454
rect 239526 543218 239568 543454
rect 239248 543134 239568 543218
rect 239248 542898 239290 543134
rect 239526 542898 239568 543134
rect 239248 542866 239568 542898
rect 269968 543454 270288 543486
rect 269968 543218 270010 543454
rect 270246 543218 270288 543454
rect 269968 543134 270288 543218
rect 269968 542898 270010 543134
rect 270246 542898 270288 543134
rect 269968 542866 270288 542898
rect 300688 543454 301008 543486
rect 300688 543218 300730 543454
rect 300966 543218 301008 543454
rect 300688 543134 301008 543218
rect 300688 542898 300730 543134
rect 300966 542898 301008 543134
rect 300688 542866 301008 542898
rect 331408 543454 331728 543486
rect 331408 543218 331450 543454
rect 331686 543218 331728 543454
rect 331408 543134 331728 543218
rect 331408 542898 331450 543134
rect 331686 542898 331728 543134
rect 331408 542866 331728 542898
rect 361794 543454 362414 578898
rect 361794 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 362414 543454
rect 361794 543134 362414 543218
rect 361794 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 362414 543134
rect 27834 533258 27866 533494
rect 28102 533258 28186 533494
rect 28422 533258 28454 533494
rect 27834 533174 28454 533258
rect 27834 532938 27866 533174
rect 28102 532938 28186 533174
rect 28422 532938 28454 533174
rect 24208 507454 24528 507486
rect 24208 507218 24250 507454
rect 24486 507218 24528 507454
rect 24208 507134 24528 507218
rect 24208 506898 24250 507134
rect 24486 506898 24528 507134
rect 24208 506866 24528 506898
rect 20394 489818 20426 490054
rect 20662 489818 20746 490054
rect 20982 489818 21014 490054
rect 20394 489734 21014 489818
rect 20394 489498 20426 489734
rect 20662 489498 20746 489734
rect 20982 489498 21014 489734
rect 20394 454054 21014 489498
rect 27834 497494 28454 532938
rect 39568 511174 39888 511206
rect 39568 510938 39610 511174
rect 39846 510938 39888 511174
rect 39568 510854 39888 510938
rect 39568 510618 39610 510854
rect 39846 510618 39888 510854
rect 39568 510586 39888 510618
rect 70288 511174 70608 511206
rect 70288 510938 70330 511174
rect 70566 510938 70608 511174
rect 70288 510854 70608 510938
rect 70288 510618 70330 510854
rect 70566 510618 70608 510854
rect 70288 510586 70608 510618
rect 101008 511174 101328 511206
rect 101008 510938 101050 511174
rect 101286 510938 101328 511174
rect 101008 510854 101328 510938
rect 101008 510618 101050 510854
rect 101286 510618 101328 510854
rect 101008 510586 101328 510618
rect 131728 511174 132048 511206
rect 131728 510938 131770 511174
rect 132006 510938 132048 511174
rect 131728 510854 132048 510938
rect 131728 510618 131770 510854
rect 132006 510618 132048 510854
rect 131728 510586 132048 510618
rect 162448 511174 162768 511206
rect 162448 510938 162490 511174
rect 162726 510938 162768 511174
rect 162448 510854 162768 510938
rect 162448 510618 162490 510854
rect 162726 510618 162768 510854
rect 162448 510586 162768 510618
rect 193168 511174 193488 511206
rect 193168 510938 193210 511174
rect 193446 510938 193488 511174
rect 193168 510854 193488 510938
rect 193168 510618 193210 510854
rect 193446 510618 193488 510854
rect 193168 510586 193488 510618
rect 223888 511174 224208 511206
rect 223888 510938 223930 511174
rect 224166 510938 224208 511174
rect 223888 510854 224208 510938
rect 223888 510618 223930 510854
rect 224166 510618 224208 510854
rect 223888 510586 224208 510618
rect 254608 511174 254928 511206
rect 254608 510938 254650 511174
rect 254886 510938 254928 511174
rect 254608 510854 254928 510938
rect 254608 510618 254650 510854
rect 254886 510618 254928 510854
rect 254608 510586 254928 510618
rect 285328 511174 285648 511206
rect 285328 510938 285370 511174
rect 285606 510938 285648 511174
rect 285328 510854 285648 510938
rect 285328 510618 285370 510854
rect 285606 510618 285648 510854
rect 285328 510586 285648 510618
rect 316048 511174 316368 511206
rect 316048 510938 316090 511174
rect 316326 510938 316368 511174
rect 316048 510854 316368 510938
rect 316048 510618 316090 510854
rect 316326 510618 316368 510854
rect 316048 510586 316368 510618
rect 346768 511174 347088 511206
rect 346768 510938 346810 511174
rect 347046 510938 347088 511174
rect 346768 510854 347088 510938
rect 346768 510618 346810 510854
rect 347046 510618 347088 510854
rect 346768 510586 347088 510618
rect 54928 507454 55248 507486
rect 54928 507218 54970 507454
rect 55206 507218 55248 507454
rect 54928 507134 55248 507218
rect 54928 506898 54970 507134
rect 55206 506898 55248 507134
rect 54928 506866 55248 506898
rect 85648 507454 85968 507486
rect 85648 507218 85690 507454
rect 85926 507218 85968 507454
rect 85648 507134 85968 507218
rect 85648 506898 85690 507134
rect 85926 506898 85968 507134
rect 85648 506866 85968 506898
rect 116368 507454 116688 507486
rect 116368 507218 116410 507454
rect 116646 507218 116688 507454
rect 116368 507134 116688 507218
rect 116368 506898 116410 507134
rect 116646 506898 116688 507134
rect 116368 506866 116688 506898
rect 147088 507454 147408 507486
rect 147088 507218 147130 507454
rect 147366 507218 147408 507454
rect 147088 507134 147408 507218
rect 147088 506898 147130 507134
rect 147366 506898 147408 507134
rect 147088 506866 147408 506898
rect 177808 507454 178128 507486
rect 177808 507218 177850 507454
rect 178086 507218 178128 507454
rect 177808 507134 178128 507218
rect 177808 506898 177850 507134
rect 178086 506898 178128 507134
rect 177808 506866 178128 506898
rect 208528 507454 208848 507486
rect 208528 507218 208570 507454
rect 208806 507218 208848 507454
rect 208528 507134 208848 507218
rect 208528 506898 208570 507134
rect 208806 506898 208848 507134
rect 208528 506866 208848 506898
rect 239248 507454 239568 507486
rect 239248 507218 239290 507454
rect 239526 507218 239568 507454
rect 239248 507134 239568 507218
rect 239248 506898 239290 507134
rect 239526 506898 239568 507134
rect 239248 506866 239568 506898
rect 269968 507454 270288 507486
rect 269968 507218 270010 507454
rect 270246 507218 270288 507454
rect 269968 507134 270288 507218
rect 269968 506898 270010 507134
rect 270246 506898 270288 507134
rect 269968 506866 270288 506898
rect 300688 507454 301008 507486
rect 300688 507218 300730 507454
rect 300966 507218 301008 507454
rect 300688 507134 301008 507218
rect 300688 506898 300730 507134
rect 300966 506898 301008 507134
rect 300688 506866 301008 506898
rect 331408 507454 331728 507486
rect 331408 507218 331450 507454
rect 331686 507218 331728 507454
rect 331408 507134 331728 507218
rect 331408 506898 331450 507134
rect 331686 506898 331728 507134
rect 331408 506866 331728 506898
rect 361794 507454 362414 542898
rect 361794 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 362414 507454
rect 361794 507134 362414 507218
rect 361794 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 362414 507134
rect 27834 497258 27866 497494
rect 28102 497258 28186 497494
rect 28422 497258 28454 497494
rect 27834 497174 28454 497258
rect 27834 496938 27866 497174
rect 28102 496938 28186 497174
rect 28422 496938 28454 497174
rect 24208 471454 24528 471486
rect 24208 471218 24250 471454
rect 24486 471218 24528 471454
rect 24208 471134 24528 471218
rect 24208 470898 24250 471134
rect 24486 470898 24528 471134
rect 24208 470866 24528 470898
rect 20394 453818 20426 454054
rect 20662 453818 20746 454054
rect 20982 453818 21014 454054
rect 20394 453734 21014 453818
rect 20394 453498 20426 453734
rect 20662 453498 20746 453734
rect 20982 453498 21014 453734
rect 20394 418054 21014 453498
rect 27834 461494 28454 496938
rect 39568 475174 39888 475206
rect 39568 474938 39610 475174
rect 39846 474938 39888 475174
rect 39568 474854 39888 474938
rect 39568 474618 39610 474854
rect 39846 474618 39888 474854
rect 39568 474586 39888 474618
rect 70288 475174 70608 475206
rect 70288 474938 70330 475174
rect 70566 474938 70608 475174
rect 70288 474854 70608 474938
rect 70288 474618 70330 474854
rect 70566 474618 70608 474854
rect 70288 474586 70608 474618
rect 101008 475174 101328 475206
rect 101008 474938 101050 475174
rect 101286 474938 101328 475174
rect 101008 474854 101328 474938
rect 101008 474618 101050 474854
rect 101286 474618 101328 474854
rect 101008 474586 101328 474618
rect 131728 475174 132048 475206
rect 131728 474938 131770 475174
rect 132006 474938 132048 475174
rect 131728 474854 132048 474938
rect 131728 474618 131770 474854
rect 132006 474618 132048 474854
rect 131728 474586 132048 474618
rect 162448 475174 162768 475206
rect 162448 474938 162490 475174
rect 162726 474938 162768 475174
rect 162448 474854 162768 474938
rect 162448 474618 162490 474854
rect 162726 474618 162768 474854
rect 162448 474586 162768 474618
rect 193168 475174 193488 475206
rect 193168 474938 193210 475174
rect 193446 474938 193488 475174
rect 193168 474854 193488 474938
rect 193168 474618 193210 474854
rect 193446 474618 193488 474854
rect 193168 474586 193488 474618
rect 223888 475174 224208 475206
rect 223888 474938 223930 475174
rect 224166 474938 224208 475174
rect 223888 474854 224208 474938
rect 223888 474618 223930 474854
rect 224166 474618 224208 474854
rect 223888 474586 224208 474618
rect 254608 475174 254928 475206
rect 254608 474938 254650 475174
rect 254886 474938 254928 475174
rect 254608 474854 254928 474938
rect 254608 474618 254650 474854
rect 254886 474618 254928 474854
rect 254608 474586 254928 474618
rect 285328 475174 285648 475206
rect 285328 474938 285370 475174
rect 285606 474938 285648 475174
rect 285328 474854 285648 474938
rect 285328 474618 285370 474854
rect 285606 474618 285648 474854
rect 285328 474586 285648 474618
rect 316048 475174 316368 475206
rect 316048 474938 316090 475174
rect 316326 474938 316368 475174
rect 316048 474854 316368 474938
rect 316048 474618 316090 474854
rect 316326 474618 316368 474854
rect 316048 474586 316368 474618
rect 346768 475174 347088 475206
rect 346768 474938 346810 475174
rect 347046 474938 347088 475174
rect 346768 474854 347088 474938
rect 346768 474618 346810 474854
rect 347046 474618 347088 474854
rect 346768 474586 347088 474618
rect 54928 471454 55248 471486
rect 54928 471218 54970 471454
rect 55206 471218 55248 471454
rect 54928 471134 55248 471218
rect 54928 470898 54970 471134
rect 55206 470898 55248 471134
rect 54928 470866 55248 470898
rect 85648 471454 85968 471486
rect 85648 471218 85690 471454
rect 85926 471218 85968 471454
rect 85648 471134 85968 471218
rect 85648 470898 85690 471134
rect 85926 470898 85968 471134
rect 85648 470866 85968 470898
rect 116368 471454 116688 471486
rect 116368 471218 116410 471454
rect 116646 471218 116688 471454
rect 116368 471134 116688 471218
rect 116368 470898 116410 471134
rect 116646 470898 116688 471134
rect 116368 470866 116688 470898
rect 147088 471454 147408 471486
rect 147088 471218 147130 471454
rect 147366 471218 147408 471454
rect 147088 471134 147408 471218
rect 147088 470898 147130 471134
rect 147366 470898 147408 471134
rect 147088 470866 147408 470898
rect 177808 471454 178128 471486
rect 177808 471218 177850 471454
rect 178086 471218 178128 471454
rect 177808 471134 178128 471218
rect 177808 470898 177850 471134
rect 178086 470898 178128 471134
rect 177808 470866 178128 470898
rect 208528 471454 208848 471486
rect 208528 471218 208570 471454
rect 208806 471218 208848 471454
rect 208528 471134 208848 471218
rect 208528 470898 208570 471134
rect 208806 470898 208848 471134
rect 208528 470866 208848 470898
rect 239248 471454 239568 471486
rect 239248 471218 239290 471454
rect 239526 471218 239568 471454
rect 239248 471134 239568 471218
rect 239248 470898 239290 471134
rect 239526 470898 239568 471134
rect 239248 470866 239568 470898
rect 269968 471454 270288 471486
rect 269968 471218 270010 471454
rect 270246 471218 270288 471454
rect 269968 471134 270288 471218
rect 269968 470898 270010 471134
rect 270246 470898 270288 471134
rect 269968 470866 270288 470898
rect 300688 471454 301008 471486
rect 300688 471218 300730 471454
rect 300966 471218 301008 471454
rect 300688 471134 301008 471218
rect 300688 470898 300730 471134
rect 300966 470898 301008 471134
rect 300688 470866 301008 470898
rect 331408 471454 331728 471486
rect 331408 471218 331450 471454
rect 331686 471218 331728 471454
rect 331408 471134 331728 471218
rect 331408 470898 331450 471134
rect 331686 470898 331728 471134
rect 331408 470866 331728 470898
rect 361794 471454 362414 506898
rect 361794 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 362414 471454
rect 361794 471134 362414 471218
rect 361794 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 362414 471134
rect 27834 461258 27866 461494
rect 28102 461258 28186 461494
rect 28422 461258 28454 461494
rect 27834 461174 28454 461258
rect 27834 460938 27866 461174
rect 28102 460938 28186 461174
rect 28422 460938 28454 461174
rect 24208 435454 24528 435486
rect 24208 435218 24250 435454
rect 24486 435218 24528 435454
rect 24208 435134 24528 435218
rect 24208 434898 24250 435134
rect 24486 434898 24528 435134
rect 24208 434866 24528 434898
rect 20394 417818 20426 418054
rect 20662 417818 20746 418054
rect 20982 417818 21014 418054
rect 20394 417734 21014 417818
rect 20394 417498 20426 417734
rect 20662 417498 20746 417734
rect 20982 417498 21014 417734
rect 20394 382054 21014 417498
rect 27834 425494 28454 460938
rect 39568 439174 39888 439206
rect 39568 438938 39610 439174
rect 39846 438938 39888 439174
rect 39568 438854 39888 438938
rect 39568 438618 39610 438854
rect 39846 438618 39888 438854
rect 39568 438586 39888 438618
rect 70288 439174 70608 439206
rect 70288 438938 70330 439174
rect 70566 438938 70608 439174
rect 70288 438854 70608 438938
rect 70288 438618 70330 438854
rect 70566 438618 70608 438854
rect 70288 438586 70608 438618
rect 101008 439174 101328 439206
rect 101008 438938 101050 439174
rect 101286 438938 101328 439174
rect 101008 438854 101328 438938
rect 101008 438618 101050 438854
rect 101286 438618 101328 438854
rect 101008 438586 101328 438618
rect 131728 439174 132048 439206
rect 131728 438938 131770 439174
rect 132006 438938 132048 439174
rect 131728 438854 132048 438938
rect 131728 438618 131770 438854
rect 132006 438618 132048 438854
rect 131728 438586 132048 438618
rect 162448 439174 162768 439206
rect 162448 438938 162490 439174
rect 162726 438938 162768 439174
rect 162448 438854 162768 438938
rect 162448 438618 162490 438854
rect 162726 438618 162768 438854
rect 162448 438586 162768 438618
rect 193168 439174 193488 439206
rect 193168 438938 193210 439174
rect 193446 438938 193488 439174
rect 193168 438854 193488 438938
rect 193168 438618 193210 438854
rect 193446 438618 193488 438854
rect 193168 438586 193488 438618
rect 223888 439174 224208 439206
rect 223888 438938 223930 439174
rect 224166 438938 224208 439174
rect 223888 438854 224208 438938
rect 223888 438618 223930 438854
rect 224166 438618 224208 438854
rect 223888 438586 224208 438618
rect 254608 439174 254928 439206
rect 254608 438938 254650 439174
rect 254886 438938 254928 439174
rect 254608 438854 254928 438938
rect 254608 438618 254650 438854
rect 254886 438618 254928 438854
rect 254608 438586 254928 438618
rect 285328 439174 285648 439206
rect 285328 438938 285370 439174
rect 285606 438938 285648 439174
rect 285328 438854 285648 438938
rect 285328 438618 285370 438854
rect 285606 438618 285648 438854
rect 285328 438586 285648 438618
rect 316048 439174 316368 439206
rect 316048 438938 316090 439174
rect 316326 438938 316368 439174
rect 316048 438854 316368 438938
rect 316048 438618 316090 438854
rect 316326 438618 316368 438854
rect 316048 438586 316368 438618
rect 346768 439174 347088 439206
rect 346768 438938 346810 439174
rect 347046 438938 347088 439174
rect 346768 438854 347088 438938
rect 346768 438618 346810 438854
rect 347046 438618 347088 438854
rect 346768 438586 347088 438618
rect 54928 435454 55248 435486
rect 54928 435218 54970 435454
rect 55206 435218 55248 435454
rect 54928 435134 55248 435218
rect 54928 434898 54970 435134
rect 55206 434898 55248 435134
rect 54928 434866 55248 434898
rect 85648 435454 85968 435486
rect 85648 435218 85690 435454
rect 85926 435218 85968 435454
rect 85648 435134 85968 435218
rect 85648 434898 85690 435134
rect 85926 434898 85968 435134
rect 85648 434866 85968 434898
rect 116368 435454 116688 435486
rect 116368 435218 116410 435454
rect 116646 435218 116688 435454
rect 116368 435134 116688 435218
rect 116368 434898 116410 435134
rect 116646 434898 116688 435134
rect 116368 434866 116688 434898
rect 147088 435454 147408 435486
rect 147088 435218 147130 435454
rect 147366 435218 147408 435454
rect 147088 435134 147408 435218
rect 147088 434898 147130 435134
rect 147366 434898 147408 435134
rect 147088 434866 147408 434898
rect 177808 435454 178128 435486
rect 177808 435218 177850 435454
rect 178086 435218 178128 435454
rect 177808 435134 178128 435218
rect 177808 434898 177850 435134
rect 178086 434898 178128 435134
rect 177808 434866 178128 434898
rect 208528 435454 208848 435486
rect 208528 435218 208570 435454
rect 208806 435218 208848 435454
rect 208528 435134 208848 435218
rect 208528 434898 208570 435134
rect 208806 434898 208848 435134
rect 208528 434866 208848 434898
rect 239248 435454 239568 435486
rect 239248 435218 239290 435454
rect 239526 435218 239568 435454
rect 239248 435134 239568 435218
rect 239248 434898 239290 435134
rect 239526 434898 239568 435134
rect 239248 434866 239568 434898
rect 269968 435454 270288 435486
rect 269968 435218 270010 435454
rect 270246 435218 270288 435454
rect 269968 435134 270288 435218
rect 269968 434898 270010 435134
rect 270246 434898 270288 435134
rect 269968 434866 270288 434898
rect 300688 435454 301008 435486
rect 300688 435218 300730 435454
rect 300966 435218 301008 435454
rect 300688 435134 301008 435218
rect 300688 434898 300730 435134
rect 300966 434898 301008 435134
rect 300688 434866 301008 434898
rect 331408 435454 331728 435486
rect 331408 435218 331450 435454
rect 331686 435218 331728 435454
rect 331408 435134 331728 435218
rect 331408 434898 331450 435134
rect 331686 434898 331728 435134
rect 331408 434866 331728 434898
rect 361794 435454 362414 470898
rect 361794 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 362414 435454
rect 361794 435134 362414 435218
rect 361794 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 362414 435134
rect 27834 425258 27866 425494
rect 28102 425258 28186 425494
rect 28422 425258 28454 425494
rect 27834 425174 28454 425258
rect 27834 424938 27866 425174
rect 28102 424938 28186 425174
rect 28422 424938 28454 425174
rect 24208 399454 24528 399486
rect 24208 399218 24250 399454
rect 24486 399218 24528 399454
rect 24208 399134 24528 399218
rect 24208 398898 24250 399134
rect 24486 398898 24528 399134
rect 24208 398866 24528 398898
rect 20394 381818 20426 382054
rect 20662 381818 20746 382054
rect 20982 381818 21014 382054
rect 20394 381734 21014 381818
rect 20394 381498 20426 381734
rect 20662 381498 20746 381734
rect 20982 381498 21014 381734
rect 20394 346054 21014 381498
rect 27834 389494 28454 424938
rect 39568 403174 39888 403206
rect 39568 402938 39610 403174
rect 39846 402938 39888 403174
rect 39568 402854 39888 402938
rect 39568 402618 39610 402854
rect 39846 402618 39888 402854
rect 39568 402586 39888 402618
rect 70288 403174 70608 403206
rect 70288 402938 70330 403174
rect 70566 402938 70608 403174
rect 70288 402854 70608 402938
rect 70288 402618 70330 402854
rect 70566 402618 70608 402854
rect 70288 402586 70608 402618
rect 101008 403174 101328 403206
rect 101008 402938 101050 403174
rect 101286 402938 101328 403174
rect 101008 402854 101328 402938
rect 101008 402618 101050 402854
rect 101286 402618 101328 402854
rect 101008 402586 101328 402618
rect 131728 403174 132048 403206
rect 131728 402938 131770 403174
rect 132006 402938 132048 403174
rect 131728 402854 132048 402938
rect 131728 402618 131770 402854
rect 132006 402618 132048 402854
rect 131728 402586 132048 402618
rect 162448 403174 162768 403206
rect 162448 402938 162490 403174
rect 162726 402938 162768 403174
rect 162448 402854 162768 402938
rect 162448 402618 162490 402854
rect 162726 402618 162768 402854
rect 162448 402586 162768 402618
rect 193168 403174 193488 403206
rect 193168 402938 193210 403174
rect 193446 402938 193488 403174
rect 193168 402854 193488 402938
rect 193168 402618 193210 402854
rect 193446 402618 193488 402854
rect 193168 402586 193488 402618
rect 223888 403174 224208 403206
rect 223888 402938 223930 403174
rect 224166 402938 224208 403174
rect 223888 402854 224208 402938
rect 223888 402618 223930 402854
rect 224166 402618 224208 402854
rect 223888 402586 224208 402618
rect 254608 403174 254928 403206
rect 254608 402938 254650 403174
rect 254886 402938 254928 403174
rect 254608 402854 254928 402938
rect 254608 402618 254650 402854
rect 254886 402618 254928 402854
rect 254608 402586 254928 402618
rect 285328 403174 285648 403206
rect 285328 402938 285370 403174
rect 285606 402938 285648 403174
rect 285328 402854 285648 402938
rect 285328 402618 285370 402854
rect 285606 402618 285648 402854
rect 285328 402586 285648 402618
rect 316048 403174 316368 403206
rect 316048 402938 316090 403174
rect 316326 402938 316368 403174
rect 316048 402854 316368 402938
rect 316048 402618 316090 402854
rect 316326 402618 316368 402854
rect 316048 402586 316368 402618
rect 346768 403174 347088 403206
rect 346768 402938 346810 403174
rect 347046 402938 347088 403174
rect 346768 402854 347088 402938
rect 346768 402618 346810 402854
rect 347046 402618 347088 402854
rect 346768 402586 347088 402618
rect 54928 399454 55248 399486
rect 54928 399218 54970 399454
rect 55206 399218 55248 399454
rect 54928 399134 55248 399218
rect 54928 398898 54970 399134
rect 55206 398898 55248 399134
rect 54928 398866 55248 398898
rect 85648 399454 85968 399486
rect 85648 399218 85690 399454
rect 85926 399218 85968 399454
rect 85648 399134 85968 399218
rect 85648 398898 85690 399134
rect 85926 398898 85968 399134
rect 85648 398866 85968 398898
rect 116368 399454 116688 399486
rect 116368 399218 116410 399454
rect 116646 399218 116688 399454
rect 116368 399134 116688 399218
rect 116368 398898 116410 399134
rect 116646 398898 116688 399134
rect 116368 398866 116688 398898
rect 147088 399454 147408 399486
rect 147088 399218 147130 399454
rect 147366 399218 147408 399454
rect 147088 399134 147408 399218
rect 147088 398898 147130 399134
rect 147366 398898 147408 399134
rect 147088 398866 147408 398898
rect 177808 399454 178128 399486
rect 177808 399218 177850 399454
rect 178086 399218 178128 399454
rect 177808 399134 178128 399218
rect 177808 398898 177850 399134
rect 178086 398898 178128 399134
rect 177808 398866 178128 398898
rect 208528 399454 208848 399486
rect 208528 399218 208570 399454
rect 208806 399218 208848 399454
rect 208528 399134 208848 399218
rect 208528 398898 208570 399134
rect 208806 398898 208848 399134
rect 208528 398866 208848 398898
rect 239248 399454 239568 399486
rect 239248 399218 239290 399454
rect 239526 399218 239568 399454
rect 239248 399134 239568 399218
rect 239248 398898 239290 399134
rect 239526 398898 239568 399134
rect 239248 398866 239568 398898
rect 269968 399454 270288 399486
rect 269968 399218 270010 399454
rect 270246 399218 270288 399454
rect 269968 399134 270288 399218
rect 269968 398898 270010 399134
rect 270246 398898 270288 399134
rect 269968 398866 270288 398898
rect 300688 399454 301008 399486
rect 300688 399218 300730 399454
rect 300966 399218 301008 399454
rect 300688 399134 301008 399218
rect 300688 398898 300730 399134
rect 300966 398898 301008 399134
rect 300688 398866 301008 398898
rect 331408 399454 331728 399486
rect 331408 399218 331450 399454
rect 331686 399218 331728 399454
rect 331408 399134 331728 399218
rect 331408 398898 331450 399134
rect 331686 398898 331728 399134
rect 331408 398866 331728 398898
rect 361794 399454 362414 434898
rect 361794 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 362414 399454
rect 361794 399134 362414 399218
rect 361794 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 362414 399134
rect 27834 389258 27866 389494
rect 28102 389258 28186 389494
rect 28422 389258 28454 389494
rect 27834 389174 28454 389258
rect 27834 388938 27866 389174
rect 28102 388938 28186 389174
rect 28422 388938 28454 389174
rect 24208 363454 24528 363486
rect 24208 363218 24250 363454
rect 24486 363218 24528 363454
rect 24208 363134 24528 363218
rect 24208 362898 24250 363134
rect 24486 362898 24528 363134
rect 24208 362866 24528 362898
rect 20394 345818 20426 346054
rect 20662 345818 20746 346054
rect 20982 345818 21014 346054
rect 20394 345734 21014 345818
rect 20394 345498 20426 345734
rect 20662 345498 20746 345734
rect 20982 345498 21014 345734
rect 20394 310054 21014 345498
rect 27834 353494 28454 388938
rect 39568 367174 39888 367206
rect 39568 366938 39610 367174
rect 39846 366938 39888 367174
rect 39568 366854 39888 366938
rect 39568 366618 39610 366854
rect 39846 366618 39888 366854
rect 39568 366586 39888 366618
rect 70288 367174 70608 367206
rect 70288 366938 70330 367174
rect 70566 366938 70608 367174
rect 70288 366854 70608 366938
rect 70288 366618 70330 366854
rect 70566 366618 70608 366854
rect 70288 366586 70608 366618
rect 101008 367174 101328 367206
rect 101008 366938 101050 367174
rect 101286 366938 101328 367174
rect 101008 366854 101328 366938
rect 101008 366618 101050 366854
rect 101286 366618 101328 366854
rect 101008 366586 101328 366618
rect 131728 367174 132048 367206
rect 131728 366938 131770 367174
rect 132006 366938 132048 367174
rect 131728 366854 132048 366938
rect 131728 366618 131770 366854
rect 132006 366618 132048 366854
rect 131728 366586 132048 366618
rect 162448 367174 162768 367206
rect 162448 366938 162490 367174
rect 162726 366938 162768 367174
rect 162448 366854 162768 366938
rect 162448 366618 162490 366854
rect 162726 366618 162768 366854
rect 162448 366586 162768 366618
rect 193168 367174 193488 367206
rect 193168 366938 193210 367174
rect 193446 366938 193488 367174
rect 193168 366854 193488 366938
rect 193168 366618 193210 366854
rect 193446 366618 193488 366854
rect 193168 366586 193488 366618
rect 223888 367174 224208 367206
rect 223888 366938 223930 367174
rect 224166 366938 224208 367174
rect 223888 366854 224208 366938
rect 223888 366618 223930 366854
rect 224166 366618 224208 366854
rect 223888 366586 224208 366618
rect 254608 367174 254928 367206
rect 254608 366938 254650 367174
rect 254886 366938 254928 367174
rect 254608 366854 254928 366938
rect 254608 366618 254650 366854
rect 254886 366618 254928 366854
rect 254608 366586 254928 366618
rect 285328 367174 285648 367206
rect 285328 366938 285370 367174
rect 285606 366938 285648 367174
rect 285328 366854 285648 366938
rect 285328 366618 285370 366854
rect 285606 366618 285648 366854
rect 285328 366586 285648 366618
rect 316048 367174 316368 367206
rect 316048 366938 316090 367174
rect 316326 366938 316368 367174
rect 316048 366854 316368 366938
rect 316048 366618 316090 366854
rect 316326 366618 316368 366854
rect 316048 366586 316368 366618
rect 346768 367174 347088 367206
rect 346768 366938 346810 367174
rect 347046 366938 347088 367174
rect 346768 366854 347088 366938
rect 346768 366618 346810 366854
rect 347046 366618 347088 366854
rect 346768 366586 347088 366618
rect 54928 363454 55248 363486
rect 54928 363218 54970 363454
rect 55206 363218 55248 363454
rect 54928 363134 55248 363218
rect 54928 362898 54970 363134
rect 55206 362898 55248 363134
rect 54928 362866 55248 362898
rect 85648 363454 85968 363486
rect 85648 363218 85690 363454
rect 85926 363218 85968 363454
rect 85648 363134 85968 363218
rect 85648 362898 85690 363134
rect 85926 362898 85968 363134
rect 85648 362866 85968 362898
rect 116368 363454 116688 363486
rect 116368 363218 116410 363454
rect 116646 363218 116688 363454
rect 116368 363134 116688 363218
rect 116368 362898 116410 363134
rect 116646 362898 116688 363134
rect 116368 362866 116688 362898
rect 147088 363454 147408 363486
rect 147088 363218 147130 363454
rect 147366 363218 147408 363454
rect 147088 363134 147408 363218
rect 147088 362898 147130 363134
rect 147366 362898 147408 363134
rect 147088 362866 147408 362898
rect 177808 363454 178128 363486
rect 177808 363218 177850 363454
rect 178086 363218 178128 363454
rect 177808 363134 178128 363218
rect 177808 362898 177850 363134
rect 178086 362898 178128 363134
rect 177808 362866 178128 362898
rect 208528 363454 208848 363486
rect 208528 363218 208570 363454
rect 208806 363218 208848 363454
rect 208528 363134 208848 363218
rect 208528 362898 208570 363134
rect 208806 362898 208848 363134
rect 208528 362866 208848 362898
rect 239248 363454 239568 363486
rect 239248 363218 239290 363454
rect 239526 363218 239568 363454
rect 239248 363134 239568 363218
rect 239248 362898 239290 363134
rect 239526 362898 239568 363134
rect 239248 362866 239568 362898
rect 269968 363454 270288 363486
rect 269968 363218 270010 363454
rect 270246 363218 270288 363454
rect 269968 363134 270288 363218
rect 269968 362898 270010 363134
rect 270246 362898 270288 363134
rect 269968 362866 270288 362898
rect 300688 363454 301008 363486
rect 300688 363218 300730 363454
rect 300966 363218 301008 363454
rect 300688 363134 301008 363218
rect 300688 362898 300730 363134
rect 300966 362898 301008 363134
rect 300688 362866 301008 362898
rect 331408 363454 331728 363486
rect 331408 363218 331450 363454
rect 331686 363218 331728 363454
rect 331408 363134 331728 363218
rect 331408 362898 331450 363134
rect 331686 362898 331728 363134
rect 331408 362866 331728 362898
rect 361794 363454 362414 398898
rect 361794 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 362414 363454
rect 361794 363134 362414 363218
rect 361794 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 362414 363134
rect 27834 353258 27866 353494
rect 28102 353258 28186 353494
rect 28422 353258 28454 353494
rect 27834 353174 28454 353258
rect 27834 352938 27866 353174
rect 28102 352938 28186 353174
rect 28422 352938 28454 353174
rect 24208 327454 24528 327486
rect 24208 327218 24250 327454
rect 24486 327218 24528 327454
rect 24208 327134 24528 327218
rect 24208 326898 24250 327134
rect 24486 326898 24528 327134
rect 24208 326866 24528 326898
rect 20394 309818 20426 310054
rect 20662 309818 20746 310054
rect 20982 309818 21014 310054
rect 20394 309734 21014 309818
rect 20394 309498 20426 309734
rect 20662 309498 20746 309734
rect 20982 309498 21014 309734
rect 20394 274054 21014 309498
rect 27834 317494 28454 352938
rect 39568 331174 39888 331206
rect 39568 330938 39610 331174
rect 39846 330938 39888 331174
rect 39568 330854 39888 330938
rect 39568 330618 39610 330854
rect 39846 330618 39888 330854
rect 39568 330586 39888 330618
rect 70288 331174 70608 331206
rect 70288 330938 70330 331174
rect 70566 330938 70608 331174
rect 70288 330854 70608 330938
rect 70288 330618 70330 330854
rect 70566 330618 70608 330854
rect 70288 330586 70608 330618
rect 101008 331174 101328 331206
rect 101008 330938 101050 331174
rect 101286 330938 101328 331174
rect 101008 330854 101328 330938
rect 101008 330618 101050 330854
rect 101286 330618 101328 330854
rect 101008 330586 101328 330618
rect 131728 331174 132048 331206
rect 131728 330938 131770 331174
rect 132006 330938 132048 331174
rect 131728 330854 132048 330938
rect 131728 330618 131770 330854
rect 132006 330618 132048 330854
rect 131728 330586 132048 330618
rect 162448 331174 162768 331206
rect 162448 330938 162490 331174
rect 162726 330938 162768 331174
rect 162448 330854 162768 330938
rect 162448 330618 162490 330854
rect 162726 330618 162768 330854
rect 162448 330586 162768 330618
rect 193168 331174 193488 331206
rect 193168 330938 193210 331174
rect 193446 330938 193488 331174
rect 193168 330854 193488 330938
rect 193168 330618 193210 330854
rect 193446 330618 193488 330854
rect 193168 330586 193488 330618
rect 223888 331174 224208 331206
rect 223888 330938 223930 331174
rect 224166 330938 224208 331174
rect 223888 330854 224208 330938
rect 223888 330618 223930 330854
rect 224166 330618 224208 330854
rect 223888 330586 224208 330618
rect 254608 331174 254928 331206
rect 254608 330938 254650 331174
rect 254886 330938 254928 331174
rect 254608 330854 254928 330938
rect 254608 330618 254650 330854
rect 254886 330618 254928 330854
rect 254608 330586 254928 330618
rect 285328 331174 285648 331206
rect 285328 330938 285370 331174
rect 285606 330938 285648 331174
rect 285328 330854 285648 330938
rect 285328 330618 285370 330854
rect 285606 330618 285648 330854
rect 285328 330586 285648 330618
rect 316048 331174 316368 331206
rect 316048 330938 316090 331174
rect 316326 330938 316368 331174
rect 316048 330854 316368 330938
rect 316048 330618 316090 330854
rect 316326 330618 316368 330854
rect 316048 330586 316368 330618
rect 346768 331174 347088 331206
rect 346768 330938 346810 331174
rect 347046 330938 347088 331174
rect 346768 330854 347088 330938
rect 346768 330618 346810 330854
rect 347046 330618 347088 330854
rect 346768 330586 347088 330618
rect 54928 327454 55248 327486
rect 54928 327218 54970 327454
rect 55206 327218 55248 327454
rect 54928 327134 55248 327218
rect 54928 326898 54970 327134
rect 55206 326898 55248 327134
rect 54928 326866 55248 326898
rect 85648 327454 85968 327486
rect 85648 327218 85690 327454
rect 85926 327218 85968 327454
rect 85648 327134 85968 327218
rect 85648 326898 85690 327134
rect 85926 326898 85968 327134
rect 85648 326866 85968 326898
rect 116368 327454 116688 327486
rect 116368 327218 116410 327454
rect 116646 327218 116688 327454
rect 116368 327134 116688 327218
rect 116368 326898 116410 327134
rect 116646 326898 116688 327134
rect 116368 326866 116688 326898
rect 147088 327454 147408 327486
rect 147088 327218 147130 327454
rect 147366 327218 147408 327454
rect 147088 327134 147408 327218
rect 147088 326898 147130 327134
rect 147366 326898 147408 327134
rect 147088 326866 147408 326898
rect 177808 327454 178128 327486
rect 177808 327218 177850 327454
rect 178086 327218 178128 327454
rect 177808 327134 178128 327218
rect 177808 326898 177850 327134
rect 178086 326898 178128 327134
rect 177808 326866 178128 326898
rect 208528 327454 208848 327486
rect 208528 327218 208570 327454
rect 208806 327218 208848 327454
rect 208528 327134 208848 327218
rect 208528 326898 208570 327134
rect 208806 326898 208848 327134
rect 208528 326866 208848 326898
rect 239248 327454 239568 327486
rect 239248 327218 239290 327454
rect 239526 327218 239568 327454
rect 239248 327134 239568 327218
rect 239248 326898 239290 327134
rect 239526 326898 239568 327134
rect 239248 326866 239568 326898
rect 269968 327454 270288 327486
rect 269968 327218 270010 327454
rect 270246 327218 270288 327454
rect 269968 327134 270288 327218
rect 269968 326898 270010 327134
rect 270246 326898 270288 327134
rect 269968 326866 270288 326898
rect 300688 327454 301008 327486
rect 300688 327218 300730 327454
rect 300966 327218 301008 327454
rect 300688 327134 301008 327218
rect 300688 326898 300730 327134
rect 300966 326898 301008 327134
rect 300688 326866 301008 326898
rect 331408 327454 331728 327486
rect 331408 327218 331450 327454
rect 331686 327218 331728 327454
rect 331408 327134 331728 327218
rect 331408 326898 331450 327134
rect 331686 326898 331728 327134
rect 331408 326866 331728 326898
rect 361794 327454 362414 362898
rect 361794 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 362414 327454
rect 361794 327134 362414 327218
rect 361794 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 362414 327134
rect 27834 317258 27866 317494
rect 28102 317258 28186 317494
rect 28422 317258 28454 317494
rect 27834 317174 28454 317258
rect 27834 316938 27866 317174
rect 28102 316938 28186 317174
rect 28422 316938 28454 317174
rect 24208 291454 24528 291486
rect 24208 291218 24250 291454
rect 24486 291218 24528 291454
rect 24208 291134 24528 291218
rect 24208 290898 24250 291134
rect 24486 290898 24528 291134
rect 24208 290866 24528 290898
rect 20394 273818 20426 274054
rect 20662 273818 20746 274054
rect 20982 273818 21014 274054
rect 20394 273734 21014 273818
rect 20394 273498 20426 273734
rect 20662 273498 20746 273734
rect 20982 273498 21014 273734
rect 20394 238054 21014 273498
rect 27834 281494 28454 316938
rect 39568 295174 39888 295206
rect 39568 294938 39610 295174
rect 39846 294938 39888 295174
rect 39568 294854 39888 294938
rect 39568 294618 39610 294854
rect 39846 294618 39888 294854
rect 39568 294586 39888 294618
rect 70288 295174 70608 295206
rect 70288 294938 70330 295174
rect 70566 294938 70608 295174
rect 70288 294854 70608 294938
rect 70288 294618 70330 294854
rect 70566 294618 70608 294854
rect 70288 294586 70608 294618
rect 101008 295174 101328 295206
rect 101008 294938 101050 295174
rect 101286 294938 101328 295174
rect 101008 294854 101328 294938
rect 101008 294618 101050 294854
rect 101286 294618 101328 294854
rect 101008 294586 101328 294618
rect 131728 295174 132048 295206
rect 131728 294938 131770 295174
rect 132006 294938 132048 295174
rect 131728 294854 132048 294938
rect 131728 294618 131770 294854
rect 132006 294618 132048 294854
rect 131728 294586 132048 294618
rect 162448 295174 162768 295206
rect 162448 294938 162490 295174
rect 162726 294938 162768 295174
rect 162448 294854 162768 294938
rect 162448 294618 162490 294854
rect 162726 294618 162768 294854
rect 162448 294586 162768 294618
rect 193168 295174 193488 295206
rect 193168 294938 193210 295174
rect 193446 294938 193488 295174
rect 193168 294854 193488 294938
rect 193168 294618 193210 294854
rect 193446 294618 193488 294854
rect 193168 294586 193488 294618
rect 223888 295174 224208 295206
rect 223888 294938 223930 295174
rect 224166 294938 224208 295174
rect 223888 294854 224208 294938
rect 223888 294618 223930 294854
rect 224166 294618 224208 294854
rect 223888 294586 224208 294618
rect 254608 295174 254928 295206
rect 254608 294938 254650 295174
rect 254886 294938 254928 295174
rect 254608 294854 254928 294938
rect 254608 294618 254650 294854
rect 254886 294618 254928 294854
rect 254608 294586 254928 294618
rect 285328 295174 285648 295206
rect 285328 294938 285370 295174
rect 285606 294938 285648 295174
rect 285328 294854 285648 294938
rect 285328 294618 285370 294854
rect 285606 294618 285648 294854
rect 285328 294586 285648 294618
rect 316048 295174 316368 295206
rect 316048 294938 316090 295174
rect 316326 294938 316368 295174
rect 316048 294854 316368 294938
rect 316048 294618 316090 294854
rect 316326 294618 316368 294854
rect 316048 294586 316368 294618
rect 346768 295174 347088 295206
rect 346768 294938 346810 295174
rect 347046 294938 347088 295174
rect 346768 294854 347088 294938
rect 346768 294618 346810 294854
rect 347046 294618 347088 294854
rect 346768 294586 347088 294618
rect 54928 291454 55248 291486
rect 54928 291218 54970 291454
rect 55206 291218 55248 291454
rect 54928 291134 55248 291218
rect 54928 290898 54970 291134
rect 55206 290898 55248 291134
rect 54928 290866 55248 290898
rect 85648 291454 85968 291486
rect 85648 291218 85690 291454
rect 85926 291218 85968 291454
rect 85648 291134 85968 291218
rect 85648 290898 85690 291134
rect 85926 290898 85968 291134
rect 85648 290866 85968 290898
rect 116368 291454 116688 291486
rect 116368 291218 116410 291454
rect 116646 291218 116688 291454
rect 116368 291134 116688 291218
rect 116368 290898 116410 291134
rect 116646 290898 116688 291134
rect 116368 290866 116688 290898
rect 147088 291454 147408 291486
rect 147088 291218 147130 291454
rect 147366 291218 147408 291454
rect 147088 291134 147408 291218
rect 147088 290898 147130 291134
rect 147366 290898 147408 291134
rect 147088 290866 147408 290898
rect 177808 291454 178128 291486
rect 177808 291218 177850 291454
rect 178086 291218 178128 291454
rect 177808 291134 178128 291218
rect 177808 290898 177850 291134
rect 178086 290898 178128 291134
rect 177808 290866 178128 290898
rect 208528 291454 208848 291486
rect 208528 291218 208570 291454
rect 208806 291218 208848 291454
rect 208528 291134 208848 291218
rect 208528 290898 208570 291134
rect 208806 290898 208848 291134
rect 208528 290866 208848 290898
rect 239248 291454 239568 291486
rect 239248 291218 239290 291454
rect 239526 291218 239568 291454
rect 239248 291134 239568 291218
rect 239248 290898 239290 291134
rect 239526 290898 239568 291134
rect 239248 290866 239568 290898
rect 269968 291454 270288 291486
rect 269968 291218 270010 291454
rect 270246 291218 270288 291454
rect 269968 291134 270288 291218
rect 269968 290898 270010 291134
rect 270246 290898 270288 291134
rect 269968 290866 270288 290898
rect 300688 291454 301008 291486
rect 300688 291218 300730 291454
rect 300966 291218 301008 291454
rect 300688 291134 301008 291218
rect 300688 290898 300730 291134
rect 300966 290898 301008 291134
rect 300688 290866 301008 290898
rect 331408 291454 331728 291486
rect 331408 291218 331450 291454
rect 331686 291218 331728 291454
rect 331408 291134 331728 291218
rect 331408 290898 331450 291134
rect 331686 290898 331728 291134
rect 331408 290866 331728 290898
rect 361794 291454 362414 326898
rect 361794 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 362414 291454
rect 361794 291134 362414 291218
rect 361794 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 362414 291134
rect 27834 281258 27866 281494
rect 28102 281258 28186 281494
rect 28422 281258 28454 281494
rect 27834 281174 28454 281258
rect 27834 280938 27866 281174
rect 28102 280938 28186 281174
rect 28422 280938 28454 281174
rect 24208 255454 24528 255486
rect 24208 255218 24250 255454
rect 24486 255218 24528 255454
rect 24208 255134 24528 255218
rect 24208 254898 24250 255134
rect 24486 254898 24528 255134
rect 24208 254866 24528 254898
rect 20394 237818 20426 238054
rect 20662 237818 20746 238054
rect 20982 237818 21014 238054
rect 20394 237734 21014 237818
rect 20394 237498 20426 237734
rect 20662 237498 20746 237734
rect 20982 237498 21014 237734
rect 20394 202054 21014 237498
rect 27834 245494 28454 280938
rect 39568 259174 39888 259206
rect 39568 258938 39610 259174
rect 39846 258938 39888 259174
rect 39568 258854 39888 258938
rect 39568 258618 39610 258854
rect 39846 258618 39888 258854
rect 39568 258586 39888 258618
rect 70288 259174 70608 259206
rect 70288 258938 70330 259174
rect 70566 258938 70608 259174
rect 70288 258854 70608 258938
rect 70288 258618 70330 258854
rect 70566 258618 70608 258854
rect 70288 258586 70608 258618
rect 101008 259174 101328 259206
rect 101008 258938 101050 259174
rect 101286 258938 101328 259174
rect 101008 258854 101328 258938
rect 101008 258618 101050 258854
rect 101286 258618 101328 258854
rect 101008 258586 101328 258618
rect 131728 259174 132048 259206
rect 131728 258938 131770 259174
rect 132006 258938 132048 259174
rect 131728 258854 132048 258938
rect 131728 258618 131770 258854
rect 132006 258618 132048 258854
rect 131728 258586 132048 258618
rect 162448 259174 162768 259206
rect 162448 258938 162490 259174
rect 162726 258938 162768 259174
rect 162448 258854 162768 258938
rect 162448 258618 162490 258854
rect 162726 258618 162768 258854
rect 162448 258586 162768 258618
rect 193168 259174 193488 259206
rect 193168 258938 193210 259174
rect 193446 258938 193488 259174
rect 193168 258854 193488 258938
rect 193168 258618 193210 258854
rect 193446 258618 193488 258854
rect 193168 258586 193488 258618
rect 223888 259174 224208 259206
rect 223888 258938 223930 259174
rect 224166 258938 224208 259174
rect 223888 258854 224208 258938
rect 223888 258618 223930 258854
rect 224166 258618 224208 258854
rect 223888 258586 224208 258618
rect 254608 259174 254928 259206
rect 254608 258938 254650 259174
rect 254886 258938 254928 259174
rect 254608 258854 254928 258938
rect 254608 258618 254650 258854
rect 254886 258618 254928 258854
rect 254608 258586 254928 258618
rect 285328 259174 285648 259206
rect 285328 258938 285370 259174
rect 285606 258938 285648 259174
rect 285328 258854 285648 258938
rect 285328 258618 285370 258854
rect 285606 258618 285648 258854
rect 285328 258586 285648 258618
rect 316048 259174 316368 259206
rect 316048 258938 316090 259174
rect 316326 258938 316368 259174
rect 316048 258854 316368 258938
rect 316048 258618 316090 258854
rect 316326 258618 316368 258854
rect 316048 258586 316368 258618
rect 346768 259174 347088 259206
rect 346768 258938 346810 259174
rect 347046 258938 347088 259174
rect 346768 258854 347088 258938
rect 346768 258618 346810 258854
rect 347046 258618 347088 258854
rect 346768 258586 347088 258618
rect 54928 255454 55248 255486
rect 54928 255218 54970 255454
rect 55206 255218 55248 255454
rect 54928 255134 55248 255218
rect 54928 254898 54970 255134
rect 55206 254898 55248 255134
rect 54928 254866 55248 254898
rect 85648 255454 85968 255486
rect 85648 255218 85690 255454
rect 85926 255218 85968 255454
rect 85648 255134 85968 255218
rect 85648 254898 85690 255134
rect 85926 254898 85968 255134
rect 85648 254866 85968 254898
rect 116368 255454 116688 255486
rect 116368 255218 116410 255454
rect 116646 255218 116688 255454
rect 116368 255134 116688 255218
rect 116368 254898 116410 255134
rect 116646 254898 116688 255134
rect 116368 254866 116688 254898
rect 147088 255454 147408 255486
rect 147088 255218 147130 255454
rect 147366 255218 147408 255454
rect 147088 255134 147408 255218
rect 147088 254898 147130 255134
rect 147366 254898 147408 255134
rect 147088 254866 147408 254898
rect 177808 255454 178128 255486
rect 177808 255218 177850 255454
rect 178086 255218 178128 255454
rect 177808 255134 178128 255218
rect 177808 254898 177850 255134
rect 178086 254898 178128 255134
rect 177808 254866 178128 254898
rect 208528 255454 208848 255486
rect 208528 255218 208570 255454
rect 208806 255218 208848 255454
rect 208528 255134 208848 255218
rect 208528 254898 208570 255134
rect 208806 254898 208848 255134
rect 208528 254866 208848 254898
rect 239248 255454 239568 255486
rect 239248 255218 239290 255454
rect 239526 255218 239568 255454
rect 239248 255134 239568 255218
rect 239248 254898 239290 255134
rect 239526 254898 239568 255134
rect 239248 254866 239568 254898
rect 269968 255454 270288 255486
rect 269968 255218 270010 255454
rect 270246 255218 270288 255454
rect 269968 255134 270288 255218
rect 269968 254898 270010 255134
rect 270246 254898 270288 255134
rect 269968 254866 270288 254898
rect 300688 255454 301008 255486
rect 300688 255218 300730 255454
rect 300966 255218 301008 255454
rect 300688 255134 301008 255218
rect 300688 254898 300730 255134
rect 300966 254898 301008 255134
rect 300688 254866 301008 254898
rect 331408 255454 331728 255486
rect 331408 255218 331450 255454
rect 331686 255218 331728 255454
rect 331408 255134 331728 255218
rect 331408 254898 331450 255134
rect 331686 254898 331728 255134
rect 331408 254866 331728 254898
rect 361794 255454 362414 290898
rect 361794 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 362414 255454
rect 361794 255134 362414 255218
rect 361794 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 362414 255134
rect 27834 245258 27866 245494
rect 28102 245258 28186 245494
rect 28422 245258 28454 245494
rect 27834 245174 28454 245258
rect 27834 244938 27866 245174
rect 28102 244938 28186 245174
rect 28422 244938 28454 245174
rect 24208 219454 24528 219486
rect 24208 219218 24250 219454
rect 24486 219218 24528 219454
rect 24208 219134 24528 219218
rect 24208 218898 24250 219134
rect 24486 218898 24528 219134
rect 24208 218866 24528 218898
rect 20394 201818 20426 202054
rect 20662 201818 20746 202054
rect 20982 201818 21014 202054
rect 20394 201734 21014 201818
rect 20394 201498 20426 201734
rect 20662 201498 20746 201734
rect 20982 201498 21014 201734
rect 20394 166054 21014 201498
rect 27834 209494 28454 244938
rect 39568 223174 39888 223206
rect 39568 222938 39610 223174
rect 39846 222938 39888 223174
rect 39568 222854 39888 222938
rect 39568 222618 39610 222854
rect 39846 222618 39888 222854
rect 39568 222586 39888 222618
rect 70288 223174 70608 223206
rect 70288 222938 70330 223174
rect 70566 222938 70608 223174
rect 70288 222854 70608 222938
rect 70288 222618 70330 222854
rect 70566 222618 70608 222854
rect 70288 222586 70608 222618
rect 101008 223174 101328 223206
rect 101008 222938 101050 223174
rect 101286 222938 101328 223174
rect 101008 222854 101328 222938
rect 101008 222618 101050 222854
rect 101286 222618 101328 222854
rect 101008 222586 101328 222618
rect 131728 223174 132048 223206
rect 131728 222938 131770 223174
rect 132006 222938 132048 223174
rect 131728 222854 132048 222938
rect 131728 222618 131770 222854
rect 132006 222618 132048 222854
rect 131728 222586 132048 222618
rect 162448 223174 162768 223206
rect 162448 222938 162490 223174
rect 162726 222938 162768 223174
rect 162448 222854 162768 222938
rect 162448 222618 162490 222854
rect 162726 222618 162768 222854
rect 162448 222586 162768 222618
rect 193168 223174 193488 223206
rect 193168 222938 193210 223174
rect 193446 222938 193488 223174
rect 193168 222854 193488 222938
rect 193168 222618 193210 222854
rect 193446 222618 193488 222854
rect 193168 222586 193488 222618
rect 223888 223174 224208 223206
rect 223888 222938 223930 223174
rect 224166 222938 224208 223174
rect 223888 222854 224208 222938
rect 223888 222618 223930 222854
rect 224166 222618 224208 222854
rect 223888 222586 224208 222618
rect 254608 223174 254928 223206
rect 254608 222938 254650 223174
rect 254886 222938 254928 223174
rect 254608 222854 254928 222938
rect 254608 222618 254650 222854
rect 254886 222618 254928 222854
rect 254608 222586 254928 222618
rect 285328 223174 285648 223206
rect 285328 222938 285370 223174
rect 285606 222938 285648 223174
rect 285328 222854 285648 222938
rect 285328 222618 285370 222854
rect 285606 222618 285648 222854
rect 285328 222586 285648 222618
rect 316048 223174 316368 223206
rect 316048 222938 316090 223174
rect 316326 222938 316368 223174
rect 316048 222854 316368 222938
rect 316048 222618 316090 222854
rect 316326 222618 316368 222854
rect 316048 222586 316368 222618
rect 346768 223174 347088 223206
rect 346768 222938 346810 223174
rect 347046 222938 347088 223174
rect 346768 222854 347088 222938
rect 346768 222618 346810 222854
rect 347046 222618 347088 222854
rect 346768 222586 347088 222618
rect 54928 219454 55248 219486
rect 54928 219218 54970 219454
rect 55206 219218 55248 219454
rect 54928 219134 55248 219218
rect 54928 218898 54970 219134
rect 55206 218898 55248 219134
rect 54928 218866 55248 218898
rect 85648 219454 85968 219486
rect 85648 219218 85690 219454
rect 85926 219218 85968 219454
rect 85648 219134 85968 219218
rect 85648 218898 85690 219134
rect 85926 218898 85968 219134
rect 85648 218866 85968 218898
rect 116368 219454 116688 219486
rect 116368 219218 116410 219454
rect 116646 219218 116688 219454
rect 116368 219134 116688 219218
rect 116368 218898 116410 219134
rect 116646 218898 116688 219134
rect 116368 218866 116688 218898
rect 147088 219454 147408 219486
rect 147088 219218 147130 219454
rect 147366 219218 147408 219454
rect 147088 219134 147408 219218
rect 147088 218898 147130 219134
rect 147366 218898 147408 219134
rect 147088 218866 147408 218898
rect 177808 219454 178128 219486
rect 177808 219218 177850 219454
rect 178086 219218 178128 219454
rect 177808 219134 178128 219218
rect 177808 218898 177850 219134
rect 178086 218898 178128 219134
rect 177808 218866 178128 218898
rect 208528 219454 208848 219486
rect 208528 219218 208570 219454
rect 208806 219218 208848 219454
rect 208528 219134 208848 219218
rect 208528 218898 208570 219134
rect 208806 218898 208848 219134
rect 208528 218866 208848 218898
rect 239248 219454 239568 219486
rect 239248 219218 239290 219454
rect 239526 219218 239568 219454
rect 239248 219134 239568 219218
rect 239248 218898 239290 219134
rect 239526 218898 239568 219134
rect 239248 218866 239568 218898
rect 269968 219454 270288 219486
rect 269968 219218 270010 219454
rect 270246 219218 270288 219454
rect 269968 219134 270288 219218
rect 269968 218898 270010 219134
rect 270246 218898 270288 219134
rect 269968 218866 270288 218898
rect 300688 219454 301008 219486
rect 300688 219218 300730 219454
rect 300966 219218 301008 219454
rect 300688 219134 301008 219218
rect 300688 218898 300730 219134
rect 300966 218898 301008 219134
rect 300688 218866 301008 218898
rect 331408 219454 331728 219486
rect 331408 219218 331450 219454
rect 331686 219218 331728 219454
rect 331408 219134 331728 219218
rect 331408 218898 331450 219134
rect 331686 218898 331728 219134
rect 331408 218866 331728 218898
rect 361794 219454 362414 254898
rect 361794 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 362414 219454
rect 361794 219134 362414 219218
rect 361794 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 362414 219134
rect 27834 209258 27866 209494
rect 28102 209258 28186 209494
rect 28422 209258 28454 209494
rect 27834 209174 28454 209258
rect 27834 208938 27866 209174
rect 28102 208938 28186 209174
rect 28422 208938 28454 209174
rect 24208 183454 24528 183486
rect 24208 183218 24250 183454
rect 24486 183218 24528 183454
rect 24208 183134 24528 183218
rect 24208 182898 24250 183134
rect 24486 182898 24528 183134
rect 24208 182866 24528 182898
rect 20394 165818 20426 166054
rect 20662 165818 20746 166054
rect 20982 165818 21014 166054
rect 20394 165734 21014 165818
rect 20394 165498 20426 165734
rect 20662 165498 20746 165734
rect 20982 165498 21014 165734
rect 20394 130054 21014 165498
rect 27834 173494 28454 208938
rect 39568 187174 39888 187206
rect 39568 186938 39610 187174
rect 39846 186938 39888 187174
rect 39568 186854 39888 186938
rect 39568 186618 39610 186854
rect 39846 186618 39888 186854
rect 39568 186586 39888 186618
rect 70288 187174 70608 187206
rect 70288 186938 70330 187174
rect 70566 186938 70608 187174
rect 70288 186854 70608 186938
rect 70288 186618 70330 186854
rect 70566 186618 70608 186854
rect 70288 186586 70608 186618
rect 101008 187174 101328 187206
rect 101008 186938 101050 187174
rect 101286 186938 101328 187174
rect 101008 186854 101328 186938
rect 101008 186618 101050 186854
rect 101286 186618 101328 186854
rect 101008 186586 101328 186618
rect 131728 187174 132048 187206
rect 131728 186938 131770 187174
rect 132006 186938 132048 187174
rect 131728 186854 132048 186938
rect 131728 186618 131770 186854
rect 132006 186618 132048 186854
rect 131728 186586 132048 186618
rect 162448 187174 162768 187206
rect 162448 186938 162490 187174
rect 162726 186938 162768 187174
rect 162448 186854 162768 186938
rect 162448 186618 162490 186854
rect 162726 186618 162768 186854
rect 162448 186586 162768 186618
rect 193168 187174 193488 187206
rect 193168 186938 193210 187174
rect 193446 186938 193488 187174
rect 193168 186854 193488 186938
rect 193168 186618 193210 186854
rect 193446 186618 193488 186854
rect 193168 186586 193488 186618
rect 223888 187174 224208 187206
rect 223888 186938 223930 187174
rect 224166 186938 224208 187174
rect 223888 186854 224208 186938
rect 223888 186618 223930 186854
rect 224166 186618 224208 186854
rect 223888 186586 224208 186618
rect 254608 187174 254928 187206
rect 254608 186938 254650 187174
rect 254886 186938 254928 187174
rect 254608 186854 254928 186938
rect 254608 186618 254650 186854
rect 254886 186618 254928 186854
rect 254608 186586 254928 186618
rect 285328 187174 285648 187206
rect 285328 186938 285370 187174
rect 285606 186938 285648 187174
rect 285328 186854 285648 186938
rect 285328 186618 285370 186854
rect 285606 186618 285648 186854
rect 285328 186586 285648 186618
rect 316048 187174 316368 187206
rect 316048 186938 316090 187174
rect 316326 186938 316368 187174
rect 316048 186854 316368 186938
rect 316048 186618 316090 186854
rect 316326 186618 316368 186854
rect 316048 186586 316368 186618
rect 346768 187174 347088 187206
rect 346768 186938 346810 187174
rect 347046 186938 347088 187174
rect 346768 186854 347088 186938
rect 346768 186618 346810 186854
rect 347046 186618 347088 186854
rect 346768 186586 347088 186618
rect 54928 183454 55248 183486
rect 54928 183218 54970 183454
rect 55206 183218 55248 183454
rect 54928 183134 55248 183218
rect 54928 182898 54970 183134
rect 55206 182898 55248 183134
rect 54928 182866 55248 182898
rect 85648 183454 85968 183486
rect 85648 183218 85690 183454
rect 85926 183218 85968 183454
rect 85648 183134 85968 183218
rect 85648 182898 85690 183134
rect 85926 182898 85968 183134
rect 85648 182866 85968 182898
rect 116368 183454 116688 183486
rect 116368 183218 116410 183454
rect 116646 183218 116688 183454
rect 116368 183134 116688 183218
rect 116368 182898 116410 183134
rect 116646 182898 116688 183134
rect 116368 182866 116688 182898
rect 147088 183454 147408 183486
rect 147088 183218 147130 183454
rect 147366 183218 147408 183454
rect 147088 183134 147408 183218
rect 147088 182898 147130 183134
rect 147366 182898 147408 183134
rect 147088 182866 147408 182898
rect 177808 183454 178128 183486
rect 177808 183218 177850 183454
rect 178086 183218 178128 183454
rect 177808 183134 178128 183218
rect 177808 182898 177850 183134
rect 178086 182898 178128 183134
rect 177808 182866 178128 182898
rect 208528 183454 208848 183486
rect 208528 183218 208570 183454
rect 208806 183218 208848 183454
rect 208528 183134 208848 183218
rect 208528 182898 208570 183134
rect 208806 182898 208848 183134
rect 208528 182866 208848 182898
rect 239248 183454 239568 183486
rect 239248 183218 239290 183454
rect 239526 183218 239568 183454
rect 239248 183134 239568 183218
rect 239248 182898 239290 183134
rect 239526 182898 239568 183134
rect 239248 182866 239568 182898
rect 269968 183454 270288 183486
rect 269968 183218 270010 183454
rect 270246 183218 270288 183454
rect 269968 183134 270288 183218
rect 269968 182898 270010 183134
rect 270246 182898 270288 183134
rect 269968 182866 270288 182898
rect 300688 183454 301008 183486
rect 300688 183218 300730 183454
rect 300966 183218 301008 183454
rect 300688 183134 301008 183218
rect 300688 182898 300730 183134
rect 300966 182898 301008 183134
rect 300688 182866 301008 182898
rect 331408 183454 331728 183486
rect 331408 183218 331450 183454
rect 331686 183218 331728 183454
rect 331408 183134 331728 183218
rect 331408 182898 331450 183134
rect 331686 182898 331728 183134
rect 331408 182866 331728 182898
rect 361794 183454 362414 218898
rect 361794 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 362414 183454
rect 361794 183134 362414 183218
rect 361794 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 362414 183134
rect 27834 173258 27866 173494
rect 28102 173258 28186 173494
rect 28422 173258 28454 173494
rect 27834 173174 28454 173258
rect 27834 172938 27866 173174
rect 28102 172938 28186 173174
rect 28422 172938 28454 173174
rect 24208 147454 24528 147486
rect 24208 147218 24250 147454
rect 24486 147218 24528 147454
rect 24208 147134 24528 147218
rect 24208 146898 24250 147134
rect 24486 146898 24528 147134
rect 24208 146866 24528 146898
rect 20394 129818 20426 130054
rect 20662 129818 20746 130054
rect 20982 129818 21014 130054
rect 20394 129734 21014 129818
rect 20394 129498 20426 129734
rect 20662 129498 20746 129734
rect 20982 129498 21014 129734
rect 20394 94054 21014 129498
rect 27834 137494 28454 172938
rect 39568 151174 39888 151206
rect 39568 150938 39610 151174
rect 39846 150938 39888 151174
rect 39568 150854 39888 150938
rect 39568 150618 39610 150854
rect 39846 150618 39888 150854
rect 39568 150586 39888 150618
rect 70288 151174 70608 151206
rect 70288 150938 70330 151174
rect 70566 150938 70608 151174
rect 70288 150854 70608 150938
rect 70288 150618 70330 150854
rect 70566 150618 70608 150854
rect 70288 150586 70608 150618
rect 101008 151174 101328 151206
rect 101008 150938 101050 151174
rect 101286 150938 101328 151174
rect 101008 150854 101328 150938
rect 101008 150618 101050 150854
rect 101286 150618 101328 150854
rect 101008 150586 101328 150618
rect 131728 151174 132048 151206
rect 131728 150938 131770 151174
rect 132006 150938 132048 151174
rect 131728 150854 132048 150938
rect 131728 150618 131770 150854
rect 132006 150618 132048 150854
rect 131728 150586 132048 150618
rect 162448 151174 162768 151206
rect 162448 150938 162490 151174
rect 162726 150938 162768 151174
rect 162448 150854 162768 150938
rect 162448 150618 162490 150854
rect 162726 150618 162768 150854
rect 162448 150586 162768 150618
rect 193168 151174 193488 151206
rect 193168 150938 193210 151174
rect 193446 150938 193488 151174
rect 193168 150854 193488 150938
rect 193168 150618 193210 150854
rect 193446 150618 193488 150854
rect 193168 150586 193488 150618
rect 223888 151174 224208 151206
rect 223888 150938 223930 151174
rect 224166 150938 224208 151174
rect 223888 150854 224208 150938
rect 223888 150618 223930 150854
rect 224166 150618 224208 150854
rect 223888 150586 224208 150618
rect 254608 151174 254928 151206
rect 254608 150938 254650 151174
rect 254886 150938 254928 151174
rect 254608 150854 254928 150938
rect 254608 150618 254650 150854
rect 254886 150618 254928 150854
rect 254608 150586 254928 150618
rect 285328 151174 285648 151206
rect 285328 150938 285370 151174
rect 285606 150938 285648 151174
rect 285328 150854 285648 150938
rect 285328 150618 285370 150854
rect 285606 150618 285648 150854
rect 285328 150586 285648 150618
rect 316048 151174 316368 151206
rect 316048 150938 316090 151174
rect 316326 150938 316368 151174
rect 316048 150854 316368 150938
rect 316048 150618 316090 150854
rect 316326 150618 316368 150854
rect 316048 150586 316368 150618
rect 346768 151174 347088 151206
rect 346768 150938 346810 151174
rect 347046 150938 347088 151174
rect 346768 150854 347088 150938
rect 346768 150618 346810 150854
rect 347046 150618 347088 150854
rect 346768 150586 347088 150618
rect 54928 147454 55248 147486
rect 54928 147218 54970 147454
rect 55206 147218 55248 147454
rect 54928 147134 55248 147218
rect 54928 146898 54970 147134
rect 55206 146898 55248 147134
rect 54928 146866 55248 146898
rect 85648 147454 85968 147486
rect 85648 147218 85690 147454
rect 85926 147218 85968 147454
rect 85648 147134 85968 147218
rect 85648 146898 85690 147134
rect 85926 146898 85968 147134
rect 85648 146866 85968 146898
rect 116368 147454 116688 147486
rect 116368 147218 116410 147454
rect 116646 147218 116688 147454
rect 116368 147134 116688 147218
rect 116368 146898 116410 147134
rect 116646 146898 116688 147134
rect 116368 146866 116688 146898
rect 147088 147454 147408 147486
rect 147088 147218 147130 147454
rect 147366 147218 147408 147454
rect 147088 147134 147408 147218
rect 147088 146898 147130 147134
rect 147366 146898 147408 147134
rect 147088 146866 147408 146898
rect 177808 147454 178128 147486
rect 177808 147218 177850 147454
rect 178086 147218 178128 147454
rect 177808 147134 178128 147218
rect 177808 146898 177850 147134
rect 178086 146898 178128 147134
rect 177808 146866 178128 146898
rect 208528 147454 208848 147486
rect 208528 147218 208570 147454
rect 208806 147218 208848 147454
rect 208528 147134 208848 147218
rect 208528 146898 208570 147134
rect 208806 146898 208848 147134
rect 208528 146866 208848 146898
rect 239248 147454 239568 147486
rect 239248 147218 239290 147454
rect 239526 147218 239568 147454
rect 239248 147134 239568 147218
rect 239248 146898 239290 147134
rect 239526 146898 239568 147134
rect 239248 146866 239568 146898
rect 269968 147454 270288 147486
rect 269968 147218 270010 147454
rect 270246 147218 270288 147454
rect 269968 147134 270288 147218
rect 269968 146898 270010 147134
rect 270246 146898 270288 147134
rect 269968 146866 270288 146898
rect 300688 147454 301008 147486
rect 300688 147218 300730 147454
rect 300966 147218 301008 147454
rect 300688 147134 301008 147218
rect 300688 146898 300730 147134
rect 300966 146898 301008 147134
rect 300688 146866 301008 146898
rect 331408 147454 331728 147486
rect 331408 147218 331450 147454
rect 331686 147218 331728 147454
rect 331408 147134 331728 147218
rect 331408 146898 331450 147134
rect 331686 146898 331728 147134
rect 331408 146866 331728 146898
rect 361794 147454 362414 182898
rect 361794 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 362414 147454
rect 361794 147134 362414 147218
rect 361794 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 362414 147134
rect 27834 137258 27866 137494
rect 28102 137258 28186 137494
rect 28422 137258 28454 137494
rect 27834 137174 28454 137258
rect 27834 136938 27866 137174
rect 28102 136938 28186 137174
rect 28422 136938 28454 137174
rect 24208 111454 24528 111486
rect 24208 111218 24250 111454
rect 24486 111218 24528 111454
rect 24208 111134 24528 111218
rect 24208 110898 24250 111134
rect 24486 110898 24528 111134
rect 24208 110866 24528 110898
rect 20394 93818 20426 94054
rect 20662 93818 20746 94054
rect 20982 93818 21014 94054
rect 20394 93734 21014 93818
rect 20394 93498 20426 93734
rect 20662 93498 20746 93734
rect 20982 93498 21014 93734
rect 20394 58054 21014 93498
rect 27834 101494 28454 136938
rect 39568 115174 39888 115206
rect 39568 114938 39610 115174
rect 39846 114938 39888 115174
rect 39568 114854 39888 114938
rect 39568 114618 39610 114854
rect 39846 114618 39888 114854
rect 39568 114586 39888 114618
rect 70288 115174 70608 115206
rect 70288 114938 70330 115174
rect 70566 114938 70608 115174
rect 70288 114854 70608 114938
rect 70288 114618 70330 114854
rect 70566 114618 70608 114854
rect 70288 114586 70608 114618
rect 101008 115174 101328 115206
rect 101008 114938 101050 115174
rect 101286 114938 101328 115174
rect 101008 114854 101328 114938
rect 101008 114618 101050 114854
rect 101286 114618 101328 114854
rect 101008 114586 101328 114618
rect 131728 115174 132048 115206
rect 131728 114938 131770 115174
rect 132006 114938 132048 115174
rect 131728 114854 132048 114938
rect 131728 114618 131770 114854
rect 132006 114618 132048 114854
rect 131728 114586 132048 114618
rect 162448 115174 162768 115206
rect 162448 114938 162490 115174
rect 162726 114938 162768 115174
rect 162448 114854 162768 114938
rect 162448 114618 162490 114854
rect 162726 114618 162768 114854
rect 162448 114586 162768 114618
rect 193168 115174 193488 115206
rect 193168 114938 193210 115174
rect 193446 114938 193488 115174
rect 193168 114854 193488 114938
rect 193168 114618 193210 114854
rect 193446 114618 193488 114854
rect 193168 114586 193488 114618
rect 223888 115174 224208 115206
rect 223888 114938 223930 115174
rect 224166 114938 224208 115174
rect 223888 114854 224208 114938
rect 223888 114618 223930 114854
rect 224166 114618 224208 114854
rect 223888 114586 224208 114618
rect 254608 115174 254928 115206
rect 254608 114938 254650 115174
rect 254886 114938 254928 115174
rect 254608 114854 254928 114938
rect 254608 114618 254650 114854
rect 254886 114618 254928 114854
rect 254608 114586 254928 114618
rect 285328 115174 285648 115206
rect 285328 114938 285370 115174
rect 285606 114938 285648 115174
rect 285328 114854 285648 114938
rect 285328 114618 285370 114854
rect 285606 114618 285648 114854
rect 285328 114586 285648 114618
rect 316048 115174 316368 115206
rect 316048 114938 316090 115174
rect 316326 114938 316368 115174
rect 316048 114854 316368 114938
rect 316048 114618 316090 114854
rect 316326 114618 316368 114854
rect 316048 114586 316368 114618
rect 346768 115174 347088 115206
rect 346768 114938 346810 115174
rect 347046 114938 347088 115174
rect 346768 114854 347088 114938
rect 346768 114618 346810 114854
rect 347046 114618 347088 114854
rect 346768 114586 347088 114618
rect 54928 111454 55248 111486
rect 54928 111218 54970 111454
rect 55206 111218 55248 111454
rect 54928 111134 55248 111218
rect 54928 110898 54970 111134
rect 55206 110898 55248 111134
rect 54928 110866 55248 110898
rect 85648 111454 85968 111486
rect 85648 111218 85690 111454
rect 85926 111218 85968 111454
rect 85648 111134 85968 111218
rect 85648 110898 85690 111134
rect 85926 110898 85968 111134
rect 85648 110866 85968 110898
rect 116368 111454 116688 111486
rect 116368 111218 116410 111454
rect 116646 111218 116688 111454
rect 116368 111134 116688 111218
rect 116368 110898 116410 111134
rect 116646 110898 116688 111134
rect 116368 110866 116688 110898
rect 147088 111454 147408 111486
rect 147088 111218 147130 111454
rect 147366 111218 147408 111454
rect 147088 111134 147408 111218
rect 147088 110898 147130 111134
rect 147366 110898 147408 111134
rect 147088 110866 147408 110898
rect 177808 111454 178128 111486
rect 177808 111218 177850 111454
rect 178086 111218 178128 111454
rect 177808 111134 178128 111218
rect 177808 110898 177850 111134
rect 178086 110898 178128 111134
rect 177808 110866 178128 110898
rect 208528 111454 208848 111486
rect 208528 111218 208570 111454
rect 208806 111218 208848 111454
rect 208528 111134 208848 111218
rect 208528 110898 208570 111134
rect 208806 110898 208848 111134
rect 208528 110866 208848 110898
rect 239248 111454 239568 111486
rect 239248 111218 239290 111454
rect 239526 111218 239568 111454
rect 239248 111134 239568 111218
rect 239248 110898 239290 111134
rect 239526 110898 239568 111134
rect 239248 110866 239568 110898
rect 269968 111454 270288 111486
rect 269968 111218 270010 111454
rect 270246 111218 270288 111454
rect 269968 111134 270288 111218
rect 269968 110898 270010 111134
rect 270246 110898 270288 111134
rect 269968 110866 270288 110898
rect 300688 111454 301008 111486
rect 300688 111218 300730 111454
rect 300966 111218 301008 111454
rect 300688 111134 301008 111218
rect 300688 110898 300730 111134
rect 300966 110898 301008 111134
rect 300688 110866 301008 110898
rect 331408 111454 331728 111486
rect 331408 111218 331450 111454
rect 331686 111218 331728 111454
rect 331408 111134 331728 111218
rect 331408 110898 331450 111134
rect 331686 110898 331728 111134
rect 331408 110866 331728 110898
rect 361794 111454 362414 146898
rect 361794 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 362414 111454
rect 361794 111134 362414 111218
rect 361794 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 362414 111134
rect 27834 101258 27866 101494
rect 28102 101258 28186 101494
rect 28422 101258 28454 101494
rect 27834 101174 28454 101258
rect 27834 100938 27866 101174
rect 28102 100938 28186 101174
rect 28422 100938 28454 101174
rect 24208 75454 24528 75486
rect 24208 75218 24250 75454
rect 24486 75218 24528 75454
rect 24208 75134 24528 75218
rect 24208 74898 24250 75134
rect 24486 74898 24528 75134
rect 24208 74866 24528 74898
rect 20394 57818 20426 58054
rect 20662 57818 20746 58054
rect 20982 57818 21014 58054
rect 20394 57734 21014 57818
rect 20394 57498 20426 57734
rect 20662 57498 20746 57734
rect 20982 57498 21014 57734
rect 20394 22054 21014 57498
rect 27834 65494 28454 100938
rect 39568 79174 39888 79206
rect 39568 78938 39610 79174
rect 39846 78938 39888 79174
rect 39568 78854 39888 78938
rect 39568 78618 39610 78854
rect 39846 78618 39888 78854
rect 39568 78586 39888 78618
rect 70288 79174 70608 79206
rect 70288 78938 70330 79174
rect 70566 78938 70608 79174
rect 70288 78854 70608 78938
rect 70288 78618 70330 78854
rect 70566 78618 70608 78854
rect 70288 78586 70608 78618
rect 101008 79174 101328 79206
rect 101008 78938 101050 79174
rect 101286 78938 101328 79174
rect 101008 78854 101328 78938
rect 101008 78618 101050 78854
rect 101286 78618 101328 78854
rect 101008 78586 101328 78618
rect 131728 79174 132048 79206
rect 131728 78938 131770 79174
rect 132006 78938 132048 79174
rect 131728 78854 132048 78938
rect 131728 78618 131770 78854
rect 132006 78618 132048 78854
rect 131728 78586 132048 78618
rect 162448 79174 162768 79206
rect 162448 78938 162490 79174
rect 162726 78938 162768 79174
rect 162448 78854 162768 78938
rect 162448 78618 162490 78854
rect 162726 78618 162768 78854
rect 162448 78586 162768 78618
rect 193168 79174 193488 79206
rect 193168 78938 193210 79174
rect 193446 78938 193488 79174
rect 193168 78854 193488 78938
rect 193168 78618 193210 78854
rect 193446 78618 193488 78854
rect 193168 78586 193488 78618
rect 223888 79174 224208 79206
rect 223888 78938 223930 79174
rect 224166 78938 224208 79174
rect 223888 78854 224208 78938
rect 223888 78618 223930 78854
rect 224166 78618 224208 78854
rect 223888 78586 224208 78618
rect 254608 79174 254928 79206
rect 254608 78938 254650 79174
rect 254886 78938 254928 79174
rect 254608 78854 254928 78938
rect 254608 78618 254650 78854
rect 254886 78618 254928 78854
rect 254608 78586 254928 78618
rect 285328 79174 285648 79206
rect 285328 78938 285370 79174
rect 285606 78938 285648 79174
rect 285328 78854 285648 78938
rect 285328 78618 285370 78854
rect 285606 78618 285648 78854
rect 285328 78586 285648 78618
rect 316048 79174 316368 79206
rect 316048 78938 316090 79174
rect 316326 78938 316368 79174
rect 316048 78854 316368 78938
rect 316048 78618 316090 78854
rect 316326 78618 316368 78854
rect 316048 78586 316368 78618
rect 346768 79174 347088 79206
rect 346768 78938 346810 79174
rect 347046 78938 347088 79174
rect 346768 78854 347088 78938
rect 346768 78618 346810 78854
rect 347046 78618 347088 78854
rect 346768 78586 347088 78618
rect 54928 75454 55248 75486
rect 54928 75218 54970 75454
rect 55206 75218 55248 75454
rect 54928 75134 55248 75218
rect 54928 74898 54970 75134
rect 55206 74898 55248 75134
rect 54928 74866 55248 74898
rect 85648 75454 85968 75486
rect 85648 75218 85690 75454
rect 85926 75218 85968 75454
rect 85648 75134 85968 75218
rect 85648 74898 85690 75134
rect 85926 74898 85968 75134
rect 85648 74866 85968 74898
rect 116368 75454 116688 75486
rect 116368 75218 116410 75454
rect 116646 75218 116688 75454
rect 116368 75134 116688 75218
rect 116368 74898 116410 75134
rect 116646 74898 116688 75134
rect 116368 74866 116688 74898
rect 147088 75454 147408 75486
rect 147088 75218 147130 75454
rect 147366 75218 147408 75454
rect 147088 75134 147408 75218
rect 147088 74898 147130 75134
rect 147366 74898 147408 75134
rect 147088 74866 147408 74898
rect 177808 75454 178128 75486
rect 177808 75218 177850 75454
rect 178086 75218 178128 75454
rect 177808 75134 178128 75218
rect 177808 74898 177850 75134
rect 178086 74898 178128 75134
rect 177808 74866 178128 74898
rect 208528 75454 208848 75486
rect 208528 75218 208570 75454
rect 208806 75218 208848 75454
rect 208528 75134 208848 75218
rect 208528 74898 208570 75134
rect 208806 74898 208848 75134
rect 208528 74866 208848 74898
rect 239248 75454 239568 75486
rect 239248 75218 239290 75454
rect 239526 75218 239568 75454
rect 239248 75134 239568 75218
rect 239248 74898 239290 75134
rect 239526 74898 239568 75134
rect 239248 74866 239568 74898
rect 269968 75454 270288 75486
rect 269968 75218 270010 75454
rect 270246 75218 270288 75454
rect 269968 75134 270288 75218
rect 269968 74898 270010 75134
rect 270246 74898 270288 75134
rect 269968 74866 270288 74898
rect 300688 75454 301008 75486
rect 300688 75218 300730 75454
rect 300966 75218 301008 75454
rect 300688 75134 301008 75218
rect 300688 74898 300730 75134
rect 300966 74898 301008 75134
rect 300688 74866 301008 74898
rect 331408 75454 331728 75486
rect 331408 75218 331450 75454
rect 331686 75218 331728 75454
rect 331408 75134 331728 75218
rect 331408 74898 331450 75134
rect 331686 74898 331728 75134
rect 331408 74866 331728 74898
rect 361794 75454 362414 110898
rect 361794 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 362414 75454
rect 361794 75134 362414 75218
rect 361794 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 362414 75134
rect 27834 65258 27866 65494
rect 28102 65258 28186 65494
rect 28422 65258 28454 65494
rect 27834 65174 28454 65258
rect 27834 64938 27866 65174
rect 28102 64938 28186 65174
rect 28422 64938 28454 65174
rect 22139 49604 22205 49605
rect 22139 49540 22140 49604
rect 22204 49540 22205 49604
rect 22139 49539 22205 49540
rect 22142 46613 22202 49539
rect 22323 48924 22389 48925
rect 22323 48860 22324 48924
rect 22388 48860 22389 48924
rect 22323 48859 22389 48860
rect 22139 46612 22205 46613
rect 22139 46548 22140 46612
rect 22204 46548 22205 46612
rect 22139 46547 22205 46548
rect 22326 46477 22386 48859
rect 22323 46476 22389 46477
rect 22323 46412 22324 46476
rect 22388 46412 22389 46476
rect 22323 46411 22389 46412
rect 20394 21818 20426 22054
rect 20662 21818 20746 22054
rect 20982 21818 21014 22054
rect 20394 21734 21014 21818
rect 20394 21498 20426 21734
rect 20662 21498 20746 21734
rect 20982 21498 21014 21734
rect 20394 -5146 21014 21498
rect 20394 -5382 20426 -5146
rect 20662 -5382 20746 -5146
rect 20982 -5382 21014 -5146
rect 20394 -5466 21014 -5382
rect 20394 -5702 20426 -5466
rect 20662 -5702 20746 -5466
rect 20982 -5702 21014 -5466
rect 20394 -7654 21014 -5702
rect 24114 25774 24734 45068
rect 24114 25538 24146 25774
rect 24382 25538 24466 25774
rect 24702 25538 24734 25774
rect 24114 25454 24734 25538
rect 24114 25218 24146 25454
rect 24382 25218 24466 25454
rect 24702 25218 24734 25454
rect 24114 -6106 24734 25218
rect 24114 -6342 24146 -6106
rect 24382 -6342 24466 -6106
rect 24702 -6342 24734 -6106
rect 24114 -6426 24734 -6342
rect 24114 -6662 24146 -6426
rect 24382 -6662 24466 -6426
rect 24702 -6662 24734 -6426
rect 24114 -7654 24734 -6662
rect 27834 29494 28454 64938
rect 27834 29258 27866 29494
rect 28102 29258 28186 29494
rect 28422 29258 28454 29494
rect 27834 29174 28454 29258
rect 27834 28938 27866 29174
rect 28102 28938 28186 29174
rect 28422 28938 28454 29174
rect 27834 -7066 28454 28938
rect 27834 -7302 27866 -7066
rect 28102 -7302 28186 -7066
rect 28422 -7302 28454 -7066
rect 27834 -7386 28454 -7302
rect 27834 -7622 27866 -7386
rect 28102 -7622 28186 -7386
rect 28422 -7622 28454 -7386
rect 27834 -7654 28454 -7622
rect 37794 39454 38414 49367
rect 37794 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 38414 39454
rect 37794 39134 38414 39218
rect 37794 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 38414 39134
rect 37794 3454 38414 38898
rect 37794 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 38414 3454
rect 37794 3134 38414 3218
rect 37794 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 38414 3134
rect 37794 -346 38414 2898
rect 37794 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 38414 -346
rect 37794 -666 38414 -582
rect 37794 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 38414 -666
rect 37794 -7654 38414 -902
rect 41514 43174 42134 49367
rect 41514 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 42134 43174
rect 41514 42854 42134 42938
rect 41514 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 42134 42854
rect 41514 7174 42134 42618
rect 41514 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 42134 7174
rect 41514 6854 42134 6938
rect 41514 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 42134 6854
rect 41514 -1306 42134 6618
rect 41514 -1542 41546 -1306
rect 41782 -1542 41866 -1306
rect 42102 -1542 42134 -1306
rect 41514 -1626 42134 -1542
rect 41514 -1862 41546 -1626
rect 41782 -1862 41866 -1626
rect 42102 -1862 42134 -1626
rect 41514 -7654 42134 -1862
rect 45234 46894 45854 49367
rect 45234 46658 45266 46894
rect 45502 46658 45586 46894
rect 45822 46658 45854 46894
rect 45234 46574 45854 46658
rect 45234 46338 45266 46574
rect 45502 46338 45586 46574
rect 45822 46338 45854 46574
rect 45234 10894 45854 46338
rect 45234 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 45854 10894
rect 45234 10574 45854 10658
rect 45234 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 45854 10574
rect 45234 -2266 45854 10338
rect 45234 -2502 45266 -2266
rect 45502 -2502 45586 -2266
rect 45822 -2502 45854 -2266
rect 45234 -2586 45854 -2502
rect 45234 -2822 45266 -2586
rect 45502 -2822 45586 -2586
rect 45822 -2822 45854 -2586
rect 45234 -7654 45854 -2822
rect 48954 14614 49574 49367
rect 48954 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 49574 14614
rect 48954 14294 49574 14378
rect 48954 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 49574 14294
rect 48954 -3226 49574 14058
rect 48954 -3462 48986 -3226
rect 49222 -3462 49306 -3226
rect 49542 -3462 49574 -3226
rect 48954 -3546 49574 -3462
rect 48954 -3782 48986 -3546
rect 49222 -3782 49306 -3546
rect 49542 -3782 49574 -3546
rect 48954 -7654 49574 -3782
rect 52674 18334 53294 49367
rect 52674 18098 52706 18334
rect 52942 18098 53026 18334
rect 53262 18098 53294 18334
rect 52674 18014 53294 18098
rect 52674 17778 52706 18014
rect 52942 17778 53026 18014
rect 53262 17778 53294 18014
rect 52674 -4186 53294 17778
rect 52674 -4422 52706 -4186
rect 52942 -4422 53026 -4186
rect 53262 -4422 53294 -4186
rect 52674 -4506 53294 -4422
rect 52674 -4742 52706 -4506
rect 52942 -4742 53026 -4506
rect 53262 -4742 53294 -4506
rect 52674 -7654 53294 -4742
rect 56394 22054 57014 49367
rect 56394 21818 56426 22054
rect 56662 21818 56746 22054
rect 56982 21818 57014 22054
rect 56394 21734 57014 21818
rect 56394 21498 56426 21734
rect 56662 21498 56746 21734
rect 56982 21498 57014 21734
rect 56394 -5146 57014 21498
rect 56394 -5382 56426 -5146
rect 56662 -5382 56746 -5146
rect 56982 -5382 57014 -5146
rect 56394 -5466 57014 -5382
rect 56394 -5702 56426 -5466
rect 56662 -5702 56746 -5466
rect 56982 -5702 57014 -5466
rect 56394 -7654 57014 -5702
rect 60114 25774 60734 49367
rect 60114 25538 60146 25774
rect 60382 25538 60466 25774
rect 60702 25538 60734 25774
rect 60114 25454 60734 25538
rect 60114 25218 60146 25454
rect 60382 25218 60466 25454
rect 60702 25218 60734 25454
rect 60114 -6106 60734 25218
rect 60114 -6342 60146 -6106
rect 60382 -6342 60466 -6106
rect 60702 -6342 60734 -6106
rect 60114 -6426 60734 -6342
rect 60114 -6662 60146 -6426
rect 60382 -6662 60466 -6426
rect 60702 -6662 60734 -6426
rect 60114 -7654 60734 -6662
rect 63834 29494 64454 49367
rect 63834 29258 63866 29494
rect 64102 29258 64186 29494
rect 64422 29258 64454 29494
rect 63834 29174 64454 29258
rect 63834 28938 63866 29174
rect 64102 28938 64186 29174
rect 64422 28938 64454 29174
rect 63834 -7066 64454 28938
rect 63834 -7302 63866 -7066
rect 64102 -7302 64186 -7066
rect 64422 -7302 64454 -7066
rect 63834 -7386 64454 -7302
rect 63834 -7622 63866 -7386
rect 64102 -7622 64186 -7386
rect 64422 -7622 64454 -7386
rect 63834 -7654 64454 -7622
rect 73794 39454 74414 49367
rect 73794 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 74414 39454
rect 73794 39134 74414 39218
rect 73794 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 74414 39134
rect 73794 3454 74414 38898
rect 73794 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 74414 3454
rect 73794 3134 74414 3218
rect 73794 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 74414 3134
rect 73794 -346 74414 2898
rect 73794 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 74414 -346
rect 73794 -666 74414 -582
rect 73794 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 74414 -666
rect 73794 -7654 74414 -902
rect 77514 43174 78134 49367
rect 77514 42938 77546 43174
rect 77782 42938 77866 43174
rect 78102 42938 78134 43174
rect 77514 42854 78134 42938
rect 77514 42618 77546 42854
rect 77782 42618 77866 42854
rect 78102 42618 78134 42854
rect 77514 7174 78134 42618
rect 77514 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 78134 7174
rect 77514 6854 78134 6938
rect 77514 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 78134 6854
rect 77514 -1306 78134 6618
rect 77514 -1542 77546 -1306
rect 77782 -1542 77866 -1306
rect 78102 -1542 78134 -1306
rect 77514 -1626 78134 -1542
rect 77514 -1862 77546 -1626
rect 77782 -1862 77866 -1626
rect 78102 -1862 78134 -1626
rect 77514 -7654 78134 -1862
rect 81234 46894 81854 49367
rect 81234 46658 81266 46894
rect 81502 46658 81586 46894
rect 81822 46658 81854 46894
rect 81234 46574 81854 46658
rect 81234 46338 81266 46574
rect 81502 46338 81586 46574
rect 81822 46338 81854 46574
rect 81234 10894 81854 46338
rect 81234 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 81854 10894
rect 81234 10574 81854 10658
rect 81234 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 81854 10574
rect 81234 -2266 81854 10338
rect 81234 -2502 81266 -2266
rect 81502 -2502 81586 -2266
rect 81822 -2502 81854 -2266
rect 81234 -2586 81854 -2502
rect 81234 -2822 81266 -2586
rect 81502 -2822 81586 -2586
rect 81822 -2822 81854 -2586
rect 81234 -7654 81854 -2822
rect 84954 14614 85574 49367
rect 84954 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 85574 14614
rect 84954 14294 85574 14378
rect 84954 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 85574 14294
rect 84954 -3226 85574 14058
rect 84954 -3462 84986 -3226
rect 85222 -3462 85306 -3226
rect 85542 -3462 85574 -3226
rect 84954 -3546 85574 -3462
rect 84954 -3782 84986 -3546
rect 85222 -3782 85306 -3546
rect 85542 -3782 85574 -3546
rect 84954 -7654 85574 -3782
rect 88674 18334 89294 49367
rect 88674 18098 88706 18334
rect 88942 18098 89026 18334
rect 89262 18098 89294 18334
rect 88674 18014 89294 18098
rect 88674 17778 88706 18014
rect 88942 17778 89026 18014
rect 89262 17778 89294 18014
rect 88674 -4186 89294 17778
rect 88674 -4422 88706 -4186
rect 88942 -4422 89026 -4186
rect 89262 -4422 89294 -4186
rect 88674 -4506 89294 -4422
rect 88674 -4742 88706 -4506
rect 88942 -4742 89026 -4506
rect 89262 -4742 89294 -4506
rect 88674 -7654 89294 -4742
rect 92394 22054 93014 49367
rect 92394 21818 92426 22054
rect 92662 21818 92746 22054
rect 92982 21818 93014 22054
rect 92394 21734 93014 21818
rect 92394 21498 92426 21734
rect 92662 21498 92746 21734
rect 92982 21498 93014 21734
rect 92394 -5146 93014 21498
rect 92394 -5382 92426 -5146
rect 92662 -5382 92746 -5146
rect 92982 -5382 93014 -5146
rect 92394 -5466 93014 -5382
rect 92394 -5702 92426 -5466
rect 92662 -5702 92746 -5466
rect 92982 -5702 93014 -5466
rect 92394 -7654 93014 -5702
rect 96114 25774 96734 49367
rect 96114 25538 96146 25774
rect 96382 25538 96466 25774
rect 96702 25538 96734 25774
rect 96114 25454 96734 25538
rect 96114 25218 96146 25454
rect 96382 25218 96466 25454
rect 96702 25218 96734 25454
rect 96114 -6106 96734 25218
rect 96114 -6342 96146 -6106
rect 96382 -6342 96466 -6106
rect 96702 -6342 96734 -6106
rect 96114 -6426 96734 -6342
rect 96114 -6662 96146 -6426
rect 96382 -6662 96466 -6426
rect 96702 -6662 96734 -6426
rect 96114 -7654 96734 -6662
rect 99834 29494 100454 49367
rect 99834 29258 99866 29494
rect 100102 29258 100186 29494
rect 100422 29258 100454 29494
rect 99834 29174 100454 29258
rect 99834 28938 99866 29174
rect 100102 28938 100186 29174
rect 100422 28938 100454 29174
rect 99834 -7066 100454 28938
rect 99834 -7302 99866 -7066
rect 100102 -7302 100186 -7066
rect 100422 -7302 100454 -7066
rect 99834 -7386 100454 -7302
rect 99834 -7622 99866 -7386
rect 100102 -7622 100186 -7386
rect 100422 -7622 100454 -7386
rect 99834 -7654 100454 -7622
rect 109794 39454 110414 49367
rect 109794 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 110414 39454
rect 109794 39134 110414 39218
rect 109794 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 110414 39134
rect 109794 3454 110414 38898
rect 109794 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 110414 3454
rect 109794 3134 110414 3218
rect 109794 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 110414 3134
rect 109794 -346 110414 2898
rect 109794 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 110414 -346
rect 109794 -666 110414 -582
rect 109794 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 110414 -666
rect 109794 -7654 110414 -902
rect 113514 43174 114134 49367
rect 113514 42938 113546 43174
rect 113782 42938 113866 43174
rect 114102 42938 114134 43174
rect 113514 42854 114134 42938
rect 113514 42618 113546 42854
rect 113782 42618 113866 42854
rect 114102 42618 114134 42854
rect 113514 7174 114134 42618
rect 113514 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 114134 7174
rect 113514 6854 114134 6938
rect 113514 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 114134 6854
rect 113514 -1306 114134 6618
rect 113514 -1542 113546 -1306
rect 113782 -1542 113866 -1306
rect 114102 -1542 114134 -1306
rect 113514 -1626 114134 -1542
rect 113514 -1862 113546 -1626
rect 113782 -1862 113866 -1626
rect 114102 -1862 114134 -1626
rect 113514 -7654 114134 -1862
rect 117234 46894 117854 49367
rect 117234 46658 117266 46894
rect 117502 46658 117586 46894
rect 117822 46658 117854 46894
rect 117234 46574 117854 46658
rect 117234 46338 117266 46574
rect 117502 46338 117586 46574
rect 117822 46338 117854 46574
rect 117234 10894 117854 46338
rect 117234 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 117854 10894
rect 117234 10574 117854 10658
rect 117234 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 117854 10574
rect 117234 -2266 117854 10338
rect 117234 -2502 117266 -2266
rect 117502 -2502 117586 -2266
rect 117822 -2502 117854 -2266
rect 117234 -2586 117854 -2502
rect 117234 -2822 117266 -2586
rect 117502 -2822 117586 -2586
rect 117822 -2822 117854 -2586
rect 117234 -7654 117854 -2822
rect 120954 14614 121574 49367
rect 120954 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 121574 14614
rect 120954 14294 121574 14378
rect 120954 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 121574 14294
rect 120954 -3226 121574 14058
rect 120954 -3462 120986 -3226
rect 121222 -3462 121306 -3226
rect 121542 -3462 121574 -3226
rect 120954 -3546 121574 -3462
rect 120954 -3782 120986 -3546
rect 121222 -3782 121306 -3546
rect 121542 -3782 121574 -3546
rect 120954 -7654 121574 -3782
rect 124674 18334 125294 49367
rect 124674 18098 124706 18334
rect 124942 18098 125026 18334
rect 125262 18098 125294 18334
rect 124674 18014 125294 18098
rect 124674 17778 124706 18014
rect 124942 17778 125026 18014
rect 125262 17778 125294 18014
rect 124674 -4186 125294 17778
rect 124674 -4422 124706 -4186
rect 124942 -4422 125026 -4186
rect 125262 -4422 125294 -4186
rect 124674 -4506 125294 -4422
rect 124674 -4742 124706 -4506
rect 124942 -4742 125026 -4506
rect 125262 -4742 125294 -4506
rect 124674 -7654 125294 -4742
rect 128394 22054 129014 49367
rect 128394 21818 128426 22054
rect 128662 21818 128746 22054
rect 128982 21818 129014 22054
rect 128394 21734 129014 21818
rect 128394 21498 128426 21734
rect 128662 21498 128746 21734
rect 128982 21498 129014 21734
rect 128394 -5146 129014 21498
rect 128394 -5382 128426 -5146
rect 128662 -5382 128746 -5146
rect 128982 -5382 129014 -5146
rect 128394 -5466 129014 -5382
rect 128394 -5702 128426 -5466
rect 128662 -5702 128746 -5466
rect 128982 -5702 129014 -5466
rect 128394 -7654 129014 -5702
rect 132114 25774 132734 49367
rect 132114 25538 132146 25774
rect 132382 25538 132466 25774
rect 132702 25538 132734 25774
rect 132114 25454 132734 25538
rect 132114 25218 132146 25454
rect 132382 25218 132466 25454
rect 132702 25218 132734 25454
rect 132114 -6106 132734 25218
rect 132114 -6342 132146 -6106
rect 132382 -6342 132466 -6106
rect 132702 -6342 132734 -6106
rect 132114 -6426 132734 -6342
rect 132114 -6662 132146 -6426
rect 132382 -6662 132466 -6426
rect 132702 -6662 132734 -6426
rect 132114 -7654 132734 -6662
rect 135834 29494 136454 49367
rect 135834 29258 135866 29494
rect 136102 29258 136186 29494
rect 136422 29258 136454 29494
rect 135834 29174 136454 29258
rect 135834 28938 135866 29174
rect 136102 28938 136186 29174
rect 136422 28938 136454 29174
rect 135834 -7066 136454 28938
rect 135834 -7302 135866 -7066
rect 136102 -7302 136186 -7066
rect 136422 -7302 136454 -7066
rect 135834 -7386 136454 -7302
rect 135834 -7622 135866 -7386
rect 136102 -7622 136186 -7386
rect 136422 -7622 136454 -7386
rect 135834 -7654 136454 -7622
rect 145794 39454 146414 49367
rect 145794 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 146414 39454
rect 145794 39134 146414 39218
rect 145794 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 146414 39134
rect 145794 3454 146414 38898
rect 145794 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 146414 3454
rect 145794 3134 146414 3218
rect 145794 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 146414 3134
rect 145794 -346 146414 2898
rect 145794 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 146414 -346
rect 145794 -666 146414 -582
rect 145794 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 146414 -666
rect 145794 -7654 146414 -902
rect 149514 43174 150134 49367
rect 149514 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 150134 43174
rect 149514 42854 150134 42938
rect 149514 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 150134 42854
rect 149514 7174 150134 42618
rect 149514 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 150134 7174
rect 149514 6854 150134 6938
rect 149514 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 150134 6854
rect 149514 -1306 150134 6618
rect 149514 -1542 149546 -1306
rect 149782 -1542 149866 -1306
rect 150102 -1542 150134 -1306
rect 149514 -1626 150134 -1542
rect 149514 -1862 149546 -1626
rect 149782 -1862 149866 -1626
rect 150102 -1862 150134 -1626
rect 149514 -7654 150134 -1862
rect 153234 46894 153854 49367
rect 153234 46658 153266 46894
rect 153502 46658 153586 46894
rect 153822 46658 153854 46894
rect 153234 46574 153854 46658
rect 153234 46338 153266 46574
rect 153502 46338 153586 46574
rect 153822 46338 153854 46574
rect 153234 10894 153854 46338
rect 153234 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 153854 10894
rect 153234 10574 153854 10658
rect 153234 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 153854 10574
rect 153234 -2266 153854 10338
rect 153234 -2502 153266 -2266
rect 153502 -2502 153586 -2266
rect 153822 -2502 153854 -2266
rect 153234 -2586 153854 -2502
rect 153234 -2822 153266 -2586
rect 153502 -2822 153586 -2586
rect 153822 -2822 153854 -2586
rect 153234 -7654 153854 -2822
rect 156954 14614 157574 49367
rect 156954 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 157574 14614
rect 156954 14294 157574 14378
rect 156954 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 157574 14294
rect 156954 -3226 157574 14058
rect 156954 -3462 156986 -3226
rect 157222 -3462 157306 -3226
rect 157542 -3462 157574 -3226
rect 156954 -3546 157574 -3462
rect 156954 -3782 156986 -3546
rect 157222 -3782 157306 -3546
rect 157542 -3782 157574 -3546
rect 156954 -7654 157574 -3782
rect 160674 18334 161294 49367
rect 160674 18098 160706 18334
rect 160942 18098 161026 18334
rect 161262 18098 161294 18334
rect 160674 18014 161294 18098
rect 160674 17778 160706 18014
rect 160942 17778 161026 18014
rect 161262 17778 161294 18014
rect 160674 -4186 161294 17778
rect 160674 -4422 160706 -4186
rect 160942 -4422 161026 -4186
rect 161262 -4422 161294 -4186
rect 160674 -4506 161294 -4422
rect 160674 -4742 160706 -4506
rect 160942 -4742 161026 -4506
rect 161262 -4742 161294 -4506
rect 160674 -7654 161294 -4742
rect 164394 22054 165014 49367
rect 164394 21818 164426 22054
rect 164662 21818 164746 22054
rect 164982 21818 165014 22054
rect 164394 21734 165014 21818
rect 164394 21498 164426 21734
rect 164662 21498 164746 21734
rect 164982 21498 165014 21734
rect 164394 -5146 165014 21498
rect 164394 -5382 164426 -5146
rect 164662 -5382 164746 -5146
rect 164982 -5382 165014 -5146
rect 164394 -5466 165014 -5382
rect 164394 -5702 164426 -5466
rect 164662 -5702 164746 -5466
rect 164982 -5702 165014 -5466
rect 164394 -7654 165014 -5702
rect 168114 25774 168734 49367
rect 168114 25538 168146 25774
rect 168382 25538 168466 25774
rect 168702 25538 168734 25774
rect 168114 25454 168734 25538
rect 168114 25218 168146 25454
rect 168382 25218 168466 25454
rect 168702 25218 168734 25454
rect 168114 -6106 168734 25218
rect 168114 -6342 168146 -6106
rect 168382 -6342 168466 -6106
rect 168702 -6342 168734 -6106
rect 168114 -6426 168734 -6342
rect 168114 -6662 168146 -6426
rect 168382 -6662 168466 -6426
rect 168702 -6662 168734 -6426
rect 168114 -7654 168734 -6662
rect 171834 29494 172454 49367
rect 171834 29258 171866 29494
rect 172102 29258 172186 29494
rect 172422 29258 172454 29494
rect 171834 29174 172454 29258
rect 171834 28938 171866 29174
rect 172102 28938 172186 29174
rect 172422 28938 172454 29174
rect 171834 -7066 172454 28938
rect 171834 -7302 171866 -7066
rect 172102 -7302 172186 -7066
rect 172422 -7302 172454 -7066
rect 171834 -7386 172454 -7302
rect 171834 -7622 171866 -7386
rect 172102 -7622 172186 -7386
rect 172422 -7622 172454 -7386
rect 171834 -7654 172454 -7622
rect 181794 39454 182414 49367
rect 181794 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 182414 39454
rect 181794 39134 182414 39218
rect 181794 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 182414 39134
rect 181794 3454 182414 38898
rect 181794 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 182414 3454
rect 181794 3134 182414 3218
rect 181794 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 182414 3134
rect 181794 -346 182414 2898
rect 181794 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 182414 -346
rect 181794 -666 182414 -582
rect 181794 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 182414 -666
rect 181794 -7654 182414 -902
rect 185514 43174 186134 49367
rect 185514 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 186134 43174
rect 185514 42854 186134 42938
rect 185514 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 186134 42854
rect 185514 7174 186134 42618
rect 185514 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 186134 7174
rect 185514 6854 186134 6938
rect 185514 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 186134 6854
rect 185514 -1306 186134 6618
rect 185514 -1542 185546 -1306
rect 185782 -1542 185866 -1306
rect 186102 -1542 186134 -1306
rect 185514 -1626 186134 -1542
rect 185514 -1862 185546 -1626
rect 185782 -1862 185866 -1626
rect 186102 -1862 186134 -1626
rect 185514 -7654 186134 -1862
rect 189234 46894 189854 49367
rect 189234 46658 189266 46894
rect 189502 46658 189586 46894
rect 189822 46658 189854 46894
rect 189234 46574 189854 46658
rect 189234 46338 189266 46574
rect 189502 46338 189586 46574
rect 189822 46338 189854 46574
rect 189234 10894 189854 46338
rect 189234 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 189854 10894
rect 189234 10574 189854 10658
rect 189234 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 189854 10574
rect 189234 -2266 189854 10338
rect 189234 -2502 189266 -2266
rect 189502 -2502 189586 -2266
rect 189822 -2502 189854 -2266
rect 189234 -2586 189854 -2502
rect 189234 -2822 189266 -2586
rect 189502 -2822 189586 -2586
rect 189822 -2822 189854 -2586
rect 189234 -7654 189854 -2822
rect 192954 14614 193574 45068
rect 192954 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 193574 14614
rect 192954 14294 193574 14378
rect 192954 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 193574 14294
rect 192954 -3226 193574 14058
rect 192954 -3462 192986 -3226
rect 193222 -3462 193306 -3226
rect 193542 -3462 193574 -3226
rect 192954 -3546 193574 -3462
rect 192954 -3782 192986 -3546
rect 193222 -3782 193306 -3546
rect 193542 -3782 193574 -3546
rect 192954 -7654 193574 -3782
rect 196674 18334 197294 49367
rect 196674 18098 196706 18334
rect 196942 18098 197026 18334
rect 197262 18098 197294 18334
rect 196674 18014 197294 18098
rect 196674 17778 196706 18014
rect 196942 17778 197026 18014
rect 197262 17778 197294 18014
rect 196674 -4186 197294 17778
rect 196674 -4422 196706 -4186
rect 196942 -4422 197026 -4186
rect 197262 -4422 197294 -4186
rect 196674 -4506 197294 -4422
rect 196674 -4742 196706 -4506
rect 196942 -4742 197026 -4506
rect 197262 -4742 197294 -4506
rect 196674 -7654 197294 -4742
rect 200394 22054 201014 49367
rect 200394 21818 200426 22054
rect 200662 21818 200746 22054
rect 200982 21818 201014 22054
rect 200394 21734 201014 21818
rect 200394 21498 200426 21734
rect 200662 21498 200746 21734
rect 200982 21498 201014 21734
rect 200394 -5146 201014 21498
rect 200394 -5382 200426 -5146
rect 200662 -5382 200746 -5146
rect 200982 -5382 201014 -5146
rect 200394 -5466 201014 -5382
rect 200394 -5702 200426 -5466
rect 200662 -5702 200746 -5466
rect 200982 -5702 201014 -5466
rect 200394 -7654 201014 -5702
rect 204114 25774 204734 49367
rect 204114 25538 204146 25774
rect 204382 25538 204466 25774
rect 204702 25538 204734 25774
rect 204114 25454 204734 25538
rect 204114 25218 204146 25454
rect 204382 25218 204466 25454
rect 204702 25218 204734 25454
rect 204114 -6106 204734 25218
rect 204114 -6342 204146 -6106
rect 204382 -6342 204466 -6106
rect 204702 -6342 204734 -6106
rect 204114 -6426 204734 -6342
rect 204114 -6662 204146 -6426
rect 204382 -6662 204466 -6426
rect 204702 -6662 204734 -6426
rect 204114 -7654 204734 -6662
rect 207834 29494 208454 49367
rect 207834 29258 207866 29494
rect 208102 29258 208186 29494
rect 208422 29258 208454 29494
rect 207834 29174 208454 29258
rect 207834 28938 207866 29174
rect 208102 28938 208186 29174
rect 208422 28938 208454 29174
rect 207834 -7066 208454 28938
rect 207834 -7302 207866 -7066
rect 208102 -7302 208186 -7066
rect 208422 -7302 208454 -7066
rect 207834 -7386 208454 -7302
rect 207834 -7622 207866 -7386
rect 208102 -7622 208186 -7386
rect 208422 -7622 208454 -7386
rect 207834 -7654 208454 -7622
rect 217794 39454 218414 49367
rect 217794 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 218414 39454
rect 217794 39134 218414 39218
rect 217794 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 218414 39134
rect 217794 3454 218414 38898
rect 217794 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 218414 3454
rect 217794 3134 218414 3218
rect 217794 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 218414 3134
rect 217794 -346 218414 2898
rect 217794 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 218414 -346
rect 217794 -666 218414 -582
rect 217794 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 218414 -666
rect 217794 -7654 218414 -902
rect 221514 43174 222134 49367
rect 221514 42938 221546 43174
rect 221782 42938 221866 43174
rect 222102 42938 222134 43174
rect 221514 42854 222134 42938
rect 221514 42618 221546 42854
rect 221782 42618 221866 42854
rect 222102 42618 222134 42854
rect 221514 7174 222134 42618
rect 221514 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 222134 7174
rect 221514 6854 222134 6938
rect 221514 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 222134 6854
rect 221514 -1306 222134 6618
rect 221514 -1542 221546 -1306
rect 221782 -1542 221866 -1306
rect 222102 -1542 222134 -1306
rect 221514 -1626 222134 -1542
rect 221514 -1862 221546 -1626
rect 221782 -1862 221866 -1626
rect 222102 -1862 222134 -1626
rect 221514 -7654 222134 -1862
rect 225234 46894 225854 49367
rect 225234 46658 225266 46894
rect 225502 46658 225586 46894
rect 225822 46658 225854 46894
rect 225234 46574 225854 46658
rect 225234 46338 225266 46574
rect 225502 46338 225586 46574
rect 225822 46338 225854 46574
rect 225234 10894 225854 46338
rect 225234 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 225854 10894
rect 225234 10574 225854 10658
rect 225234 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 225854 10574
rect 225234 -2266 225854 10338
rect 225234 -2502 225266 -2266
rect 225502 -2502 225586 -2266
rect 225822 -2502 225854 -2266
rect 225234 -2586 225854 -2502
rect 225234 -2822 225266 -2586
rect 225502 -2822 225586 -2586
rect 225822 -2822 225854 -2586
rect 225234 -7654 225854 -2822
rect 228954 14614 229574 49367
rect 228954 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 229574 14614
rect 228954 14294 229574 14378
rect 228954 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 229574 14294
rect 228954 -3226 229574 14058
rect 228954 -3462 228986 -3226
rect 229222 -3462 229306 -3226
rect 229542 -3462 229574 -3226
rect 228954 -3546 229574 -3462
rect 228954 -3782 228986 -3546
rect 229222 -3782 229306 -3546
rect 229542 -3782 229574 -3546
rect 228954 -7654 229574 -3782
rect 232674 18334 233294 49367
rect 232674 18098 232706 18334
rect 232942 18098 233026 18334
rect 233262 18098 233294 18334
rect 232674 18014 233294 18098
rect 232674 17778 232706 18014
rect 232942 17778 233026 18014
rect 233262 17778 233294 18014
rect 232674 -4186 233294 17778
rect 232674 -4422 232706 -4186
rect 232942 -4422 233026 -4186
rect 233262 -4422 233294 -4186
rect 232674 -4506 233294 -4422
rect 232674 -4742 232706 -4506
rect 232942 -4742 233026 -4506
rect 233262 -4742 233294 -4506
rect 232674 -7654 233294 -4742
rect 236394 22054 237014 49367
rect 236394 21818 236426 22054
rect 236662 21818 236746 22054
rect 236982 21818 237014 22054
rect 236394 21734 237014 21818
rect 236394 21498 236426 21734
rect 236662 21498 236746 21734
rect 236982 21498 237014 21734
rect 236394 -5146 237014 21498
rect 236394 -5382 236426 -5146
rect 236662 -5382 236746 -5146
rect 236982 -5382 237014 -5146
rect 236394 -5466 237014 -5382
rect 236394 -5702 236426 -5466
rect 236662 -5702 236746 -5466
rect 236982 -5702 237014 -5466
rect 236394 -7654 237014 -5702
rect 240114 25774 240734 49367
rect 240114 25538 240146 25774
rect 240382 25538 240466 25774
rect 240702 25538 240734 25774
rect 240114 25454 240734 25538
rect 240114 25218 240146 25454
rect 240382 25218 240466 25454
rect 240702 25218 240734 25454
rect 240114 -6106 240734 25218
rect 240114 -6342 240146 -6106
rect 240382 -6342 240466 -6106
rect 240702 -6342 240734 -6106
rect 240114 -6426 240734 -6342
rect 240114 -6662 240146 -6426
rect 240382 -6662 240466 -6426
rect 240702 -6662 240734 -6426
rect 240114 -7654 240734 -6662
rect 243834 29494 244454 49367
rect 243834 29258 243866 29494
rect 244102 29258 244186 29494
rect 244422 29258 244454 29494
rect 243834 29174 244454 29258
rect 243834 28938 243866 29174
rect 244102 28938 244186 29174
rect 244422 28938 244454 29174
rect 243834 -7066 244454 28938
rect 243834 -7302 243866 -7066
rect 244102 -7302 244186 -7066
rect 244422 -7302 244454 -7066
rect 243834 -7386 244454 -7302
rect 243834 -7622 243866 -7386
rect 244102 -7622 244186 -7386
rect 244422 -7622 244454 -7386
rect 243834 -7654 244454 -7622
rect 253794 39454 254414 49367
rect 253794 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 254414 39454
rect 253794 39134 254414 39218
rect 253794 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 254414 39134
rect 253794 3454 254414 38898
rect 253794 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 254414 3454
rect 253794 3134 254414 3218
rect 253794 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 254414 3134
rect 253794 -346 254414 2898
rect 253794 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 254414 -346
rect 253794 -666 254414 -582
rect 253794 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 254414 -666
rect 253794 -7654 254414 -902
rect 257514 43174 258134 49367
rect 257514 42938 257546 43174
rect 257782 42938 257866 43174
rect 258102 42938 258134 43174
rect 257514 42854 258134 42938
rect 257514 42618 257546 42854
rect 257782 42618 257866 42854
rect 258102 42618 258134 42854
rect 257514 7174 258134 42618
rect 257514 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 258134 7174
rect 257514 6854 258134 6938
rect 257514 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 258134 6854
rect 257514 -1306 258134 6618
rect 257514 -1542 257546 -1306
rect 257782 -1542 257866 -1306
rect 258102 -1542 258134 -1306
rect 257514 -1626 258134 -1542
rect 257514 -1862 257546 -1626
rect 257782 -1862 257866 -1626
rect 258102 -1862 258134 -1626
rect 257514 -7654 258134 -1862
rect 261234 46894 261854 49367
rect 261234 46658 261266 46894
rect 261502 46658 261586 46894
rect 261822 46658 261854 46894
rect 261234 46574 261854 46658
rect 261234 46338 261266 46574
rect 261502 46338 261586 46574
rect 261822 46338 261854 46574
rect 261234 10894 261854 46338
rect 261234 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 261854 10894
rect 261234 10574 261854 10658
rect 261234 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 261854 10574
rect 261234 -2266 261854 10338
rect 261234 -2502 261266 -2266
rect 261502 -2502 261586 -2266
rect 261822 -2502 261854 -2266
rect 261234 -2586 261854 -2502
rect 261234 -2822 261266 -2586
rect 261502 -2822 261586 -2586
rect 261822 -2822 261854 -2586
rect 261234 -7654 261854 -2822
rect 264954 14614 265574 49367
rect 264954 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 265574 14614
rect 264954 14294 265574 14378
rect 264954 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 265574 14294
rect 264954 -3226 265574 14058
rect 264954 -3462 264986 -3226
rect 265222 -3462 265306 -3226
rect 265542 -3462 265574 -3226
rect 264954 -3546 265574 -3462
rect 264954 -3782 264986 -3546
rect 265222 -3782 265306 -3546
rect 265542 -3782 265574 -3546
rect 264954 -7654 265574 -3782
rect 268674 18334 269294 49367
rect 268674 18098 268706 18334
rect 268942 18098 269026 18334
rect 269262 18098 269294 18334
rect 268674 18014 269294 18098
rect 268674 17778 268706 18014
rect 268942 17778 269026 18014
rect 269262 17778 269294 18014
rect 268674 -4186 269294 17778
rect 268674 -4422 268706 -4186
rect 268942 -4422 269026 -4186
rect 269262 -4422 269294 -4186
rect 268674 -4506 269294 -4422
rect 268674 -4742 268706 -4506
rect 268942 -4742 269026 -4506
rect 269262 -4742 269294 -4506
rect 268674 -7654 269294 -4742
rect 272394 22054 273014 49367
rect 272394 21818 272426 22054
rect 272662 21818 272746 22054
rect 272982 21818 273014 22054
rect 272394 21734 273014 21818
rect 272394 21498 272426 21734
rect 272662 21498 272746 21734
rect 272982 21498 273014 21734
rect 272394 -5146 273014 21498
rect 272394 -5382 272426 -5146
rect 272662 -5382 272746 -5146
rect 272982 -5382 273014 -5146
rect 272394 -5466 273014 -5382
rect 272394 -5702 272426 -5466
rect 272662 -5702 272746 -5466
rect 272982 -5702 273014 -5466
rect 272394 -7654 273014 -5702
rect 276114 25774 276734 49367
rect 276114 25538 276146 25774
rect 276382 25538 276466 25774
rect 276702 25538 276734 25774
rect 276114 25454 276734 25538
rect 276114 25218 276146 25454
rect 276382 25218 276466 25454
rect 276702 25218 276734 25454
rect 276114 -6106 276734 25218
rect 276114 -6342 276146 -6106
rect 276382 -6342 276466 -6106
rect 276702 -6342 276734 -6106
rect 276114 -6426 276734 -6342
rect 276114 -6662 276146 -6426
rect 276382 -6662 276466 -6426
rect 276702 -6662 276734 -6426
rect 276114 -7654 276734 -6662
rect 279834 29494 280454 49367
rect 279834 29258 279866 29494
rect 280102 29258 280186 29494
rect 280422 29258 280454 29494
rect 279834 29174 280454 29258
rect 279834 28938 279866 29174
rect 280102 28938 280186 29174
rect 280422 28938 280454 29174
rect 279834 -7066 280454 28938
rect 279834 -7302 279866 -7066
rect 280102 -7302 280186 -7066
rect 280422 -7302 280454 -7066
rect 279834 -7386 280454 -7302
rect 279834 -7622 279866 -7386
rect 280102 -7622 280186 -7386
rect 280422 -7622 280454 -7386
rect 279834 -7654 280454 -7622
rect 289794 39454 290414 49367
rect 289794 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 290414 39454
rect 289794 39134 290414 39218
rect 289794 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 290414 39134
rect 289794 3454 290414 38898
rect 289794 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 290414 3454
rect 289794 3134 290414 3218
rect 289794 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 290414 3134
rect 289794 -346 290414 2898
rect 289794 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 290414 -346
rect 289794 -666 290414 -582
rect 289794 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 290414 -666
rect 289794 -7654 290414 -902
rect 293514 43174 294134 49367
rect 293514 42938 293546 43174
rect 293782 42938 293866 43174
rect 294102 42938 294134 43174
rect 293514 42854 294134 42938
rect 293514 42618 293546 42854
rect 293782 42618 293866 42854
rect 294102 42618 294134 42854
rect 293514 7174 294134 42618
rect 293514 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 294134 7174
rect 293514 6854 294134 6938
rect 293514 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 294134 6854
rect 293514 -1306 294134 6618
rect 293514 -1542 293546 -1306
rect 293782 -1542 293866 -1306
rect 294102 -1542 294134 -1306
rect 293514 -1626 294134 -1542
rect 293514 -1862 293546 -1626
rect 293782 -1862 293866 -1626
rect 294102 -1862 294134 -1626
rect 293514 -7654 294134 -1862
rect 297234 46894 297854 49367
rect 297234 46658 297266 46894
rect 297502 46658 297586 46894
rect 297822 46658 297854 46894
rect 297234 46574 297854 46658
rect 297234 46338 297266 46574
rect 297502 46338 297586 46574
rect 297822 46338 297854 46574
rect 297234 10894 297854 46338
rect 297234 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 297854 10894
rect 297234 10574 297854 10658
rect 297234 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 297854 10574
rect 297234 -2266 297854 10338
rect 297234 -2502 297266 -2266
rect 297502 -2502 297586 -2266
rect 297822 -2502 297854 -2266
rect 297234 -2586 297854 -2502
rect 297234 -2822 297266 -2586
rect 297502 -2822 297586 -2586
rect 297822 -2822 297854 -2586
rect 297234 -7654 297854 -2822
rect 300954 14614 301574 45068
rect 300954 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 301574 14614
rect 300954 14294 301574 14378
rect 300954 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 301574 14294
rect 300954 -3226 301574 14058
rect 300954 -3462 300986 -3226
rect 301222 -3462 301306 -3226
rect 301542 -3462 301574 -3226
rect 300954 -3546 301574 -3462
rect 300954 -3782 300986 -3546
rect 301222 -3782 301306 -3546
rect 301542 -3782 301574 -3546
rect 300954 -7654 301574 -3782
rect 304674 18334 305294 49367
rect 304674 18098 304706 18334
rect 304942 18098 305026 18334
rect 305262 18098 305294 18334
rect 304674 18014 305294 18098
rect 304674 17778 304706 18014
rect 304942 17778 305026 18014
rect 305262 17778 305294 18014
rect 304674 -4186 305294 17778
rect 304674 -4422 304706 -4186
rect 304942 -4422 305026 -4186
rect 305262 -4422 305294 -4186
rect 304674 -4506 305294 -4422
rect 304674 -4742 304706 -4506
rect 304942 -4742 305026 -4506
rect 305262 -4742 305294 -4506
rect 304674 -7654 305294 -4742
rect 308394 22054 309014 49367
rect 308394 21818 308426 22054
rect 308662 21818 308746 22054
rect 308982 21818 309014 22054
rect 308394 21734 309014 21818
rect 308394 21498 308426 21734
rect 308662 21498 308746 21734
rect 308982 21498 309014 21734
rect 308394 -5146 309014 21498
rect 308394 -5382 308426 -5146
rect 308662 -5382 308746 -5146
rect 308982 -5382 309014 -5146
rect 308394 -5466 309014 -5382
rect 308394 -5702 308426 -5466
rect 308662 -5702 308746 -5466
rect 308982 -5702 309014 -5466
rect 308394 -7654 309014 -5702
rect 312114 25774 312734 49367
rect 312114 25538 312146 25774
rect 312382 25538 312466 25774
rect 312702 25538 312734 25774
rect 312114 25454 312734 25538
rect 312114 25218 312146 25454
rect 312382 25218 312466 25454
rect 312702 25218 312734 25454
rect 312114 -6106 312734 25218
rect 312114 -6342 312146 -6106
rect 312382 -6342 312466 -6106
rect 312702 -6342 312734 -6106
rect 312114 -6426 312734 -6342
rect 312114 -6662 312146 -6426
rect 312382 -6662 312466 -6426
rect 312702 -6662 312734 -6426
rect 312114 -7654 312734 -6662
rect 315834 29494 316454 45068
rect 315834 29258 315866 29494
rect 316102 29258 316186 29494
rect 316422 29258 316454 29494
rect 315834 29174 316454 29258
rect 315834 28938 315866 29174
rect 316102 28938 316186 29174
rect 316422 28938 316454 29174
rect 315834 -7066 316454 28938
rect 315834 -7302 315866 -7066
rect 316102 -7302 316186 -7066
rect 316422 -7302 316454 -7066
rect 315834 -7386 316454 -7302
rect 315834 -7622 315866 -7386
rect 316102 -7622 316186 -7386
rect 316422 -7622 316454 -7386
rect 315834 -7654 316454 -7622
rect 325794 39454 326414 49367
rect 325794 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 326414 39454
rect 325794 39134 326414 39218
rect 325794 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 326414 39134
rect 325794 3454 326414 38898
rect 325794 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 326414 3454
rect 325794 3134 326414 3218
rect 325794 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 326414 3134
rect 325794 -346 326414 2898
rect 325794 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 326414 -346
rect 325794 -666 326414 -582
rect 325794 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 326414 -666
rect 325794 -7654 326414 -902
rect 329514 43174 330134 49367
rect 329514 42938 329546 43174
rect 329782 42938 329866 43174
rect 330102 42938 330134 43174
rect 329514 42854 330134 42938
rect 329514 42618 329546 42854
rect 329782 42618 329866 42854
rect 330102 42618 330134 42854
rect 329514 7174 330134 42618
rect 329514 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 330134 7174
rect 329514 6854 330134 6938
rect 329514 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 330134 6854
rect 329514 -1306 330134 6618
rect 329514 -1542 329546 -1306
rect 329782 -1542 329866 -1306
rect 330102 -1542 330134 -1306
rect 329514 -1626 330134 -1542
rect 329514 -1862 329546 -1626
rect 329782 -1862 329866 -1626
rect 330102 -1862 330134 -1626
rect 329514 -7654 330134 -1862
rect 333234 46894 333854 49367
rect 333234 46658 333266 46894
rect 333502 46658 333586 46894
rect 333822 46658 333854 46894
rect 333234 46574 333854 46658
rect 333234 46338 333266 46574
rect 333502 46338 333586 46574
rect 333822 46338 333854 46574
rect 333234 10894 333854 46338
rect 333234 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 333854 10894
rect 333234 10574 333854 10658
rect 333234 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 333854 10574
rect 333234 -2266 333854 10338
rect 333234 -2502 333266 -2266
rect 333502 -2502 333586 -2266
rect 333822 -2502 333854 -2266
rect 333234 -2586 333854 -2502
rect 333234 -2822 333266 -2586
rect 333502 -2822 333586 -2586
rect 333822 -2822 333854 -2586
rect 333234 -7654 333854 -2822
rect 336954 14614 337574 49367
rect 336954 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 337574 14614
rect 336954 14294 337574 14378
rect 336954 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 337574 14294
rect 336954 -3226 337574 14058
rect 336954 -3462 336986 -3226
rect 337222 -3462 337306 -3226
rect 337542 -3462 337574 -3226
rect 336954 -3546 337574 -3462
rect 336954 -3782 336986 -3546
rect 337222 -3782 337306 -3546
rect 337542 -3782 337574 -3546
rect 336954 -7654 337574 -3782
rect 340674 18334 341294 49367
rect 340674 18098 340706 18334
rect 340942 18098 341026 18334
rect 341262 18098 341294 18334
rect 340674 18014 341294 18098
rect 340674 17778 340706 18014
rect 340942 17778 341026 18014
rect 341262 17778 341294 18014
rect 340674 -4186 341294 17778
rect 340674 -4422 340706 -4186
rect 340942 -4422 341026 -4186
rect 341262 -4422 341294 -4186
rect 340674 -4506 341294 -4422
rect 340674 -4742 340706 -4506
rect 340942 -4742 341026 -4506
rect 341262 -4742 341294 -4506
rect 340674 -7654 341294 -4742
rect 344394 22054 345014 49367
rect 344394 21818 344426 22054
rect 344662 21818 344746 22054
rect 344982 21818 345014 22054
rect 344394 21734 345014 21818
rect 344394 21498 344426 21734
rect 344662 21498 344746 21734
rect 344982 21498 345014 21734
rect 344394 -5146 345014 21498
rect 344394 -5382 344426 -5146
rect 344662 -5382 344746 -5146
rect 344982 -5382 345014 -5146
rect 344394 -5466 345014 -5382
rect 344394 -5702 344426 -5466
rect 344662 -5702 344746 -5466
rect 344982 -5702 345014 -5466
rect 344394 -7654 345014 -5702
rect 348114 25774 348734 49367
rect 348114 25538 348146 25774
rect 348382 25538 348466 25774
rect 348702 25538 348734 25774
rect 348114 25454 348734 25538
rect 348114 25218 348146 25454
rect 348382 25218 348466 25454
rect 348702 25218 348734 25454
rect 348114 -6106 348734 25218
rect 348114 -6342 348146 -6106
rect 348382 -6342 348466 -6106
rect 348702 -6342 348734 -6106
rect 348114 -6426 348734 -6342
rect 348114 -6662 348146 -6426
rect 348382 -6662 348466 -6426
rect 348702 -6662 348734 -6426
rect 348114 -7654 348734 -6662
rect 351834 29494 352454 49367
rect 351834 29258 351866 29494
rect 352102 29258 352186 29494
rect 352422 29258 352454 29494
rect 351834 29174 352454 29258
rect 351834 28938 351866 29174
rect 352102 28938 352186 29174
rect 352422 28938 352454 29174
rect 351834 -7066 352454 28938
rect 351834 -7302 351866 -7066
rect 352102 -7302 352186 -7066
rect 352422 -7302 352454 -7066
rect 351834 -7386 352454 -7302
rect 351834 -7622 351866 -7386
rect 352102 -7622 352186 -7386
rect 352422 -7622 352454 -7386
rect 351834 -7654 352454 -7622
rect 361794 39454 362414 74898
rect 361794 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 362414 39454
rect 361794 39134 362414 39218
rect 361794 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 362414 39134
rect 361794 3454 362414 38898
rect 361794 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 362414 3454
rect 361794 3134 362414 3218
rect 361794 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 362414 3134
rect 361794 -346 362414 2898
rect 361794 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 362414 -346
rect 361794 -666 362414 -582
rect 361794 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 362414 -666
rect 361794 -7654 362414 -902
rect 365514 705798 366134 711590
rect 365514 705562 365546 705798
rect 365782 705562 365866 705798
rect 366102 705562 366134 705798
rect 365514 705478 366134 705562
rect 365514 705242 365546 705478
rect 365782 705242 365866 705478
rect 366102 705242 366134 705478
rect 365514 691174 366134 705242
rect 365514 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 366134 691174
rect 365514 690854 366134 690938
rect 365514 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 366134 690854
rect 365514 655174 366134 690618
rect 365514 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 366134 655174
rect 365514 654854 366134 654938
rect 365514 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 366134 654854
rect 365514 619174 366134 654618
rect 365514 618938 365546 619174
rect 365782 618938 365866 619174
rect 366102 618938 366134 619174
rect 365514 618854 366134 618938
rect 365514 618618 365546 618854
rect 365782 618618 365866 618854
rect 366102 618618 366134 618854
rect 365514 583174 366134 618618
rect 365514 582938 365546 583174
rect 365782 582938 365866 583174
rect 366102 582938 366134 583174
rect 365514 582854 366134 582938
rect 365514 582618 365546 582854
rect 365782 582618 365866 582854
rect 366102 582618 366134 582854
rect 365514 547174 366134 582618
rect 365514 546938 365546 547174
rect 365782 546938 365866 547174
rect 366102 546938 366134 547174
rect 365514 546854 366134 546938
rect 365514 546618 365546 546854
rect 365782 546618 365866 546854
rect 366102 546618 366134 546854
rect 365514 511174 366134 546618
rect 365514 510938 365546 511174
rect 365782 510938 365866 511174
rect 366102 510938 366134 511174
rect 365514 510854 366134 510938
rect 365514 510618 365546 510854
rect 365782 510618 365866 510854
rect 366102 510618 366134 510854
rect 365514 475174 366134 510618
rect 365514 474938 365546 475174
rect 365782 474938 365866 475174
rect 366102 474938 366134 475174
rect 365514 474854 366134 474938
rect 365514 474618 365546 474854
rect 365782 474618 365866 474854
rect 366102 474618 366134 474854
rect 365514 439174 366134 474618
rect 365514 438938 365546 439174
rect 365782 438938 365866 439174
rect 366102 438938 366134 439174
rect 365514 438854 366134 438938
rect 365514 438618 365546 438854
rect 365782 438618 365866 438854
rect 366102 438618 366134 438854
rect 365514 403174 366134 438618
rect 365514 402938 365546 403174
rect 365782 402938 365866 403174
rect 366102 402938 366134 403174
rect 365514 402854 366134 402938
rect 365514 402618 365546 402854
rect 365782 402618 365866 402854
rect 366102 402618 366134 402854
rect 365514 367174 366134 402618
rect 365514 366938 365546 367174
rect 365782 366938 365866 367174
rect 366102 366938 366134 367174
rect 365514 366854 366134 366938
rect 365514 366618 365546 366854
rect 365782 366618 365866 366854
rect 366102 366618 366134 366854
rect 365514 331174 366134 366618
rect 365514 330938 365546 331174
rect 365782 330938 365866 331174
rect 366102 330938 366134 331174
rect 365514 330854 366134 330938
rect 365514 330618 365546 330854
rect 365782 330618 365866 330854
rect 366102 330618 366134 330854
rect 365514 295174 366134 330618
rect 365514 294938 365546 295174
rect 365782 294938 365866 295174
rect 366102 294938 366134 295174
rect 365514 294854 366134 294938
rect 365514 294618 365546 294854
rect 365782 294618 365866 294854
rect 366102 294618 366134 294854
rect 365514 259174 366134 294618
rect 365514 258938 365546 259174
rect 365782 258938 365866 259174
rect 366102 258938 366134 259174
rect 365514 258854 366134 258938
rect 365514 258618 365546 258854
rect 365782 258618 365866 258854
rect 366102 258618 366134 258854
rect 365514 223174 366134 258618
rect 365514 222938 365546 223174
rect 365782 222938 365866 223174
rect 366102 222938 366134 223174
rect 365514 222854 366134 222938
rect 365514 222618 365546 222854
rect 365782 222618 365866 222854
rect 366102 222618 366134 222854
rect 365514 187174 366134 222618
rect 365514 186938 365546 187174
rect 365782 186938 365866 187174
rect 366102 186938 366134 187174
rect 365514 186854 366134 186938
rect 365514 186618 365546 186854
rect 365782 186618 365866 186854
rect 366102 186618 366134 186854
rect 365514 151174 366134 186618
rect 365514 150938 365546 151174
rect 365782 150938 365866 151174
rect 366102 150938 366134 151174
rect 365514 150854 366134 150938
rect 365514 150618 365546 150854
rect 365782 150618 365866 150854
rect 366102 150618 366134 150854
rect 365514 115174 366134 150618
rect 365514 114938 365546 115174
rect 365782 114938 365866 115174
rect 366102 114938 366134 115174
rect 365514 114854 366134 114938
rect 365514 114618 365546 114854
rect 365782 114618 365866 114854
rect 366102 114618 366134 114854
rect 365514 79174 366134 114618
rect 365514 78938 365546 79174
rect 365782 78938 365866 79174
rect 366102 78938 366134 79174
rect 365514 78854 366134 78938
rect 365514 78618 365546 78854
rect 365782 78618 365866 78854
rect 366102 78618 366134 78854
rect 365514 43174 366134 78618
rect 365514 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 366134 43174
rect 365514 42854 366134 42938
rect 365514 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 366134 42854
rect 365514 7174 366134 42618
rect 365514 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 366134 7174
rect 365514 6854 366134 6938
rect 365514 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 366134 6854
rect 365514 -1306 366134 6618
rect 365514 -1542 365546 -1306
rect 365782 -1542 365866 -1306
rect 366102 -1542 366134 -1306
rect 365514 -1626 366134 -1542
rect 365514 -1862 365546 -1626
rect 365782 -1862 365866 -1626
rect 366102 -1862 366134 -1626
rect 365514 -7654 366134 -1862
rect 369234 706758 369854 711590
rect 369234 706522 369266 706758
rect 369502 706522 369586 706758
rect 369822 706522 369854 706758
rect 369234 706438 369854 706522
rect 369234 706202 369266 706438
rect 369502 706202 369586 706438
rect 369822 706202 369854 706438
rect 369234 694894 369854 706202
rect 369234 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 369854 694894
rect 369234 694574 369854 694658
rect 369234 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 369854 694574
rect 369234 658894 369854 694338
rect 369234 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 369854 658894
rect 369234 658574 369854 658658
rect 369234 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 369854 658574
rect 369234 622894 369854 658338
rect 369234 622658 369266 622894
rect 369502 622658 369586 622894
rect 369822 622658 369854 622894
rect 369234 622574 369854 622658
rect 369234 622338 369266 622574
rect 369502 622338 369586 622574
rect 369822 622338 369854 622574
rect 369234 586894 369854 622338
rect 369234 586658 369266 586894
rect 369502 586658 369586 586894
rect 369822 586658 369854 586894
rect 369234 586574 369854 586658
rect 369234 586338 369266 586574
rect 369502 586338 369586 586574
rect 369822 586338 369854 586574
rect 369234 550894 369854 586338
rect 369234 550658 369266 550894
rect 369502 550658 369586 550894
rect 369822 550658 369854 550894
rect 369234 550574 369854 550658
rect 369234 550338 369266 550574
rect 369502 550338 369586 550574
rect 369822 550338 369854 550574
rect 369234 514894 369854 550338
rect 369234 514658 369266 514894
rect 369502 514658 369586 514894
rect 369822 514658 369854 514894
rect 369234 514574 369854 514658
rect 369234 514338 369266 514574
rect 369502 514338 369586 514574
rect 369822 514338 369854 514574
rect 369234 478894 369854 514338
rect 369234 478658 369266 478894
rect 369502 478658 369586 478894
rect 369822 478658 369854 478894
rect 369234 478574 369854 478658
rect 369234 478338 369266 478574
rect 369502 478338 369586 478574
rect 369822 478338 369854 478574
rect 369234 442894 369854 478338
rect 369234 442658 369266 442894
rect 369502 442658 369586 442894
rect 369822 442658 369854 442894
rect 369234 442574 369854 442658
rect 369234 442338 369266 442574
rect 369502 442338 369586 442574
rect 369822 442338 369854 442574
rect 369234 406894 369854 442338
rect 369234 406658 369266 406894
rect 369502 406658 369586 406894
rect 369822 406658 369854 406894
rect 369234 406574 369854 406658
rect 369234 406338 369266 406574
rect 369502 406338 369586 406574
rect 369822 406338 369854 406574
rect 369234 370894 369854 406338
rect 369234 370658 369266 370894
rect 369502 370658 369586 370894
rect 369822 370658 369854 370894
rect 369234 370574 369854 370658
rect 369234 370338 369266 370574
rect 369502 370338 369586 370574
rect 369822 370338 369854 370574
rect 369234 334894 369854 370338
rect 369234 334658 369266 334894
rect 369502 334658 369586 334894
rect 369822 334658 369854 334894
rect 369234 334574 369854 334658
rect 369234 334338 369266 334574
rect 369502 334338 369586 334574
rect 369822 334338 369854 334574
rect 369234 298894 369854 334338
rect 369234 298658 369266 298894
rect 369502 298658 369586 298894
rect 369822 298658 369854 298894
rect 369234 298574 369854 298658
rect 369234 298338 369266 298574
rect 369502 298338 369586 298574
rect 369822 298338 369854 298574
rect 369234 262894 369854 298338
rect 369234 262658 369266 262894
rect 369502 262658 369586 262894
rect 369822 262658 369854 262894
rect 369234 262574 369854 262658
rect 369234 262338 369266 262574
rect 369502 262338 369586 262574
rect 369822 262338 369854 262574
rect 369234 226894 369854 262338
rect 369234 226658 369266 226894
rect 369502 226658 369586 226894
rect 369822 226658 369854 226894
rect 369234 226574 369854 226658
rect 369234 226338 369266 226574
rect 369502 226338 369586 226574
rect 369822 226338 369854 226574
rect 369234 190894 369854 226338
rect 369234 190658 369266 190894
rect 369502 190658 369586 190894
rect 369822 190658 369854 190894
rect 369234 190574 369854 190658
rect 369234 190338 369266 190574
rect 369502 190338 369586 190574
rect 369822 190338 369854 190574
rect 369234 154894 369854 190338
rect 369234 154658 369266 154894
rect 369502 154658 369586 154894
rect 369822 154658 369854 154894
rect 369234 154574 369854 154658
rect 369234 154338 369266 154574
rect 369502 154338 369586 154574
rect 369822 154338 369854 154574
rect 369234 118894 369854 154338
rect 369234 118658 369266 118894
rect 369502 118658 369586 118894
rect 369822 118658 369854 118894
rect 369234 118574 369854 118658
rect 369234 118338 369266 118574
rect 369502 118338 369586 118574
rect 369822 118338 369854 118574
rect 369234 82894 369854 118338
rect 369234 82658 369266 82894
rect 369502 82658 369586 82894
rect 369822 82658 369854 82894
rect 369234 82574 369854 82658
rect 369234 82338 369266 82574
rect 369502 82338 369586 82574
rect 369822 82338 369854 82574
rect 369234 46894 369854 82338
rect 369234 46658 369266 46894
rect 369502 46658 369586 46894
rect 369822 46658 369854 46894
rect 369234 46574 369854 46658
rect 369234 46338 369266 46574
rect 369502 46338 369586 46574
rect 369822 46338 369854 46574
rect 369234 10894 369854 46338
rect 369234 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 369854 10894
rect 369234 10574 369854 10658
rect 369234 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 369854 10574
rect 369234 -2266 369854 10338
rect 369234 -2502 369266 -2266
rect 369502 -2502 369586 -2266
rect 369822 -2502 369854 -2266
rect 369234 -2586 369854 -2502
rect 369234 -2822 369266 -2586
rect 369502 -2822 369586 -2586
rect 369822 -2822 369854 -2586
rect 369234 -7654 369854 -2822
rect 372954 707718 373574 711590
rect 372954 707482 372986 707718
rect 373222 707482 373306 707718
rect 373542 707482 373574 707718
rect 372954 707398 373574 707482
rect 372954 707162 372986 707398
rect 373222 707162 373306 707398
rect 373542 707162 373574 707398
rect 372954 698614 373574 707162
rect 372954 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 373574 698614
rect 372954 698294 373574 698378
rect 372954 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 373574 698294
rect 372954 662614 373574 698058
rect 372954 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 373574 662614
rect 372954 662294 373574 662378
rect 372954 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 373574 662294
rect 372954 626614 373574 662058
rect 372954 626378 372986 626614
rect 373222 626378 373306 626614
rect 373542 626378 373574 626614
rect 372954 626294 373574 626378
rect 372954 626058 372986 626294
rect 373222 626058 373306 626294
rect 373542 626058 373574 626294
rect 372954 590614 373574 626058
rect 372954 590378 372986 590614
rect 373222 590378 373306 590614
rect 373542 590378 373574 590614
rect 372954 590294 373574 590378
rect 372954 590058 372986 590294
rect 373222 590058 373306 590294
rect 373542 590058 373574 590294
rect 372954 554614 373574 590058
rect 372954 554378 372986 554614
rect 373222 554378 373306 554614
rect 373542 554378 373574 554614
rect 372954 554294 373574 554378
rect 372954 554058 372986 554294
rect 373222 554058 373306 554294
rect 373542 554058 373574 554294
rect 372954 518614 373574 554058
rect 372954 518378 372986 518614
rect 373222 518378 373306 518614
rect 373542 518378 373574 518614
rect 372954 518294 373574 518378
rect 372954 518058 372986 518294
rect 373222 518058 373306 518294
rect 373542 518058 373574 518294
rect 372954 482614 373574 518058
rect 372954 482378 372986 482614
rect 373222 482378 373306 482614
rect 373542 482378 373574 482614
rect 372954 482294 373574 482378
rect 372954 482058 372986 482294
rect 373222 482058 373306 482294
rect 373542 482058 373574 482294
rect 372954 446614 373574 482058
rect 372954 446378 372986 446614
rect 373222 446378 373306 446614
rect 373542 446378 373574 446614
rect 372954 446294 373574 446378
rect 372954 446058 372986 446294
rect 373222 446058 373306 446294
rect 373542 446058 373574 446294
rect 372954 410614 373574 446058
rect 372954 410378 372986 410614
rect 373222 410378 373306 410614
rect 373542 410378 373574 410614
rect 372954 410294 373574 410378
rect 372954 410058 372986 410294
rect 373222 410058 373306 410294
rect 373542 410058 373574 410294
rect 372954 374614 373574 410058
rect 372954 374378 372986 374614
rect 373222 374378 373306 374614
rect 373542 374378 373574 374614
rect 372954 374294 373574 374378
rect 372954 374058 372986 374294
rect 373222 374058 373306 374294
rect 373542 374058 373574 374294
rect 372954 338614 373574 374058
rect 372954 338378 372986 338614
rect 373222 338378 373306 338614
rect 373542 338378 373574 338614
rect 372954 338294 373574 338378
rect 372954 338058 372986 338294
rect 373222 338058 373306 338294
rect 373542 338058 373574 338294
rect 372954 302614 373574 338058
rect 372954 302378 372986 302614
rect 373222 302378 373306 302614
rect 373542 302378 373574 302614
rect 372954 302294 373574 302378
rect 372954 302058 372986 302294
rect 373222 302058 373306 302294
rect 373542 302058 373574 302294
rect 372954 266614 373574 302058
rect 372954 266378 372986 266614
rect 373222 266378 373306 266614
rect 373542 266378 373574 266614
rect 372954 266294 373574 266378
rect 372954 266058 372986 266294
rect 373222 266058 373306 266294
rect 373542 266058 373574 266294
rect 372954 230614 373574 266058
rect 372954 230378 372986 230614
rect 373222 230378 373306 230614
rect 373542 230378 373574 230614
rect 372954 230294 373574 230378
rect 372954 230058 372986 230294
rect 373222 230058 373306 230294
rect 373542 230058 373574 230294
rect 372954 194614 373574 230058
rect 372954 194378 372986 194614
rect 373222 194378 373306 194614
rect 373542 194378 373574 194614
rect 372954 194294 373574 194378
rect 372954 194058 372986 194294
rect 373222 194058 373306 194294
rect 373542 194058 373574 194294
rect 372954 158614 373574 194058
rect 372954 158378 372986 158614
rect 373222 158378 373306 158614
rect 373542 158378 373574 158614
rect 372954 158294 373574 158378
rect 372954 158058 372986 158294
rect 373222 158058 373306 158294
rect 373542 158058 373574 158294
rect 372954 122614 373574 158058
rect 372954 122378 372986 122614
rect 373222 122378 373306 122614
rect 373542 122378 373574 122614
rect 372954 122294 373574 122378
rect 372954 122058 372986 122294
rect 373222 122058 373306 122294
rect 373542 122058 373574 122294
rect 372954 86614 373574 122058
rect 372954 86378 372986 86614
rect 373222 86378 373306 86614
rect 373542 86378 373574 86614
rect 372954 86294 373574 86378
rect 372954 86058 372986 86294
rect 373222 86058 373306 86294
rect 373542 86058 373574 86294
rect 372954 50614 373574 86058
rect 372954 50378 372986 50614
rect 373222 50378 373306 50614
rect 373542 50378 373574 50614
rect 372954 50294 373574 50378
rect 372954 50058 372986 50294
rect 373222 50058 373306 50294
rect 373542 50058 373574 50294
rect 372954 14614 373574 50058
rect 372954 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 373574 14614
rect 372954 14294 373574 14378
rect 372954 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 373574 14294
rect 372954 -3226 373574 14058
rect 372954 -3462 372986 -3226
rect 373222 -3462 373306 -3226
rect 373542 -3462 373574 -3226
rect 372954 -3546 373574 -3462
rect 372954 -3782 372986 -3546
rect 373222 -3782 373306 -3546
rect 373542 -3782 373574 -3546
rect 372954 -7654 373574 -3782
rect 376674 708678 377294 711590
rect 376674 708442 376706 708678
rect 376942 708442 377026 708678
rect 377262 708442 377294 708678
rect 376674 708358 377294 708442
rect 376674 708122 376706 708358
rect 376942 708122 377026 708358
rect 377262 708122 377294 708358
rect 376674 666334 377294 708122
rect 376674 666098 376706 666334
rect 376942 666098 377026 666334
rect 377262 666098 377294 666334
rect 376674 666014 377294 666098
rect 376674 665778 376706 666014
rect 376942 665778 377026 666014
rect 377262 665778 377294 666014
rect 376674 630334 377294 665778
rect 376674 630098 376706 630334
rect 376942 630098 377026 630334
rect 377262 630098 377294 630334
rect 376674 630014 377294 630098
rect 376674 629778 376706 630014
rect 376942 629778 377026 630014
rect 377262 629778 377294 630014
rect 376674 594334 377294 629778
rect 376674 594098 376706 594334
rect 376942 594098 377026 594334
rect 377262 594098 377294 594334
rect 376674 594014 377294 594098
rect 376674 593778 376706 594014
rect 376942 593778 377026 594014
rect 377262 593778 377294 594014
rect 376674 558334 377294 593778
rect 376674 558098 376706 558334
rect 376942 558098 377026 558334
rect 377262 558098 377294 558334
rect 376674 558014 377294 558098
rect 376674 557778 376706 558014
rect 376942 557778 377026 558014
rect 377262 557778 377294 558014
rect 376674 522334 377294 557778
rect 376674 522098 376706 522334
rect 376942 522098 377026 522334
rect 377262 522098 377294 522334
rect 376674 522014 377294 522098
rect 376674 521778 376706 522014
rect 376942 521778 377026 522014
rect 377262 521778 377294 522014
rect 376674 486334 377294 521778
rect 376674 486098 376706 486334
rect 376942 486098 377026 486334
rect 377262 486098 377294 486334
rect 376674 486014 377294 486098
rect 376674 485778 376706 486014
rect 376942 485778 377026 486014
rect 377262 485778 377294 486014
rect 376674 450334 377294 485778
rect 376674 450098 376706 450334
rect 376942 450098 377026 450334
rect 377262 450098 377294 450334
rect 376674 450014 377294 450098
rect 376674 449778 376706 450014
rect 376942 449778 377026 450014
rect 377262 449778 377294 450014
rect 376674 414334 377294 449778
rect 376674 414098 376706 414334
rect 376942 414098 377026 414334
rect 377262 414098 377294 414334
rect 376674 414014 377294 414098
rect 376674 413778 376706 414014
rect 376942 413778 377026 414014
rect 377262 413778 377294 414014
rect 376674 378334 377294 413778
rect 376674 378098 376706 378334
rect 376942 378098 377026 378334
rect 377262 378098 377294 378334
rect 376674 378014 377294 378098
rect 376674 377778 376706 378014
rect 376942 377778 377026 378014
rect 377262 377778 377294 378014
rect 376674 342334 377294 377778
rect 376674 342098 376706 342334
rect 376942 342098 377026 342334
rect 377262 342098 377294 342334
rect 376674 342014 377294 342098
rect 376674 341778 376706 342014
rect 376942 341778 377026 342014
rect 377262 341778 377294 342014
rect 376674 306334 377294 341778
rect 376674 306098 376706 306334
rect 376942 306098 377026 306334
rect 377262 306098 377294 306334
rect 376674 306014 377294 306098
rect 376674 305778 376706 306014
rect 376942 305778 377026 306014
rect 377262 305778 377294 306014
rect 376674 270334 377294 305778
rect 376674 270098 376706 270334
rect 376942 270098 377026 270334
rect 377262 270098 377294 270334
rect 376674 270014 377294 270098
rect 376674 269778 376706 270014
rect 376942 269778 377026 270014
rect 377262 269778 377294 270014
rect 376674 234334 377294 269778
rect 376674 234098 376706 234334
rect 376942 234098 377026 234334
rect 377262 234098 377294 234334
rect 376674 234014 377294 234098
rect 376674 233778 376706 234014
rect 376942 233778 377026 234014
rect 377262 233778 377294 234014
rect 376674 198334 377294 233778
rect 376674 198098 376706 198334
rect 376942 198098 377026 198334
rect 377262 198098 377294 198334
rect 376674 198014 377294 198098
rect 376674 197778 376706 198014
rect 376942 197778 377026 198014
rect 377262 197778 377294 198014
rect 376674 162334 377294 197778
rect 376674 162098 376706 162334
rect 376942 162098 377026 162334
rect 377262 162098 377294 162334
rect 376674 162014 377294 162098
rect 376674 161778 376706 162014
rect 376942 161778 377026 162014
rect 377262 161778 377294 162014
rect 376674 126334 377294 161778
rect 376674 126098 376706 126334
rect 376942 126098 377026 126334
rect 377262 126098 377294 126334
rect 376674 126014 377294 126098
rect 376674 125778 376706 126014
rect 376942 125778 377026 126014
rect 377262 125778 377294 126014
rect 376674 90334 377294 125778
rect 376674 90098 376706 90334
rect 376942 90098 377026 90334
rect 377262 90098 377294 90334
rect 376674 90014 377294 90098
rect 376674 89778 376706 90014
rect 376942 89778 377026 90014
rect 377262 89778 377294 90014
rect 376674 54334 377294 89778
rect 376674 54098 376706 54334
rect 376942 54098 377026 54334
rect 377262 54098 377294 54334
rect 376674 54014 377294 54098
rect 376674 53778 376706 54014
rect 376942 53778 377026 54014
rect 377262 53778 377294 54014
rect 376674 18334 377294 53778
rect 376674 18098 376706 18334
rect 376942 18098 377026 18334
rect 377262 18098 377294 18334
rect 376674 18014 377294 18098
rect 376674 17778 376706 18014
rect 376942 17778 377026 18014
rect 377262 17778 377294 18014
rect 376674 -4186 377294 17778
rect 376674 -4422 376706 -4186
rect 376942 -4422 377026 -4186
rect 377262 -4422 377294 -4186
rect 376674 -4506 377294 -4422
rect 376674 -4742 376706 -4506
rect 376942 -4742 377026 -4506
rect 377262 -4742 377294 -4506
rect 376674 -7654 377294 -4742
rect 380394 709638 381014 711590
rect 380394 709402 380426 709638
rect 380662 709402 380746 709638
rect 380982 709402 381014 709638
rect 380394 709318 381014 709402
rect 380394 709082 380426 709318
rect 380662 709082 380746 709318
rect 380982 709082 381014 709318
rect 380394 670054 381014 709082
rect 380394 669818 380426 670054
rect 380662 669818 380746 670054
rect 380982 669818 381014 670054
rect 380394 669734 381014 669818
rect 380394 669498 380426 669734
rect 380662 669498 380746 669734
rect 380982 669498 381014 669734
rect 380394 634054 381014 669498
rect 380394 633818 380426 634054
rect 380662 633818 380746 634054
rect 380982 633818 381014 634054
rect 380394 633734 381014 633818
rect 380394 633498 380426 633734
rect 380662 633498 380746 633734
rect 380982 633498 381014 633734
rect 380394 598054 381014 633498
rect 380394 597818 380426 598054
rect 380662 597818 380746 598054
rect 380982 597818 381014 598054
rect 380394 597734 381014 597818
rect 380394 597498 380426 597734
rect 380662 597498 380746 597734
rect 380982 597498 381014 597734
rect 380394 562054 381014 597498
rect 380394 561818 380426 562054
rect 380662 561818 380746 562054
rect 380982 561818 381014 562054
rect 380394 561734 381014 561818
rect 380394 561498 380426 561734
rect 380662 561498 380746 561734
rect 380982 561498 381014 561734
rect 380394 526054 381014 561498
rect 380394 525818 380426 526054
rect 380662 525818 380746 526054
rect 380982 525818 381014 526054
rect 380394 525734 381014 525818
rect 380394 525498 380426 525734
rect 380662 525498 380746 525734
rect 380982 525498 381014 525734
rect 380394 490054 381014 525498
rect 380394 489818 380426 490054
rect 380662 489818 380746 490054
rect 380982 489818 381014 490054
rect 380394 489734 381014 489818
rect 380394 489498 380426 489734
rect 380662 489498 380746 489734
rect 380982 489498 381014 489734
rect 380394 454054 381014 489498
rect 380394 453818 380426 454054
rect 380662 453818 380746 454054
rect 380982 453818 381014 454054
rect 380394 453734 381014 453818
rect 380394 453498 380426 453734
rect 380662 453498 380746 453734
rect 380982 453498 381014 453734
rect 380394 418054 381014 453498
rect 380394 417818 380426 418054
rect 380662 417818 380746 418054
rect 380982 417818 381014 418054
rect 380394 417734 381014 417818
rect 380394 417498 380426 417734
rect 380662 417498 380746 417734
rect 380982 417498 381014 417734
rect 380394 382054 381014 417498
rect 380394 381818 380426 382054
rect 380662 381818 380746 382054
rect 380982 381818 381014 382054
rect 380394 381734 381014 381818
rect 380394 381498 380426 381734
rect 380662 381498 380746 381734
rect 380982 381498 381014 381734
rect 380394 346054 381014 381498
rect 380394 345818 380426 346054
rect 380662 345818 380746 346054
rect 380982 345818 381014 346054
rect 380394 345734 381014 345818
rect 380394 345498 380426 345734
rect 380662 345498 380746 345734
rect 380982 345498 381014 345734
rect 380394 310054 381014 345498
rect 380394 309818 380426 310054
rect 380662 309818 380746 310054
rect 380982 309818 381014 310054
rect 380394 309734 381014 309818
rect 380394 309498 380426 309734
rect 380662 309498 380746 309734
rect 380982 309498 381014 309734
rect 380394 274054 381014 309498
rect 380394 273818 380426 274054
rect 380662 273818 380746 274054
rect 380982 273818 381014 274054
rect 380394 273734 381014 273818
rect 380394 273498 380426 273734
rect 380662 273498 380746 273734
rect 380982 273498 381014 273734
rect 380394 238054 381014 273498
rect 380394 237818 380426 238054
rect 380662 237818 380746 238054
rect 380982 237818 381014 238054
rect 380394 237734 381014 237818
rect 380394 237498 380426 237734
rect 380662 237498 380746 237734
rect 380982 237498 381014 237734
rect 380394 202054 381014 237498
rect 380394 201818 380426 202054
rect 380662 201818 380746 202054
rect 380982 201818 381014 202054
rect 380394 201734 381014 201818
rect 380394 201498 380426 201734
rect 380662 201498 380746 201734
rect 380982 201498 381014 201734
rect 380394 166054 381014 201498
rect 380394 165818 380426 166054
rect 380662 165818 380746 166054
rect 380982 165818 381014 166054
rect 380394 165734 381014 165818
rect 380394 165498 380426 165734
rect 380662 165498 380746 165734
rect 380982 165498 381014 165734
rect 380394 130054 381014 165498
rect 380394 129818 380426 130054
rect 380662 129818 380746 130054
rect 380982 129818 381014 130054
rect 380394 129734 381014 129818
rect 380394 129498 380426 129734
rect 380662 129498 380746 129734
rect 380982 129498 381014 129734
rect 380394 94054 381014 129498
rect 380394 93818 380426 94054
rect 380662 93818 380746 94054
rect 380982 93818 381014 94054
rect 380394 93734 381014 93818
rect 380394 93498 380426 93734
rect 380662 93498 380746 93734
rect 380982 93498 381014 93734
rect 380394 58054 381014 93498
rect 380394 57818 380426 58054
rect 380662 57818 380746 58054
rect 380982 57818 381014 58054
rect 380394 57734 381014 57818
rect 380394 57498 380426 57734
rect 380662 57498 380746 57734
rect 380982 57498 381014 57734
rect 380394 22054 381014 57498
rect 380394 21818 380426 22054
rect 380662 21818 380746 22054
rect 380982 21818 381014 22054
rect 380394 21734 381014 21818
rect 380394 21498 380426 21734
rect 380662 21498 380746 21734
rect 380982 21498 381014 21734
rect 380394 -5146 381014 21498
rect 380394 -5382 380426 -5146
rect 380662 -5382 380746 -5146
rect 380982 -5382 381014 -5146
rect 380394 -5466 381014 -5382
rect 380394 -5702 380426 -5466
rect 380662 -5702 380746 -5466
rect 380982 -5702 381014 -5466
rect 380394 -7654 381014 -5702
rect 384114 710598 384734 711590
rect 384114 710362 384146 710598
rect 384382 710362 384466 710598
rect 384702 710362 384734 710598
rect 384114 710278 384734 710362
rect 384114 710042 384146 710278
rect 384382 710042 384466 710278
rect 384702 710042 384734 710278
rect 384114 673774 384734 710042
rect 384114 673538 384146 673774
rect 384382 673538 384466 673774
rect 384702 673538 384734 673774
rect 384114 673454 384734 673538
rect 384114 673218 384146 673454
rect 384382 673218 384466 673454
rect 384702 673218 384734 673454
rect 384114 637774 384734 673218
rect 384114 637538 384146 637774
rect 384382 637538 384466 637774
rect 384702 637538 384734 637774
rect 384114 637454 384734 637538
rect 384114 637218 384146 637454
rect 384382 637218 384466 637454
rect 384702 637218 384734 637454
rect 384114 601774 384734 637218
rect 384114 601538 384146 601774
rect 384382 601538 384466 601774
rect 384702 601538 384734 601774
rect 384114 601454 384734 601538
rect 384114 601218 384146 601454
rect 384382 601218 384466 601454
rect 384702 601218 384734 601454
rect 384114 565774 384734 601218
rect 384114 565538 384146 565774
rect 384382 565538 384466 565774
rect 384702 565538 384734 565774
rect 384114 565454 384734 565538
rect 384114 565218 384146 565454
rect 384382 565218 384466 565454
rect 384702 565218 384734 565454
rect 384114 529774 384734 565218
rect 384114 529538 384146 529774
rect 384382 529538 384466 529774
rect 384702 529538 384734 529774
rect 384114 529454 384734 529538
rect 384114 529218 384146 529454
rect 384382 529218 384466 529454
rect 384702 529218 384734 529454
rect 384114 493774 384734 529218
rect 384114 493538 384146 493774
rect 384382 493538 384466 493774
rect 384702 493538 384734 493774
rect 384114 493454 384734 493538
rect 384114 493218 384146 493454
rect 384382 493218 384466 493454
rect 384702 493218 384734 493454
rect 384114 457774 384734 493218
rect 384114 457538 384146 457774
rect 384382 457538 384466 457774
rect 384702 457538 384734 457774
rect 384114 457454 384734 457538
rect 384114 457218 384146 457454
rect 384382 457218 384466 457454
rect 384702 457218 384734 457454
rect 384114 421774 384734 457218
rect 384114 421538 384146 421774
rect 384382 421538 384466 421774
rect 384702 421538 384734 421774
rect 384114 421454 384734 421538
rect 384114 421218 384146 421454
rect 384382 421218 384466 421454
rect 384702 421218 384734 421454
rect 384114 385774 384734 421218
rect 384114 385538 384146 385774
rect 384382 385538 384466 385774
rect 384702 385538 384734 385774
rect 384114 385454 384734 385538
rect 384114 385218 384146 385454
rect 384382 385218 384466 385454
rect 384702 385218 384734 385454
rect 384114 349774 384734 385218
rect 384114 349538 384146 349774
rect 384382 349538 384466 349774
rect 384702 349538 384734 349774
rect 384114 349454 384734 349538
rect 384114 349218 384146 349454
rect 384382 349218 384466 349454
rect 384702 349218 384734 349454
rect 384114 313774 384734 349218
rect 384114 313538 384146 313774
rect 384382 313538 384466 313774
rect 384702 313538 384734 313774
rect 384114 313454 384734 313538
rect 384114 313218 384146 313454
rect 384382 313218 384466 313454
rect 384702 313218 384734 313454
rect 384114 277774 384734 313218
rect 384114 277538 384146 277774
rect 384382 277538 384466 277774
rect 384702 277538 384734 277774
rect 384114 277454 384734 277538
rect 384114 277218 384146 277454
rect 384382 277218 384466 277454
rect 384702 277218 384734 277454
rect 384114 241774 384734 277218
rect 384114 241538 384146 241774
rect 384382 241538 384466 241774
rect 384702 241538 384734 241774
rect 384114 241454 384734 241538
rect 384114 241218 384146 241454
rect 384382 241218 384466 241454
rect 384702 241218 384734 241454
rect 384114 205774 384734 241218
rect 384114 205538 384146 205774
rect 384382 205538 384466 205774
rect 384702 205538 384734 205774
rect 384114 205454 384734 205538
rect 384114 205218 384146 205454
rect 384382 205218 384466 205454
rect 384702 205218 384734 205454
rect 384114 169774 384734 205218
rect 384114 169538 384146 169774
rect 384382 169538 384466 169774
rect 384702 169538 384734 169774
rect 384114 169454 384734 169538
rect 384114 169218 384146 169454
rect 384382 169218 384466 169454
rect 384702 169218 384734 169454
rect 384114 133774 384734 169218
rect 384114 133538 384146 133774
rect 384382 133538 384466 133774
rect 384702 133538 384734 133774
rect 384114 133454 384734 133538
rect 384114 133218 384146 133454
rect 384382 133218 384466 133454
rect 384702 133218 384734 133454
rect 384114 97774 384734 133218
rect 384114 97538 384146 97774
rect 384382 97538 384466 97774
rect 384702 97538 384734 97774
rect 384114 97454 384734 97538
rect 384114 97218 384146 97454
rect 384382 97218 384466 97454
rect 384702 97218 384734 97454
rect 384114 61774 384734 97218
rect 387834 711558 388454 711590
rect 387834 711322 387866 711558
rect 388102 711322 388186 711558
rect 388422 711322 388454 711558
rect 387834 711238 388454 711322
rect 387834 711002 387866 711238
rect 388102 711002 388186 711238
rect 388422 711002 388454 711238
rect 387834 677494 388454 711002
rect 387834 677258 387866 677494
rect 388102 677258 388186 677494
rect 388422 677258 388454 677494
rect 387834 677174 388454 677258
rect 387834 676938 387866 677174
rect 388102 676938 388186 677174
rect 388422 676938 388454 677174
rect 387834 641494 388454 676938
rect 387834 641258 387866 641494
rect 388102 641258 388186 641494
rect 388422 641258 388454 641494
rect 387834 641174 388454 641258
rect 387834 640938 387866 641174
rect 388102 640938 388186 641174
rect 388422 640938 388454 641174
rect 387834 605494 388454 640938
rect 387834 605258 387866 605494
rect 388102 605258 388186 605494
rect 388422 605258 388454 605494
rect 387834 605174 388454 605258
rect 387834 604938 387866 605174
rect 388102 604938 388186 605174
rect 388422 604938 388454 605174
rect 387834 569494 388454 604938
rect 387834 569258 387866 569494
rect 388102 569258 388186 569494
rect 388422 569258 388454 569494
rect 387834 569174 388454 569258
rect 387834 568938 387866 569174
rect 388102 568938 388186 569174
rect 388422 568938 388454 569174
rect 387834 533494 388454 568938
rect 387834 533258 387866 533494
rect 388102 533258 388186 533494
rect 388422 533258 388454 533494
rect 387834 533174 388454 533258
rect 387834 532938 387866 533174
rect 388102 532938 388186 533174
rect 388422 532938 388454 533174
rect 387834 497494 388454 532938
rect 387834 497258 387866 497494
rect 388102 497258 388186 497494
rect 388422 497258 388454 497494
rect 387834 497174 388454 497258
rect 387834 496938 387866 497174
rect 388102 496938 388186 497174
rect 388422 496938 388454 497174
rect 387834 461494 388454 496938
rect 387834 461258 387866 461494
rect 388102 461258 388186 461494
rect 388422 461258 388454 461494
rect 387834 461174 388454 461258
rect 387834 460938 387866 461174
rect 388102 460938 388186 461174
rect 388422 460938 388454 461174
rect 387834 425494 388454 460938
rect 387834 425258 387866 425494
rect 388102 425258 388186 425494
rect 388422 425258 388454 425494
rect 387834 425174 388454 425258
rect 387834 424938 387866 425174
rect 388102 424938 388186 425174
rect 388422 424938 388454 425174
rect 387834 389494 388454 424938
rect 387834 389258 387866 389494
rect 388102 389258 388186 389494
rect 388422 389258 388454 389494
rect 387834 389174 388454 389258
rect 387834 388938 387866 389174
rect 388102 388938 388186 389174
rect 388422 388938 388454 389174
rect 387834 353494 388454 388938
rect 387834 353258 387866 353494
rect 388102 353258 388186 353494
rect 388422 353258 388454 353494
rect 387834 353174 388454 353258
rect 387834 352938 387866 353174
rect 388102 352938 388186 353174
rect 388422 352938 388454 353174
rect 387834 317494 388454 352938
rect 387834 317258 387866 317494
rect 388102 317258 388186 317494
rect 388422 317258 388454 317494
rect 387834 317174 388454 317258
rect 387834 316938 387866 317174
rect 388102 316938 388186 317174
rect 388422 316938 388454 317174
rect 387834 281494 388454 316938
rect 387834 281258 387866 281494
rect 388102 281258 388186 281494
rect 388422 281258 388454 281494
rect 387834 281174 388454 281258
rect 387834 280938 387866 281174
rect 388102 280938 388186 281174
rect 388422 280938 388454 281174
rect 387834 245494 388454 280938
rect 387834 245258 387866 245494
rect 388102 245258 388186 245494
rect 388422 245258 388454 245494
rect 387834 245174 388454 245258
rect 387834 244938 387866 245174
rect 388102 244938 388186 245174
rect 388422 244938 388454 245174
rect 387834 209494 388454 244938
rect 387834 209258 387866 209494
rect 388102 209258 388186 209494
rect 388422 209258 388454 209494
rect 387834 209174 388454 209258
rect 387834 208938 387866 209174
rect 388102 208938 388186 209174
rect 388422 208938 388454 209174
rect 387834 173494 388454 208938
rect 387834 173258 387866 173494
rect 388102 173258 388186 173494
rect 388422 173258 388454 173494
rect 387834 173174 388454 173258
rect 387834 172938 387866 173174
rect 388102 172938 388186 173174
rect 388422 172938 388454 173174
rect 387834 137494 388454 172938
rect 387834 137258 387866 137494
rect 388102 137258 388186 137494
rect 388422 137258 388454 137494
rect 387834 137174 388454 137258
rect 387834 136938 387866 137174
rect 388102 136938 388186 137174
rect 388422 136938 388454 137174
rect 387834 101494 388454 136938
rect 387834 101258 387866 101494
rect 388102 101258 388186 101494
rect 388422 101258 388454 101494
rect 387834 101174 388454 101258
rect 387834 100938 387866 101174
rect 388102 100938 388186 101174
rect 388422 100938 388454 101174
rect 387834 92137 388454 100938
rect 397794 704838 398414 711590
rect 397794 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 398414 704838
rect 397794 704518 398414 704602
rect 397794 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 398414 704518
rect 397794 687454 398414 704282
rect 397794 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 398414 687454
rect 397794 687134 398414 687218
rect 397794 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 398414 687134
rect 397794 651454 398414 686898
rect 397794 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 398414 651454
rect 397794 651134 398414 651218
rect 397794 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 398414 651134
rect 397794 615454 398414 650898
rect 397794 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 398414 615454
rect 397794 615134 398414 615218
rect 397794 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 398414 615134
rect 397794 579454 398414 614898
rect 397794 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 398414 579454
rect 397794 579134 398414 579218
rect 397794 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 398414 579134
rect 397794 543454 398414 578898
rect 397794 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 398414 543454
rect 397794 543134 398414 543218
rect 397794 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 398414 543134
rect 397794 507454 398414 542898
rect 397794 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 398414 507454
rect 397794 507134 398414 507218
rect 397794 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 398414 507134
rect 397794 471454 398414 506898
rect 397794 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 398414 471454
rect 397794 471134 398414 471218
rect 397794 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 398414 471134
rect 397794 435454 398414 470898
rect 397794 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 398414 435454
rect 397794 435134 398414 435218
rect 397794 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 398414 435134
rect 397794 399454 398414 434898
rect 397794 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 398414 399454
rect 397794 399134 398414 399218
rect 397794 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 398414 399134
rect 397794 363454 398414 398898
rect 397794 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 398414 363454
rect 397794 363134 398414 363218
rect 397794 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 398414 363134
rect 397794 327454 398414 362898
rect 397794 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 398414 327454
rect 397794 327134 398414 327218
rect 397794 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 398414 327134
rect 397794 291454 398414 326898
rect 397794 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 398414 291454
rect 397794 291134 398414 291218
rect 397794 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 398414 291134
rect 397794 255454 398414 290898
rect 397794 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 398414 255454
rect 397794 255134 398414 255218
rect 397794 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 398414 255134
rect 397794 219454 398414 254898
rect 397794 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 398414 219454
rect 397794 219134 398414 219218
rect 397794 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 398414 219134
rect 397794 183454 398414 218898
rect 397794 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 398414 183454
rect 397794 183134 398414 183218
rect 397794 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 398414 183134
rect 397794 147454 398414 182898
rect 397794 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 398414 147454
rect 397794 147134 398414 147218
rect 397794 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 398414 147134
rect 397794 111454 398414 146898
rect 397794 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 398414 111454
rect 397794 111134 398414 111218
rect 397794 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 398414 111134
rect 397794 92137 398414 110898
rect 401514 705798 402134 711590
rect 401514 705562 401546 705798
rect 401782 705562 401866 705798
rect 402102 705562 402134 705798
rect 401514 705478 402134 705562
rect 401514 705242 401546 705478
rect 401782 705242 401866 705478
rect 402102 705242 402134 705478
rect 401514 691174 402134 705242
rect 401514 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 402134 691174
rect 401514 690854 402134 690938
rect 401514 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 402134 690854
rect 401514 655174 402134 690618
rect 401514 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 402134 655174
rect 401514 654854 402134 654938
rect 401514 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 402134 654854
rect 401514 619174 402134 654618
rect 401514 618938 401546 619174
rect 401782 618938 401866 619174
rect 402102 618938 402134 619174
rect 401514 618854 402134 618938
rect 401514 618618 401546 618854
rect 401782 618618 401866 618854
rect 402102 618618 402134 618854
rect 401514 583174 402134 618618
rect 401514 582938 401546 583174
rect 401782 582938 401866 583174
rect 402102 582938 402134 583174
rect 401514 582854 402134 582938
rect 401514 582618 401546 582854
rect 401782 582618 401866 582854
rect 402102 582618 402134 582854
rect 401514 547174 402134 582618
rect 401514 546938 401546 547174
rect 401782 546938 401866 547174
rect 402102 546938 402134 547174
rect 401514 546854 402134 546938
rect 401514 546618 401546 546854
rect 401782 546618 401866 546854
rect 402102 546618 402134 546854
rect 401514 511174 402134 546618
rect 401514 510938 401546 511174
rect 401782 510938 401866 511174
rect 402102 510938 402134 511174
rect 401514 510854 402134 510938
rect 401514 510618 401546 510854
rect 401782 510618 401866 510854
rect 402102 510618 402134 510854
rect 401514 475174 402134 510618
rect 401514 474938 401546 475174
rect 401782 474938 401866 475174
rect 402102 474938 402134 475174
rect 401514 474854 402134 474938
rect 401514 474618 401546 474854
rect 401782 474618 401866 474854
rect 402102 474618 402134 474854
rect 401514 439174 402134 474618
rect 401514 438938 401546 439174
rect 401782 438938 401866 439174
rect 402102 438938 402134 439174
rect 401514 438854 402134 438938
rect 401514 438618 401546 438854
rect 401782 438618 401866 438854
rect 402102 438618 402134 438854
rect 401514 403174 402134 438618
rect 401514 402938 401546 403174
rect 401782 402938 401866 403174
rect 402102 402938 402134 403174
rect 401514 402854 402134 402938
rect 401514 402618 401546 402854
rect 401782 402618 401866 402854
rect 402102 402618 402134 402854
rect 401514 367174 402134 402618
rect 401514 366938 401546 367174
rect 401782 366938 401866 367174
rect 402102 366938 402134 367174
rect 401514 366854 402134 366938
rect 401514 366618 401546 366854
rect 401782 366618 401866 366854
rect 402102 366618 402134 366854
rect 401514 331174 402134 366618
rect 401514 330938 401546 331174
rect 401782 330938 401866 331174
rect 402102 330938 402134 331174
rect 401514 330854 402134 330938
rect 401514 330618 401546 330854
rect 401782 330618 401866 330854
rect 402102 330618 402134 330854
rect 401514 295174 402134 330618
rect 405234 706758 405854 711590
rect 405234 706522 405266 706758
rect 405502 706522 405586 706758
rect 405822 706522 405854 706758
rect 405234 706438 405854 706522
rect 405234 706202 405266 706438
rect 405502 706202 405586 706438
rect 405822 706202 405854 706438
rect 405234 694894 405854 706202
rect 405234 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 405854 694894
rect 405234 694574 405854 694658
rect 405234 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 405854 694574
rect 405234 658894 405854 694338
rect 405234 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 405854 658894
rect 405234 658574 405854 658658
rect 405234 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 405854 658574
rect 405234 622894 405854 658338
rect 405234 622658 405266 622894
rect 405502 622658 405586 622894
rect 405822 622658 405854 622894
rect 405234 622574 405854 622658
rect 405234 622338 405266 622574
rect 405502 622338 405586 622574
rect 405822 622338 405854 622574
rect 405234 586894 405854 622338
rect 405234 586658 405266 586894
rect 405502 586658 405586 586894
rect 405822 586658 405854 586894
rect 405234 586574 405854 586658
rect 405234 586338 405266 586574
rect 405502 586338 405586 586574
rect 405822 586338 405854 586574
rect 405234 550894 405854 586338
rect 405234 550658 405266 550894
rect 405502 550658 405586 550894
rect 405822 550658 405854 550894
rect 405234 550574 405854 550658
rect 405234 550338 405266 550574
rect 405502 550338 405586 550574
rect 405822 550338 405854 550574
rect 405234 514894 405854 550338
rect 405234 514658 405266 514894
rect 405502 514658 405586 514894
rect 405822 514658 405854 514894
rect 405234 514574 405854 514658
rect 405234 514338 405266 514574
rect 405502 514338 405586 514574
rect 405822 514338 405854 514574
rect 405234 478894 405854 514338
rect 405234 478658 405266 478894
rect 405502 478658 405586 478894
rect 405822 478658 405854 478894
rect 405234 478574 405854 478658
rect 405234 478338 405266 478574
rect 405502 478338 405586 478574
rect 405822 478338 405854 478574
rect 405234 442894 405854 478338
rect 405234 442658 405266 442894
rect 405502 442658 405586 442894
rect 405822 442658 405854 442894
rect 405234 442574 405854 442658
rect 405234 442338 405266 442574
rect 405502 442338 405586 442574
rect 405822 442338 405854 442574
rect 405234 406894 405854 442338
rect 405234 406658 405266 406894
rect 405502 406658 405586 406894
rect 405822 406658 405854 406894
rect 405234 406574 405854 406658
rect 405234 406338 405266 406574
rect 405502 406338 405586 406574
rect 405822 406338 405854 406574
rect 405234 370894 405854 406338
rect 405234 370658 405266 370894
rect 405502 370658 405586 370894
rect 405822 370658 405854 370894
rect 405234 370574 405854 370658
rect 405234 370338 405266 370574
rect 405502 370338 405586 370574
rect 405822 370338 405854 370574
rect 405234 334894 405854 370338
rect 405234 334658 405266 334894
rect 405502 334658 405586 334894
rect 405822 334658 405854 334894
rect 405234 334574 405854 334658
rect 405234 334338 405266 334574
rect 405502 334338 405586 334574
rect 405822 334338 405854 334574
rect 404417 327454 404737 327486
rect 404417 327218 404459 327454
rect 404695 327218 404737 327454
rect 404417 327134 404737 327218
rect 404417 326898 404459 327134
rect 404695 326898 404737 327134
rect 404417 326866 404737 326898
rect 401514 294938 401546 295174
rect 401782 294938 401866 295174
rect 402102 294938 402134 295174
rect 401514 294854 402134 294938
rect 401514 294618 401546 294854
rect 401782 294618 401866 294854
rect 402102 294618 402134 294854
rect 401514 259174 402134 294618
rect 401514 258938 401546 259174
rect 401782 258938 401866 259174
rect 402102 258938 402134 259174
rect 401514 258854 402134 258938
rect 401514 258618 401546 258854
rect 401782 258618 401866 258854
rect 402102 258618 402134 258854
rect 401514 223174 402134 258618
rect 401514 222938 401546 223174
rect 401782 222938 401866 223174
rect 402102 222938 402134 223174
rect 401514 222854 402134 222938
rect 401514 222618 401546 222854
rect 401782 222618 401866 222854
rect 402102 222618 402134 222854
rect 401514 187174 402134 222618
rect 401514 186938 401546 187174
rect 401782 186938 401866 187174
rect 402102 186938 402134 187174
rect 401514 186854 402134 186938
rect 401514 186618 401546 186854
rect 401782 186618 401866 186854
rect 402102 186618 402134 186854
rect 401514 151174 402134 186618
rect 401514 150938 401546 151174
rect 401782 150938 401866 151174
rect 402102 150938 402134 151174
rect 401514 150854 402134 150938
rect 401514 150618 401546 150854
rect 401782 150618 401866 150854
rect 402102 150618 402134 150854
rect 401514 115174 402134 150618
rect 401514 114938 401546 115174
rect 401782 114938 401866 115174
rect 402102 114938 402134 115174
rect 401514 114854 402134 114938
rect 401514 114618 401546 114854
rect 401782 114618 401866 114854
rect 402102 114618 402134 114854
rect 401514 92137 402134 114618
rect 405234 298894 405854 334338
rect 408954 707718 409574 711590
rect 408954 707482 408986 707718
rect 409222 707482 409306 707718
rect 409542 707482 409574 707718
rect 408954 707398 409574 707482
rect 408954 707162 408986 707398
rect 409222 707162 409306 707398
rect 409542 707162 409574 707398
rect 408954 698614 409574 707162
rect 408954 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 409574 698614
rect 408954 698294 409574 698378
rect 408954 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 409574 698294
rect 408954 662614 409574 698058
rect 408954 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 409574 662614
rect 408954 662294 409574 662378
rect 408954 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 409574 662294
rect 408954 626614 409574 662058
rect 408954 626378 408986 626614
rect 409222 626378 409306 626614
rect 409542 626378 409574 626614
rect 408954 626294 409574 626378
rect 408954 626058 408986 626294
rect 409222 626058 409306 626294
rect 409542 626058 409574 626294
rect 408954 590614 409574 626058
rect 408954 590378 408986 590614
rect 409222 590378 409306 590614
rect 409542 590378 409574 590614
rect 408954 590294 409574 590378
rect 408954 590058 408986 590294
rect 409222 590058 409306 590294
rect 409542 590058 409574 590294
rect 408954 554614 409574 590058
rect 408954 554378 408986 554614
rect 409222 554378 409306 554614
rect 409542 554378 409574 554614
rect 408954 554294 409574 554378
rect 408954 554058 408986 554294
rect 409222 554058 409306 554294
rect 409542 554058 409574 554294
rect 408954 518614 409574 554058
rect 408954 518378 408986 518614
rect 409222 518378 409306 518614
rect 409542 518378 409574 518614
rect 408954 518294 409574 518378
rect 408954 518058 408986 518294
rect 409222 518058 409306 518294
rect 409542 518058 409574 518294
rect 408954 482614 409574 518058
rect 408954 482378 408986 482614
rect 409222 482378 409306 482614
rect 409542 482378 409574 482614
rect 408954 482294 409574 482378
rect 408954 482058 408986 482294
rect 409222 482058 409306 482294
rect 409542 482058 409574 482294
rect 408954 446614 409574 482058
rect 408954 446378 408986 446614
rect 409222 446378 409306 446614
rect 409542 446378 409574 446614
rect 408954 446294 409574 446378
rect 408954 446058 408986 446294
rect 409222 446058 409306 446294
rect 409542 446058 409574 446294
rect 408954 410614 409574 446058
rect 408954 410378 408986 410614
rect 409222 410378 409306 410614
rect 409542 410378 409574 410614
rect 408954 410294 409574 410378
rect 408954 410058 408986 410294
rect 409222 410058 409306 410294
rect 409542 410058 409574 410294
rect 408954 374614 409574 410058
rect 408954 374378 408986 374614
rect 409222 374378 409306 374614
rect 409542 374378 409574 374614
rect 408954 374294 409574 374378
rect 408954 374058 408986 374294
rect 409222 374058 409306 374294
rect 409542 374058 409574 374294
rect 408954 338614 409574 374058
rect 408954 338378 408986 338614
rect 409222 338378 409306 338614
rect 409542 338378 409574 338614
rect 408954 338294 409574 338378
rect 408954 338058 408986 338294
rect 409222 338058 409306 338294
rect 409542 338058 409574 338294
rect 407890 331174 408210 331206
rect 407890 330938 407932 331174
rect 408168 330938 408210 331174
rect 407890 330854 408210 330938
rect 407890 330618 407932 330854
rect 408168 330618 408210 330854
rect 407890 330586 408210 330618
rect 405234 298658 405266 298894
rect 405502 298658 405586 298894
rect 405822 298658 405854 298894
rect 405234 298574 405854 298658
rect 405234 298338 405266 298574
rect 405502 298338 405586 298574
rect 405822 298338 405854 298574
rect 405234 262894 405854 298338
rect 405234 262658 405266 262894
rect 405502 262658 405586 262894
rect 405822 262658 405854 262894
rect 405234 262574 405854 262658
rect 405234 262338 405266 262574
rect 405502 262338 405586 262574
rect 405822 262338 405854 262574
rect 405234 226894 405854 262338
rect 405234 226658 405266 226894
rect 405502 226658 405586 226894
rect 405822 226658 405854 226894
rect 405234 226574 405854 226658
rect 405234 226338 405266 226574
rect 405502 226338 405586 226574
rect 405822 226338 405854 226574
rect 405234 190894 405854 226338
rect 405234 190658 405266 190894
rect 405502 190658 405586 190894
rect 405822 190658 405854 190894
rect 405234 190574 405854 190658
rect 405234 190338 405266 190574
rect 405502 190338 405586 190574
rect 405822 190338 405854 190574
rect 405234 154894 405854 190338
rect 405234 154658 405266 154894
rect 405502 154658 405586 154894
rect 405822 154658 405854 154894
rect 405234 154574 405854 154658
rect 405234 154338 405266 154574
rect 405502 154338 405586 154574
rect 405822 154338 405854 154574
rect 405234 118894 405854 154338
rect 405234 118658 405266 118894
rect 405502 118658 405586 118894
rect 405822 118658 405854 118894
rect 405234 118574 405854 118658
rect 405234 118338 405266 118574
rect 405502 118338 405586 118574
rect 405822 118338 405854 118574
rect 405234 104460 405854 118338
rect 408954 302614 409574 338058
rect 412674 708678 413294 711590
rect 412674 708442 412706 708678
rect 412942 708442 413026 708678
rect 413262 708442 413294 708678
rect 412674 708358 413294 708442
rect 412674 708122 412706 708358
rect 412942 708122 413026 708358
rect 413262 708122 413294 708358
rect 412674 666334 413294 708122
rect 412674 666098 412706 666334
rect 412942 666098 413026 666334
rect 413262 666098 413294 666334
rect 412674 666014 413294 666098
rect 412674 665778 412706 666014
rect 412942 665778 413026 666014
rect 413262 665778 413294 666014
rect 412674 630334 413294 665778
rect 412674 630098 412706 630334
rect 412942 630098 413026 630334
rect 413262 630098 413294 630334
rect 412674 630014 413294 630098
rect 412674 629778 412706 630014
rect 412942 629778 413026 630014
rect 413262 629778 413294 630014
rect 412674 594334 413294 629778
rect 412674 594098 412706 594334
rect 412942 594098 413026 594334
rect 413262 594098 413294 594334
rect 412674 594014 413294 594098
rect 412674 593778 412706 594014
rect 412942 593778 413026 594014
rect 413262 593778 413294 594014
rect 412674 558334 413294 593778
rect 412674 558098 412706 558334
rect 412942 558098 413026 558334
rect 413262 558098 413294 558334
rect 412674 558014 413294 558098
rect 412674 557778 412706 558014
rect 412942 557778 413026 558014
rect 413262 557778 413294 558014
rect 412674 522334 413294 557778
rect 412674 522098 412706 522334
rect 412942 522098 413026 522334
rect 413262 522098 413294 522334
rect 412674 522014 413294 522098
rect 412674 521778 412706 522014
rect 412942 521778 413026 522014
rect 413262 521778 413294 522014
rect 412674 486334 413294 521778
rect 412674 486098 412706 486334
rect 412942 486098 413026 486334
rect 413262 486098 413294 486334
rect 412674 486014 413294 486098
rect 412674 485778 412706 486014
rect 412942 485778 413026 486014
rect 413262 485778 413294 486014
rect 412674 450334 413294 485778
rect 412674 450098 412706 450334
rect 412942 450098 413026 450334
rect 413262 450098 413294 450334
rect 412674 450014 413294 450098
rect 412674 449778 412706 450014
rect 412942 449778 413026 450014
rect 413262 449778 413294 450014
rect 412674 414334 413294 449778
rect 412674 414098 412706 414334
rect 412942 414098 413026 414334
rect 413262 414098 413294 414334
rect 412674 414014 413294 414098
rect 412674 413778 412706 414014
rect 412942 413778 413026 414014
rect 413262 413778 413294 414014
rect 412674 378334 413294 413778
rect 412674 378098 412706 378334
rect 412942 378098 413026 378334
rect 413262 378098 413294 378334
rect 412674 378014 413294 378098
rect 412674 377778 412706 378014
rect 412942 377778 413026 378014
rect 413262 377778 413294 378014
rect 412674 342334 413294 377778
rect 412674 342098 412706 342334
rect 412942 342098 413026 342334
rect 413262 342098 413294 342334
rect 412674 342014 413294 342098
rect 412674 341778 412706 342014
rect 412942 341778 413026 342014
rect 413262 341778 413294 342014
rect 411363 327454 411683 327486
rect 411363 327218 411405 327454
rect 411641 327218 411683 327454
rect 411363 327134 411683 327218
rect 411363 326898 411405 327134
rect 411641 326898 411683 327134
rect 411363 326866 411683 326898
rect 408954 302378 408986 302614
rect 409222 302378 409306 302614
rect 409542 302378 409574 302614
rect 408954 302294 409574 302378
rect 408954 302058 408986 302294
rect 409222 302058 409306 302294
rect 409542 302058 409574 302294
rect 408954 266614 409574 302058
rect 408954 266378 408986 266614
rect 409222 266378 409306 266614
rect 409542 266378 409574 266614
rect 408954 266294 409574 266378
rect 408954 266058 408986 266294
rect 409222 266058 409306 266294
rect 409542 266058 409574 266294
rect 408954 230614 409574 266058
rect 408954 230378 408986 230614
rect 409222 230378 409306 230614
rect 409542 230378 409574 230614
rect 408954 230294 409574 230378
rect 408954 230058 408986 230294
rect 409222 230058 409306 230294
rect 409542 230058 409574 230294
rect 408954 194614 409574 230058
rect 408954 194378 408986 194614
rect 409222 194378 409306 194614
rect 409542 194378 409574 194614
rect 408954 194294 409574 194378
rect 408954 194058 408986 194294
rect 409222 194058 409306 194294
rect 409542 194058 409574 194294
rect 408954 158614 409574 194058
rect 408954 158378 408986 158614
rect 409222 158378 409306 158614
rect 409542 158378 409574 158614
rect 408954 158294 409574 158378
rect 408954 158058 408986 158294
rect 409222 158058 409306 158294
rect 409542 158058 409574 158294
rect 408954 122614 409574 158058
rect 408954 122378 408986 122614
rect 409222 122378 409306 122614
rect 409542 122378 409574 122614
rect 408954 122294 409574 122378
rect 408954 122058 408986 122294
rect 409222 122058 409306 122294
rect 409542 122058 409574 122294
rect 408954 92137 409574 122058
rect 412674 306334 413294 341778
rect 416394 709638 417014 711590
rect 416394 709402 416426 709638
rect 416662 709402 416746 709638
rect 416982 709402 417014 709638
rect 416394 709318 417014 709402
rect 416394 709082 416426 709318
rect 416662 709082 416746 709318
rect 416982 709082 417014 709318
rect 416394 670054 417014 709082
rect 416394 669818 416426 670054
rect 416662 669818 416746 670054
rect 416982 669818 417014 670054
rect 416394 669734 417014 669818
rect 416394 669498 416426 669734
rect 416662 669498 416746 669734
rect 416982 669498 417014 669734
rect 416394 634054 417014 669498
rect 416394 633818 416426 634054
rect 416662 633818 416746 634054
rect 416982 633818 417014 634054
rect 416394 633734 417014 633818
rect 416394 633498 416426 633734
rect 416662 633498 416746 633734
rect 416982 633498 417014 633734
rect 416394 598054 417014 633498
rect 416394 597818 416426 598054
rect 416662 597818 416746 598054
rect 416982 597818 417014 598054
rect 416394 597734 417014 597818
rect 416394 597498 416426 597734
rect 416662 597498 416746 597734
rect 416982 597498 417014 597734
rect 416394 562054 417014 597498
rect 416394 561818 416426 562054
rect 416662 561818 416746 562054
rect 416982 561818 417014 562054
rect 416394 561734 417014 561818
rect 416394 561498 416426 561734
rect 416662 561498 416746 561734
rect 416982 561498 417014 561734
rect 416394 526054 417014 561498
rect 416394 525818 416426 526054
rect 416662 525818 416746 526054
rect 416982 525818 417014 526054
rect 416394 525734 417014 525818
rect 416394 525498 416426 525734
rect 416662 525498 416746 525734
rect 416982 525498 417014 525734
rect 416394 490054 417014 525498
rect 416394 489818 416426 490054
rect 416662 489818 416746 490054
rect 416982 489818 417014 490054
rect 416394 489734 417014 489818
rect 416394 489498 416426 489734
rect 416662 489498 416746 489734
rect 416982 489498 417014 489734
rect 416394 454054 417014 489498
rect 416394 453818 416426 454054
rect 416662 453818 416746 454054
rect 416982 453818 417014 454054
rect 416394 453734 417014 453818
rect 416394 453498 416426 453734
rect 416662 453498 416746 453734
rect 416982 453498 417014 453734
rect 416394 418054 417014 453498
rect 416394 417818 416426 418054
rect 416662 417818 416746 418054
rect 416982 417818 417014 418054
rect 416394 417734 417014 417818
rect 416394 417498 416426 417734
rect 416662 417498 416746 417734
rect 416982 417498 417014 417734
rect 416394 382054 417014 417498
rect 416394 381818 416426 382054
rect 416662 381818 416746 382054
rect 416982 381818 417014 382054
rect 416394 381734 417014 381818
rect 416394 381498 416426 381734
rect 416662 381498 416746 381734
rect 416982 381498 417014 381734
rect 416394 346054 417014 381498
rect 416394 345818 416426 346054
rect 416662 345818 416746 346054
rect 416982 345818 417014 346054
rect 416394 345734 417014 345818
rect 416394 345498 416426 345734
rect 416662 345498 416746 345734
rect 416982 345498 417014 345734
rect 414836 331174 415156 331206
rect 414836 330938 414878 331174
rect 415114 330938 415156 331174
rect 414836 330854 415156 330938
rect 414836 330618 414878 330854
rect 415114 330618 415156 330854
rect 414836 330586 415156 330618
rect 412674 306098 412706 306334
rect 412942 306098 413026 306334
rect 413262 306098 413294 306334
rect 412674 306014 413294 306098
rect 412674 305778 412706 306014
rect 412942 305778 413026 306014
rect 413262 305778 413294 306014
rect 412674 270334 413294 305778
rect 412674 270098 412706 270334
rect 412942 270098 413026 270334
rect 413262 270098 413294 270334
rect 412674 270014 413294 270098
rect 412674 269778 412706 270014
rect 412942 269778 413026 270014
rect 413262 269778 413294 270014
rect 412674 234334 413294 269778
rect 412674 234098 412706 234334
rect 412942 234098 413026 234334
rect 413262 234098 413294 234334
rect 412674 234014 413294 234098
rect 412674 233778 412706 234014
rect 412942 233778 413026 234014
rect 413262 233778 413294 234014
rect 412674 198334 413294 233778
rect 412674 198098 412706 198334
rect 412942 198098 413026 198334
rect 413262 198098 413294 198334
rect 412674 198014 413294 198098
rect 412674 197778 412706 198014
rect 412942 197778 413026 198014
rect 413262 197778 413294 198014
rect 412674 162334 413294 197778
rect 412674 162098 412706 162334
rect 412942 162098 413026 162334
rect 413262 162098 413294 162334
rect 412674 162014 413294 162098
rect 412674 161778 412706 162014
rect 412942 161778 413026 162014
rect 413262 161778 413294 162014
rect 412674 126334 413294 161778
rect 416394 310054 417014 345498
rect 420114 710598 420734 711590
rect 420114 710362 420146 710598
rect 420382 710362 420466 710598
rect 420702 710362 420734 710598
rect 420114 710278 420734 710362
rect 420114 710042 420146 710278
rect 420382 710042 420466 710278
rect 420702 710042 420734 710278
rect 420114 673774 420734 710042
rect 420114 673538 420146 673774
rect 420382 673538 420466 673774
rect 420702 673538 420734 673774
rect 420114 673454 420734 673538
rect 420114 673218 420146 673454
rect 420382 673218 420466 673454
rect 420702 673218 420734 673454
rect 420114 637774 420734 673218
rect 420114 637538 420146 637774
rect 420382 637538 420466 637774
rect 420702 637538 420734 637774
rect 420114 637454 420734 637538
rect 420114 637218 420146 637454
rect 420382 637218 420466 637454
rect 420702 637218 420734 637454
rect 420114 601774 420734 637218
rect 420114 601538 420146 601774
rect 420382 601538 420466 601774
rect 420702 601538 420734 601774
rect 420114 601454 420734 601538
rect 420114 601218 420146 601454
rect 420382 601218 420466 601454
rect 420702 601218 420734 601454
rect 420114 565774 420734 601218
rect 420114 565538 420146 565774
rect 420382 565538 420466 565774
rect 420702 565538 420734 565774
rect 420114 565454 420734 565538
rect 420114 565218 420146 565454
rect 420382 565218 420466 565454
rect 420702 565218 420734 565454
rect 420114 529774 420734 565218
rect 420114 529538 420146 529774
rect 420382 529538 420466 529774
rect 420702 529538 420734 529774
rect 420114 529454 420734 529538
rect 420114 529218 420146 529454
rect 420382 529218 420466 529454
rect 420702 529218 420734 529454
rect 420114 493774 420734 529218
rect 420114 493538 420146 493774
rect 420382 493538 420466 493774
rect 420702 493538 420734 493774
rect 420114 493454 420734 493538
rect 420114 493218 420146 493454
rect 420382 493218 420466 493454
rect 420702 493218 420734 493454
rect 420114 457774 420734 493218
rect 420114 457538 420146 457774
rect 420382 457538 420466 457774
rect 420702 457538 420734 457774
rect 420114 457454 420734 457538
rect 420114 457218 420146 457454
rect 420382 457218 420466 457454
rect 420702 457218 420734 457454
rect 420114 421774 420734 457218
rect 423834 711558 424454 711590
rect 423834 711322 423866 711558
rect 424102 711322 424186 711558
rect 424422 711322 424454 711558
rect 423834 711238 424454 711322
rect 423834 711002 423866 711238
rect 424102 711002 424186 711238
rect 424422 711002 424454 711238
rect 423834 677494 424454 711002
rect 423834 677258 423866 677494
rect 424102 677258 424186 677494
rect 424422 677258 424454 677494
rect 423834 677174 424454 677258
rect 423834 676938 423866 677174
rect 424102 676938 424186 677174
rect 424422 676938 424454 677174
rect 423834 641494 424454 676938
rect 423834 641258 423866 641494
rect 424102 641258 424186 641494
rect 424422 641258 424454 641494
rect 423834 641174 424454 641258
rect 423834 640938 423866 641174
rect 424102 640938 424186 641174
rect 424422 640938 424454 641174
rect 423834 605494 424454 640938
rect 423834 605258 423866 605494
rect 424102 605258 424186 605494
rect 424422 605258 424454 605494
rect 423834 605174 424454 605258
rect 423834 604938 423866 605174
rect 424102 604938 424186 605174
rect 424422 604938 424454 605174
rect 423834 569494 424454 604938
rect 423834 569258 423866 569494
rect 424102 569258 424186 569494
rect 424422 569258 424454 569494
rect 423834 569174 424454 569258
rect 423834 568938 423866 569174
rect 424102 568938 424186 569174
rect 424422 568938 424454 569174
rect 423834 533494 424454 568938
rect 423834 533258 423866 533494
rect 424102 533258 424186 533494
rect 424422 533258 424454 533494
rect 423834 533174 424454 533258
rect 423834 532938 423866 533174
rect 424102 532938 424186 533174
rect 424422 532938 424454 533174
rect 423834 497494 424454 532938
rect 423834 497258 423866 497494
rect 424102 497258 424186 497494
rect 424422 497258 424454 497494
rect 423834 497174 424454 497258
rect 423834 496938 423866 497174
rect 424102 496938 424186 497174
rect 424422 496938 424454 497174
rect 423834 461494 424454 496938
rect 423834 461258 423866 461494
rect 424102 461258 424186 461494
rect 424422 461258 424454 461494
rect 423834 461174 424454 461258
rect 423834 460938 423866 461174
rect 424102 460938 424186 461174
rect 424422 460938 424454 461174
rect 423834 444412 424454 460938
rect 433794 704838 434414 711590
rect 433794 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 434414 704838
rect 433794 704518 434414 704602
rect 433794 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 434414 704518
rect 433794 687454 434414 704282
rect 433794 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 434414 687454
rect 433794 687134 434414 687218
rect 433794 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 434414 687134
rect 433794 651454 434414 686898
rect 433794 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 434414 651454
rect 433794 651134 434414 651218
rect 433794 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 434414 651134
rect 433794 615454 434414 650898
rect 433794 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 434414 615454
rect 433794 615134 434414 615218
rect 433794 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 434414 615134
rect 433794 579454 434414 614898
rect 433794 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 434414 579454
rect 433794 579134 434414 579218
rect 433794 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 434414 579134
rect 433794 543454 434414 578898
rect 433794 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 434414 543454
rect 433794 543134 434414 543218
rect 433794 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 434414 543134
rect 433794 507454 434414 542898
rect 433794 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 434414 507454
rect 433794 507134 434414 507218
rect 433794 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 434414 507134
rect 433794 471454 434414 506898
rect 433794 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 434414 471454
rect 433794 471134 434414 471218
rect 433794 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 434414 471134
rect 433794 442833 434414 470898
rect 437514 705798 438134 711590
rect 437514 705562 437546 705798
rect 437782 705562 437866 705798
rect 438102 705562 438134 705798
rect 437514 705478 438134 705562
rect 437514 705242 437546 705478
rect 437782 705242 437866 705478
rect 438102 705242 438134 705478
rect 437514 691174 438134 705242
rect 437514 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 438134 691174
rect 437514 690854 438134 690938
rect 437514 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 438134 690854
rect 437514 655174 438134 690618
rect 437514 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 438134 655174
rect 437514 654854 438134 654938
rect 437514 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 438134 654854
rect 437514 619174 438134 654618
rect 437514 618938 437546 619174
rect 437782 618938 437866 619174
rect 438102 618938 438134 619174
rect 437514 618854 438134 618938
rect 437514 618618 437546 618854
rect 437782 618618 437866 618854
rect 438102 618618 438134 618854
rect 437514 583174 438134 618618
rect 437514 582938 437546 583174
rect 437782 582938 437866 583174
rect 438102 582938 438134 583174
rect 437514 582854 438134 582938
rect 437514 582618 437546 582854
rect 437782 582618 437866 582854
rect 438102 582618 438134 582854
rect 437514 547174 438134 582618
rect 437514 546938 437546 547174
rect 437782 546938 437866 547174
rect 438102 546938 438134 547174
rect 437514 546854 438134 546938
rect 437514 546618 437546 546854
rect 437782 546618 437866 546854
rect 438102 546618 438134 546854
rect 437514 511174 438134 546618
rect 437514 510938 437546 511174
rect 437782 510938 437866 511174
rect 438102 510938 438134 511174
rect 437514 510854 438134 510938
rect 437514 510618 437546 510854
rect 437782 510618 437866 510854
rect 438102 510618 438134 510854
rect 437514 475174 438134 510618
rect 437514 474938 437546 475174
rect 437782 474938 437866 475174
rect 438102 474938 438134 475174
rect 437514 474854 438134 474938
rect 437514 474618 437546 474854
rect 437782 474618 437866 474854
rect 438102 474618 438134 474854
rect 437514 444412 438134 474618
rect 441234 706758 441854 711590
rect 441234 706522 441266 706758
rect 441502 706522 441586 706758
rect 441822 706522 441854 706758
rect 441234 706438 441854 706522
rect 441234 706202 441266 706438
rect 441502 706202 441586 706438
rect 441822 706202 441854 706438
rect 441234 694894 441854 706202
rect 441234 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 441854 694894
rect 441234 694574 441854 694658
rect 441234 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 441854 694574
rect 441234 658894 441854 694338
rect 444954 707718 445574 711590
rect 444954 707482 444986 707718
rect 445222 707482 445306 707718
rect 445542 707482 445574 707718
rect 444954 707398 445574 707482
rect 444954 707162 444986 707398
rect 445222 707162 445306 707398
rect 445542 707162 445574 707398
rect 444954 698614 445574 707162
rect 448674 708678 449294 711590
rect 448674 708442 448706 708678
rect 448942 708442 449026 708678
rect 449262 708442 449294 708678
rect 448674 708358 449294 708442
rect 448674 708122 448706 708358
rect 448942 708122 449026 708358
rect 449262 708122 449294 708358
rect 447915 700636 447981 700637
rect 447915 700572 447916 700636
rect 447980 700572 447981 700636
rect 447915 700571 447981 700572
rect 447731 700364 447797 700365
rect 447731 700300 447732 700364
rect 447796 700300 447797 700364
rect 447731 700299 447797 700300
rect 444954 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 445574 698614
rect 444954 698294 445574 698378
rect 444954 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 445574 698294
rect 444235 689348 444301 689349
rect 444235 689284 444236 689348
rect 444300 689284 444301 689348
rect 444235 689283 444301 689284
rect 441234 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 441854 658894
rect 441234 658574 441854 658658
rect 441234 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 441854 658574
rect 441234 622894 441854 658338
rect 441234 622658 441266 622894
rect 441502 622658 441586 622894
rect 441822 622658 441854 622894
rect 441234 622574 441854 622658
rect 441234 622338 441266 622574
rect 441502 622338 441586 622574
rect 441822 622338 441854 622574
rect 441234 586894 441854 622338
rect 441234 586658 441266 586894
rect 441502 586658 441586 586894
rect 441822 586658 441854 586894
rect 441234 586574 441854 586658
rect 441234 586338 441266 586574
rect 441502 586338 441586 586574
rect 441822 586338 441854 586574
rect 441234 550894 441854 586338
rect 441234 550658 441266 550894
rect 441502 550658 441586 550894
rect 441822 550658 441854 550894
rect 441234 550574 441854 550658
rect 441234 550338 441266 550574
rect 441502 550338 441586 550574
rect 441822 550338 441854 550574
rect 441234 514894 441854 550338
rect 441234 514658 441266 514894
rect 441502 514658 441586 514894
rect 441822 514658 441854 514894
rect 441234 514574 441854 514658
rect 441234 514338 441266 514574
rect 441502 514338 441586 514574
rect 441822 514338 441854 514574
rect 441234 478894 441854 514338
rect 441234 478658 441266 478894
rect 441502 478658 441586 478894
rect 441822 478658 441854 478894
rect 441234 478574 441854 478658
rect 441234 478338 441266 478574
rect 441502 478338 441586 478574
rect 441822 478338 441854 478574
rect 441234 442833 441854 478338
rect 426624 439174 426944 439206
rect 426624 438938 426666 439174
rect 426902 438938 426944 439174
rect 426624 438854 426944 438938
rect 426624 438618 426666 438854
rect 426902 438618 426944 438854
rect 426624 438586 426944 438618
rect 432305 439174 432625 439206
rect 432305 438938 432347 439174
rect 432583 438938 432625 439174
rect 432305 438854 432625 438938
rect 432305 438618 432347 438854
rect 432583 438618 432625 438854
rect 432305 438586 432625 438618
rect 437986 439174 438306 439206
rect 437986 438938 438028 439174
rect 438264 438938 438306 439174
rect 437986 438854 438306 438938
rect 437986 438618 438028 438854
rect 438264 438618 438306 438854
rect 437986 438586 438306 438618
rect 443667 439174 443987 439206
rect 443667 438938 443709 439174
rect 443945 438938 443987 439174
rect 443667 438854 443987 438938
rect 443667 438618 443709 438854
rect 443945 438618 443987 438854
rect 443667 438586 443987 438618
rect 423784 435454 424104 435486
rect 423784 435218 423826 435454
rect 424062 435218 424104 435454
rect 423784 435134 424104 435218
rect 423784 434898 423826 435134
rect 424062 434898 424104 435134
rect 423784 434866 424104 434898
rect 429465 435454 429785 435486
rect 429465 435218 429507 435454
rect 429743 435218 429785 435454
rect 429465 435134 429785 435218
rect 429465 434898 429507 435134
rect 429743 434898 429785 435134
rect 429465 434866 429785 434898
rect 435146 435454 435466 435486
rect 435146 435218 435188 435454
rect 435424 435218 435466 435454
rect 435146 435134 435466 435218
rect 435146 434898 435188 435134
rect 435424 434898 435466 435134
rect 435146 434866 435466 434898
rect 440827 435454 441147 435486
rect 440827 435218 440869 435454
rect 441105 435218 441147 435454
rect 440827 435134 441147 435218
rect 440827 434898 440869 435134
rect 441105 434898 441147 435134
rect 440827 434866 441147 434898
rect 420114 421538 420146 421774
rect 420382 421538 420466 421774
rect 420702 421538 420734 421774
rect 420114 421454 420734 421538
rect 420114 421218 420146 421454
rect 420382 421218 420466 421454
rect 420702 421218 420734 421454
rect 420114 385774 420734 421218
rect 420114 385538 420146 385774
rect 420382 385538 420466 385774
rect 420702 385538 420734 385774
rect 420114 385454 420734 385538
rect 420114 385218 420146 385454
rect 420382 385218 420466 385454
rect 420702 385218 420734 385454
rect 420114 349774 420734 385218
rect 420114 349538 420146 349774
rect 420382 349538 420466 349774
rect 420702 349538 420734 349774
rect 420114 349454 420734 349538
rect 420114 349218 420146 349454
rect 420382 349218 420466 349454
rect 420702 349218 420734 349454
rect 418309 327454 418629 327486
rect 418309 327218 418351 327454
rect 418587 327218 418629 327454
rect 418309 327134 418629 327218
rect 418309 326898 418351 327134
rect 418587 326898 418629 327134
rect 418309 326866 418629 326898
rect 416394 309818 416426 310054
rect 416662 309818 416746 310054
rect 416982 309818 417014 310054
rect 416394 309734 417014 309818
rect 416394 309498 416426 309734
rect 416662 309498 416746 309734
rect 416982 309498 417014 309734
rect 416394 274054 417014 309498
rect 416394 273818 416426 274054
rect 416662 273818 416746 274054
rect 416982 273818 417014 274054
rect 416394 273734 417014 273818
rect 416394 273498 416426 273734
rect 416662 273498 416746 273734
rect 416982 273498 417014 273734
rect 416394 238054 417014 273498
rect 416394 237818 416426 238054
rect 416662 237818 416746 238054
rect 416982 237818 417014 238054
rect 416394 237734 417014 237818
rect 416394 237498 416426 237734
rect 416662 237498 416746 237734
rect 416982 237498 417014 237734
rect 416394 202054 417014 237498
rect 416394 201818 416426 202054
rect 416662 201818 416746 202054
rect 416982 201818 417014 202054
rect 416394 201734 417014 201818
rect 416394 201498 416426 201734
rect 416662 201498 416746 201734
rect 416982 201498 417014 201734
rect 416394 166054 417014 201498
rect 416394 165818 416426 166054
rect 416662 165818 416746 166054
rect 416982 165818 417014 166054
rect 416394 165734 417014 165818
rect 416394 165498 416426 165734
rect 416662 165498 416746 165734
rect 416982 165498 417014 165734
rect 416394 157249 417014 165498
rect 420114 313774 420734 349218
rect 423834 389494 424454 420068
rect 423834 389258 423866 389494
rect 424102 389258 424186 389494
rect 424422 389258 424454 389494
rect 423834 389174 424454 389258
rect 423834 388938 423866 389174
rect 424102 388938 424186 389174
rect 424422 388938 424454 389174
rect 423834 353494 424454 388938
rect 423834 353258 423866 353494
rect 424102 353258 424186 353494
rect 424422 353258 424454 353494
rect 423834 353174 424454 353258
rect 423834 352938 423866 353174
rect 424102 352938 424186 353174
rect 424422 352938 424454 353174
rect 421419 334116 421485 334117
rect 421419 334052 421420 334116
rect 421484 334052 421485 334116
rect 421419 334051 421485 334052
rect 420114 313538 420146 313774
rect 420382 313538 420466 313774
rect 420702 313538 420734 313774
rect 420114 313454 420734 313538
rect 420114 313218 420146 313454
rect 420382 313218 420466 313454
rect 420702 313218 420734 313454
rect 420114 277774 420734 313218
rect 420114 277538 420146 277774
rect 420382 277538 420466 277774
rect 420702 277538 420734 277774
rect 420114 277454 420734 277538
rect 420114 277218 420146 277454
rect 420382 277218 420466 277454
rect 420702 277218 420734 277454
rect 420114 241774 420734 277218
rect 420114 241538 420146 241774
rect 420382 241538 420466 241774
rect 420702 241538 420734 241774
rect 420114 241454 420734 241538
rect 420114 241218 420146 241454
rect 420382 241218 420466 241454
rect 420702 241218 420734 241454
rect 420114 205774 420734 241218
rect 420114 205538 420146 205774
rect 420382 205538 420466 205774
rect 420702 205538 420734 205774
rect 420114 205454 420734 205538
rect 420114 205218 420146 205454
rect 420382 205218 420466 205454
rect 420702 205218 420734 205454
rect 420114 169774 420734 205218
rect 420114 169538 420146 169774
rect 420382 169538 420466 169774
rect 420702 169538 420734 169774
rect 420114 169454 420734 169538
rect 420114 169218 420146 169454
rect 420382 169218 420466 169454
rect 420702 169218 420734 169454
rect 420114 157249 420734 169218
rect 421422 162757 421482 334051
rect 421782 331174 422102 331206
rect 421782 330938 421824 331174
rect 422060 330938 422102 331174
rect 421782 330854 422102 330938
rect 421782 330618 421824 330854
rect 422060 330618 422102 330854
rect 421782 330586 422102 330618
rect 423834 317494 424454 352938
rect 433794 399454 434414 422599
rect 433794 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 434414 399454
rect 433794 399134 434414 399218
rect 433794 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 434414 399134
rect 433794 363454 434414 398898
rect 433794 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 434414 363454
rect 433794 363134 434414 363218
rect 433794 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 434414 363134
rect 428411 334524 428477 334525
rect 428411 334460 428412 334524
rect 428476 334460 428477 334524
rect 428411 334459 428477 334460
rect 425835 334388 425901 334389
rect 425835 334324 425836 334388
rect 425900 334324 425901 334388
rect 425835 334323 425901 334324
rect 425255 327454 425575 327486
rect 425255 327218 425297 327454
rect 425533 327218 425575 327454
rect 425255 327134 425575 327218
rect 425255 326898 425297 327134
rect 425533 326898 425575 327134
rect 425255 326866 425575 326898
rect 423834 317258 423866 317494
rect 424102 317258 424186 317494
rect 424422 317258 424454 317494
rect 423834 317174 424454 317258
rect 423834 316938 423866 317174
rect 424102 316938 424186 317174
rect 424422 316938 424454 317174
rect 423834 281494 424454 316938
rect 423834 281258 423866 281494
rect 424102 281258 424186 281494
rect 424422 281258 424454 281494
rect 423834 281174 424454 281258
rect 423834 280938 423866 281174
rect 424102 280938 424186 281174
rect 424422 280938 424454 281174
rect 423834 245494 424454 280938
rect 423834 245258 423866 245494
rect 424102 245258 424186 245494
rect 424422 245258 424454 245494
rect 423834 245174 424454 245258
rect 423834 244938 423866 245174
rect 424102 244938 424186 245174
rect 424422 244938 424454 245174
rect 423834 209494 424454 244938
rect 423834 209258 423866 209494
rect 424102 209258 424186 209494
rect 424422 209258 424454 209494
rect 423834 209174 424454 209258
rect 423834 208938 423866 209174
rect 424102 208938 424186 209174
rect 424422 208938 424454 209174
rect 423834 173494 424454 208938
rect 423834 173258 423866 173494
rect 424102 173258 424186 173494
rect 424422 173258 424454 173494
rect 423834 173174 424454 173258
rect 423834 172938 423866 173174
rect 424102 172938 424186 173174
rect 424422 172938 424454 173174
rect 421419 162756 421485 162757
rect 421419 162692 421420 162756
rect 421484 162692 421485 162756
rect 421419 162691 421485 162692
rect 423834 157249 424454 172938
rect 425838 162757 425898 334323
rect 428414 162757 428474 334459
rect 428728 331174 429048 331206
rect 428728 330938 428770 331174
rect 429006 330938 429048 331174
rect 428728 330854 429048 330938
rect 428728 330618 428770 330854
rect 429006 330618 429048 330854
rect 428728 330586 429048 330618
rect 433794 327454 434414 362898
rect 433794 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 434414 327454
rect 433794 327134 434414 327218
rect 433794 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 434414 327134
rect 433794 291454 434414 326898
rect 433794 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 434414 291454
rect 433794 291134 434414 291218
rect 433794 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 434414 291134
rect 433794 255454 434414 290898
rect 433794 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 434414 255454
rect 433794 255134 434414 255218
rect 433794 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 434414 255134
rect 433794 219454 434414 254898
rect 433794 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 434414 219454
rect 433794 219134 434414 219218
rect 433794 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 434414 219134
rect 433794 183454 434414 218898
rect 433794 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 434414 183454
rect 433794 183134 434414 183218
rect 433794 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 434414 183134
rect 425835 162756 425901 162757
rect 425835 162692 425836 162756
rect 425900 162692 425901 162756
rect 425835 162691 425901 162692
rect 428411 162756 428477 162757
rect 428411 162692 428412 162756
rect 428476 162692 428477 162756
rect 428411 162691 428477 162692
rect 433794 157249 434414 182898
rect 437514 403174 438134 420068
rect 437514 402938 437546 403174
rect 437782 402938 437866 403174
rect 438102 402938 438134 403174
rect 437514 402854 438134 402938
rect 437514 402618 437546 402854
rect 437782 402618 437866 402854
rect 438102 402618 438134 402854
rect 437514 367174 438134 402618
rect 437514 366938 437546 367174
rect 437782 366938 437866 367174
rect 438102 366938 438134 367174
rect 437514 366854 438134 366938
rect 437514 366618 437546 366854
rect 437782 366618 437866 366854
rect 438102 366618 438134 366854
rect 437514 331174 438134 366618
rect 437514 330938 437546 331174
rect 437782 330938 437866 331174
rect 438102 330938 438134 331174
rect 437514 330854 438134 330938
rect 437514 330618 437546 330854
rect 437782 330618 437866 330854
rect 438102 330618 438134 330854
rect 437514 295174 438134 330618
rect 437514 294938 437546 295174
rect 437782 294938 437866 295174
rect 438102 294938 438134 295174
rect 437514 294854 438134 294938
rect 437514 294618 437546 294854
rect 437782 294618 437866 294854
rect 438102 294618 438134 294854
rect 437514 259174 438134 294618
rect 437514 258938 437546 259174
rect 437782 258938 437866 259174
rect 438102 258938 438134 259174
rect 437514 258854 438134 258938
rect 437514 258618 437546 258854
rect 437782 258618 437866 258854
rect 438102 258618 438134 258854
rect 437514 223174 438134 258618
rect 437514 222938 437546 223174
rect 437782 222938 437866 223174
rect 438102 222938 438134 223174
rect 437514 222854 438134 222938
rect 437514 222618 437546 222854
rect 437782 222618 437866 222854
rect 438102 222618 438134 222854
rect 437514 187174 438134 222618
rect 437514 186938 437546 187174
rect 437782 186938 437866 187174
rect 438102 186938 438134 187174
rect 437514 186854 438134 186938
rect 437514 186618 437546 186854
rect 437782 186618 437866 186854
rect 438102 186618 438134 186854
rect 437514 157249 438134 186618
rect 441234 406894 441854 422599
rect 444051 421972 444117 421973
rect 444051 421908 444052 421972
rect 444116 421908 444117 421972
rect 444051 421907 444117 421908
rect 441234 406658 441266 406894
rect 441502 406658 441586 406894
rect 441822 406658 441854 406894
rect 441234 406574 441854 406658
rect 441234 406338 441266 406574
rect 441502 406338 441586 406574
rect 441822 406338 441854 406574
rect 441234 370894 441854 406338
rect 441234 370658 441266 370894
rect 441502 370658 441586 370894
rect 441822 370658 441854 370894
rect 441234 370574 441854 370658
rect 441234 370338 441266 370574
rect 441502 370338 441586 370574
rect 441822 370338 441854 370574
rect 441234 334894 441854 370338
rect 441234 334658 441266 334894
rect 441502 334658 441586 334894
rect 441822 334658 441854 334894
rect 441234 334574 441854 334658
rect 441234 334338 441266 334574
rect 441502 334338 441586 334574
rect 441822 334338 441854 334574
rect 441234 298894 441854 334338
rect 444054 321469 444114 421907
rect 444051 321468 444117 321469
rect 444051 321404 444052 321468
rect 444116 321404 444117 321468
rect 444051 321403 444117 321404
rect 444238 319837 444298 689283
rect 444954 662614 445574 698058
rect 446259 686492 446325 686493
rect 446259 686428 446260 686492
rect 446324 686428 446325 686492
rect 446259 686427 446325 686428
rect 444954 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 445574 662614
rect 444954 662294 445574 662378
rect 444954 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 445574 662294
rect 444954 626614 445574 662058
rect 444954 626378 444986 626614
rect 445222 626378 445306 626614
rect 445542 626378 445574 626614
rect 444954 626294 445574 626378
rect 444954 626058 444986 626294
rect 445222 626058 445306 626294
rect 445542 626058 445574 626294
rect 444954 590614 445574 626058
rect 444954 590378 444986 590614
rect 445222 590378 445306 590614
rect 445542 590378 445574 590614
rect 444954 590294 445574 590378
rect 444954 590058 444986 590294
rect 445222 590058 445306 590294
rect 445542 590058 445574 590294
rect 444954 554614 445574 590058
rect 444954 554378 444986 554614
rect 445222 554378 445306 554614
rect 445542 554378 445574 554614
rect 444954 554294 445574 554378
rect 444954 554058 444986 554294
rect 445222 554058 445306 554294
rect 445542 554058 445574 554294
rect 444954 518614 445574 554058
rect 444954 518378 444986 518614
rect 445222 518378 445306 518614
rect 445542 518378 445574 518614
rect 444954 518294 445574 518378
rect 444954 518058 444986 518294
rect 445222 518058 445306 518294
rect 445542 518058 445574 518294
rect 444954 482614 445574 518058
rect 444954 482378 444986 482614
rect 445222 482378 445306 482614
rect 445542 482378 445574 482614
rect 444954 482294 445574 482378
rect 444954 482058 444986 482294
rect 445222 482058 445306 482294
rect 445542 482058 445574 482294
rect 444954 446614 445574 482058
rect 444954 446378 444986 446614
rect 445222 446378 445306 446614
rect 445542 446378 445574 446614
rect 444954 446294 445574 446378
rect 444954 446058 444986 446294
rect 445222 446058 445306 446294
rect 445542 446058 445574 446294
rect 444954 410614 445574 446058
rect 444954 410378 444986 410614
rect 445222 410378 445306 410614
rect 445542 410378 445574 410614
rect 444954 410294 445574 410378
rect 444954 410058 444986 410294
rect 445222 410058 445306 410294
rect 445542 410058 445574 410294
rect 444954 374614 445574 410058
rect 444954 374378 444986 374614
rect 445222 374378 445306 374614
rect 445542 374378 445574 374614
rect 444954 374294 445574 374378
rect 444954 374058 444986 374294
rect 445222 374058 445306 374294
rect 445542 374058 445574 374294
rect 444954 338614 445574 374058
rect 444954 338378 444986 338614
rect 445222 338378 445306 338614
rect 445542 338378 445574 338614
rect 444954 338294 445574 338378
rect 444954 338058 444986 338294
rect 445222 338058 445306 338294
rect 445542 338058 445574 338294
rect 444235 319836 444301 319837
rect 444235 319772 444236 319836
rect 444300 319772 444301 319836
rect 444235 319771 444301 319772
rect 441234 298658 441266 298894
rect 441502 298658 441586 298894
rect 441822 298658 441854 298894
rect 441234 298574 441854 298658
rect 441234 298338 441266 298574
rect 441502 298338 441586 298574
rect 441822 298338 441854 298574
rect 441234 262894 441854 298338
rect 441234 262658 441266 262894
rect 441502 262658 441586 262894
rect 441822 262658 441854 262894
rect 441234 262574 441854 262658
rect 441234 262338 441266 262574
rect 441502 262338 441586 262574
rect 441822 262338 441854 262574
rect 441234 226894 441854 262338
rect 441234 226658 441266 226894
rect 441502 226658 441586 226894
rect 441822 226658 441854 226894
rect 441234 226574 441854 226658
rect 441234 226338 441266 226574
rect 441502 226338 441586 226574
rect 441822 226338 441854 226574
rect 441234 190894 441854 226338
rect 441234 190658 441266 190894
rect 441502 190658 441586 190894
rect 441822 190658 441854 190894
rect 441234 190574 441854 190658
rect 441234 190338 441266 190574
rect 441502 190338 441586 190574
rect 441822 190338 441854 190574
rect 441234 157249 441854 190338
rect 444954 302614 445574 338058
rect 446262 319973 446322 686427
rect 447734 321333 447794 700299
rect 447918 322421 447978 700571
rect 448674 666334 449294 708122
rect 452394 709638 453014 711590
rect 452394 709402 452426 709638
rect 452662 709402 452746 709638
rect 452982 709402 453014 709638
rect 452394 709318 453014 709402
rect 452394 709082 452426 709318
rect 452662 709082 452746 709318
rect 452982 709082 453014 709318
rect 449571 700500 449637 700501
rect 449571 700436 449572 700500
rect 449636 700436 449637 700500
rect 449571 700435 449637 700436
rect 448674 666098 448706 666334
rect 448942 666098 449026 666334
rect 449262 666098 449294 666334
rect 448674 666014 449294 666098
rect 448674 665778 448706 666014
rect 448942 665778 449026 666014
rect 449262 665778 449294 666014
rect 448674 630334 449294 665778
rect 448674 630098 448706 630334
rect 448942 630098 449026 630334
rect 449262 630098 449294 630334
rect 448674 630014 449294 630098
rect 448674 629778 448706 630014
rect 448942 629778 449026 630014
rect 449262 629778 449294 630014
rect 448674 594334 449294 629778
rect 448674 594098 448706 594334
rect 448942 594098 449026 594334
rect 449262 594098 449294 594334
rect 448674 594014 449294 594098
rect 448674 593778 448706 594014
rect 448942 593778 449026 594014
rect 449262 593778 449294 594014
rect 448674 558334 449294 593778
rect 448674 558098 448706 558334
rect 448942 558098 449026 558334
rect 449262 558098 449294 558334
rect 448674 558014 449294 558098
rect 448674 557778 448706 558014
rect 448942 557778 449026 558014
rect 449262 557778 449294 558014
rect 448674 522334 449294 557778
rect 448674 522098 448706 522334
rect 448942 522098 449026 522334
rect 449262 522098 449294 522334
rect 448674 522014 449294 522098
rect 448674 521778 448706 522014
rect 448942 521778 449026 522014
rect 449262 521778 449294 522014
rect 448674 486334 449294 521778
rect 448674 486098 448706 486334
rect 448942 486098 449026 486334
rect 449262 486098 449294 486334
rect 448674 486014 449294 486098
rect 448674 485778 448706 486014
rect 448942 485778 449026 486014
rect 449262 485778 449294 486014
rect 448674 450334 449294 485778
rect 448674 450098 448706 450334
rect 448942 450098 449026 450334
rect 449262 450098 449294 450334
rect 448674 450014 449294 450098
rect 448674 449778 448706 450014
rect 448942 449778 449026 450014
rect 449262 449778 449294 450014
rect 448674 414334 449294 449778
rect 448674 414098 448706 414334
rect 448942 414098 449026 414334
rect 449262 414098 449294 414334
rect 448674 414014 449294 414098
rect 448674 413778 448706 414014
rect 448942 413778 449026 414014
rect 449262 413778 449294 414014
rect 448283 388380 448349 388381
rect 448283 388316 448284 388380
rect 448348 388316 448349 388380
rect 448283 388315 448349 388316
rect 448286 349213 448346 388315
rect 448674 378334 449294 413778
rect 448674 378098 448706 378334
rect 448942 378098 449026 378334
rect 449262 378098 449294 378334
rect 448674 378014 449294 378098
rect 448674 377778 448706 378014
rect 448942 377778 449026 378014
rect 449262 377778 449294 378014
rect 448283 349212 448349 349213
rect 448283 349148 448284 349212
rect 448348 349148 448349 349212
rect 448283 349147 448349 349148
rect 448674 342334 449294 377778
rect 448674 342098 448706 342334
rect 448942 342098 449026 342334
rect 449262 342098 449294 342334
rect 448674 342014 449294 342098
rect 448674 341778 448706 342014
rect 448942 341778 449026 342014
rect 449262 341778 449294 342014
rect 447915 322420 447981 322421
rect 447915 322356 447916 322420
rect 447980 322356 447981 322420
rect 447915 322355 447981 322356
rect 447731 321332 447797 321333
rect 447731 321268 447732 321332
rect 447796 321268 447797 321332
rect 447731 321267 447797 321268
rect 446259 319972 446325 319973
rect 446259 319908 446260 319972
rect 446324 319908 446325 319972
rect 446259 319907 446325 319908
rect 444954 302378 444986 302614
rect 445222 302378 445306 302614
rect 445542 302378 445574 302614
rect 444954 302294 445574 302378
rect 444954 302058 444986 302294
rect 445222 302058 445306 302294
rect 445542 302058 445574 302294
rect 444954 266614 445574 302058
rect 444954 266378 444986 266614
rect 445222 266378 445306 266614
rect 445542 266378 445574 266614
rect 444954 266294 445574 266378
rect 444954 266058 444986 266294
rect 445222 266058 445306 266294
rect 445542 266058 445574 266294
rect 444954 230614 445574 266058
rect 444954 230378 444986 230614
rect 445222 230378 445306 230614
rect 445542 230378 445574 230614
rect 444954 230294 445574 230378
rect 444954 230058 444986 230294
rect 445222 230058 445306 230294
rect 445542 230058 445574 230294
rect 444954 194614 445574 230058
rect 444954 194378 444986 194614
rect 445222 194378 445306 194614
rect 445542 194378 445574 194614
rect 444954 194294 445574 194378
rect 444954 194058 444986 194294
rect 445222 194058 445306 194294
rect 445542 194058 445574 194294
rect 444954 159644 445574 194058
rect 448674 306334 449294 341778
rect 449574 321061 449634 700435
rect 452394 670054 453014 709082
rect 452394 669818 452426 670054
rect 452662 669818 452746 670054
rect 452982 669818 453014 670054
rect 452394 669734 453014 669818
rect 452394 669498 452426 669734
rect 452662 669498 452746 669734
rect 452982 669498 453014 669734
rect 452394 634054 453014 669498
rect 452394 633818 452426 634054
rect 452662 633818 452746 634054
rect 452982 633818 453014 634054
rect 452394 633734 453014 633818
rect 452394 633498 452426 633734
rect 452662 633498 452746 633734
rect 452982 633498 453014 633734
rect 452394 598054 453014 633498
rect 452394 597818 452426 598054
rect 452662 597818 452746 598054
rect 452982 597818 453014 598054
rect 452394 597734 453014 597818
rect 452394 597498 452426 597734
rect 452662 597498 452746 597734
rect 452982 597498 453014 597734
rect 452394 562054 453014 597498
rect 452394 561818 452426 562054
rect 452662 561818 452746 562054
rect 452982 561818 453014 562054
rect 452394 561734 453014 561818
rect 452394 561498 452426 561734
rect 452662 561498 452746 561734
rect 452982 561498 453014 561734
rect 452394 526054 453014 561498
rect 452394 525818 452426 526054
rect 452662 525818 452746 526054
rect 452982 525818 453014 526054
rect 452394 525734 453014 525818
rect 452394 525498 452426 525734
rect 452662 525498 452746 525734
rect 452982 525498 453014 525734
rect 452394 517884 453014 525498
rect 456114 710598 456734 711590
rect 456114 710362 456146 710598
rect 456382 710362 456466 710598
rect 456702 710362 456734 710598
rect 456114 710278 456734 710362
rect 456114 710042 456146 710278
rect 456382 710042 456466 710278
rect 456702 710042 456734 710278
rect 456114 673774 456734 710042
rect 456114 673538 456146 673774
rect 456382 673538 456466 673774
rect 456702 673538 456734 673774
rect 456114 673454 456734 673538
rect 456114 673218 456146 673454
rect 456382 673218 456466 673454
rect 456702 673218 456734 673454
rect 456114 637774 456734 673218
rect 459834 711558 460454 711590
rect 459834 711322 459866 711558
rect 460102 711322 460186 711558
rect 460422 711322 460454 711558
rect 459834 711238 460454 711322
rect 459834 711002 459866 711238
rect 460102 711002 460186 711238
rect 460422 711002 460454 711238
rect 459834 677494 460454 711002
rect 459834 677258 459866 677494
rect 460102 677258 460186 677494
rect 460422 677258 460454 677494
rect 459834 677174 460454 677258
rect 459834 676938 459866 677174
rect 460102 676938 460186 677174
rect 460422 676938 460454 677174
rect 459834 669073 460454 676938
rect 469794 704838 470414 711590
rect 469794 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 470414 704838
rect 469794 704518 470414 704602
rect 469794 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 470414 704518
rect 469794 687454 470414 704282
rect 469794 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 470414 687454
rect 469794 687134 470414 687218
rect 469794 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 470414 687134
rect 469794 669073 470414 686898
rect 473514 705798 474134 711590
rect 473514 705562 473546 705798
rect 473782 705562 473866 705798
rect 474102 705562 474134 705798
rect 473514 705478 474134 705562
rect 473514 705242 473546 705478
rect 473782 705242 473866 705478
rect 474102 705242 474134 705478
rect 473514 691174 474134 705242
rect 473514 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 474134 691174
rect 473514 690854 474134 690938
rect 473514 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 474134 690854
rect 473514 669073 474134 690618
rect 477234 706758 477854 711590
rect 477234 706522 477266 706758
rect 477502 706522 477586 706758
rect 477822 706522 477854 706758
rect 477234 706438 477854 706522
rect 477234 706202 477266 706438
rect 477502 706202 477586 706438
rect 477822 706202 477854 706438
rect 477234 694894 477854 706202
rect 477234 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 477854 694894
rect 477234 694574 477854 694658
rect 477234 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 477854 694574
rect 477234 669073 477854 694338
rect 480954 707718 481574 711590
rect 480954 707482 480986 707718
rect 481222 707482 481306 707718
rect 481542 707482 481574 707718
rect 480954 707398 481574 707482
rect 480954 707162 480986 707398
rect 481222 707162 481306 707398
rect 481542 707162 481574 707398
rect 480954 698614 481574 707162
rect 480954 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 481574 698614
rect 480954 698294 481574 698378
rect 480954 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 481574 698294
rect 480954 669073 481574 698058
rect 488394 709638 489014 711590
rect 488394 709402 488426 709638
rect 488662 709402 488746 709638
rect 488982 709402 489014 709638
rect 488394 709318 489014 709402
rect 488394 709082 488426 709318
rect 488662 709082 488746 709318
rect 488982 709082 489014 709318
rect 488394 670054 489014 709082
rect 488394 669818 488426 670054
rect 488662 669818 488746 670054
rect 488982 669818 489014 670054
rect 488394 669734 489014 669818
rect 488394 669498 488426 669734
rect 488662 669498 488746 669734
rect 488982 669498 489014 669734
rect 488394 669073 489014 669498
rect 492114 710598 492734 711590
rect 492114 710362 492146 710598
rect 492382 710362 492466 710598
rect 492702 710362 492734 710598
rect 492114 710278 492734 710362
rect 492114 710042 492146 710278
rect 492382 710042 492466 710278
rect 492702 710042 492734 710278
rect 492114 673774 492734 710042
rect 492114 673538 492146 673774
rect 492382 673538 492466 673774
rect 492702 673538 492734 673774
rect 492114 673454 492734 673538
rect 492114 673218 492146 673454
rect 492382 673218 492466 673454
rect 492702 673218 492734 673454
rect 492114 669073 492734 673218
rect 495834 711558 496454 711590
rect 495834 711322 495866 711558
rect 496102 711322 496186 711558
rect 496422 711322 496454 711558
rect 495834 711238 496454 711322
rect 495834 711002 495866 711238
rect 496102 711002 496186 711238
rect 496422 711002 496454 711238
rect 495834 677494 496454 711002
rect 495834 677258 495866 677494
rect 496102 677258 496186 677494
rect 496422 677258 496454 677494
rect 495834 677174 496454 677258
rect 495834 676938 495866 677174
rect 496102 676938 496186 677174
rect 496422 676938 496454 677174
rect 495834 669073 496454 676938
rect 505794 704838 506414 711590
rect 505794 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 506414 704838
rect 505794 704518 506414 704602
rect 505794 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 506414 704518
rect 505794 687454 506414 704282
rect 505794 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 506414 687454
rect 505794 687134 506414 687218
rect 505794 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 506414 687134
rect 505794 669073 506414 686898
rect 509514 705798 510134 711590
rect 509514 705562 509546 705798
rect 509782 705562 509866 705798
rect 510102 705562 510134 705798
rect 509514 705478 510134 705562
rect 509514 705242 509546 705478
rect 509782 705242 509866 705478
rect 510102 705242 510134 705478
rect 509514 691174 510134 705242
rect 509514 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 510134 691174
rect 509514 690854 510134 690938
rect 509514 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 510134 690854
rect 509514 669073 510134 690618
rect 513234 706758 513854 711590
rect 513234 706522 513266 706758
rect 513502 706522 513586 706758
rect 513822 706522 513854 706758
rect 513234 706438 513854 706522
rect 513234 706202 513266 706438
rect 513502 706202 513586 706438
rect 513822 706202 513854 706438
rect 513234 694894 513854 706202
rect 513234 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 513854 694894
rect 513234 694574 513854 694658
rect 513234 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 513854 694574
rect 513234 669073 513854 694338
rect 516954 707718 517574 711590
rect 516954 707482 516986 707718
rect 517222 707482 517306 707718
rect 517542 707482 517574 707718
rect 516954 707398 517574 707482
rect 516954 707162 516986 707398
rect 517222 707162 517306 707398
rect 517542 707162 517574 707398
rect 516954 698614 517574 707162
rect 516954 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 517574 698614
rect 516954 698294 517574 698378
rect 516954 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 517574 698294
rect 516954 669073 517574 698058
rect 520674 708678 521294 711590
rect 520674 708442 520706 708678
rect 520942 708442 521026 708678
rect 521262 708442 521294 708678
rect 520674 708358 521294 708442
rect 520674 708122 520706 708358
rect 520942 708122 521026 708358
rect 521262 708122 521294 708358
rect 520674 666334 521294 708122
rect 520674 666098 520706 666334
rect 520942 666098 521026 666334
rect 521262 666098 521294 666334
rect 520674 666014 521294 666098
rect 520674 665778 520706 666014
rect 520942 665778 521026 666014
rect 521262 665778 521294 666014
rect 457851 665276 457917 665277
rect 457851 665212 457852 665276
rect 457916 665212 457917 665276
rect 457851 665211 457917 665212
rect 456114 637538 456146 637774
rect 456382 637538 456466 637774
rect 456702 637538 456734 637774
rect 456114 637454 456734 637538
rect 456114 637218 456146 637454
rect 456382 637218 456466 637454
rect 456702 637218 456734 637454
rect 456114 601774 456734 637218
rect 456114 601538 456146 601774
rect 456382 601538 456466 601774
rect 456702 601538 456734 601774
rect 456114 601454 456734 601538
rect 456114 601218 456146 601454
rect 456382 601218 456466 601454
rect 456702 601218 456734 601454
rect 456114 565774 456734 601218
rect 457854 597685 457914 665211
rect 458035 662556 458101 662557
rect 458035 662492 458036 662556
rect 458100 662492 458101 662556
rect 458035 662491 458101 662492
rect 457851 597684 457917 597685
rect 457851 597620 457852 597684
rect 457916 597620 457917 597684
rect 457851 597619 457917 597620
rect 456114 565538 456146 565774
rect 456382 565538 456466 565774
rect 456702 565538 456734 565774
rect 456114 565454 456734 565538
rect 456114 565218 456146 565454
rect 456382 565218 456466 565454
rect 456702 565218 456734 565454
rect 456114 529774 456734 565218
rect 456114 529538 456146 529774
rect 456382 529538 456466 529774
rect 456702 529538 456734 529774
rect 456114 529454 456734 529538
rect 456114 529218 456146 529454
rect 456382 529218 456466 529454
rect 456702 529218 456734 529454
rect 456114 517884 456734 529218
rect 458038 518125 458098 662491
rect 459507 655688 459573 655689
rect 459507 655624 459508 655688
rect 459572 655624 459573 655688
rect 459507 655623 459573 655624
rect 459510 595509 459570 655623
rect 479568 655174 479888 655206
rect 479568 654938 479610 655174
rect 479846 654938 479888 655174
rect 479568 654854 479888 654938
rect 479568 654618 479610 654854
rect 479846 654618 479888 654854
rect 479568 654586 479888 654618
rect 510288 655174 510608 655206
rect 510288 654938 510330 655174
rect 510566 654938 510608 655174
rect 510288 654854 510608 654938
rect 510288 654618 510330 654854
rect 510566 654618 510608 654854
rect 510288 654586 510608 654618
rect 464208 651454 464528 651486
rect 464208 651218 464250 651454
rect 464486 651218 464528 651454
rect 464208 651134 464528 651218
rect 464208 650898 464250 651134
rect 464486 650898 464528 651134
rect 464208 650866 464528 650898
rect 494928 651454 495248 651486
rect 494928 651218 494970 651454
rect 495206 651218 495248 651454
rect 494928 651134 495248 651218
rect 494928 650898 494970 651134
rect 495206 650898 495248 651134
rect 494928 650866 495248 650898
rect 520674 630334 521294 665778
rect 520674 630098 520706 630334
rect 520942 630098 521026 630334
rect 521262 630098 521294 630334
rect 520674 630014 521294 630098
rect 520674 629778 520706 630014
rect 520942 629778 521026 630014
rect 521262 629778 521294 630014
rect 479568 619174 479888 619206
rect 479568 618938 479610 619174
rect 479846 618938 479888 619174
rect 479568 618854 479888 618938
rect 479568 618618 479610 618854
rect 479846 618618 479888 618854
rect 479568 618586 479888 618618
rect 510288 619174 510608 619206
rect 510288 618938 510330 619174
rect 510566 618938 510608 619174
rect 510288 618854 510608 618938
rect 510288 618618 510330 618854
rect 510566 618618 510608 618854
rect 510288 618586 510608 618618
rect 464208 615454 464528 615486
rect 464208 615218 464250 615454
rect 464486 615218 464528 615454
rect 464208 615134 464528 615218
rect 464208 614898 464250 615134
rect 464486 614898 464528 615134
rect 464208 614866 464528 614898
rect 494928 615454 495248 615486
rect 494928 615218 494970 615454
rect 495206 615218 495248 615454
rect 494928 615134 495248 615218
rect 494928 614898 494970 615134
rect 495206 614898 495248 615134
rect 494928 614866 495248 614898
rect 459507 595508 459573 595509
rect 459507 595444 459508 595508
rect 459572 595444 459573 595508
rect 459507 595443 459573 595444
rect 459834 569494 460454 601103
rect 459834 569258 459866 569494
rect 460102 569258 460186 569494
rect 460422 569258 460454 569494
rect 459834 569174 460454 569258
rect 459834 568938 459866 569174
rect 460102 568938 460186 569174
rect 460422 568938 460454 569174
rect 459834 533494 460454 568938
rect 459834 533258 459866 533494
rect 460102 533258 460186 533494
rect 460422 533258 460454 533494
rect 459834 533174 460454 533258
rect 459834 532938 459866 533174
rect 460102 532938 460186 533174
rect 460422 532938 460454 533174
rect 458035 518124 458101 518125
rect 458035 518060 458036 518124
rect 458100 518060 458101 518124
rect 458035 518059 458101 518060
rect 459834 517884 460454 532938
rect 469794 579454 470414 601103
rect 472019 598228 472085 598229
rect 472019 598164 472020 598228
rect 472084 598164 472085 598228
rect 472019 598163 472085 598164
rect 469794 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 470414 579454
rect 469794 579134 470414 579218
rect 469794 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 470414 579134
rect 469794 543454 470414 578898
rect 469794 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 470414 543454
rect 469794 543134 470414 543218
rect 469794 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 470414 543134
rect 451043 516764 451109 516765
rect 451043 516700 451044 516764
rect 451108 516700 451109 516764
rect 451043 516699 451109 516700
rect 450491 514384 450557 514385
rect 450491 514320 450492 514384
rect 450556 514320 450557 514384
rect 450491 514319 450557 514320
rect 450494 328405 450554 514319
rect 451046 335370 451106 516699
rect 453382 511174 453702 511206
rect 453382 510938 453424 511174
rect 453660 510938 453702 511174
rect 453382 510854 453702 510938
rect 453382 510618 453424 510854
rect 453660 510618 453702 510854
rect 453382 510586 453702 510618
rect 455820 511174 456140 511206
rect 455820 510938 455862 511174
rect 456098 510938 456140 511174
rect 455820 510854 456140 510938
rect 455820 510618 455862 510854
rect 456098 510618 456140 510854
rect 455820 510586 456140 510618
rect 458258 511174 458578 511206
rect 458258 510938 458300 511174
rect 458536 510938 458578 511174
rect 458258 510854 458578 510938
rect 458258 510618 458300 510854
rect 458536 510618 458578 510854
rect 458258 510586 458578 510618
rect 460696 511174 461016 511206
rect 460696 510938 460738 511174
rect 460974 510938 461016 511174
rect 460696 510854 461016 510938
rect 460696 510618 460738 510854
rect 460974 510618 461016 510854
rect 460696 510586 461016 510618
rect 452163 507454 452483 507486
rect 452163 507218 452205 507454
rect 452441 507218 452483 507454
rect 452163 507134 452483 507218
rect 452163 506898 452205 507134
rect 452441 506898 452483 507134
rect 452163 506866 452483 506898
rect 454601 507454 454921 507486
rect 454601 507218 454643 507454
rect 454879 507218 454921 507454
rect 454601 507134 454921 507218
rect 454601 506898 454643 507134
rect 454879 506898 454921 507134
rect 454601 506866 454921 506898
rect 457039 507454 457359 507486
rect 457039 507218 457081 507454
rect 457317 507218 457359 507454
rect 457039 507134 457359 507218
rect 457039 506898 457081 507134
rect 457317 506898 457359 507134
rect 457039 506866 457359 506898
rect 459477 507454 459797 507486
rect 459477 507218 459519 507454
rect 459755 507218 459797 507454
rect 459477 507134 459797 507218
rect 459477 506898 459519 507134
rect 459755 506898 459797 507134
rect 459477 506866 459797 506898
rect 469794 507454 470414 542898
rect 469794 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 470414 507454
rect 469794 507134 470414 507218
rect 469794 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 470414 507134
rect 450678 335310 451106 335370
rect 452394 490054 453014 500068
rect 452394 489818 452426 490054
rect 452662 489818 452746 490054
rect 452982 489818 453014 490054
rect 452394 489734 453014 489818
rect 452394 489498 452426 489734
rect 452662 489498 452746 489734
rect 452982 489498 453014 489734
rect 452394 454054 453014 489498
rect 452394 453818 452426 454054
rect 452662 453818 452746 454054
rect 452982 453818 453014 454054
rect 452394 453734 453014 453818
rect 452394 453498 452426 453734
rect 452662 453498 452746 453734
rect 452982 453498 453014 453734
rect 452394 418054 453014 453498
rect 452394 417818 452426 418054
rect 452662 417818 452746 418054
rect 452982 417818 453014 418054
rect 452394 417734 453014 417818
rect 452394 417498 452426 417734
rect 452662 417498 452746 417734
rect 452982 417498 453014 417734
rect 452394 382054 453014 417498
rect 452394 381818 452426 382054
rect 452662 381818 452746 382054
rect 452982 381818 453014 382054
rect 452394 381734 453014 381818
rect 452394 381498 452426 381734
rect 452662 381498 452746 381734
rect 452982 381498 453014 381734
rect 452394 346054 453014 381498
rect 456114 493774 456734 500068
rect 456114 493538 456146 493774
rect 456382 493538 456466 493774
rect 456702 493538 456734 493774
rect 456114 493454 456734 493538
rect 456114 493218 456146 493454
rect 456382 493218 456466 493454
rect 456702 493218 456734 493454
rect 456114 457774 456734 493218
rect 456114 457538 456146 457774
rect 456382 457538 456466 457774
rect 456702 457538 456734 457774
rect 456114 457454 456734 457538
rect 456114 457218 456146 457454
rect 456382 457218 456466 457454
rect 456702 457218 456734 457454
rect 456114 421774 456734 457218
rect 456114 421538 456146 421774
rect 456382 421538 456466 421774
rect 456702 421538 456734 421774
rect 456114 421454 456734 421538
rect 456114 421218 456146 421454
rect 456382 421218 456466 421454
rect 456702 421218 456734 421454
rect 456114 385774 456734 421218
rect 456114 385538 456146 385774
rect 456382 385538 456466 385774
rect 456702 385538 456734 385774
rect 456114 385454 456734 385538
rect 456114 385218 456146 385454
rect 456382 385218 456466 385454
rect 456702 385218 456734 385454
rect 454208 363454 454528 363486
rect 454208 363218 454250 363454
rect 454486 363218 454528 363454
rect 454208 363134 454528 363218
rect 454208 362898 454250 363134
rect 454486 362898 454528 363134
rect 454208 362866 454528 362898
rect 452394 345818 452426 346054
rect 452662 345818 452746 346054
rect 452982 345818 453014 346054
rect 452394 345734 453014 345818
rect 452394 345498 452426 345734
rect 452662 345498 452746 345734
rect 452982 345498 453014 345734
rect 450678 328813 450738 335310
rect 450675 328812 450741 328813
rect 450675 328748 450676 328812
rect 450740 328748 450741 328812
rect 450675 328747 450741 328748
rect 450491 328404 450557 328405
rect 450491 328340 450492 328404
rect 450556 328340 450557 328404
rect 450491 328339 450557 328340
rect 449571 321060 449637 321061
rect 449571 320996 449572 321060
rect 449636 320996 449637 321060
rect 449571 320995 449637 320996
rect 448674 306098 448706 306334
rect 448942 306098 449026 306334
rect 449262 306098 449294 306334
rect 448674 306014 449294 306098
rect 448674 305778 448706 306014
rect 448942 305778 449026 306014
rect 449262 305778 449294 306014
rect 448674 270334 449294 305778
rect 448674 270098 448706 270334
rect 448942 270098 449026 270334
rect 449262 270098 449294 270334
rect 448674 270014 449294 270098
rect 448674 269778 448706 270014
rect 448942 269778 449026 270014
rect 449262 269778 449294 270014
rect 448674 234334 449294 269778
rect 448674 234098 448706 234334
rect 448942 234098 449026 234334
rect 449262 234098 449294 234334
rect 448674 234014 449294 234098
rect 448674 233778 448706 234014
rect 448942 233778 449026 234014
rect 449262 233778 449294 234014
rect 448674 198334 449294 233778
rect 448674 198098 448706 198334
rect 448942 198098 449026 198334
rect 449262 198098 449294 198334
rect 448674 198014 449294 198098
rect 448674 197778 448706 198014
rect 448942 197778 449026 198014
rect 449262 197778 449294 198014
rect 448674 162334 449294 197778
rect 448674 162098 448706 162334
rect 448942 162098 449026 162334
rect 449262 162098 449294 162334
rect 448674 162014 449294 162098
rect 448674 161778 448706 162014
rect 448942 161778 449026 162014
rect 449262 161778 449294 162014
rect 429568 151174 429888 151206
rect 429568 150938 429610 151174
rect 429846 150938 429888 151174
rect 429568 150854 429888 150938
rect 429568 150618 429610 150854
rect 429846 150618 429888 150854
rect 429568 150586 429888 150618
rect 414208 147454 414528 147486
rect 414208 147218 414250 147454
rect 414486 147218 414528 147454
rect 414208 147134 414528 147218
rect 414208 146898 414250 147134
rect 414486 146898 414528 147134
rect 414208 146866 414528 146898
rect 444928 147454 445248 147486
rect 444928 147218 444970 147454
rect 445206 147218 445248 147454
rect 444928 147134 445248 147218
rect 444928 146898 444970 147134
rect 445206 146898 445248 147134
rect 444928 146866 445248 146898
rect 412674 126098 412706 126334
rect 412942 126098 413026 126334
rect 413262 126098 413294 126334
rect 412674 126014 413294 126098
rect 412674 125778 412706 126014
rect 412942 125778 413026 126014
rect 413262 125778 413294 126014
rect 412674 92137 413294 125778
rect 416394 94054 417014 127767
rect 416394 93818 416426 94054
rect 416662 93818 416746 94054
rect 416982 93818 417014 94054
rect 416394 93734 417014 93818
rect 416394 93498 416426 93734
rect 416662 93498 416746 93734
rect 416982 93498 417014 93734
rect 416394 92137 417014 93498
rect 420114 97774 420734 127767
rect 420114 97538 420146 97774
rect 420382 97538 420466 97774
rect 420702 97538 420734 97774
rect 420114 97454 420734 97538
rect 420114 97218 420146 97454
rect 420382 97218 420466 97454
rect 420702 97218 420734 97454
rect 420114 92137 420734 97218
rect 423834 101494 424454 127767
rect 423834 101258 423866 101494
rect 424102 101258 424186 101494
rect 424422 101258 424454 101494
rect 423834 101174 424454 101258
rect 423834 100938 423866 101174
rect 424102 100938 424186 101174
rect 424422 100938 424454 101174
rect 423834 92137 424454 100938
rect 448674 126334 449294 161778
rect 448674 126098 448706 126334
rect 448942 126098 449026 126334
rect 449262 126098 449294 126334
rect 448674 126014 449294 126098
rect 448674 125778 448706 126014
rect 448942 125778 449026 126014
rect 449262 125778 449294 126014
rect 448674 92137 449294 125778
rect 452394 310054 453014 345498
rect 456114 349774 456734 385218
rect 456114 349538 456146 349774
rect 456382 349538 456466 349774
rect 456702 349538 456734 349774
rect 456114 349454 456734 349538
rect 456114 349218 456146 349454
rect 456382 349218 456466 349454
rect 456702 349218 456734 349454
rect 454208 327454 454528 327486
rect 454208 327218 454250 327454
rect 454486 327218 454528 327454
rect 454208 327134 454528 327218
rect 454208 326898 454250 327134
rect 454486 326898 454528 327134
rect 454208 326866 454528 326898
rect 452394 309818 452426 310054
rect 452662 309818 452746 310054
rect 452982 309818 453014 310054
rect 452394 309734 453014 309818
rect 452394 309498 452426 309734
rect 452662 309498 452746 309734
rect 452982 309498 453014 309734
rect 452394 274054 453014 309498
rect 452394 273818 452426 274054
rect 452662 273818 452746 274054
rect 452982 273818 453014 274054
rect 452394 273734 453014 273818
rect 452394 273498 452426 273734
rect 452662 273498 452746 273734
rect 452982 273498 453014 273734
rect 452394 238054 453014 273498
rect 452394 237818 452426 238054
rect 452662 237818 452746 238054
rect 452982 237818 453014 238054
rect 452394 237734 453014 237818
rect 452394 237498 452426 237734
rect 452662 237498 452746 237734
rect 452982 237498 453014 237734
rect 452394 202054 453014 237498
rect 452394 201818 452426 202054
rect 452662 201818 452746 202054
rect 452982 201818 453014 202054
rect 452394 201734 453014 201818
rect 452394 201498 452426 201734
rect 452662 201498 452746 201734
rect 452982 201498 453014 201734
rect 452394 166054 453014 201498
rect 452394 165818 452426 166054
rect 452662 165818 452746 166054
rect 452982 165818 453014 166054
rect 452394 165734 453014 165818
rect 452394 165498 452426 165734
rect 452662 165498 452746 165734
rect 452982 165498 453014 165734
rect 452394 130054 453014 165498
rect 452394 129818 452426 130054
rect 452662 129818 452746 130054
rect 452982 129818 453014 130054
rect 452394 129734 453014 129818
rect 452394 129498 452426 129734
rect 452662 129498 452746 129734
rect 452982 129498 453014 129734
rect 452394 94054 453014 129498
rect 452394 93818 452426 94054
rect 452662 93818 452746 94054
rect 452982 93818 453014 94054
rect 452394 93734 453014 93818
rect 452394 93498 452426 93734
rect 452662 93498 452746 93734
rect 452982 93498 453014 93734
rect 452394 92137 453014 93498
rect 456114 313774 456734 349218
rect 456114 313538 456146 313774
rect 456382 313538 456466 313774
rect 456702 313538 456734 313774
rect 456114 313454 456734 313538
rect 456114 313218 456146 313454
rect 456382 313218 456466 313454
rect 456702 313218 456734 313454
rect 456114 277774 456734 313218
rect 456114 277538 456146 277774
rect 456382 277538 456466 277774
rect 456702 277538 456734 277774
rect 456114 277454 456734 277538
rect 456114 277218 456146 277454
rect 456382 277218 456466 277454
rect 456702 277218 456734 277454
rect 456114 241774 456734 277218
rect 456114 241538 456146 241774
rect 456382 241538 456466 241774
rect 456702 241538 456734 241774
rect 456114 241454 456734 241538
rect 456114 241218 456146 241454
rect 456382 241218 456466 241454
rect 456702 241218 456734 241454
rect 456114 205774 456734 241218
rect 456114 205538 456146 205774
rect 456382 205538 456466 205774
rect 456702 205538 456734 205774
rect 456114 205454 456734 205538
rect 456114 205218 456146 205454
rect 456382 205218 456466 205454
rect 456702 205218 456734 205454
rect 456114 169774 456734 205218
rect 456114 169538 456146 169774
rect 456382 169538 456466 169774
rect 456702 169538 456734 169774
rect 456114 169454 456734 169538
rect 456114 169218 456146 169454
rect 456382 169218 456466 169454
rect 456702 169218 456734 169454
rect 456114 133774 456734 169218
rect 456114 133538 456146 133774
rect 456382 133538 456466 133774
rect 456702 133538 456734 133774
rect 456114 133454 456734 133538
rect 456114 133218 456146 133454
rect 456382 133218 456466 133454
rect 456702 133218 456734 133454
rect 456114 97774 456734 133218
rect 456114 97538 456146 97774
rect 456382 97538 456466 97774
rect 456702 97538 456734 97774
rect 456114 97454 456734 97538
rect 456114 97218 456146 97454
rect 456382 97218 456466 97454
rect 456702 97218 456734 97454
rect 456114 92137 456734 97218
rect 459834 497494 460454 500068
rect 459834 497258 459866 497494
rect 460102 497258 460186 497494
rect 460422 497258 460454 497494
rect 459834 497174 460454 497258
rect 459834 496938 459866 497174
rect 460102 496938 460186 497174
rect 460422 496938 460454 497174
rect 459834 461494 460454 496938
rect 459834 461258 459866 461494
rect 460102 461258 460186 461494
rect 460422 461258 460454 461494
rect 459834 461174 460454 461258
rect 459834 460938 459866 461174
rect 460102 460938 460186 461174
rect 460422 460938 460454 461174
rect 459834 425494 460454 460938
rect 459834 425258 459866 425494
rect 460102 425258 460186 425494
rect 460422 425258 460454 425494
rect 459834 425174 460454 425258
rect 459834 424938 459866 425174
rect 460102 424938 460186 425174
rect 460422 424938 460454 425174
rect 459834 389494 460454 424938
rect 459834 389258 459866 389494
rect 460102 389258 460186 389494
rect 460422 389258 460454 389494
rect 459834 389174 460454 389258
rect 459834 388938 459866 389174
rect 460102 388938 460186 389174
rect 460422 388938 460454 389174
rect 459834 353494 460454 388938
rect 469794 471454 470414 506898
rect 469794 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 470414 471454
rect 469794 471134 470414 471218
rect 469794 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 470414 471134
rect 469794 435454 470414 470898
rect 469794 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 470414 435454
rect 469794 435134 470414 435218
rect 469794 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 470414 435134
rect 469794 399454 470414 434898
rect 469794 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 470414 399454
rect 469794 399134 470414 399218
rect 469794 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 470414 399134
rect 469794 385580 470414 398898
rect 472022 388925 472082 598163
rect 472203 595644 472269 595645
rect 472203 595580 472204 595644
rect 472268 595580 472269 595644
rect 472203 595579 472269 595580
rect 472206 389061 472266 595579
rect 473514 583174 474134 601103
rect 474411 599588 474477 599589
rect 474411 599524 474412 599588
rect 474476 599524 474477 599588
rect 474411 599523 474477 599524
rect 473514 582938 473546 583174
rect 473782 582938 473866 583174
rect 474102 582938 474134 583174
rect 473514 582854 474134 582938
rect 473514 582618 473546 582854
rect 473782 582618 473866 582854
rect 474102 582618 474134 582854
rect 473514 547174 474134 582618
rect 473514 546938 473546 547174
rect 473782 546938 473866 547174
rect 474102 546938 474134 547174
rect 473514 546854 474134 546938
rect 473514 546618 473546 546854
rect 473782 546618 473866 546854
rect 474102 546618 474134 546854
rect 473514 511174 474134 546618
rect 473514 510938 473546 511174
rect 473782 510938 473866 511174
rect 474102 510938 474134 511174
rect 473514 510854 474134 510938
rect 473514 510618 473546 510854
rect 473782 510618 473866 510854
rect 474102 510618 474134 510854
rect 473514 475174 474134 510618
rect 473514 474938 473546 475174
rect 473782 474938 473866 475174
rect 474102 474938 474134 475174
rect 473514 474854 474134 474938
rect 473514 474618 473546 474854
rect 473782 474618 473866 474854
rect 474102 474618 474134 474854
rect 473514 453692 474134 474618
rect 473416 435454 473736 435486
rect 473416 435218 473458 435454
rect 473694 435218 473736 435454
rect 473416 435134 473736 435218
rect 473416 434898 473458 435134
rect 473694 434898 473736 435134
rect 473416 434866 473736 434898
rect 474414 389061 474474 599523
rect 476435 591292 476501 591293
rect 476435 591228 476436 591292
rect 476500 591228 476501 591292
rect 476435 591227 476501 591228
rect 474779 589932 474845 589933
rect 474779 589868 474780 589932
rect 474844 589868 474845 589932
rect 474779 589867 474845 589868
rect 474782 389061 474842 589867
rect 475888 439174 476208 439206
rect 475888 438938 475930 439174
rect 476166 438938 476208 439174
rect 475888 438854 476208 438938
rect 475888 438618 475930 438854
rect 476166 438618 476208 438854
rect 475888 438586 476208 438618
rect 476438 389061 476498 591227
rect 477234 586894 477854 601103
rect 478827 595508 478893 595509
rect 478827 595444 478828 595508
rect 478892 595444 478893 595508
rect 478827 595443 478893 595444
rect 477234 586658 477266 586894
rect 477502 586658 477586 586894
rect 477822 586658 477854 586894
rect 477234 586574 477854 586658
rect 477234 586338 477266 586574
rect 477502 586338 477586 586574
rect 477822 586338 477854 586574
rect 477234 550894 477854 586338
rect 477234 550658 477266 550894
rect 477502 550658 477586 550894
rect 477822 550658 477854 550894
rect 477234 550574 477854 550658
rect 477234 550338 477266 550574
rect 477502 550338 477586 550574
rect 477822 550338 477854 550574
rect 477234 514894 477854 550338
rect 477234 514658 477266 514894
rect 477502 514658 477586 514894
rect 477822 514658 477854 514894
rect 477234 514574 477854 514658
rect 477234 514338 477266 514574
rect 477502 514338 477586 514574
rect 477822 514338 477854 514574
rect 477234 478894 477854 514338
rect 477234 478658 477266 478894
rect 477502 478658 477586 478894
rect 477822 478658 477854 478894
rect 477234 478574 477854 478658
rect 477234 478338 477266 478574
rect 477502 478338 477586 478574
rect 477822 478338 477854 478574
rect 477234 442894 477854 478338
rect 477234 442658 477266 442894
rect 477502 442658 477586 442894
rect 477822 442658 477854 442894
rect 477234 442574 477854 442658
rect 477234 442338 477266 442574
rect 477502 442338 477586 442574
rect 477822 442338 477854 442574
rect 477234 406894 477854 442338
rect 478361 435454 478681 435486
rect 478361 435218 478403 435454
rect 478639 435218 478681 435454
rect 478361 435134 478681 435218
rect 478361 434898 478403 435134
rect 478639 434898 478681 435134
rect 478361 434866 478681 434898
rect 477234 406658 477266 406894
rect 477502 406658 477586 406894
rect 477822 406658 477854 406894
rect 477234 406574 477854 406658
rect 477234 406338 477266 406574
rect 477502 406338 477586 406574
rect 477822 406338 477854 406574
rect 472203 389060 472269 389061
rect 472203 388996 472204 389060
rect 472268 388996 472269 389060
rect 472203 388995 472269 388996
rect 474411 389060 474477 389061
rect 474411 388996 474412 389060
rect 474476 388996 474477 389060
rect 474411 388995 474477 388996
rect 474779 389060 474845 389061
rect 474779 388996 474780 389060
rect 474844 388996 474845 389060
rect 474779 388995 474845 388996
rect 476435 389060 476501 389061
rect 476435 388996 476436 389060
rect 476500 388996 476501 389060
rect 476435 388995 476501 388996
rect 472019 388924 472085 388925
rect 472019 388860 472020 388924
rect 472084 388860 472085 388924
rect 472019 388859 472085 388860
rect 477234 384817 477854 406338
rect 478830 389061 478890 595443
rect 480954 590614 481574 601103
rect 480954 590378 480986 590614
rect 481222 590378 481306 590614
rect 481542 590378 481574 590614
rect 480954 590294 481574 590378
rect 480954 590058 480986 590294
rect 481222 590058 481306 590294
rect 481542 590058 481574 590294
rect 480954 554614 481574 590058
rect 480954 554378 480986 554614
rect 481222 554378 481306 554614
rect 481542 554378 481574 554614
rect 480954 554294 481574 554378
rect 480954 554058 480986 554294
rect 481222 554058 481306 554294
rect 481542 554058 481574 554294
rect 480954 518614 481574 554058
rect 480954 518378 480986 518614
rect 481222 518378 481306 518614
rect 481542 518378 481574 518614
rect 480954 518294 481574 518378
rect 480954 518058 480986 518294
rect 481222 518058 481306 518294
rect 481542 518058 481574 518294
rect 480954 482614 481574 518058
rect 484674 594334 485294 601103
rect 484674 594098 484706 594334
rect 484942 594098 485026 594334
rect 485262 594098 485294 594334
rect 484674 594014 485294 594098
rect 484674 593778 484706 594014
rect 484942 593778 485026 594014
rect 485262 593778 485294 594014
rect 484674 558334 485294 593778
rect 484674 558098 484706 558334
rect 484942 558098 485026 558334
rect 485262 558098 485294 558334
rect 484674 558014 485294 558098
rect 484674 557778 484706 558014
rect 484942 557778 485026 558014
rect 485262 557778 485294 558014
rect 484674 522334 485294 557778
rect 484674 522098 484706 522334
rect 484942 522098 485026 522334
rect 485262 522098 485294 522334
rect 484674 522014 485294 522098
rect 484674 521778 484706 522014
rect 484942 521778 485026 522014
rect 485262 521778 485294 522014
rect 484674 517884 485294 521778
rect 488394 598054 489014 601103
rect 488394 597818 488426 598054
rect 488662 597818 488746 598054
rect 488982 597818 489014 598054
rect 488394 597734 489014 597818
rect 488394 597498 488426 597734
rect 488662 597498 488746 597734
rect 488982 597498 489014 597734
rect 488394 562054 489014 597498
rect 488394 561818 488426 562054
rect 488662 561818 488746 562054
rect 488982 561818 489014 562054
rect 488394 561734 489014 561818
rect 488394 561498 488426 561734
rect 488662 561498 488746 561734
rect 488982 561498 489014 561734
rect 488394 526054 489014 561498
rect 488394 525818 488426 526054
rect 488662 525818 488746 526054
rect 488982 525818 489014 526054
rect 488394 525734 489014 525818
rect 488394 525498 488426 525734
rect 488662 525498 488746 525734
rect 488982 525498 489014 525734
rect 488394 517884 489014 525498
rect 492114 565774 492734 601103
rect 492114 565538 492146 565774
rect 492382 565538 492466 565774
rect 492702 565538 492734 565774
rect 492114 565454 492734 565538
rect 492114 565218 492146 565454
rect 492382 565218 492466 565454
rect 492702 565218 492734 565454
rect 492114 529774 492734 565218
rect 492114 529538 492146 529774
rect 492382 529538 492466 529774
rect 492702 529538 492734 529774
rect 492114 529454 492734 529538
rect 492114 529218 492146 529454
rect 492382 529218 492466 529454
rect 492702 529218 492734 529454
rect 482691 517580 482757 517581
rect 482691 517516 482692 517580
rect 482756 517516 482757 517580
rect 482691 517515 482757 517516
rect 482163 507454 482483 507486
rect 482163 507218 482205 507454
rect 482441 507218 482483 507454
rect 482163 507134 482483 507218
rect 482163 506898 482205 507134
rect 482441 506898 482483 507134
rect 482163 506866 482483 506898
rect 480954 482378 480986 482614
rect 481222 482378 481306 482614
rect 481542 482378 481574 482614
rect 480954 482294 481574 482378
rect 480954 482058 480986 482294
rect 481222 482058 481306 482294
rect 481542 482058 481574 482294
rect 480954 453692 481574 482058
rect 482694 462909 482754 517515
rect 483382 511174 483702 511206
rect 483382 510938 483424 511174
rect 483660 510938 483702 511174
rect 483382 510854 483702 510938
rect 483382 510618 483424 510854
rect 483660 510618 483702 510854
rect 483382 510586 483702 510618
rect 485820 511174 486140 511206
rect 485820 510938 485862 511174
rect 486098 510938 486140 511174
rect 485820 510854 486140 510938
rect 485820 510618 485862 510854
rect 486098 510618 486140 510854
rect 485820 510586 486140 510618
rect 488258 511174 488578 511206
rect 488258 510938 488300 511174
rect 488536 510938 488578 511174
rect 488258 510854 488578 510938
rect 488258 510618 488300 510854
rect 488536 510618 488578 510854
rect 488258 510586 488578 510618
rect 490696 511174 491016 511206
rect 490696 510938 490738 511174
rect 490974 510938 491016 511174
rect 490696 510854 491016 510938
rect 490696 510618 490738 510854
rect 490974 510618 491016 510854
rect 490696 510586 491016 510618
rect 484601 507454 484921 507486
rect 484601 507218 484643 507454
rect 484879 507218 484921 507454
rect 484601 507134 484921 507218
rect 484601 506898 484643 507134
rect 484879 506898 484921 507134
rect 484601 506866 484921 506898
rect 487039 507454 487359 507486
rect 487039 507218 487081 507454
rect 487317 507218 487359 507454
rect 487039 507134 487359 507218
rect 487039 506898 487081 507134
rect 487317 506898 487359 507134
rect 487039 506866 487359 506898
rect 489477 507454 489797 507486
rect 489477 507218 489519 507454
rect 489755 507218 489797 507454
rect 489477 507134 489797 507218
rect 489477 506898 489519 507134
rect 489755 506898 489797 507134
rect 489477 506866 489797 506898
rect 484674 486334 485294 500068
rect 484674 486098 484706 486334
rect 484942 486098 485026 486334
rect 485262 486098 485294 486334
rect 484674 486014 485294 486098
rect 484674 485778 484706 486014
rect 484942 485778 485026 486014
rect 485262 485778 485294 486014
rect 482691 462908 482757 462909
rect 482691 462844 482692 462908
rect 482756 462844 482757 462908
rect 482691 462843 482757 462844
rect 484674 450334 485294 485778
rect 488394 490054 489014 500068
rect 489315 496908 489381 496909
rect 489315 496844 489316 496908
rect 489380 496844 489381 496908
rect 489315 496843 489381 496844
rect 488394 489818 488426 490054
rect 488662 489818 488746 490054
rect 488982 489818 489014 490054
rect 488394 489734 489014 489818
rect 488394 489498 488426 489734
rect 488662 489498 488746 489734
rect 488982 489498 489014 489734
rect 488394 454007 489014 489498
rect 488394 453771 488426 454007
rect 488662 453771 488746 454007
rect 488982 453771 489014 454007
rect 488394 453692 489014 453771
rect 484674 450098 484706 450334
rect 484942 450098 485026 450334
rect 485262 450098 485294 450334
rect 484674 450014 485294 450098
rect 484674 449778 484706 450014
rect 484942 449778 485026 450014
rect 485262 449778 485294 450014
rect 480833 439174 481153 439206
rect 480833 438938 480875 439174
rect 481111 438938 481153 439174
rect 480833 438854 481153 438938
rect 480833 438618 480875 438854
rect 481111 438618 481153 438854
rect 480833 438586 481153 438618
rect 483306 435454 483626 435486
rect 483306 435218 483348 435454
rect 483584 435218 483626 435454
rect 483306 435134 483626 435218
rect 483306 434898 483348 435134
rect 483584 434898 483626 435134
rect 483306 434866 483626 434898
rect 484674 414334 485294 449778
rect 485778 439174 486098 439206
rect 485778 438938 485820 439174
rect 486056 438938 486098 439174
rect 485778 438854 486098 438938
rect 485778 438618 485820 438854
rect 486056 438618 486098 438854
rect 485778 438586 486098 438618
rect 488251 435454 488571 435486
rect 488251 435218 488293 435454
rect 488529 435218 488571 435454
rect 488251 435134 488571 435218
rect 488251 434898 488293 435134
rect 488529 434898 488571 435134
rect 488251 434866 488571 434898
rect 484674 414098 484706 414334
rect 484942 414098 485026 414334
rect 485262 414098 485294 414334
rect 484674 414014 485294 414098
rect 484674 413778 484706 414014
rect 484942 413778 485026 414014
rect 485262 413778 485294 414014
rect 478827 389060 478893 389061
rect 478827 388996 478828 389060
rect 478892 388996 478893 389060
rect 478827 388995 478893 388996
rect 484674 385580 485294 413778
rect 489318 387021 489378 496843
rect 492114 493774 492734 529218
rect 492114 493538 492146 493774
rect 492382 493538 492466 493774
rect 492702 493538 492734 493774
rect 492114 493454 492734 493538
rect 492114 493218 492146 493454
rect 492382 493218 492466 493454
rect 492702 493218 492734 493454
rect 492114 457774 492734 493218
rect 492114 457538 492146 457774
rect 492382 457538 492466 457774
rect 492702 457538 492734 457774
rect 492114 457454 492734 457538
rect 492114 457218 492146 457454
rect 492382 457218 492466 457454
rect 492702 457218 492734 457454
rect 490723 439174 491043 439206
rect 490723 438938 490765 439174
rect 491001 438938 491043 439174
rect 490723 438854 491043 438938
rect 490723 438618 490765 438854
rect 491001 438618 491043 438854
rect 490723 438586 491043 438618
rect 492114 421774 492734 457218
rect 492114 421538 492146 421774
rect 492382 421538 492466 421774
rect 492702 421538 492734 421774
rect 492114 421454 492734 421538
rect 492114 421218 492146 421454
rect 492382 421218 492466 421454
rect 492702 421218 492734 421454
rect 489315 387020 489381 387021
rect 489315 386956 489316 387020
rect 489380 386956 489381 387020
rect 489315 386955 489381 386956
rect 492114 385774 492734 421218
rect 492114 385538 492146 385774
rect 492382 385538 492466 385774
rect 492702 385538 492734 385774
rect 492114 385454 492734 385538
rect 492114 385218 492146 385454
rect 492382 385218 492466 385454
rect 492702 385218 492734 385454
rect 492114 384817 492734 385218
rect 495834 569494 496454 601103
rect 495834 569258 495866 569494
rect 496102 569258 496186 569494
rect 496422 569258 496454 569494
rect 495834 569174 496454 569258
rect 495834 568938 495866 569174
rect 496102 568938 496186 569174
rect 496422 568938 496454 569174
rect 495834 533494 496454 568938
rect 495834 533258 495866 533494
rect 496102 533258 496186 533494
rect 496422 533258 496454 533494
rect 495834 533174 496454 533258
rect 495834 532938 495866 533174
rect 496102 532938 496186 533174
rect 496422 532938 496454 533174
rect 495834 497494 496454 532938
rect 495834 497258 495866 497494
rect 496102 497258 496186 497494
rect 496422 497258 496454 497494
rect 495834 497174 496454 497258
rect 495834 496938 495866 497174
rect 496102 496938 496186 497174
rect 496422 496938 496454 497174
rect 495834 461494 496454 496938
rect 495834 461258 495866 461494
rect 496102 461258 496186 461494
rect 496422 461258 496454 461494
rect 495834 461174 496454 461258
rect 495834 460938 495866 461174
rect 496102 460938 496186 461174
rect 496422 460938 496454 461174
rect 495834 425494 496454 460938
rect 495834 425258 495866 425494
rect 496102 425258 496186 425494
rect 496422 425258 496454 425494
rect 495834 425174 496454 425258
rect 495834 424938 495866 425174
rect 496102 424938 496186 425174
rect 496422 424938 496454 425174
rect 495834 389494 496454 424938
rect 495834 389258 495866 389494
rect 496102 389258 496186 389494
rect 496422 389258 496454 389494
rect 495834 389174 496454 389258
rect 495834 388938 495866 389174
rect 496102 388938 496186 389174
rect 496422 388938 496454 389174
rect 495834 384817 496454 388938
rect 505794 579454 506414 601103
rect 505794 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 506414 579454
rect 505794 579134 506414 579218
rect 505794 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 506414 579134
rect 505794 543454 506414 578898
rect 505794 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 506414 543454
rect 505794 543134 506414 543218
rect 505794 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 506414 543134
rect 505794 507454 506414 542898
rect 505794 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 506414 507454
rect 505794 507134 506414 507218
rect 505794 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 506414 507134
rect 505794 471454 506414 506898
rect 505794 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 506414 471454
rect 505794 471134 506414 471218
rect 505794 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 506414 471134
rect 505794 435454 506414 470898
rect 505794 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 506414 435454
rect 505794 435134 506414 435218
rect 505794 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 506414 435134
rect 505794 399454 506414 434898
rect 505794 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 506414 399454
rect 505794 399134 506414 399218
rect 505794 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 506414 399134
rect 469568 367174 469888 367206
rect 469568 366938 469610 367174
rect 469846 366938 469888 367174
rect 469568 366854 469888 366938
rect 469568 366618 469610 366854
rect 469846 366618 469888 366854
rect 469568 366586 469888 366618
rect 500288 367174 500608 367206
rect 500288 366938 500330 367174
rect 500566 366938 500608 367174
rect 500288 366854 500608 366938
rect 500288 366618 500330 366854
rect 500566 366618 500608 366854
rect 500288 366586 500608 366618
rect 484928 363454 485248 363486
rect 484928 363218 484970 363454
rect 485206 363218 485248 363454
rect 484928 363134 485248 363218
rect 484928 362898 484970 363134
rect 485206 362898 485248 363134
rect 484928 362866 485248 362898
rect 505794 363454 506414 398898
rect 505794 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 506414 363454
rect 505794 363134 506414 363218
rect 505794 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 506414 363134
rect 459834 353258 459866 353494
rect 460102 353258 460186 353494
rect 460422 353258 460454 353494
rect 459834 353174 460454 353258
rect 459834 352938 459866 353174
rect 460102 352938 460186 353174
rect 460422 352938 460454 353174
rect 459834 317494 460454 352938
rect 469568 331174 469888 331206
rect 469568 330938 469610 331174
rect 469846 330938 469888 331174
rect 469568 330854 469888 330938
rect 469568 330618 469610 330854
rect 469846 330618 469888 330854
rect 469568 330586 469888 330618
rect 500288 331174 500608 331206
rect 500288 330938 500330 331174
rect 500566 330938 500608 331174
rect 500288 330854 500608 330938
rect 500288 330618 500330 330854
rect 500566 330618 500608 330854
rect 500288 330586 500608 330618
rect 484928 327454 485248 327486
rect 484928 327218 484970 327454
rect 485206 327218 485248 327454
rect 484928 327134 485248 327218
rect 484928 326898 484970 327134
rect 485206 326898 485248 327134
rect 484928 326866 485248 326898
rect 505794 327454 506414 362898
rect 505794 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 506414 327454
rect 505794 327134 506414 327218
rect 505794 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 506414 327134
rect 460795 320788 460861 320789
rect 460795 320724 460796 320788
rect 460860 320724 460861 320788
rect 460795 320723 460861 320724
rect 459834 317258 459866 317494
rect 460102 317258 460186 317494
rect 460422 317258 460454 317494
rect 459834 317174 460454 317258
rect 459834 316938 459866 317174
rect 460102 316938 460186 317174
rect 460422 316938 460454 317174
rect 459834 281494 460454 316938
rect 459834 281258 459866 281494
rect 460102 281258 460186 281494
rect 460422 281258 460454 281494
rect 459834 281174 460454 281258
rect 459834 280938 459866 281174
rect 460102 280938 460186 281174
rect 460422 280938 460454 281174
rect 459834 245494 460454 280938
rect 459834 245258 459866 245494
rect 460102 245258 460186 245494
rect 460422 245258 460454 245494
rect 459834 245174 460454 245258
rect 459834 244938 459866 245174
rect 460102 244938 460186 245174
rect 460422 244938 460454 245174
rect 459834 209494 460454 244938
rect 459834 209258 459866 209494
rect 460102 209258 460186 209494
rect 460422 209258 460454 209494
rect 459834 209174 460454 209258
rect 459834 208938 459866 209174
rect 460102 208938 460186 209174
rect 460422 208938 460454 209174
rect 459834 173494 460454 208938
rect 459834 173258 459866 173494
rect 460102 173258 460186 173494
rect 460422 173258 460454 173494
rect 459834 173174 460454 173258
rect 459834 172938 459866 173174
rect 460102 172938 460186 173174
rect 460422 172938 460454 173174
rect 459834 137494 460454 172938
rect 459834 137258 459866 137494
rect 460102 137258 460186 137494
rect 460422 137258 460454 137494
rect 459834 137174 460454 137258
rect 459834 136938 459866 137174
rect 460102 136938 460186 137174
rect 460422 136938 460454 137174
rect 459834 101494 460454 136938
rect 459834 101258 459866 101494
rect 460102 101258 460186 101494
rect 460422 101258 460454 101494
rect 459834 101174 460454 101258
rect 459834 100938 459866 101174
rect 460102 100938 460186 101174
rect 460422 100938 460454 101174
rect 405568 79174 405888 79206
rect 405568 78938 405610 79174
rect 405846 78938 405888 79174
rect 405568 78854 405888 78938
rect 405568 78618 405610 78854
rect 405846 78618 405888 78854
rect 405568 78586 405888 78618
rect 436288 79174 436608 79206
rect 436288 78938 436330 79174
rect 436566 78938 436608 79174
rect 436288 78854 436608 78938
rect 436288 78618 436330 78854
rect 436566 78618 436608 78854
rect 436288 78586 436608 78618
rect 390208 75454 390528 75486
rect 390208 75218 390250 75454
rect 390486 75218 390528 75454
rect 390208 75134 390528 75218
rect 390208 74898 390250 75134
rect 390486 74898 390528 75134
rect 390208 74866 390528 74898
rect 420928 75454 421248 75486
rect 420928 75218 420970 75454
rect 421206 75218 421248 75454
rect 420928 75134 421248 75218
rect 420928 74898 420970 75134
rect 421206 74898 421248 75134
rect 420928 74866 421248 74898
rect 451648 75454 451968 75486
rect 451648 75218 451690 75454
rect 451926 75218 451968 75454
rect 451648 75134 451968 75218
rect 451648 74898 451690 75134
rect 451926 74898 451968 75134
rect 451648 74866 451968 74898
rect 384114 61538 384146 61774
rect 384382 61538 384466 61774
rect 384702 61538 384734 61774
rect 384114 61454 384734 61538
rect 384114 61218 384146 61454
rect 384382 61218 384466 61454
rect 384702 61218 384734 61454
rect 384114 25774 384734 61218
rect 459834 65494 460454 100938
rect 459834 65258 459866 65494
rect 460102 65258 460186 65494
rect 460422 65258 460454 65494
rect 459834 65174 460454 65258
rect 459834 64938 459866 65174
rect 460102 64938 460186 65174
rect 460422 64938 460454 65174
rect 405568 43174 405888 43206
rect 405568 42938 405610 43174
rect 405846 42938 405888 43174
rect 405568 42854 405888 42938
rect 405568 42618 405610 42854
rect 405846 42618 405888 42854
rect 405568 42586 405888 42618
rect 436288 43174 436608 43206
rect 436288 42938 436330 43174
rect 436566 42938 436608 43174
rect 436288 42854 436608 42938
rect 436288 42618 436330 42854
rect 436566 42618 436608 42854
rect 436288 42586 436608 42618
rect 390208 39454 390528 39486
rect 390208 39218 390250 39454
rect 390486 39218 390528 39454
rect 390208 39134 390528 39218
rect 390208 38898 390250 39134
rect 390486 38898 390528 39134
rect 390208 38866 390528 38898
rect 420928 39454 421248 39486
rect 420928 39218 420970 39454
rect 421206 39218 421248 39454
rect 420928 39134 421248 39218
rect 420928 38898 420970 39134
rect 421206 38898 421248 39134
rect 420928 38866 421248 38898
rect 451648 39454 451968 39486
rect 451648 39218 451690 39454
rect 451926 39218 451968 39454
rect 451648 39134 451968 39218
rect 451648 38898 451690 39134
rect 451926 38898 451968 39134
rect 451648 38866 451968 38898
rect 384114 25538 384146 25774
rect 384382 25538 384466 25774
rect 384702 25538 384734 25774
rect 384114 25454 384734 25538
rect 384114 25218 384146 25454
rect 384382 25218 384466 25454
rect 384702 25218 384734 25454
rect 384114 -6106 384734 25218
rect 384114 -6342 384146 -6106
rect 384382 -6342 384466 -6106
rect 384702 -6342 384734 -6106
rect 384114 -6426 384734 -6342
rect 384114 -6662 384146 -6426
rect 384382 -6662 384466 -6426
rect 384702 -6662 384734 -6426
rect 384114 -7654 384734 -6662
rect 387834 29494 388454 31919
rect 387834 29258 387866 29494
rect 388102 29258 388186 29494
rect 388422 29258 388454 29494
rect 387834 29174 388454 29258
rect 387834 28938 387866 29174
rect 388102 28938 388186 29174
rect 388422 28938 388454 29174
rect 387834 -7066 388454 28938
rect 387834 -7302 387866 -7066
rect 388102 -7302 388186 -7066
rect 388422 -7302 388454 -7066
rect 387834 -7386 388454 -7302
rect 387834 -7622 387866 -7386
rect 388102 -7622 388186 -7386
rect 388422 -7622 388454 -7386
rect 387834 -7654 388454 -7622
rect 397794 3454 398414 31919
rect 397794 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 398414 3454
rect 397794 3134 398414 3218
rect 397794 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 398414 3134
rect 397794 -346 398414 2898
rect 397794 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 398414 -346
rect 397794 -666 398414 -582
rect 397794 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 398414 -666
rect 397794 -7654 398414 -902
rect 401514 7174 402134 31919
rect 401514 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 402134 7174
rect 401514 6854 402134 6938
rect 401514 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 402134 6854
rect 401514 -1306 402134 6618
rect 401514 -1542 401546 -1306
rect 401782 -1542 401866 -1306
rect 402102 -1542 402134 -1306
rect 401514 -1626 402134 -1542
rect 401514 -1862 401546 -1626
rect 401782 -1862 401866 -1626
rect 402102 -1862 402134 -1626
rect 401514 -7654 402134 -1862
rect 405234 10894 405854 30068
rect 405234 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 405854 10894
rect 405234 10574 405854 10658
rect 405234 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 405854 10574
rect 405234 -2266 405854 10338
rect 405234 -2502 405266 -2266
rect 405502 -2502 405586 -2266
rect 405822 -2502 405854 -2266
rect 405234 -2586 405854 -2502
rect 405234 -2822 405266 -2586
rect 405502 -2822 405586 -2586
rect 405822 -2822 405854 -2586
rect 405234 -7654 405854 -2822
rect 408954 14614 409574 31919
rect 408954 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 409574 14614
rect 408954 14294 409574 14378
rect 408954 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 409574 14294
rect 408954 -3226 409574 14058
rect 408954 -3462 408986 -3226
rect 409222 -3462 409306 -3226
rect 409542 -3462 409574 -3226
rect 408954 -3546 409574 -3462
rect 408954 -3782 408986 -3546
rect 409222 -3782 409306 -3546
rect 409542 -3782 409574 -3546
rect 408954 -7654 409574 -3782
rect 412674 18334 413294 31919
rect 412674 18098 412706 18334
rect 412942 18098 413026 18334
rect 413262 18098 413294 18334
rect 412674 18014 413294 18098
rect 412674 17778 412706 18014
rect 412942 17778 413026 18014
rect 413262 17778 413294 18014
rect 412674 -4186 413294 17778
rect 412674 -4422 412706 -4186
rect 412942 -4422 413026 -4186
rect 413262 -4422 413294 -4186
rect 412674 -4506 413294 -4422
rect 412674 -4742 412706 -4506
rect 412942 -4742 413026 -4506
rect 413262 -4742 413294 -4506
rect 412674 -7654 413294 -4742
rect 416394 22054 417014 31919
rect 416394 21818 416426 22054
rect 416662 21818 416746 22054
rect 416982 21818 417014 22054
rect 416394 21734 417014 21818
rect 416394 21498 416426 21734
rect 416662 21498 416746 21734
rect 416982 21498 417014 21734
rect 416394 -5146 417014 21498
rect 416394 -5382 416426 -5146
rect 416662 -5382 416746 -5146
rect 416982 -5382 417014 -5146
rect 416394 -5466 417014 -5382
rect 416394 -5702 416426 -5466
rect 416662 -5702 416746 -5466
rect 416982 -5702 417014 -5466
rect 416394 -7654 417014 -5702
rect 420114 25774 420734 31919
rect 420114 25538 420146 25774
rect 420382 25538 420466 25774
rect 420702 25538 420734 25774
rect 420114 25454 420734 25538
rect 420114 25218 420146 25454
rect 420382 25218 420466 25454
rect 420702 25218 420734 25454
rect 420114 -6106 420734 25218
rect 420114 -6342 420146 -6106
rect 420382 -6342 420466 -6106
rect 420702 -6342 420734 -6106
rect 420114 -6426 420734 -6342
rect 420114 -6662 420146 -6426
rect 420382 -6662 420466 -6426
rect 420702 -6662 420734 -6426
rect 420114 -7654 420734 -6662
rect 423834 29494 424454 31919
rect 423834 29258 423866 29494
rect 424102 29258 424186 29494
rect 424422 29258 424454 29494
rect 423834 29174 424454 29258
rect 423834 28938 423866 29174
rect 424102 28938 424186 29174
rect 424422 28938 424454 29174
rect 423834 -7066 424454 28938
rect 423834 -7302 423866 -7066
rect 424102 -7302 424186 -7066
rect 424422 -7302 424454 -7066
rect 423834 -7386 424454 -7302
rect 423834 -7622 423866 -7386
rect 424102 -7622 424186 -7386
rect 424422 -7622 424454 -7386
rect 423834 -7654 424454 -7622
rect 433794 3454 434414 31919
rect 433794 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 434414 3454
rect 433794 3134 434414 3218
rect 433794 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 434414 3134
rect 433794 -346 434414 2898
rect 433794 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 434414 -346
rect 433794 -666 434414 -582
rect 433794 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 434414 -666
rect 433794 -7654 434414 -902
rect 437514 7174 438134 31919
rect 437514 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 438134 7174
rect 437514 6854 438134 6938
rect 437514 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 438134 6854
rect 437514 -1306 438134 6618
rect 437514 -1542 437546 -1306
rect 437782 -1542 437866 -1306
rect 438102 -1542 438134 -1306
rect 437514 -1626 438134 -1542
rect 437514 -1862 437546 -1626
rect 437782 -1862 437866 -1626
rect 438102 -1862 438134 -1626
rect 437514 -7654 438134 -1862
rect 441234 10894 441854 31919
rect 441234 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 441854 10894
rect 441234 10574 441854 10658
rect 441234 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 441854 10574
rect 441234 -2266 441854 10338
rect 441234 -2502 441266 -2266
rect 441502 -2502 441586 -2266
rect 441822 -2502 441854 -2266
rect 441234 -2586 441854 -2502
rect 441234 -2822 441266 -2586
rect 441502 -2822 441586 -2586
rect 441822 -2822 441854 -2586
rect 441234 -7654 441854 -2822
rect 444954 14614 445574 31919
rect 444954 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 445574 14614
rect 444954 14294 445574 14378
rect 444954 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 445574 14294
rect 444954 -3226 445574 14058
rect 444954 -3462 444986 -3226
rect 445222 -3462 445306 -3226
rect 445542 -3462 445574 -3226
rect 444954 -3546 445574 -3462
rect 444954 -3782 444986 -3546
rect 445222 -3782 445306 -3546
rect 445542 -3782 445574 -3546
rect 444954 -7654 445574 -3782
rect 448674 18334 449294 31919
rect 448674 18098 448706 18334
rect 448942 18098 449026 18334
rect 449262 18098 449294 18334
rect 448674 18014 449294 18098
rect 448674 17778 448706 18014
rect 448942 17778 449026 18014
rect 449262 17778 449294 18014
rect 448674 -4186 449294 17778
rect 448674 -4422 448706 -4186
rect 448942 -4422 449026 -4186
rect 449262 -4422 449294 -4186
rect 448674 -4506 449294 -4422
rect 448674 -4742 448706 -4506
rect 448942 -4742 449026 -4506
rect 449262 -4742 449294 -4506
rect 448674 -7654 449294 -4742
rect 452394 22054 453014 31919
rect 452394 21818 452426 22054
rect 452662 21818 452746 22054
rect 452982 21818 453014 22054
rect 452394 21734 453014 21818
rect 452394 21498 452426 21734
rect 452662 21498 452746 21734
rect 452982 21498 453014 21734
rect 452394 -5146 453014 21498
rect 452394 -5382 452426 -5146
rect 452662 -5382 452746 -5146
rect 452982 -5382 453014 -5146
rect 452394 -5466 453014 -5382
rect 452394 -5702 452426 -5466
rect 452662 -5702 452746 -5466
rect 452982 -5702 453014 -5466
rect 452394 -7654 453014 -5702
rect 456114 25774 456734 31919
rect 456114 25538 456146 25774
rect 456382 25538 456466 25774
rect 456702 25538 456734 25774
rect 456114 25454 456734 25538
rect 456114 25218 456146 25454
rect 456382 25218 456466 25454
rect 456702 25218 456734 25454
rect 456114 -6106 456734 25218
rect 456114 -6342 456146 -6106
rect 456382 -6342 456466 -6106
rect 456702 -6342 456734 -6106
rect 456114 -6426 456734 -6342
rect 456114 -6662 456146 -6426
rect 456382 -6662 456466 -6426
rect 456702 -6662 456734 -6426
rect 456114 -7654 456734 -6662
rect 459834 29494 460454 64938
rect 459834 29258 459866 29494
rect 460102 29258 460186 29494
rect 460422 29258 460454 29494
rect 459834 29174 460454 29258
rect 459834 28938 459866 29174
rect 460102 28938 460186 29174
rect 460422 28938 460454 29174
rect 459834 -7066 460454 28938
rect 460798 3365 460858 320723
rect 477234 298894 477854 322287
rect 477234 298658 477266 298894
rect 477502 298658 477586 298894
rect 477822 298658 477854 298894
rect 477234 298574 477854 298658
rect 477234 298338 477266 298574
rect 477502 298338 477586 298574
rect 477822 298338 477854 298574
rect 477234 262894 477854 298338
rect 477234 262658 477266 262894
rect 477502 262658 477586 262894
rect 477822 262658 477854 262894
rect 477234 262574 477854 262658
rect 477234 262338 477266 262574
rect 477502 262338 477586 262574
rect 477822 262338 477854 262574
rect 477234 259417 477854 262338
rect 480954 302614 481574 322287
rect 480954 302378 480986 302614
rect 481222 302378 481306 302614
rect 481542 302378 481574 302614
rect 480954 302294 481574 302378
rect 480954 302058 480986 302294
rect 481222 302058 481306 302294
rect 481542 302058 481574 302294
rect 480954 266614 481574 302058
rect 480954 266378 480986 266614
rect 481222 266378 481306 266614
rect 481542 266378 481574 266614
rect 480954 266294 481574 266378
rect 480954 266058 480986 266294
rect 481222 266058 481306 266294
rect 481542 266058 481574 266294
rect 480954 259417 481574 266058
rect 484674 306334 485294 322068
rect 484674 306098 484706 306334
rect 484942 306098 485026 306334
rect 485262 306098 485294 306334
rect 484674 306014 485294 306098
rect 484674 305778 484706 306014
rect 484942 305778 485026 306014
rect 485262 305778 485294 306014
rect 484674 270334 485294 305778
rect 484674 270098 484706 270334
rect 484942 270098 485026 270334
rect 485262 270098 485294 270334
rect 484674 270014 485294 270098
rect 484674 269778 484706 270014
rect 484942 269778 485026 270014
rect 485262 269778 485294 270014
rect 484674 259417 485294 269778
rect 488394 310054 489014 322287
rect 488394 309818 488426 310054
rect 488662 309818 488746 310054
rect 488982 309818 489014 310054
rect 488394 309734 489014 309818
rect 488394 309498 488426 309734
rect 488662 309498 488746 309734
rect 488982 309498 489014 309734
rect 488394 274054 489014 309498
rect 488394 273818 488426 274054
rect 488662 273818 488746 274054
rect 488982 273818 489014 274054
rect 488394 273734 489014 273818
rect 488394 273498 488426 273734
rect 488662 273498 488746 273734
rect 488982 273498 489014 273734
rect 488394 259417 489014 273498
rect 492114 313774 492734 322287
rect 492114 313538 492146 313774
rect 492382 313538 492466 313774
rect 492702 313538 492734 313774
rect 492114 313454 492734 313538
rect 492114 313218 492146 313454
rect 492382 313218 492466 313454
rect 492702 313218 492734 313454
rect 492114 277774 492734 313218
rect 492114 277538 492146 277774
rect 492382 277538 492466 277774
rect 492702 277538 492734 277774
rect 492114 277454 492734 277538
rect 492114 277218 492146 277454
rect 492382 277218 492466 277454
rect 492702 277218 492734 277454
rect 492114 259417 492734 277218
rect 495834 317494 496454 322287
rect 495834 317258 495866 317494
rect 496102 317258 496186 317494
rect 496422 317258 496454 317494
rect 495834 317174 496454 317258
rect 495834 316938 495866 317174
rect 496102 316938 496186 317174
rect 496422 316938 496454 317174
rect 495834 281494 496454 316938
rect 495834 281258 495866 281494
rect 496102 281258 496186 281494
rect 496422 281258 496454 281494
rect 495834 281174 496454 281258
rect 495834 280938 495866 281174
rect 496102 280938 496186 281174
rect 496422 280938 496454 281174
rect 495834 259417 496454 280938
rect 505794 291454 506414 326898
rect 509514 583174 510134 601103
rect 509514 582938 509546 583174
rect 509782 582938 509866 583174
rect 510102 582938 510134 583174
rect 509514 582854 510134 582938
rect 509514 582618 509546 582854
rect 509782 582618 509866 582854
rect 510102 582618 510134 582854
rect 509514 547174 510134 582618
rect 509514 546938 509546 547174
rect 509782 546938 509866 547174
rect 510102 546938 510134 547174
rect 509514 546854 510134 546938
rect 509514 546618 509546 546854
rect 509782 546618 509866 546854
rect 510102 546618 510134 546854
rect 509514 511174 510134 546618
rect 509514 510938 509546 511174
rect 509782 510938 509866 511174
rect 510102 510938 510134 511174
rect 509514 510854 510134 510938
rect 509514 510618 509546 510854
rect 509782 510618 509866 510854
rect 510102 510618 510134 510854
rect 509514 475174 510134 510618
rect 509514 474938 509546 475174
rect 509782 474938 509866 475174
rect 510102 474938 510134 475174
rect 509514 474854 510134 474938
rect 509514 474618 509546 474854
rect 509782 474618 509866 474854
rect 510102 474618 510134 474854
rect 509514 439174 510134 474618
rect 509514 438938 509546 439174
rect 509782 438938 509866 439174
rect 510102 438938 510134 439174
rect 509514 438854 510134 438938
rect 509514 438618 509546 438854
rect 509782 438618 509866 438854
rect 510102 438618 510134 438854
rect 509514 403174 510134 438618
rect 509514 402938 509546 403174
rect 509782 402938 509866 403174
rect 510102 402938 510134 403174
rect 509514 402854 510134 402938
rect 509514 402618 509546 402854
rect 509782 402618 509866 402854
rect 510102 402618 510134 402854
rect 509514 367174 510134 402618
rect 509514 366938 509546 367174
rect 509782 366938 509866 367174
rect 510102 366938 510134 367174
rect 509514 366854 510134 366938
rect 509514 366618 509546 366854
rect 509782 366618 509866 366854
rect 510102 366618 510134 366854
rect 509514 331174 510134 366618
rect 513234 586894 513854 601103
rect 513234 586658 513266 586894
rect 513502 586658 513586 586894
rect 513822 586658 513854 586894
rect 513234 586574 513854 586658
rect 513234 586338 513266 586574
rect 513502 586338 513586 586574
rect 513822 586338 513854 586574
rect 513234 550894 513854 586338
rect 513234 550658 513266 550894
rect 513502 550658 513586 550894
rect 513822 550658 513854 550894
rect 513234 550574 513854 550658
rect 513234 550338 513266 550574
rect 513502 550338 513586 550574
rect 513822 550338 513854 550574
rect 513234 514894 513854 550338
rect 513234 514658 513266 514894
rect 513502 514658 513586 514894
rect 513822 514658 513854 514894
rect 513234 514574 513854 514658
rect 513234 514338 513266 514574
rect 513502 514338 513586 514574
rect 513822 514338 513854 514574
rect 513234 478894 513854 514338
rect 513234 478658 513266 478894
rect 513502 478658 513586 478894
rect 513822 478658 513854 478894
rect 513234 478574 513854 478658
rect 513234 478338 513266 478574
rect 513502 478338 513586 478574
rect 513822 478338 513854 478574
rect 513234 442894 513854 478338
rect 513234 442658 513266 442894
rect 513502 442658 513586 442894
rect 513822 442658 513854 442894
rect 513234 442574 513854 442658
rect 513234 442338 513266 442574
rect 513502 442338 513586 442574
rect 513822 442338 513854 442574
rect 513234 406894 513854 442338
rect 513234 406658 513266 406894
rect 513502 406658 513586 406894
rect 513822 406658 513854 406894
rect 513234 406574 513854 406658
rect 513234 406338 513266 406574
rect 513502 406338 513586 406574
rect 513822 406338 513854 406574
rect 513234 370894 513854 406338
rect 513234 370658 513266 370894
rect 513502 370658 513586 370894
rect 513822 370658 513854 370894
rect 513234 370574 513854 370658
rect 513234 370338 513266 370574
rect 513502 370338 513586 370574
rect 513822 370338 513854 370574
rect 511211 335748 511277 335749
rect 511211 335684 511212 335748
rect 511276 335684 511277 335748
rect 511211 335683 511277 335684
rect 510659 333028 510725 333029
rect 510659 332964 510660 333028
rect 510724 332964 510725 333028
rect 510659 332963 510725 332964
rect 509514 330938 509546 331174
rect 509782 330938 509866 331174
rect 510102 330938 510134 331174
rect 509514 330854 510134 330938
rect 509514 330618 509546 330854
rect 509782 330618 509866 330854
rect 510102 330618 510134 330854
rect 509187 316708 509253 316709
rect 509187 316644 509188 316708
rect 509252 316644 509253 316708
rect 509187 316643 509253 316644
rect 509190 311910 509250 316643
rect 509006 311850 509250 311910
rect 509006 306101 509066 311850
rect 509003 306100 509069 306101
rect 509003 306036 509004 306100
rect 509068 306036 509069 306100
rect 509003 306035 509069 306036
rect 505794 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 506414 291454
rect 505794 291134 506414 291218
rect 505794 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 506414 291134
rect 505794 259417 506414 290898
rect 509514 295174 510134 330618
rect 510475 327588 510541 327589
rect 510475 327524 510476 327588
rect 510540 327524 510541 327588
rect 510475 327523 510541 327524
rect 510291 324324 510357 324325
rect 510291 324260 510292 324324
rect 510356 324260 510357 324324
rect 510291 324259 510357 324260
rect 510294 316709 510354 324259
rect 510478 321877 510538 327523
rect 510475 321876 510541 321877
rect 510475 321812 510476 321876
rect 510540 321812 510541 321876
rect 510475 321811 510541 321812
rect 510291 316708 510357 316709
rect 510291 316644 510292 316708
rect 510356 316644 510357 316708
rect 510291 316643 510357 316644
rect 510662 297669 510722 332963
rect 510843 326500 510909 326501
rect 510843 326436 510844 326500
rect 510908 326436 510909 326500
rect 510843 326435 510909 326436
rect 510846 303109 510906 326435
rect 511027 323780 511093 323781
rect 511027 323716 511028 323780
rect 511092 323716 511093 323780
rect 511027 323715 511093 323716
rect 511030 305965 511090 323715
rect 511214 318341 511274 335683
rect 513234 334894 513854 370338
rect 513234 334658 513266 334894
rect 513502 334658 513586 334894
rect 513822 334658 513854 334894
rect 513234 334574 513854 334658
rect 513234 334338 513266 334574
rect 513502 334338 513586 334574
rect 513822 334338 513854 334574
rect 511211 318340 511277 318341
rect 511211 318276 511212 318340
rect 511276 318276 511277 318340
rect 511211 318275 511277 318276
rect 511027 305964 511093 305965
rect 511027 305900 511028 305964
rect 511092 305900 511093 305964
rect 511027 305899 511093 305900
rect 510843 303108 510909 303109
rect 510843 303044 510844 303108
rect 510908 303044 510909 303108
rect 510843 303043 510909 303044
rect 513234 298894 513854 334338
rect 516954 590614 517574 601103
rect 516954 590378 516986 590614
rect 517222 590378 517306 590614
rect 517542 590378 517574 590614
rect 516954 590294 517574 590378
rect 516954 590058 516986 590294
rect 517222 590058 517306 590294
rect 517542 590058 517574 590294
rect 516954 554614 517574 590058
rect 516954 554378 516986 554614
rect 517222 554378 517306 554614
rect 517542 554378 517574 554614
rect 516954 554294 517574 554378
rect 516954 554058 516986 554294
rect 517222 554058 517306 554294
rect 517542 554058 517574 554294
rect 516954 518614 517574 554058
rect 516954 518378 516986 518614
rect 517222 518378 517306 518614
rect 517542 518378 517574 518614
rect 516954 518294 517574 518378
rect 516954 518058 516986 518294
rect 517222 518058 517306 518294
rect 517542 518058 517574 518294
rect 516954 482614 517574 518058
rect 516954 482378 516986 482614
rect 517222 482378 517306 482614
rect 517542 482378 517574 482614
rect 516954 482294 517574 482378
rect 516954 482058 516986 482294
rect 517222 482058 517306 482294
rect 517542 482058 517574 482294
rect 516954 446614 517574 482058
rect 516954 446378 516986 446614
rect 517222 446378 517306 446614
rect 517542 446378 517574 446614
rect 516954 446294 517574 446378
rect 516954 446058 516986 446294
rect 517222 446058 517306 446294
rect 517542 446058 517574 446294
rect 516954 410614 517574 446058
rect 516954 410378 516986 410614
rect 517222 410378 517306 410614
rect 517542 410378 517574 410614
rect 516954 410294 517574 410378
rect 516954 410058 516986 410294
rect 517222 410058 517306 410294
rect 517542 410058 517574 410294
rect 516954 374614 517574 410058
rect 516954 374378 516986 374614
rect 517222 374378 517306 374614
rect 517542 374378 517574 374614
rect 516954 374294 517574 374378
rect 516954 374058 516986 374294
rect 517222 374058 517306 374294
rect 517542 374058 517574 374294
rect 516954 338614 517574 374058
rect 516954 338378 516986 338614
rect 517222 338378 517306 338614
rect 517542 338378 517574 338614
rect 516954 338294 517574 338378
rect 516954 338058 516986 338294
rect 517222 338058 517306 338294
rect 517542 338058 517574 338294
rect 514707 331940 514773 331941
rect 514707 331876 514708 331940
rect 514772 331876 514773 331940
rect 514707 331875 514773 331876
rect 514710 331230 514770 331875
rect 514891 331396 514957 331397
rect 514891 331332 514892 331396
rect 514956 331332 514957 331396
rect 514891 331331 514957 331332
rect 514526 331170 514770 331230
rect 514339 328676 514405 328677
rect 514339 328612 514340 328676
rect 514404 328612 514405 328676
rect 514339 328611 514405 328612
rect 514155 324868 514221 324869
rect 514155 324804 514156 324868
rect 514220 324804 514221 324868
rect 514155 324803 514221 324804
rect 513234 298658 513266 298894
rect 513502 298658 513586 298894
rect 513822 298658 513854 298894
rect 513234 298574 513854 298658
rect 513234 298338 513266 298574
rect 513502 298338 513586 298574
rect 513822 298338 513854 298574
rect 510659 297668 510725 297669
rect 510659 297604 510660 297668
rect 510724 297604 510725 297668
rect 510659 297603 510725 297604
rect 509514 294938 509546 295174
rect 509782 294938 509866 295174
rect 510102 294938 510134 295174
rect 509514 294854 510134 294938
rect 509514 294618 509546 294854
rect 509782 294618 509866 294854
rect 510102 294618 510134 294854
rect 509514 259417 510134 294618
rect 513234 262894 513854 298338
rect 514158 297533 514218 324803
rect 514342 320245 514402 328611
rect 514339 320244 514405 320245
rect 514339 320180 514340 320244
rect 514404 320180 514405 320244
rect 514339 320179 514405 320180
rect 514526 311910 514586 331170
rect 514526 311850 514770 311910
rect 514155 297532 514221 297533
rect 514155 297468 514156 297532
rect 514220 297468 514221 297532
rect 514155 297467 514221 297468
rect 514710 291821 514770 311850
rect 514894 297397 514954 331331
rect 515075 329220 515141 329221
rect 515075 329156 515076 329220
rect 515140 329156 515141 329220
rect 515075 329155 515141 329156
rect 515078 321741 515138 329155
rect 515075 321740 515141 321741
rect 515075 321676 515076 321740
rect 515140 321676 515141 321740
rect 515075 321675 515141 321676
rect 516954 302614 517574 338058
rect 520674 594334 521294 629778
rect 520674 594098 520706 594334
rect 520942 594098 521026 594334
rect 521262 594098 521294 594334
rect 520674 594014 521294 594098
rect 520674 593778 520706 594014
rect 520942 593778 521026 594014
rect 521262 593778 521294 594014
rect 520674 558334 521294 593778
rect 520674 558098 520706 558334
rect 520942 558098 521026 558334
rect 521262 558098 521294 558334
rect 520674 558014 521294 558098
rect 520674 557778 520706 558014
rect 520942 557778 521026 558014
rect 521262 557778 521294 558014
rect 520674 522334 521294 557778
rect 520674 522098 520706 522334
rect 520942 522098 521026 522334
rect 521262 522098 521294 522334
rect 520674 522014 521294 522098
rect 520674 521778 520706 522014
rect 520942 521778 521026 522014
rect 521262 521778 521294 522014
rect 520674 486334 521294 521778
rect 520674 486098 520706 486334
rect 520942 486098 521026 486334
rect 521262 486098 521294 486334
rect 520674 486014 521294 486098
rect 520674 485778 520706 486014
rect 520942 485778 521026 486014
rect 521262 485778 521294 486014
rect 520674 450334 521294 485778
rect 520674 450098 520706 450334
rect 520942 450098 521026 450334
rect 521262 450098 521294 450334
rect 520674 450014 521294 450098
rect 520674 449778 520706 450014
rect 520942 449778 521026 450014
rect 521262 449778 521294 450014
rect 520674 414334 521294 449778
rect 520674 414098 520706 414334
rect 520942 414098 521026 414334
rect 521262 414098 521294 414334
rect 520674 414014 521294 414098
rect 520674 413778 520706 414014
rect 520942 413778 521026 414014
rect 521262 413778 521294 414014
rect 520674 378334 521294 413778
rect 520674 378098 520706 378334
rect 520942 378098 521026 378334
rect 521262 378098 521294 378334
rect 520674 378014 521294 378098
rect 520674 377778 520706 378014
rect 520942 377778 521026 378014
rect 521262 377778 521294 378014
rect 520674 342334 521294 377778
rect 520674 342098 520706 342334
rect 520942 342098 521026 342334
rect 521262 342098 521294 342334
rect 520674 342014 521294 342098
rect 520674 341778 520706 342014
rect 520942 341778 521026 342014
rect 521262 341778 521294 342014
rect 517835 330852 517901 330853
rect 517835 330788 517836 330852
rect 517900 330788 517901 330852
rect 517835 330787 517901 330788
rect 516954 302378 516986 302614
rect 517222 302378 517306 302614
rect 517542 302378 517574 302614
rect 516954 302294 517574 302378
rect 516954 302058 516986 302294
rect 517222 302058 517306 302294
rect 517542 302058 517574 302294
rect 514891 297396 514957 297397
rect 514891 297332 514892 297396
rect 514956 297332 514957 297396
rect 514891 297331 514957 297332
rect 514707 291820 514773 291821
rect 514707 291756 514708 291820
rect 514772 291756 514773 291820
rect 514707 291755 514773 291756
rect 513234 262658 513266 262894
rect 513502 262658 513586 262894
rect 513822 262658 513854 262894
rect 513234 262574 513854 262658
rect 513234 262338 513266 262574
rect 513502 262338 513586 262574
rect 513822 262338 513854 262574
rect 513234 259417 513854 262338
rect 516954 266614 517574 302058
rect 517838 286381 517898 330787
rect 518939 325820 519005 325821
rect 518939 325756 518940 325820
rect 519004 325756 519005 325820
rect 518939 325755 519005 325756
rect 518942 318069 519002 325755
rect 518939 318068 519005 318069
rect 518939 318004 518940 318068
rect 519004 318004 519005 318068
rect 518939 318003 519005 318004
rect 520674 306334 521294 341778
rect 520674 306098 520706 306334
rect 520942 306098 521026 306334
rect 521262 306098 521294 306334
rect 520674 306014 521294 306098
rect 520674 305778 520706 306014
rect 520942 305778 521026 306014
rect 521262 305778 521294 306014
rect 517835 286380 517901 286381
rect 517835 286316 517836 286380
rect 517900 286316 517901 286380
rect 517835 286315 517901 286316
rect 516954 266378 516986 266614
rect 517222 266378 517306 266614
rect 517542 266378 517574 266614
rect 516954 266294 517574 266378
rect 516954 266058 516986 266294
rect 517222 266058 517306 266294
rect 517542 266058 517574 266294
rect 516954 259417 517574 266058
rect 520674 270334 521294 305778
rect 520674 270098 520706 270334
rect 520942 270098 521026 270334
rect 521262 270098 521294 270334
rect 520674 270014 521294 270098
rect 520674 269778 520706 270014
rect 520942 269778 521026 270014
rect 521262 269778 521294 270014
rect 520674 259417 521294 269778
rect 524394 709638 525014 711590
rect 524394 709402 524426 709638
rect 524662 709402 524746 709638
rect 524982 709402 525014 709638
rect 524394 709318 525014 709402
rect 524394 709082 524426 709318
rect 524662 709082 524746 709318
rect 524982 709082 525014 709318
rect 524394 670054 525014 709082
rect 528114 710598 528734 711590
rect 528114 710362 528146 710598
rect 528382 710362 528466 710598
rect 528702 710362 528734 710598
rect 528114 710278 528734 710362
rect 528114 710042 528146 710278
rect 528382 710042 528466 710278
rect 528702 710042 528734 710278
rect 527219 699820 527285 699821
rect 527219 699756 527220 699820
rect 527284 699756 527285 699820
rect 527219 699755 527285 699756
rect 524394 669818 524426 670054
rect 524662 669818 524746 670054
rect 524982 669818 525014 670054
rect 524394 669734 525014 669818
rect 524394 669498 524426 669734
rect 524662 669498 524746 669734
rect 524982 669498 525014 669734
rect 524394 634054 525014 669498
rect 525648 651454 525968 651486
rect 525648 651218 525690 651454
rect 525926 651218 525968 651454
rect 525648 651134 525968 651218
rect 525648 650898 525690 651134
rect 525926 650898 525968 651134
rect 525648 650866 525968 650898
rect 524394 633818 524426 634054
rect 524662 633818 524746 634054
rect 524982 633818 525014 634054
rect 524394 633734 525014 633818
rect 524394 633498 524426 633734
rect 524662 633498 524746 633734
rect 524982 633498 525014 633734
rect 524394 598054 525014 633498
rect 525648 615454 525968 615486
rect 525648 615218 525690 615454
rect 525926 615218 525968 615454
rect 525648 615134 525968 615218
rect 525648 614898 525690 615134
rect 525926 614898 525968 615134
rect 525648 614866 525968 614898
rect 524394 597818 524426 598054
rect 524662 597818 524746 598054
rect 524982 597818 525014 598054
rect 524394 597734 525014 597818
rect 524394 597498 524426 597734
rect 524662 597498 524746 597734
rect 524982 597498 525014 597734
rect 524394 562054 525014 597498
rect 524394 561818 524426 562054
rect 524662 561818 524746 562054
rect 524982 561818 525014 562054
rect 524394 561734 525014 561818
rect 524394 561498 524426 561734
rect 524662 561498 524746 561734
rect 524982 561498 525014 561734
rect 524394 526054 525014 561498
rect 524394 525818 524426 526054
rect 524662 525818 524746 526054
rect 524982 525818 525014 526054
rect 524394 525734 525014 525818
rect 524394 525498 524426 525734
rect 524662 525498 524746 525734
rect 524982 525498 525014 525734
rect 524394 490054 525014 525498
rect 527222 502349 527282 699755
rect 528114 673774 528734 710042
rect 531834 711558 532454 711590
rect 531834 711322 531866 711558
rect 532102 711322 532186 711558
rect 532422 711322 532454 711558
rect 531834 711238 532454 711322
rect 531834 711002 531866 711238
rect 532102 711002 532186 711238
rect 532422 711002 532454 711238
rect 530531 700364 530597 700365
rect 530531 700300 530532 700364
rect 530596 700300 530597 700364
rect 530531 700299 530597 700300
rect 528114 673538 528146 673774
rect 528382 673538 528466 673774
rect 528702 673538 528734 673774
rect 528114 673454 528734 673538
rect 528114 673218 528146 673454
rect 528382 673218 528466 673454
rect 528702 673218 528734 673454
rect 528114 637774 528734 673218
rect 528114 637538 528146 637774
rect 528382 637538 528466 637774
rect 528702 637538 528734 637774
rect 528114 637454 528734 637538
rect 528114 637218 528146 637454
rect 528382 637218 528466 637454
rect 528702 637218 528734 637454
rect 528114 601774 528734 637218
rect 528114 601538 528146 601774
rect 528382 601538 528466 601774
rect 528702 601538 528734 601774
rect 528114 601454 528734 601538
rect 528114 601218 528146 601454
rect 528382 601218 528466 601454
rect 528702 601218 528734 601454
rect 528114 565774 528734 601218
rect 528114 565538 528146 565774
rect 528382 565538 528466 565774
rect 528702 565538 528734 565774
rect 528114 565454 528734 565538
rect 528114 565218 528146 565454
rect 528382 565218 528466 565454
rect 528702 565218 528734 565454
rect 528114 529774 528734 565218
rect 528114 529538 528146 529774
rect 528382 529538 528466 529774
rect 528702 529538 528734 529774
rect 528114 529454 528734 529538
rect 528114 529218 528146 529454
rect 528382 529218 528466 529454
rect 528702 529218 528734 529454
rect 527219 502348 527285 502349
rect 527219 502284 527220 502348
rect 527284 502284 527285 502348
rect 527219 502283 527285 502284
rect 524394 489818 524426 490054
rect 524662 489818 524746 490054
rect 524982 489818 525014 490054
rect 524394 489734 525014 489818
rect 524394 489498 524426 489734
rect 524662 489498 524746 489734
rect 524982 489498 525014 489734
rect 524394 454054 525014 489498
rect 524394 453818 524426 454054
rect 524662 453818 524746 454054
rect 524982 453818 525014 454054
rect 524394 453734 525014 453818
rect 524394 453498 524426 453734
rect 524662 453498 524746 453734
rect 524982 453498 525014 453734
rect 524394 418054 525014 453498
rect 528114 493774 528734 529218
rect 528114 493538 528146 493774
rect 528382 493538 528466 493774
rect 528702 493538 528734 493774
rect 528114 493454 528734 493538
rect 528114 493218 528146 493454
rect 528382 493218 528466 493454
rect 528702 493218 528734 493454
rect 528114 457774 528734 493218
rect 528114 457538 528146 457774
rect 528382 457538 528466 457774
rect 528702 457538 528734 457774
rect 528114 457454 528734 457538
rect 528114 457218 528146 457454
rect 528382 457218 528466 457454
rect 528702 457218 528734 457454
rect 525164 435454 525484 435486
rect 525164 435218 525206 435454
rect 525442 435218 525484 435454
rect 525164 435134 525484 435218
rect 525164 434898 525206 435134
rect 525442 434898 525484 435134
rect 525164 434866 525484 434898
rect 524394 417818 524426 418054
rect 524662 417818 524746 418054
rect 524982 417818 525014 418054
rect 524394 417734 525014 417818
rect 524394 417498 524426 417734
rect 524662 417498 524746 417734
rect 524982 417498 525014 417734
rect 524394 382054 525014 417498
rect 524394 381818 524426 382054
rect 524662 381818 524746 382054
rect 524982 381818 525014 382054
rect 524394 381734 525014 381818
rect 524394 381498 524426 381734
rect 524662 381498 524746 381734
rect 524982 381498 525014 381734
rect 524394 346054 525014 381498
rect 524394 345818 524426 346054
rect 524662 345818 524746 346054
rect 524982 345818 525014 346054
rect 524394 345734 525014 345818
rect 524394 345498 524426 345734
rect 524662 345498 524746 345734
rect 524982 345498 525014 345734
rect 524394 310054 525014 345498
rect 524394 309818 524426 310054
rect 524662 309818 524746 310054
rect 524982 309818 525014 310054
rect 524394 309734 525014 309818
rect 524394 309498 524426 309734
rect 524662 309498 524746 309734
rect 524982 309498 525014 309734
rect 524394 274054 525014 309498
rect 524394 273818 524426 274054
rect 524662 273818 524746 274054
rect 524982 273818 525014 274054
rect 524394 273734 525014 273818
rect 524394 273498 524426 273734
rect 524662 273498 524746 273734
rect 524982 273498 525014 273734
rect 524394 259417 525014 273498
rect 528114 421774 528734 457218
rect 529384 439174 529704 439206
rect 529384 438938 529426 439174
rect 529662 438938 529704 439174
rect 529384 438854 529704 438938
rect 529384 438618 529426 438854
rect 529662 438618 529704 438854
rect 529384 438586 529704 438618
rect 528114 421538 528146 421774
rect 528382 421538 528466 421774
rect 528702 421538 528734 421774
rect 528114 421454 528734 421538
rect 528114 421218 528146 421454
rect 528382 421218 528466 421454
rect 528702 421218 528734 421454
rect 528114 385774 528734 421218
rect 528114 385538 528146 385774
rect 528382 385538 528466 385774
rect 528702 385538 528734 385774
rect 528114 385454 528734 385538
rect 528114 385218 528146 385454
rect 528382 385218 528466 385454
rect 528702 385218 528734 385454
rect 528114 349774 528734 385218
rect 528114 349538 528146 349774
rect 528382 349538 528466 349774
rect 528702 349538 528734 349774
rect 528114 349454 528734 349538
rect 528114 349218 528146 349454
rect 528382 349218 528466 349454
rect 528702 349218 528734 349454
rect 528114 313774 528734 349218
rect 530534 321333 530594 700299
rect 531834 677494 532454 711002
rect 531834 677258 531866 677494
rect 532102 677258 532186 677494
rect 532422 677258 532454 677494
rect 531834 677174 532454 677258
rect 531834 676938 531866 677174
rect 532102 676938 532186 677174
rect 532422 676938 532454 677174
rect 531834 641494 532454 676938
rect 531834 641258 531866 641494
rect 532102 641258 532186 641494
rect 532422 641258 532454 641494
rect 531834 641174 532454 641258
rect 531834 640938 531866 641174
rect 532102 640938 532186 641174
rect 532422 640938 532454 641174
rect 531834 605494 532454 640938
rect 531834 605258 531866 605494
rect 532102 605258 532186 605494
rect 532422 605258 532454 605494
rect 531834 605174 532454 605258
rect 531834 604938 531866 605174
rect 532102 604938 532186 605174
rect 532422 604938 532454 605174
rect 531834 569494 532454 604938
rect 531834 569258 531866 569494
rect 532102 569258 532186 569494
rect 532422 569258 532454 569494
rect 531834 569174 532454 569258
rect 531834 568938 531866 569174
rect 532102 568938 532186 569174
rect 532422 568938 532454 569174
rect 531834 533494 532454 568938
rect 531834 533258 531866 533494
rect 532102 533258 532186 533494
rect 532422 533258 532454 533494
rect 531834 533174 532454 533258
rect 531834 532938 531866 533174
rect 532102 532938 532186 533174
rect 532422 532938 532454 533174
rect 531834 497494 532454 532938
rect 531834 497258 531866 497494
rect 532102 497258 532186 497494
rect 532422 497258 532454 497494
rect 531834 497174 532454 497258
rect 531834 496938 531866 497174
rect 532102 496938 532186 497174
rect 532422 496938 532454 497174
rect 531834 461494 532454 496938
rect 531834 461258 531866 461494
rect 532102 461258 532186 461494
rect 532422 461258 532454 461494
rect 531834 461174 532454 461258
rect 531834 460938 531866 461174
rect 532102 460938 532186 461174
rect 532422 460938 532454 461174
rect 531834 425494 532454 460938
rect 541794 704838 542414 711590
rect 541794 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 542414 704838
rect 541794 704518 542414 704602
rect 541794 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 542414 704518
rect 541794 687454 542414 704282
rect 541794 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 542414 687454
rect 541794 687134 542414 687218
rect 541794 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 542414 687134
rect 541794 651454 542414 686898
rect 541794 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 542414 651454
rect 541794 651134 542414 651218
rect 541794 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 542414 651134
rect 541794 615454 542414 650898
rect 541794 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 542414 615454
rect 541794 615134 542414 615218
rect 541794 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 542414 615134
rect 541794 579454 542414 614898
rect 541794 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 542414 579454
rect 541794 579134 542414 579218
rect 541794 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 542414 579134
rect 541794 543454 542414 578898
rect 541794 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 542414 543454
rect 541794 543134 542414 543218
rect 541794 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 542414 543134
rect 541794 507454 542414 542898
rect 541794 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 542414 507454
rect 541794 507134 542414 507218
rect 541794 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 542414 507134
rect 541794 471454 542414 506898
rect 541794 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 542414 471454
rect 541794 471134 542414 471218
rect 541794 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 542414 471134
rect 541794 460836 542414 470898
rect 545514 705798 546134 711590
rect 545514 705562 545546 705798
rect 545782 705562 545866 705798
rect 546102 705562 546134 705798
rect 545514 705478 546134 705562
rect 545514 705242 545546 705478
rect 545782 705242 545866 705478
rect 546102 705242 546134 705478
rect 545514 691174 546134 705242
rect 545514 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 546134 691174
rect 545514 690854 546134 690938
rect 545514 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 546134 690854
rect 545514 655174 546134 690618
rect 545514 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 546134 655174
rect 545514 654854 546134 654938
rect 545514 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 546134 654854
rect 545514 619174 546134 654618
rect 545514 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 546134 619174
rect 545514 618854 546134 618938
rect 545514 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 546134 618854
rect 545514 583174 546134 618618
rect 545514 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 546134 583174
rect 545514 582854 546134 582938
rect 545514 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 546134 582854
rect 545514 547174 546134 582618
rect 545514 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 546134 547174
rect 545514 546854 546134 546938
rect 545514 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 546134 546854
rect 545514 511174 546134 546618
rect 545514 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 546134 511174
rect 545514 510854 546134 510938
rect 545514 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 546134 510854
rect 545514 475174 546134 510618
rect 545514 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 546134 475174
rect 545514 474854 546134 474938
rect 545514 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 546134 474854
rect 537825 439174 538145 439206
rect 537825 438938 537867 439174
rect 538103 438938 538145 439174
rect 537825 438854 538145 438938
rect 537825 438618 537867 438854
rect 538103 438618 538145 438854
rect 537825 438586 538145 438618
rect 545514 439174 546134 474618
rect 549234 706758 549854 711590
rect 549234 706522 549266 706758
rect 549502 706522 549586 706758
rect 549822 706522 549854 706758
rect 549234 706438 549854 706522
rect 549234 706202 549266 706438
rect 549502 706202 549586 706438
rect 549822 706202 549854 706438
rect 549234 694894 549854 706202
rect 549234 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 549854 694894
rect 549234 694574 549854 694658
rect 549234 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 549854 694574
rect 549234 658894 549854 694338
rect 549234 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 549854 658894
rect 549234 658574 549854 658658
rect 549234 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 549854 658574
rect 549234 622894 549854 658338
rect 549234 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 549854 622894
rect 549234 622574 549854 622658
rect 549234 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 549854 622574
rect 549234 586894 549854 622338
rect 549234 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 549854 586894
rect 549234 586574 549854 586658
rect 549234 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 549854 586574
rect 549234 550894 549854 586338
rect 549234 550658 549266 550894
rect 549502 550658 549586 550894
rect 549822 550658 549854 550894
rect 549234 550574 549854 550658
rect 549234 550338 549266 550574
rect 549502 550338 549586 550574
rect 549822 550338 549854 550574
rect 549234 514894 549854 550338
rect 549234 514658 549266 514894
rect 549502 514658 549586 514894
rect 549822 514658 549854 514894
rect 549234 514574 549854 514658
rect 549234 514338 549266 514574
rect 549502 514338 549586 514574
rect 549822 514338 549854 514574
rect 549234 478894 549854 514338
rect 549234 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 549854 478894
rect 549234 478574 549854 478658
rect 549234 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 549854 478574
rect 549234 442894 549854 478338
rect 549234 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 549854 442894
rect 549234 442574 549854 442658
rect 549234 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 549854 442574
rect 545514 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 546134 439174
rect 545514 438854 546134 438938
rect 545514 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 546134 438854
rect 533605 435454 533925 435486
rect 533605 435218 533647 435454
rect 533883 435218 533925 435454
rect 533605 435134 533925 435218
rect 533605 434898 533647 435134
rect 533883 434898 533925 435134
rect 533605 434866 533925 434898
rect 542046 435454 542366 435486
rect 542046 435218 542088 435454
rect 542324 435218 542366 435454
rect 542046 435134 542366 435218
rect 542046 434898 542088 435134
rect 542324 434898 542366 435134
rect 542046 434866 542366 434898
rect 531834 425258 531866 425494
rect 532102 425258 532186 425494
rect 532422 425258 532454 425494
rect 531834 425174 532454 425258
rect 531834 424938 531866 425174
rect 532102 424938 532186 425174
rect 532422 424938 532454 425174
rect 531834 389494 532454 424938
rect 531834 389258 531866 389494
rect 532102 389258 532186 389494
rect 532422 389258 532454 389494
rect 531834 389174 532454 389258
rect 531834 388938 531866 389174
rect 532102 388938 532186 389174
rect 532422 388938 532454 389174
rect 531834 353494 532454 388938
rect 531834 353258 531866 353494
rect 532102 353258 532186 353494
rect 532422 353258 532454 353494
rect 531834 353174 532454 353258
rect 531834 352938 531866 353174
rect 532102 352938 532186 353174
rect 532422 352938 532454 353174
rect 530531 321332 530597 321333
rect 530531 321268 530532 321332
rect 530596 321268 530597 321332
rect 530531 321267 530597 321268
rect 528114 313538 528146 313774
rect 528382 313538 528466 313774
rect 528702 313538 528734 313774
rect 528114 313454 528734 313538
rect 528114 313218 528146 313454
rect 528382 313218 528466 313454
rect 528702 313218 528734 313454
rect 528114 277774 528734 313218
rect 528114 277538 528146 277774
rect 528382 277538 528466 277774
rect 528702 277538 528734 277774
rect 528114 277454 528734 277538
rect 528114 277218 528146 277454
rect 528382 277218 528466 277454
rect 528702 277218 528734 277454
rect 528114 259417 528734 277218
rect 531834 317494 532454 352938
rect 531834 317258 531866 317494
rect 532102 317258 532186 317494
rect 532422 317258 532454 317494
rect 531834 317174 532454 317258
rect 531834 316938 531866 317174
rect 532102 316938 532186 317174
rect 532422 316938 532454 317174
rect 531834 281494 532454 316938
rect 541794 399454 542414 425068
rect 541794 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 542414 399454
rect 541794 399134 542414 399218
rect 541794 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 542414 399134
rect 541794 363454 542414 398898
rect 541794 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 542414 363454
rect 541794 363134 542414 363218
rect 541794 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 542414 363134
rect 541794 327454 542414 362898
rect 541794 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 542414 327454
rect 541794 327134 542414 327218
rect 541794 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 542414 327134
rect 538443 315348 538509 315349
rect 538443 315284 538444 315348
rect 538508 315284 538509 315348
rect 538443 315283 538509 315284
rect 538259 313988 538325 313989
rect 538259 313924 538260 313988
rect 538324 313924 538325 313988
rect 538259 313923 538325 313924
rect 531834 281258 531866 281494
rect 532102 281258 532186 281494
rect 532422 281258 532454 281494
rect 531834 281174 532454 281258
rect 531834 280938 531866 281174
rect 532102 280938 532186 281174
rect 532422 280938 532454 281174
rect 479568 259174 479888 259206
rect 479568 258938 479610 259174
rect 479846 258938 479888 259174
rect 479568 258854 479888 258938
rect 479568 258618 479610 258854
rect 479846 258618 479888 258854
rect 479568 258586 479888 258618
rect 510288 259174 510608 259206
rect 510288 258938 510330 259174
rect 510566 258938 510608 259174
rect 510288 258854 510608 258938
rect 510288 258618 510330 258854
rect 510566 258618 510608 258854
rect 510288 258586 510608 258618
rect 464208 255454 464528 255486
rect 464208 255218 464250 255454
rect 464486 255218 464528 255454
rect 464208 255134 464528 255218
rect 464208 254898 464250 255134
rect 464486 254898 464528 255134
rect 464208 254866 464528 254898
rect 494928 255454 495248 255486
rect 494928 255218 494970 255454
rect 495206 255218 495248 255454
rect 494928 255134 495248 255218
rect 494928 254898 494970 255134
rect 495206 254898 495248 255134
rect 494928 254866 495248 254898
rect 525648 255454 525968 255486
rect 525648 255218 525690 255454
rect 525926 255218 525968 255454
rect 525648 255134 525968 255218
rect 525648 254898 525690 255134
rect 525926 254898 525968 255134
rect 525648 254866 525968 254898
rect 531834 245494 532454 280938
rect 531834 245258 531866 245494
rect 532102 245258 532186 245494
rect 532422 245258 532454 245494
rect 531834 245174 532454 245258
rect 531834 244938 531866 245174
rect 532102 244938 532186 245174
rect 532422 244938 532454 245174
rect 479568 223174 479888 223206
rect 479568 222938 479610 223174
rect 479846 222938 479888 223174
rect 479568 222854 479888 222938
rect 479568 222618 479610 222854
rect 479846 222618 479888 222854
rect 479568 222586 479888 222618
rect 510288 223174 510608 223206
rect 510288 222938 510330 223174
rect 510566 222938 510608 223174
rect 510288 222854 510608 222938
rect 510288 222618 510330 222854
rect 510566 222618 510608 222854
rect 510288 222586 510608 222618
rect 464208 219454 464528 219486
rect 464208 219218 464250 219454
rect 464486 219218 464528 219454
rect 464208 219134 464528 219218
rect 464208 218898 464250 219134
rect 464486 218898 464528 219134
rect 464208 218866 464528 218898
rect 494928 219454 495248 219486
rect 494928 219218 494970 219454
rect 495206 219218 495248 219454
rect 494928 219134 495248 219218
rect 494928 218898 494970 219134
rect 495206 218898 495248 219134
rect 494928 218866 495248 218898
rect 525648 219454 525968 219486
rect 525648 219218 525690 219454
rect 525926 219218 525968 219454
rect 525648 219134 525968 219218
rect 525648 218898 525690 219134
rect 525926 218898 525968 219134
rect 525648 218866 525968 218898
rect 531834 209494 532454 244938
rect 531834 209258 531866 209494
rect 532102 209258 532186 209494
rect 532422 209258 532454 209494
rect 531834 209174 532454 209258
rect 531834 208938 531866 209174
rect 532102 208938 532186 209174
rect 532422 208938 532454 209174
rect 469794 183454 470414 201919
rect 469794 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 470414 183454
rect 469794 183134 470414 183218
rect 469794 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 470414 183134
rect 469794 147454 470414 182898
rect 469794 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 470414 147454
rect 469794 147134 470414 147218
rect 469794 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 470414 147134
rect 469794 111454 470414 146898
rect 469794 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 470414 111454
rect 469794 111134 470414 111218
rect 469794 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 470414 111134
rect 469794 75454 470414 110898
rect 469794 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 470414 75454
rect 469794 75134 470414 75218
rect 469794 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 470414 75134
rect 469794 39454 470414 74898
rect 469794 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 470414 39454
rect 469794 39134 470414 39218
rect 469794 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 470414 39134
rect 469794 3454 470414 38898
rect 460795 3364 460861 3365
rect 460795 3300 460796 3364
rect 460860 3300 460861 3364
rect 460795 3299 460861 3300
rect 459834 -7302 459866 -7066
rect 460102 -7302 460186 -7066
rect 460422 -7302 460454 -7066
rect 459834 -7386 460454 -7302
rect 459834 -7622 459866 -7386
rect 460102 -7622 460186 -7386
rect 460422 -7622 460454 -7386
rect 459834 -7654 460454 -7622
rect 469794 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 470414 3454
rect 469794 3134 470414 3218
rect 469794 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 470414 3134
rect 469794 -346 470414 2898
rect 469794 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 470414 -346
rect 469794 -666 470414 -582
rect 469794 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 470414 -666
rect 469794 -7654 470414 -902
rect 473514 187174 474134 201919
rect 473514 186938 473546 187174
rect 473782 186938 473866 187174
rect 474102 186938 474134 187174
rect 473514 186854 474134 186938
rect 473514 186618 473546 186854
rect 473782 186618 473866 186854
rect 474102 186618 474134 186854
rect 473514 151174 474134 186618
rect 473514 150938 473546 151174
rect 473782 150938 473866 151174
rect 474102 150938 474134 151174
rect 473514 150854 474134 150938
rect 473514 150618 473546 150854
rect 473782 150618 473866 150854
rect 474102 150618 474134 150854
rect 473514 115174 474134 150618
rect 473514 114938 473546 115174
rect 473782 114938 473866 115174
rect 474102 114938 474134 115174
rect 473514 114854 474134 114938
rect 473514 114618 473546 114854
rect 473782 114618 473866 114854
rect 474102 114618 474134 114854
rect 473514 79174 474134 114618
rect 473514 78938 473546 79174
rect 473782 78938 473866 79174
rect 474102 78938 474134 79174
rect 473514 78854 474134 78938
rect 473514 78618 473546 78854
rect 473782 78618 473866 78854
rect 474102 78618 474134 78854
rect 473514 43174 474134 78618
rect 473514 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 474134 43174
rect 473514 42854 474134 42938
rect 473514 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 474134 42854
rect 473514 7174 474134 42618
rect 473514 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 474134 7174
rect 473514 6854 474134 6938
rect 473514 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 474134 6854
rect 473514 -1306 474134 6618
rect 473514 -1542 473546 -1306
rect 473782 -1542 473866 -1306
rect 474102 -1542 474134 -1306
rect 473514 -1626 474134 -1542
rect 473514 -1862 473546 -1626
rect 473782 -1862 473866 -1626
rect 474102 -1862 474134 -1626
rect 473514 -7654 474134 -1862
rect 477234 190894 477854 201919
rect 477234 190658 477266 190894
rect 477502 190658 477586 190894
rect 477822 190658 477854 190894
rect 477234 190574 477854 190658
rect 477234 190338 477266 190574
rect 477502 190338 477586 190574
rect 477822 190338 477854 190574
rect 477234 154894 477854 190338
rect 477234 154658 477266 154894
rect 477502 154658 477586 154894
rect 477822 154658 477854 154894
rect 477234 154574 477854 154658
rect 477234 154338 477266 154574
rect 477502 154338 477586 154574
rect 477822 154338 477854 154574
rect 477234 118894 477854 154338
rect 477234 118658 477266 118894
rect 477502 118658 477586 118894
rect 477822 118658 477854 118894
rect 477234 118574 477854 118658
rect 477234 118338 477266 118574
rect 477502 118338 477586 118574
rect 477822 118338 477854 118574
rect 477234 82894 477854 118338
rect 477234 82658 477266 82894
rect 477502 82658 477586 82894
rect 477822 82658 477854 82894
rect 477234 82574 477854 82658
rect 477234 82338 477266 82574
rect 477502 82338 477586 82574
rect 477822 82338 477854 82574
rect 477234 46894 477854 82338
rect 477234 46658 477266 46894
rect 477502 46658 477586 46894
rect 477822 46658 477854 46894
rect 477234 46574 477854 46658
rect 477234 46338 477266 46574
rect 477502 46338 477586 46574
rect 477822 46338 477854 46574
rect 477234 10894 477854 46338
rect 477234 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 477854 10894
rect 477234 10574 477854 10658
rect 477234 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 477854 10574
rect 477234 -2266 477854 10338
rect 477234 -2502 477266 -2266
rect 477502 -2502 477586 -2266
rect 477822 -2502 477854 -2266
rect 477234 -2586 477854 -2502
rect 477234 -2822 477266 -2586
rect 477502 -2822 477586 -2586
rect 477822 -2822 477854 -2586
rect 477234 -7654 477854 -2822
rect 480954 194614 481574 201919
rect 480954 194378 480986 194614
rect 481222 194378 481306 194614
rect 481542 194378 481574 194614
rect 480954 194294 481574 194378
rect 480954 194058 480986 194294
rect 481222 194058 481306 194294
rect 481542 194058 481574 194294
rect 480954 158614 481574 194058
rect 480954 158378 480986 158614
rect 481222 158378 481306 158614
rect 481542 158378 481574 158614
rect 480954 158294 481574 158378
rect 480954 158058 480986 158294
rect 481222 158058 481306 158294
rect 481542 158058 481574 158294
rect 480954 122614 481574 158058
rect 480954 122378 480986 122614
rect 481222 122378 481306 122614
rect 481542 122378 481574 122614
rect 480954 122294 481574 122378
rect 480954 122058 480986 122294
rect 481222 122058 481306 122294
rect 481542 122058 481574 122294
rect 480954 86614 481574 122058
rect 484674 198334 485294 201919
rect 484674 198098 484706 198334
rect 484942 198098 485026 198334
rect 485262 198098 485294 198334
rect 484674 198014 485294 198098
rect 484674 197778 484706 198014
rect 484942 197778 485026 198014
rect 485262 197778 485294 198014
rect 484674 162334 485294 197778
rect 484674 162098 484706 162334
rect 484942 162098 485026 162334
rect 485262 162098 485294 162334
rect 484674 162014 485294 162098
rect 484674 161778 484706 162014
rect 484942 161778 485026 162014
rect 485262 161778 485294 162014
rect 484674 126334 485294 161778
rect 488394 166054 489014 201919
rect 488394 165818 488426 166054
rect 488662 165818 488746 166054
rect 488982 165818 489014 166054
rect 488394 165734 489014 165818
rect 488394 165498 488426 165734
rect 488662 165498 488746 165734
rect 488982 165498 489014 165734
rect 488394 139281 489014 165498
rect 505794 183454 506414 201919
rect 505794 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 506414 183454
rect 505794 183134 506414 183218
rect 505794 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 506414 183134
rect 505794 147454 506414 182898
rect 505794 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 506414 147454
rect 505794 147134 506414 147218
rect 505794 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 506414 147134
rect 505794 139281 506414 146898
rect 509514 187174 510134 201919
rect 509514 186938 509546 187174
rect 509782 186938 509866 187174
rect 510102 186938 510134 187174
rect 509514 186854 510134 186938
rect 509514 186618 509546 186854
rect 509782 186618 509866 186854
rect 510102 186618 510134 186854
rect 509514 151174 510134 186618
rect 509514 150938 509546 151174
rect 509782 150938 509866 151174
rect 510102 150938 510134 151174
rect 509514 150854 510134 150938
rect 509514 150618 509546 150854
rect 509782 150618 509866 150854
rect 510102 150618 510134 150854
rect 509514 139281 510134 150618
rect 513234 190894 513854 201919
rect 513234 190658 513266 190894
rect 513502 190658 513586 190894
rect 513822 190658 513854 190894
rect 513234 190574 513854 190658
rect 513234 190338 513266 190574
rect 513502 190338 513586 190574
rect 513822 190338 513854 190574
rect 513234 154894 513854 190338
rect 513234 154658 513266 154894
rect 513502 154658 513586 154894
rect 513822 154658 513854 154894
rect 513234 154574 513854 154658
rect 513234 154338 513266 154574
rect 513502 154338 513586 154574
rect 513822 154338 513854 154574
rect 513234 139281 513854 154338
rect 516954 194614 517574 201919
rect 516954 194378 516986 194614
rect 517222 194378 517306 194614
rect 517542 194378 517574 194614
rect 516954 194294 517574 194378
rect 516954 194058 516986 194294
rect 517222 194058 517306 194294
rect 517542 194058 517574 194294
rect 516954 158614 517574 194058
rect 516954 158378 516986 158614
rect 517222 158378 517306 158614
rect 517542 158378 517574 158614
rect 516954 158294 517574 158378
rect 516954 158058 516986 158294
rect 517222 158058 517306 158294
rect 517542 158058 517574 158294
rect 516954 139281 517574 158058
rect 520674 198334 521294 201919
rect 520674 198098 520706 198334
rect 520942 198098 521026 198334
rect 521262 198098 521294 198334
rect 520674 198014 521294 198098
rect 520674 197778 520706 198014
rect 520942 197778 521026 198014
rect 521262 197778 521294 198014
rect 520674 162334 521294 197778
rect 520674 162098 520706 162334
rect 520942 162098 521026 162334
rect 521262 162098 521294 162334
rect 520674 162014 521294 162098
rect 520674 161778 520706 162014
rect 520942 161778 521026 162014
rect 521262 161778 521294 162014
rect 520674 139281 521294 161778
rect 524394 166054 525014 201919
rect 524394 165818 524426 166054
rect 524662 165818 524746 166054
rect 524982 165818 525014 166054
rect 524394 165734 525014 165818
rect 524394 165498 524426 165734
rect 524662 165498 524746 165734
rect 524982 165498 525014 165734
rect 524394 139281 525014 165498
rect 531834 173494 532454 208938
rect 531834 173258 531866 173494
rect 532102 173258 532186 173494
rect 532422 173258 532454 173494
rect 531834 173174 532454 173258
rect 531834 172938 531866 173174
rect 532102 172938 532186 173174
rect 532422 172938 532454 173174
rect 531834 139281 532454 172938
rect 538262 137730 538322 313923
rect 538446 137869 538506 315283
rect 541794 291454 542414 326898
rect 541794 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 542414 291454
rect 541794 291134 542414 291218
rect 541794 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 542414 291134
rect 541794 255454 542414 290898
rect 541794 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 542414 255454
rect 541794 255134 542414 255218
rect 541794 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 542414 255134
rect 541794 219454 542414 254898
rect 541794 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 542414 219454
rect 541794 219134 542414 219218
rect 541794 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 542414 219134
rect 541794 183454 542414 218898
rect 541794 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 542414 183454
rect 541794 183134 542414 183218
rect 541794 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 542414 183134
rect 541794 147454 542414 182898
rect 541794 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 542414 147454
rect 541794 147134 542414 147218
rect 541794 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 542414 147134
rect 538443 137868 538509 137869
rect 538443 137804 538444 137868
rect 538508 137804 538509 137868
rect 538443 137803 538509 137804
rect 538262 137670 539426 137730
rect 539366 133381 539426 137670
rect 539363 133380 539429 133381
rect 539363 133316 539364 133380
rect 539428 133316 539429 133380
rect 539363 133315 539429 133316
rect 484674 126098 484706 126334
rect 484942 126098 485026 126334
rect 485262 126098 485294 126334
rect 484674 126014 485294 126098
rect 484674 125778 484706 126014
rect 484942 125778 485026 126014
rect 485262 125778 485294 126014
rect 484208 111454 484528 111486
rect 484208 111218 484250 111454
rect 484486 111218 484528 111454
rect 484208 111134 484528 111218
rect 484208 110898 484250 111134
rect 484486 110898 484528 111134
rect 484208 110866 484528 110898
rect 480954 86378 480986 86614
rect 481222 86378 481306 86614
rect 481542 86378 481574 86614
rect 480954 86294 481574 86378
rect 480954 86058 480986 86294
rect 481222 86058 481306 86294
rect 481542 86058 481574 86294
rect 480954 50614 481574 86058
rect 480954 50378 480986 50614
rect 481222 50378 481306 50614
rect 481542 50378 481574 50614
rect 480954 50294 481574 50378
rect 480954 50058 480986 50294
rect 481222 50058 481306 50294
rect 481542 50058 481574 50294
rect 480954 14614 481574 50058
rect 480954 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 481574 14614
rect 480954 14294 481574 14378
rect 480954 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 481574 14294
rect 480954 -3226 481574 14058
rect 480954 -3462 480986 -3226
rect 481222 -3462 481306 -3226
rect 481542 -3462 481574 -3226
rect 480954 -3546 481574 -3462
rect 480954 -3782 480986 -3546
rect 481222 -3782 481306 -3546
rect 481542 -3782 481574 -3546
rect 480954 -7654 481574 -3782
rect 484674 90334 485294 125778
rect 499568 115174 499888 115206
rect 499568 114938 499610 115174
rect 499846 114938 499888 115174
rect 499568 114854 499888 114938
rect 499568 114618 499610 114854
rect 499846 114618 499888 114854
rect 499568 114586 499888 114618
rect 530288 115174 530608 115206
rect 530288 114938 530330 115174
rect 530566 114938 530608 115174
rect 530288 114854 530608 114938
rect 530288 114618 530330 114854
rect 530566 114618 530608 114854
rect 530288 114586 530608 114618
rect 514928 111454 515248 111486
rect 514928 111218 514970 111454
rect 515206 111218 515248 111454
rect 514928 111134 515248 111218
rect 514928 110898 514970 111134
rect 515206 110898 515248 111134
rect 514928 110866 515248 110898
rect 541794 111454 542414 146898
rect 541794 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 542414 111454
rect 541794 111134 542414 111218
rect 541794 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 542414 111134
rect 484674 90098 484706 90334
rect 484942 90098 485026 90334
rect 485262 90098 485294 90334
rect 484674 90014 485294 90098
rect 484674 89778 484706 90014
rect 484942 89778 485026 90014
rect 485262 89778 485294 90014
rect 484674 54334 485294 89778
rect 484674 54098 484706 54334
rect 484942 54098 485026 54334
rect 485262 54098 485294 54334
rect 484674 54014 485294 54098
rect 484674 53778 484706 54014
rect 484942 53778 485026 54014
rect 485262 53778 485294 54014
rect 484674 18334 485294 53778
rect 484674 18098 484706 18334
rect 484942 18098 485026 18334
rect 485262 18098 485294 18334
rect 484674 18014 485294 18098
rect 484674 17778 484706 18014
rect 484942 17778 485026 18014
rect 485262 17778 485294 18014
rect 484674 -4186 485294 17778
rect 484674 -4422 484706 -4186
rect 484942 -4422 485026 -4186
rect 485262 -4422 485294 -4186
rect 484674 -4506 485294 -4422
rect 484674 -4742 484706 -4506
rect 484942 -4742 485026 -4506
rect 485262 -4742 485294 -4506
rect 484674 -7654 485294 -4742
rect 488394 58054 489014 82599
rect 488394 57818 488426 58054
rect 488662 57818 488746 58054
rect 488982 57818 489014 58054
rect 488394 57734 489014 57818
rect 488394 57498 488426 57734
rect 488662 57498 488746 57734
rect 488982 57498 489014 57734
rect 488394 22054 489014 57498
rect 488394 21818 488426 22054
rect 488662 21818 488746 22054
rect 488982 21818 489014 22054
rect 488394 21734 489014 21818
rect 488394 21498 488426 21734
rect 488662 21498 488746 21734
rect 488982 21498 489014 21734
rect 488394 -5146 489014 21498
rect 488394 -5382 488426 -5146
rect 488662 -5382 488746 -5146
rect 488982 -5382 489014 -5146
rect 488394 -5466 489014 -5382
rect 488394 -5702 488426 -5466
rect 488662 -5702 488746 -5466
rect 488982 -5702 489014 -5466
rect 488394 -7654 489014 -5702
rect 492114 61774 492734 82599
rect 492114 61538 492146 61774
rect 492382 61538 492466 61774
rect 492702 61538 492734 61774
rect 492114 61454 492734 61538
rect 492114 61218 492146 61454
rect 492382 61218 492466 61454
rect 492702 61218 492734 61454
rect 492114 25774 492734 61218
rect 492114 25538 492146 25774
rect 492382 25538 492466 25774
rect 492702 25538 492734 25774
rect 492114 25454 492734 25538
rect 492114 25218 492146 25454
rect 492382 25218 492466 25454
rect 492702 25218 492734 25454
rect 492114 -6106 492734 25218
rect 492114 -6342 492146 -6106
rect 492382 -6342 492466 -6106
rect 492702 -6342 492734 -6106
rect 492114 -6426 492734 -6342
rect 492114 -6662 492146 -6426
rect 492382 -6662 492466 -6426
rect 492702 -6662 492734 -6426
rect 492114 -7654 492734 -6662
rect 495834 65494 496454 82599
rect 495834 65258 495866 65494
rect 496102 65258 496186 65494
rect 496422 65258 496454 65494
rect 495834 65174 496454 65258
rect 495834 64938 495866 65174
rect 496102 64938 496186 65174
rect 496422 64938 496454 65174
rect 495834 29494 496454 64938
rect 495834 29258 495866 29494
rect 496102 29258 496186 29494
rect 496422 29258 496454 29494
rect 495834 29174 496454 29258
rect 495834 28938 495866 29174
rect 496102 28938 496186 29174
rect 496422 28938 496454 29174
rect 495834 -7066 496454 28938
rect 495834 -7302 495866 -7066
rect 496102 -7302 496186 -7066
rect 496422 -7302 496454 -7066
rect 495834 -7386 496454 -7302
rect 495834 -7622 495866 -7386
rect 496102 -7622 496186 -7386
rect 496422 -7622 496454 -7386
rect 495834 -7654 496454 -7622
rect 505794 75454 506414 82599
rect 505794 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 506414 75454
rect 505794 75134 506414 75218
rect 505794 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 506414 75134
rect 505794 39454 506414 74898
rect 505794 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 506414 39454
rect 505794 39134 506414 39218
rect 505794 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 506414 39134
rect 505794 3454 506414 38898
rect 505794 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 506414 3454
rect 505794 3134 506414 3218
rect 505794 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 506414 3134
rect 505794 -346 506414 2898
rect 505794 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 506414 -346
rect 505794 -666 506414 -582
rect 505794 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 506414 -666
rect 505794 -7654 506414 -902
rect 509514 79174 510134 82599
rect 509514 78938 509546 79174
rect 509782 78938 509866 79174
rect 510102 78938 510134 79174
rect 509514 78854 510134 78938
rect 509514 78618 509546 78854
rect 509782 78618 509866 78854
rect 510102 78618 510134 78854
rect 509514 43174 510134 78618
rect 509514 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 510134 43174
rect 509514 42854 510134 42938
rect 509514 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 510134 42854
rect 509514 7174 510134 42618
rect 509514 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 510134 7174
rect 509514 6854 510134 6938
rect 509514 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 510134 6854
rect 509514 -1306 510134 6618
rect 509514 -1542 509546 -1306
rect 509782 -1542 509866 -1306
rect 510102 -1542 510134 -1306
rect 509514 -1626 510134 -1542
rect 509514 -1862 509546 -1626
rect 509782 -1862 509866 -1626
rect 510102 -1862 510134 -1626
rect 509514 -7654 510134 -1862
rect 513234 46894 513854 82599
rect 513234 46658 513266 46894
rect 513502 46658 513586 46894
rect 513822 46658 513854 46894
rect 513234 46574 513854 46658
rect 513234 46338 513266 46574
rect 513502 46338 513586 46574
rect 513822 46338 513854 46574
rect 513234 10894 513854 46338
rect 513234 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 513854 10894
rect 513234 10574 513854 10658
rect 513234 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 513854 10574
rect 513234 -2266 513854 10338
rect 513234 -2502 513266 -2266
rect 513502 -2502 513586 -2266
rect 513822 -2502 513854 -2266
rect 513234 -2586 513854 -2502
rect 513234 -2822 513266 -2586
rect 513502 -2822 513586 -2586
rect 513822 -2822 513854 -2586
rect 513234 -7654 513854 -2822
rect 516954 50614 517574 82599
rect 516954 50378 516986 50614
rect 517222 50378 517306 50614
rect 517542 50378 517574 50614
rect 516954 50294 517574 50378
rect 516954 50058 516986 50294
rect 517222 50058 517306 50294
rect 517542 50058 517574 50294
rect 516954 14614 517574 50058
rect 516954 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 517574 14614
rect 516954 14294 517574 14378
rect 516954 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 517574 14294
rect 516954 -3226 517574 14058
rect 516954 -3462 516986 -3226
rect 517222 -3462 517306 -3226
rect 517542 -3462 517574 -3226
rect 516954 -3546 517574 -3462
rect 516954 -3782 516986 -3546
rect 517222 -3782 517306 -3546
rect 517542 -3782 517574 -3546
rect 516954 -7654 517574 -3782
rect 520674 54334 521294 82599
rect 520674 54098 520706 54334
rect 520942 54098 521026 54334
rect 521262 54098 521294 54334
rect 520674 54014 521294 54098
rect 520674 53778 520706 54014
rect 520942 53778 521026 54014
rect 521262 53778 521294 54014
rect 520674 18334 521294 53778
rect 520674 18098 520706 18334
rect 520942 18098 521026 18334
rect 521262 18098 521294 18334
rect 520674 18014 521294 18098
rect 520674 17778 520706 18014
rect 520942 17778 521026 18014
rect 521262 17778 521294 18014
rect 520674 -4186 521294 17778
rect 520674 -4422 520706 -4186
rect 520942 -4422 521026 -4186
rect 521262 -4422 521294 -4186
rect 520674 -4506 521294 -4422
rect 520674 -4742 520706 -4506
rect 520942 -4742 521026 -4506
rect 521262 -4742 521294 -4506
rect 520674 -7654 521294 -4742
rect 524394 58054 525014 82599
rect 524394 57818 524426 58054
rect 524662 57818 524746 58054
rect 524982 57818 525014 58054
rect 524394 57734 525014 57818
rect 524394 57498 524426 57734
rect 524662 57498 524746 57734
rect 524982 57498 525014 57734
rect 524394 22054 525014 57498
rect 524394 21818 524426 22054
rect 524662 21818 524746 22054
rect 524982 21818 525014 22054
rect 524394 21734 525014 21818
rect 524394 21498 524426 21734
rect 524662 21498 524746 21734
rect 524982 21498 525014 21734
rect 524394 -5146 525014 21498
rect 524394 -5382 524426 -5146
rect 524662 -5382 524746 -5146
rect 524982 -5382 525014 -5146
rect 524394 -5466 525014 -5382
rect 524394 -5702 524426 -5466
rect 524662 -5702 524746 -5466
rect 524982 -5702 525014 -5466
rect 524394 -7654 525014 -5702
rect 528114 61774 528734 82599
rect 528114 61538 528146 61774
rect 528382 61538 528466 61774
rect 528702 61538 528734 61774
rect 528114 61454 528734 61538
rect 528114 61218 528146 61454
rect 528382 61218 528466 61454
rect 528702 61218 528734 61454
rect 528114 25774 528734 61218
rect 528114 25538 528146 25774
rect 528382 25538 528466 25774
rect 528702 25538 528734 25774
rect 528114 25454 528734 25538
rect 528114 25218 528146 25454
rect 528382 25218 528466 25454
rect 528702 25218 528734 25454
rect 528114 -6106 528734 25218
rect 528114 -6342 528146 -6106
rect 528382 -6342 528466 -6106
rect 528702 -6342 528734 -6106
rect 528114 -6426 528734 -6342
rect 528114 -6662 528146 -6426
rect 528382 -6662 528466 -6426
rect 528702 -6662 528734 -6426
rect 528114 -7654 528734 -6662
rect 531834 65494 532454 82599
rect 531834 65258 531866 65494
rect 532102 65258 532186 65494
rect 532422 65258 532454 65494
rect 531834 65174 532454 65258
rect 531834 64938 531866 65174
rect 532102 64938 532186 65174
rect 532422 64938 532454 65174
rect 531834 29494 532454 64938
rect 531834 29258 531866 29494
rect 532102 29258 532186 29494
rect 532422 29258 532454 29494
rect 531834 29174 532454 29258
rect 531834 28938 531866 29174
rect 532102 28938 532186 29174
rect 532422 28938 532454 29174
rect 531834 -7066 532454 28938
rect 531834 -7302 531866 -7066
rect 532102 -7302 532186 -7066
rect 532422 -7302 532454 -7066
rect 531834 -7386 532454 -7302
rect 531834 -7622 531866 -7386
rect 532102 -7622 532186 -7386
rect 532422 -7622 532454 -7386
rect 531834 -7654 532454 -7622
rect 541794 75454 542414 110898
rect 541794 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 542414 75454
rect 541794 75134 542414 75218
rect 541794 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 542414 75134
rect 541794 39454 542414 74898
rect 545514 403174 546134 438618
rect 546266 439174 546586 439206
rect 546266 438938 546308 439174
rect 546544 438938 546586 439174
rect 546266 438854 546586 438938
rect 546266 438618 546308 438854
rect 546544 438618 546586 438854
rect 546266 438586 546586 438618
rect 545514 402938 545546 403174
rect 545782 402938 545866 403174
rect 546102 402938 546134 403174
rect 545514 402854 546134 402938
rect 545514 402618 545546 402854
rect 545782 402618 545866 402854
rect 546102 402618 546134 402854
rect 545514 367174 546134 402618
rect 545514 366938 545546 367174
rect 545782 366938 545866 367174
rect 546102 366938 546134 367174
rect 545514 366854 546134 366938
rect 545514 366618 545546 366854
rect 545782 366618 545866 366854
rect 546102 366618 546134 366854
rect 545514 331174 546134 366618
rect 545514 330938 545546 331174
rect 545782 330938 545866 331174
rect 546102 330938 546134 331174
rect 545514 330854 546134 330938
rect 545514 330618 545546 330854
rect 545782 330618 545866 330854
rect 546102 330618 546134 330854
rect 545514 295174 546134 330618
rect 545514 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 546134 295174
rect 545514 294854 546134 294938
rect 545514 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 546134 294854
rect 545514 259174 546134 294618
rect 545514 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 546134 259174
rect 545514 258854 546134 258938
rect 545514 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 546134 258854
rect 545514 223174 546134 258618
rect 545514 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 546134 223174
rect 545514 222854 546134 222938
rect 545514 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 546134 222854
rect 545514 187174 546134 222618
rect 545514 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 546134 187174
rect 545514 186854 546134 186938
rect 545514 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 546134 186854
rect 545514 151174 546134 186618
rect 545514 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 546134 151174
rect 545514 150854 546134 150938
rect 545514 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 546134 150854
rect 545514 115174 546134 150618
rect 545514 114938 545546 115174
rect 545782 114938 545866 115174
rect 546102 114938 546134 115174
rect 545514 114854 546134 114938
rect 545514 114618 545546 114854
rect 545782 114618 545866 114854
rect 546102 114618 546134 114854
rect 545514 79174 546134 114618
rect 545514 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 546134 79174
rect 545514 78854 546134 78938
rect 545514 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 546134 78854
rect 545514 51692 546134 78618
rect 549234 406894 549854 442338
rect 552954 707718 553574 711590
rect 552954 707482 552986 707718
rect 553222 707482 553306 707718
rect 553542 707482 553574 707718
rect 552954 707398 553574 707482
rect 552954 707162 552986 707398
rect 553222 707162 553306 707398
rect 553542 707162 553574 707398
rect 552954 698614 553574 707162
rect 552954 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 553574 698614
rect 552954 698294 553574 698378
rect 552954 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 553574 698294
rect 552954 662614 553574 698058
rect 552954 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 553574 662614
rect 552954 662294 553574 662378
rect 552954 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 553574 662294
rect 552954 626614 553574 662058
rect 552954 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 553574 626614
rect 552954 626294 553574 626378
rect 552954 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 553574 626294
rect 552954 590614 553574 626058
rect 552954 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 553574 590614
rect 552954 590294 553574 590378
rect 552954 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 553574 590294
rect 552954 554614 553574 590058
rect 552954 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 553574 554614
rect 552954 554294 553574 554378
rect 552954 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 553574 554294
rect 552954 518614 553574 554058
rect 552954 518378 552986 518614
rect 553222 518378 553306 518614
rect 553542 518378 553574 518614
rect 552954 518294 553574 518378
rect 552954 518058 552986 518294
rect 553222 518058 553306 518294
rect 553542 518058 553574 518294
rect 552954 482614 553574 518058
rect 552954 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 553574 482614
rect 552954 482294 553574 482378
rect 552954 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 553574 482294
rect 552954 446614 553574 482058
rect 552954 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 553574 446614
rect 552954 446294 553574 446378
rect 552954 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 553574 446294
rect 550487 435454 550807 435486
rect 550487 435218 550529 435454
rect 550765 435218 550807 435454
rect 550487 435134 550807 435218
rect 550487 434898 550529 435134
rect 550765 434898 550807 435134
rect 550487 434866 550807 434898
rect 549234 406658 549266 406894
rect 549502 406658 549586 406894
rect 549822 406658 549854 406894
rect 549234 406574 549854 406658
rect 549234 406338 549266 406574
rect 549502 406338 549586 406574
rect 549822 406338 549854 406574
rect 549234 370894 549854 406338
rect 552954 410614 553574 446058
rect 556674 708678 557294 711590
rect 556674 708442 556706 708678
rect 556942 708442 557026 708678
rect 557262 708442 557294 708678
rect 556674 708358 557294 708442
rect 556674 708122 556706 708358
rect 556942 708122 557026 708358
rect 557262 708122 557294 708358
rect 556674 666334 557294 708122
rect 560394 709638 561014 711590
rect 560394 709402 560426 709638
rect 560662 709402 560746 709638
rect 560982 709402 561014 709638
rect 560394 709318 561014 709402
rect 560394 709082 560426 709318
rect 560662 709082 560746 709318
rect 560982 709082 561014 709318
rect 558131 699820 558197 699821
rect 558131 699756 558132 699820
rect 558196 699756 558197 699820
rect 558131 699755 558197 699756
rect 556674 666098 556706 666334
rect 556942 666098 557026 666334
rect 557262 666098 557294 666334
rect 556674 666014 557294 666098
rect 556674 665778 556706 666014
rect 556942 665778 557026 666014
rect 557262 665778 557294 666014
rect 556674 630334 557294 665778
rect 556674 630098 556706 630334
rect 556942 630098 557026 630334
rect 557262 630098 557294 630334
rect 556674 630014 557294 630098
rect 556674 629778 556706 630014
rect 556942 629778 557026 630014
rect 557262 629778 557294 630014
rect 556674 594334 557294 629778
rect 556674 594098 556706 594334
rect 556942 594098 557026 594334
rect 557262 594098 557294 594334
rect 556674 594014 557294 594098
rect 556674 593778 556706 594014
rect 556942 593778 557026 594014
rect 557262 593778 557294 594014
rect 556674 558334 557294 593778
rect 556674 558098 556706 558334
rect 556942 558098 557026 558334
rect 557262 558098 557294 558334
rect 556674 558014 557294 558098
rect 556674 557778 556706 558014
rect 556942 557778 557026 558014
rect 557262 557778 557294 558014
rect 556674 522334 557294 557778
rect 556674 522098 556706 522334
rect 556942 522098 557026 522334
rect 557262 522098 557294 522334
rect 556674 522014 557294 522098
rect 556674 521778 556706 522014
rect 556942 521778 557026 522014
rect 557262 521778 557294 522014
rect 556674 486334 557294 521778
rect 556674 486098 556706 486334
rect 556942 486098 557026 486334
rect 557262 486098 557294 486334
rect 556674 486014 557294 486098
rect 556674 485778 556706 486014
rect 556942 485778 557026 486014
rect 557262 485778 557294 486014
rect 556674 450334 557294 485778
rect 556674 450098 556706 450334
rect 556942 450098 557026 450334
rect 557262 450098 557294 450334
rect 556674 450014 557294 450098
rect 556674 449778 556706 450014
rect 556942 449778 557026 450014
rect 557262 449778 557294 450014
rect 554707 439174 555027 439206
rect 554707 438938 554749 439174
rect 554985 438938 555027 439174
rect 554707 438854 555027 438938
rect 554707 438618 554749 438854
rect 554985 438618 555027 438854
rect 554707 438586 555027 438618
rect 552954 410378 552986 410614
rect 553222 410378 553306 410614
rect 553542 410378 553574 410614
rect 552954 410294 553574 410378
rect 552954 410058 552986 410294
rect 553222 410058 553306 410294
rect 553542 410058 553574 410294
rect 552954 377884 553574 410058
rect 556674 414334 557294 449778
rect 556674 414098 556706 414334
rect 556942 414098 557026 414334
rect 557262 414098 557294 414334
rect 556674 414014 557294 414098
rect 556674 413778 556706 414014
rect 556942 413778 557026 414014
rect 557262 413778 557294 414014
rect 556674 378243 557294 413778
rect 556674 378007 556706 378243
rect 556942 378007 557026 378243
rect 557262 378007 557294 378243
rect 556674 377884 557294 378007
rect 549234 370658 549266 370894
rect 549502 370658 549586 370894
rect 549822 370658 549854 370894
rect 549234 370574 549854 370658
rect 549234 370338 549266 370574
rect 549502 370338 549586 370574
rect 549822 370338 549854 370574
rect 549234 334894 549854 370338
rect 554876 367174 555196 367206
rect 554876 366938 554918 367174
rect 555154 366938 555196 367174
rect 554876 366854 555196 366938
rect 554876 366618 554918 366854
rect 555154 366618 555196 366854
rect 554876 366586 555196 366618
rect 552910 363454 553230 363486
rect 552910 363218 552952 363454
rect 553188 363218 553230 363454
rect 552910 363134 553230 363218
rect 552910 362898 552952 363134
rect 553188 362898 553230 363134
rect 552910 362866 553230 362898
rect 556843 363454 557163 363486
rect 556843 363218 556885 363454
rect 557121 363218 557163 363454
rect 556843 363134 557163 363218
rect 556843 362898 556885 363134
rect 557121 362898 557163 363134
rect 556843 362866 557163 362898
rect 549234 334658 549266 334894
rect 549502 334658 549586 334894
rect 549822 334658 549854 334894
rect 549234 334574 549854 334658
rect 549234 334338 549266 334574
rect 549502 334338 549586 334574
rect 549822 334338 549854 334574
rect 549234 298894 549854 334338
rect 549234 298658 549266 298894
rect 549502 298658 549586 298894
rect 549822 298658 549854 298894
rect 549234 298574 549854 298658
rect 549234 298338 549266 298574
rect 549502 298338 549586 298574
rect 549822 298338 549854 298574
rect 549234 262894 549854 298338
rect 549234 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 549854 262894
rect 549234 262574 549854 262658
rect 549234 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 549854 262574
rect 549234 226894 549854 262338
rect 549234 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 549854 226894
rect 549234 226574 549854 226658
rect 549234 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 549854 226574
rect 549234 190894 549854 226338
rect 549234 190658 549266 190894
rect 549502 190658 549586 190894
rect 549822 190658 549854 190894
rect 549234 190574 549854 190658
rect 549234 190338 549266 190574
rect 549502 190338 549586 190574
rect 549822 190338 549854 190574
rect 549234 154894 549854 190338
rect 549234 154658 549266 154894
rect 549502 154658 549586 154894
rect 549822 154658 549854 154894
rect 549234 154574 549854 154658
rect 549234 154338 549266 154574
rect 549502 154338 549586 154574
rect 549822 154338 549854 154574
rect 549234 118894 549854 154338
rect 549234 118658 549266 118894
rect 549502 118658 549586 118894
rect 549822 118658 549854 118894
rect 549234 118574 549854 118658
rect 549234 118338 549266 118574
rect 549502 118338 549586 118574
rect 549822 118338 549854 118574
rect 549234 82894 549854 118338
rect 549234 82658 549266 82894
rect 549502 82658 549586 82894
rect 549822 82658 549854 82894
rect 549234 82574 549854 82658
rect 549234 82338 549266 82574
rect 549502 82338 549586 82574
rect 549822 82338 549854 82574
rect 549234 46894 549854 82338
rect 552954 338614 553574 360068
rect 552954 338378 552986 338614
rect 553222 338378 553306 338614
rect 553542 338378 553574 338614
rect 552954 338294 553574 338378
rect 552954 338058 552986 338294
rect 553222 338058 553306 338294
rect 553542 338058 553574 338294
rect 552954 302614 553574 338058
rect 552954 302378 552986 302614
rect 553222 302378 553306 302614
rect 553542 302378 553574 302614
rect 552954 302294 553574 302378
rect 552954 302058 552986 302294
rect 553222 302058 553306 302294
rect 553542 302058 553574 302294
rect 552954 266614 553574 302058
rect 552954 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 553574 266614
rect 552954 266294 553574 266378
rect 552954 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 553574 266294
rect 552954 230614 553574 266058
rect 552954 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 553574 230614
rect 552954 230294 553574 230378
rect 552954 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 553574 230294
rect 552954 194614 553574 230058
rect 552954 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 553574 194614
rect 552954 194294 553574 194378
rect 552954 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 553574 194294
rect 552954 158614 553574 194058
rect 552954 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 553574 158614
rect 552954 158294 553574 158378
rect 552954 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 553574 158294
rect 552954 122614 553574 158058
rect 552954 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 553574 122614
rect 552954 122294 553574 122378
rect 552954 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 553574 122294
rect 552954 86614 553574 122058
rect 552954 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 553574 86614
rect 552954 86294 553574 86378
rect 552954 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 553574 86294
rect 552954 51692 553574 86058
rect 556674 342334 557294 360068
rect 556674 342098 556706 342334
rect 556942 342098 557026 342334
rect 557262 342098 557294 342334
rect 556674 342014 557294 342098
rect 556674 341778 556706 342014
rect 556942 341778 557026 342014
rect 557262 341778 557294 342014
rect 556674 306334 557294 341778
rect 558134 320653 558194 699755
rect 560394 670054 561014 709082
rect 560394 669818 560426 670054
rect 560662 669818 560746 670054
rect 560982 669818 561014 670054
rect 560394 669734 561014 669818
rect 560394 669498 560426 669734
rect 560662 669498 560746 669734
rect 560982 669498 561014 669734
rect 560394 634054 561014 669498
rect 560394 633818 560426 634054
rect 560662 633818 560746 634054
rect 560982 633818 561014 634054
rect 560394 633734 561014 633818
rect 560394 633498 560426 633734
rect 560662 633498 560746 633734
rect 560982 633498 561014 633734
rect 560394 598054 561014 633498
rect 560394 597818 560426 598054
rect 560662 597818 560746 598054
rect 560982 597818 561014 598054
rect 560394 597734 561014 597818
rect 560394 597498 560426 597734
rect 560662 597498 560746 597734
rect 560982 597498 561014 597734
rect 560394 562054 561014 597498
rect 560394 561818 560426 562054
rect 560662 561818 560746 562054
rect 560982 561818 561014 562054
rect 560394 561734 561014 561818
rect 560394 561498 560426 561734
rect 560662 561498 560746 561734
rect 560982 561498 561014 561734
rect 560394 526054 561014 561498
rect 560394 525818 560426 526054
rect 560662 525818 560746 526054
rect 560982 525818 561014 526054
rect 560394 525734 561014 525818
rect 560394 525498 560426 525734
rect 560662 525498 560746 525734
rect 560982 525498 561014 525734
rect 560394 490054 561014 525498
rect 560394 489818 560426 490054
rect 560662 489818 560746 490054
rect 560982 489818 561014 490054
rect 560394 489734 561014 489818
rect 560394 489498 560426 489734
rect 560662 489498 560746 489734
rect 560982 489498 561014 489734
rect 560394 454054 561014 489498
rect 560394 453818 560426 454054
rect 560662 453818 560746 454054
rect 560982 453818 561014 454054
rect 560394 453734 561014 453818
rect 560394 453498 560426 453734
rect 560662 453498 560746 453734
rect 560982 453498 561014 453734
rect 560394 418054 561014 453498
rect 560394 417818 560426 418054
rect 560662 417818 560746 418054
rect 560982 417818 561014 418054
rect 560394 417734 561014 417818
rect 560394 417498 560426 417734
rect 560662 417498 560746 417734
rect 560982 417498 561014 417734
rect 560394 382054 561014 417498
rect 560394 381818 560426 382054
rect 560662 381818 560746 382054
rect 560982 381818 561014 382054
rect 560394 381734 561014 381818
rect 560394 381498 560426 381734
rect 560662 381498 560746 381734
rect 560982 381498 561014 381734
rect 560394 377884 561014 381498
rect 564114 710598 564734 711590
rect 564114 710362 564146 710598
rect 564382 710362 564466 710598
rect 564702 710362 564734 710598
rect 564114 710278 564734 710362
rect 564114 710042 564146 710278
rect 564382 710042 564466 710278
rect 564702 710042 564734 710278
rect 564114 673774 564734 710042
rect 564114 673538 564146 673774
rect 564382 673538 564466 673774
rect 564702 673538 564734 673774
rect 564114 673454 564734 673538
rect 564114 673218 564146 673454
rect 564382 673218 564466 673454
rect 564702 673218 564734 673454
rect 564114 637774 564734 673218
rect 564114 637538 564146 637774
rect 564382 637538 564466 637774
rect 564702 637538 564734 637774
rect 564114 637454 564734 637538
rect 564114 637218 564146 637454
rect 564382 637218 564466 637454
rect 564702 637218 564734 637454
rect 564114 601774 564734 637218
rect 564114 601538 564146 601774
rect 564382 601538 564466 601774
rect 564702 601538 564734 601774
rect 564114 601454 564734 601538
rect 564114 601218 564146 601454
rect 564382 601218 564466 601454
rect 564702 601218 564734 601454
rect 564114 565774 564734 601218
rect 564114 565538 564146 565774
rect 564382 565538 564466 565774
rect 564702 565538 564734 565774
rect 564114 565454 564734 565538
rect 564114 565218 564146 565454
rect 564382 565218 564466 565454
rect 564702 565218 564734 565454
rect 564114 529774 564734 565218
rect 564114 529538 564146 529774
rect 564382 529538 564466 529774
rect 564702 529538 564734 529774
rect 564114 529454 564734 529538
rect 564114 529218 564146 529454
rect 564382 529218 564466 529454
rect 564702 529218 564734 529454
rect 564114 493774 564734 529218
rect 564114 493538 564146 493774
rect 564382 493538 564466 493774
rect 564702 493538 564734 493774
rect 564114 493454 564734 493538
rect 564114 493218 564146 493454
rect 564382 493218 564466 493454
rect 564702 493218 564734 493454
rect 564114 457774 564734 493218
rect 564114 457538 564146 457774
rect 564382 457538 564466 457774
rect 564702 457538 564734 457774
rect 564114 457454 564734 457538
rect 564114 457218 564146 457454
rect 564382 457218 564466 457454
rect 564702 457218 564734 457454
rect 564114 421774 564734 457218
rect 564114 421538 564146 421774
rect 564382 421538 564466 421774
rect 564702 421538 564734 421774
rect 564114 421454 564734 421538
rect 564114 421218 564146 421454
rect 564382 421218 564466 421454
rect 564702 421218 564734 421454
rect 564114 385774 564734 421218
rect 564114 385538 564146 385774
rect 564382 385538 564466 385774
rect 564702 385538 564734 385774
rect 564114 385454 564734 385538
rect 564114 385218 564146 385454
rect 564382 385218 564466 385454
rect 564702 385218 564734 385454
rect 564114 377884 564734 385218
rect 567834 711558 568454 711590
rect 567834 711322 567866 711558
rect 568102 711322 568186 711558
rect 568422 711322 568454 711558
rect 567834 711238 568454 711322
rect 567834 711002 567866 711238
rect 568102 711002 568186 711238
rect 568422 711002 568454 711238
rect 567834 677494 568454 711002
rect 567834 677258 567866 677494
rect 568102 677258 568186 677494
rect 568422 677258 568454 677494
rect 567834 677174 568454 677258
rect 567834 676938 567866 677174
rect 568102 676938 568186 677174
rect 568422 676938 568454 677174
rect 567834 641494 568454 676938
rect 567834 641258 567866 641494
rect 568102 641258 568186 641494
rect 568422 641258 568454 641494
rect 567834 641174 568454 641258
rect 567834 640938 567866 641174
rect 568102 640938 568186 641174
rect 568422 640938 568454 641174
rect 567834 605494 568454 640938
rect 567834 605258 567866 605494
rect 568102 605258 568186 605494
rect 568422 605258 568454 605494
rect 567834 605174 568454 605258
rect 567834 604938 567866 605174
rect 568102 604938 568186 605174
rect 568422 604938 568454 605174
rect 567834 569494 568454 604938
rect 567834 569258 567866 569494
rect 568102 569258 568186 569494
rect 568422 569258 568454 569494
rect 567834 569174 568454 569258
rect 567834 568938 567866 569174
rect 568102 568938 568186 569174
rect 568422 568938 568454 569174
rect 567834 533494 568454 568938
rect 567834 533258 567866 533494
rect 568102 533258 568186 533494
rect 568422 533258 568454 533494
rect 567834 533174 568454 533258
rect 567834 532938 567866 533174
rect 568102 532938 568186 533174
rect 568422 532938 568454 533174
rect 567834 497494 568454 532938
rect 567834 497258 567866 497494
rect 568102 497258 568186 497494
rect 568422 497258 568454 497494
rect 567834 497174 568454 497258
rect 567834 496938 567866 497174
rect 568102 496938 568186 497174
rect 568422 496938 568454 497174
rect 567834 461494 568454 496938
rect 567834 461258 567866 461494
rect 568102 461258 568186 461494
rect 568422 461258 568454 461494
rect 567834 461174 568454 461258
rect 567834 460938 567866 461174
rect 568102 460938 568186 461174
rect 568422 460938 568454 461174
rect 567834 425494 568454 460938
rect 567834 425258 567866 425494
rect 568102 425258 568186 425494
rect 568422 425258 568454 425494
rect 567834 425174 568454 425258
rect 567834 424938 567866 425174
rect 568102 424938 568186 425174
rect 568422 424938 568454 425174
rect 567834 389494 568454 424938
rect 567834 389258 567866 389494
rect 568102 389258 568186 389494
rect 568422 389258 568454 389494
rect 567834 389174 568454 389258
rect 567834 388938 567866 389174
rect 568102 388938 568186 389174
rect 568422 388938 568454 389174
rect 558809 367174 559129 367206
rect 558809 366938 558851 367174
rect 559087 366938 559129 367174
rect 558809 366854 559129 366938
rect 558809 366618 558851 366854
rect 559087 366618 559129 366854
rect 558809 366586 559129 366618
rect 562742 367174 563062 367206
rect 562742 366938 562784 367174
rect 563020 366938 563062 367174
rect 562742 366854 563062 366938
rect 562742 366618 562784 366854
rect 563020 366618 563062 366854
rect 562742 366586 563062 366618
rect 566675 367174 566995 367206
rect 566675 366938 566717 367174
rect 566953 366938 566995 367174
rect 566675 366854 566995 366938
rect 566675 366618 566717 366854
rect 566953 366618 566995 366854
rect 566675 366586 566995 366618
rect 560776 363454 561096 363486
rect 560776 363218 560818 363454
rect 561054 363218 561096 363454
rect 560776 363134 561096 363218
rect 560776 362898 560818 363134
rect 561054 362898 561096 363134
rect 560776 362866 561096 362898
rect 564709 363454 565029 363486
rect 564709 363218 564751 363454
rect 564987 363218 565029 363454
rect 564709 363134 565029 363218
rect 564709 362898 564751 363134
rect 564987 362898 565029 363134
rect 564709 362866 565029 362898
rect 560394 346054 561014 360068
rect 560394 345818 560426 346054
rect 560662 345818 560746 346054
rect 560982 345818 561014 346054
rect 560394 345734 561014 345818
rect 560394 345498 560426 345734
rect 560662 345498 560746 345734
rect 560982 345498 561014 345734
rect 558131 320652 558197 320653
rect 558131 320588 558132 320652
rect 558196 320588 558197 320652
rect 558131 320587 558197 320588
rect 556674 306098 556706 306334
rect 556942 306098 557026 306334
rect 557262 306098 557294 306334
rect 556674 306014 557294 306098
rect 556674 305778 556706 306014
rect 556942 305778 557026 306014
rect 557262 305778 557294 306014
rect 556674 270334 557294 305778
rect 556674 270098 556706 270334
rect 556942 270098 557026 270334
rect 557262 270098 557294 270334
rect 556674 270014 557294 270098
rect 556674 269778 556706 270014
rect 556942 269778 557026 270014
rect 557262 269778 557294 270014
rect 556674 234334 557294 269778
rect 556674 234098 556706 234334
rect 556942 234098 557026 234334
rect 557262 234098 557294 234334
rect 556674 234014 557294 234098
rect 556674 233778 556706 234014
rect 556942 233778 557026 234014
rect 557262 233778 557294 234014
rect 556674 198334 557294 233778
rect 556674 198098 556706 198334
rect 556942 198098 557026 198334
rect 557262 198098 557294 198334
rect 556674 198014 557294 198098
rect 556674 197778 556706 198014
rect 556942 197778 557026 198014
rect 557262 197778 557294 198014
rect 556674 162334 557294 197778
rect 556674 162098 556706 162334
rect 556942 162098 557026 162334
rect 557262 162098 557294 162334
rect 556674 162014 557294 162098
rect 556674 161778 556706 162014
rect 556942 161778 557026 162014
rect 557262 161778 557294 162014
rect 556674 126334 557294 161778
rect 556674 126098 556706 126334
rect 556942 126098 557026 126334
rect 557262 126098 557294 126334
rect 556674 126014 557294 126098
rect 556674 125778 556706 126014
rect 556942 125778 557026 126014
rect 557262 125778 557294 126014
rect 556674 90334 557294 125778
rect 556674 90098 556706 90334
rect 556942 90098 557026 90334
rect 557262 90098 557294 90334
rect 556674 90014 557294 90098
rect 556674 89778 556706 90014
rect 556942 89778 557026 90014
rect 557262 89778 557294 90014
rect 556674 54334 557294 89778
rect 556674 54098 556706 54334
rect 556942 54098 557026 54334
rect 557262 54098 557294 54334
rect 556674 54014 557294 54098
rect 556674 53778 556706 54014
rect 556942 53778 557026 54014
rect 557262 53778 557294 54014
rect 549234 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 549854 46894
rect 549234 46574 549854 46658
rect 549234 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 549854 46574
rect 545888 43174 546208 43206
rect 545888 42938 545930 43174
rect 546166 42938 546208 43174
rect 545888 42854 546208 42938
rect 545888 42618 545930 42854
rect 546166 42618 546208 42854
rect 545888 42586 546208 42618
rect 541794 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 542414 39454
rect 541794 39134 542414 39218
rect 541794 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 542414 39134
rect 541794 3454 542414 38898
rect 543416 39454 543736 39486
rect 543416 39218 543458 39454
rect 543694 39218 543736 39454
rect 543416 39134 543736 39218
rect 543416 38898 543458 39134
rect 543694 38898 543736 39134
rect 543416 38866 543736 38898
rect 548361 39454 548681 39486
rect 548361 39218 548403 39454
rect 548639 39218 548681 39454
rect 548361 39134 548681 39218
rect 548361 38898 548403 39134
rect 548639 38898 548681 39134
rect 548361 38866 548681 38898
rect 541794 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 542414 3454
rect 541794 3134 542414 3218
rect 541794 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 542414 3134
rect 541794 -346 542414 2898
rect 541794 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 542414 -346
rect 541794 -666 542414 -582
rect 541794 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 542414 -666
rect 541794 -7654 542414 -902
rect 545514 7174 546134 30068
rect 545514 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 546134 7174
rect 545514 6854 546134 6938
rect 545514 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 546134 6854
rect 545514 -1306 546134 6618
rect 545514 -1542 545546 -1306
rect 545782 -1542 545866 -1306
rect 546102 -1542 546134 -1306
rect 545514 -1626 546134 -1542
rect 545514 -1862 545546 -1626
rect 545782 -1862 545866 -1626
rect 546102 -1862 546134 -1626
rect 545514 -7654 546134 -1862
rect 549234 10894 549854 46338
rect 550833 43174 551153 43206
rect 550833 42938 550875 43174
rect 551111 42938 551153 43174
rect 550833 42854 551153 42938
rect 550833 42618 550875 42854
rect 551111 42618 551153 42854
rect 550833 42586 551153 42618
rect 555778 43174 556098 43206
rect 555778 42938 555820 43174
rect 556056 42938 556098 43174
rect 555778 42854 556098 42938
rect 555778 42618 555820 42854
rect 556056 42618 556098 42854
rect 555778 42586 556098 42618
rect 553306 39454 553626 39486
rect 553306 39218 553348 39454
rect 553584 39218 553626 39454
rect 553306 39134 553626 39218
rect 553306 38898 553348 39134
rect 553584 38898 553626 39134
rect 553306 38866 553626 38898
rect 549234 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 549854 10894
rect 549234 10574 549854 10658
rect 549234 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 549854 10574
rect 549234 -2266 549854 10338
rect 549234 -2502 549266 -2266
rect 549502 -2502 549586 -2266
rect 549822 -2502 549854 -2266
rect 549234 -2586 549854 -2502
rect 549234 -2822 549266 -2586
rect 549502 -2822 549586 -2586
rect 549822 -2822 549854 -2586
rect 549234 -7654 549854 -2822
rect 552954 14614 553574 30068
rect 552954 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 553574 14614
rect 552954 14294 553574 14378
rect 552954 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 553574 14294
rect 552954 -3226 553574 14058
rect 552954 -3462 552986 -3226
rect 553222 -3462 553306 -3226
rect 553542 -3462 553574 -3226
rect 552954 -3546 553574 -3462
rect 552954 -3782 552986 -3546
rect 553222 -3782 553306 -3546
rect 553542 -3782 553574 -3546
rect 552954 -7654 553574 -3782
rect 556674 18334 557294 53778
rect 560394 310054 561014 345498
rect 560394 309818 560426 310054
rect 560662 309818 560746 310054
rect 560982 309818 561014 310054
rect 560394 309734 561014 309818
rect 560394 309498 560426 309734
rect 560662 309498 560746 309734
rect 560982 309498 561014 309734
rect 560394 274054 561014 309498
rect 560394 273818 560426 274054
rect 560662 273818 560746 274054
rect 560982 273818 561014 274054
rect 560394 273734 561014 273818
rect 560394 273498 560426 273734
rect 560662 273498 560746 273734
rect 560982 273498 561014 273734
rect 560394 238054 561014 273498
rect 560394 237818 560426 238054
rect 560662 237818 560746 238054
rect 560982 237818 561014 238054
rect 560394 237734 561014 237818
rect 560394 237498 560426 237734
rect 560662 237498 560746 237734
rect 560982 237498 561014 237734
rect 560394 202054 561014 237498
rect 560394 201818 560426 202054
rect 560662 201818 560746 202054
rect 560982 201818 561014 202054
rect 560394 201734 561014 201818
rect 560394 201498 560426 201734
rect 560662 201498 560746 201734
rect 560982 201498 561014 201734
rect 560394 166054 561014 201498
rect 560394 165818 560426 166054
rect 560662 165818 560746 166054
rect 560982 165818 561014 166054
rect 560394 165734 561014 165818
rect 560394 165498 560426 165734
rect 560662 165498 560746 165734
rect 560982 165498 561014 165734
rect 560394 130054 561014 165498
rect 560394 129818 560426 130054
rect 560662 129818 560746 130054
rect 560982 129818 561014 130054
rect 560394 129734 561014 129818
rect 560394 129498 560426 129734
rect 560662 129498 560746 129734
rect 560982 129498 561014 129734
rect 560394 94054 561014 129498
rect 560394 93818 560426 94054
rect 560662 93818 560746 94054
rect 560982 93818 561014 94054
rect 560394 93734 561014 93818
rect 560394 93498 560426 93734
rect 560662 93498 560746 93734
rect 560982 93498 561014 93734
rect 560394 58054 561014 93498
rect 560394 57818 560426 58054
rect 560662 57818 560746 58054
rect 560982 57818 561014 58054
rect 560394 57734 561014 57818
rect 560394 57498 560426 57734
rect 560662 57498 560746 57734
rect 560982 57498 561014 57734
rect 560394 51692 561014 57498
rect 564114 349774 564734 360068
rect 564114 349538 564146 349774
rect 564382 349538 564466 349774
rect 564702 349538 564734 349774
rect 564114 349454 564734 349538
rect 564114 349218 564146 349454
rect 564382 349218 564466 349454
rect 564702 349218 564734 349454
rect 564114 313774 564734 349218
rect 564114 313538 564146 313774
rect 564382 313538 564466 313774
rect 564702 313538 564734 313774
rect 564114 313454 564734 313538
rect 564114 313218 564146 313454
rect 564382 313218 564466 313454
rect 564702 313218 564734 313454
rect 564114 277774 564734 313218
rect 564114 277538 564146 277774
rect 564382 277538 564466 277774
rect 564702 277538 564734 277774
rect 564114 277454 564734 277538
rect 564114 277218 564146 277454
rect 564382 277218 564466 277454
rect 564702 277218 564734 277454
rect 564114 241774 564734 277218
rect 564114 241538 564146 241774
rect 564382 241538 564466 241774
rect 564702 241538 564734 241774
rect 564114 241454 564734 241538
rect 564114 241218 564146 241454
rect 564382 241218 564466 241454
rect 564702 241218 564734 241454
rect 564114 205774 564734 241218
rect 564114 205538 564146 205774
rect 564382 205538 564466 205774
rect 564702 205538 564734 205774
rect 564114 205454 564734 205538
rect 564114 205218 564146 205454
rect 564382 205218 564466 205454
rect 564702 205218 564734 205454
rect 564114 169774 564734 205218
rect 564114 169538 564146 169774
rect 564382 169538 564466 169774
rect 564702 169538 564734 169774
rect 564114 169454 564734 169538
rect 564114 169218 564146 169454
rect 564382 169218 564466 169454
rect 564702 169218 564734 169454
rect 564114 133774 564734 169218
rect 564114 133538 564146 133774
rect 564382 133538 564466 133774
rect 564702 133538 564734 133774
rect 564114 133454 564734 133538
rect 564114 133218 564146 133454
rect 564382 133218 564466 133454
rect 564702 133218 564734 133454
rect 564114 97774 564734 133218
rect 564114 97538 564146 97774
rect 564382 97538 564466 97774
rect 564702 97538 564734 97774
rect 564114 97454 564734 97538
rect 564114 97218 564146 97454
rect 564382 97218 564466 97454
rect 564702 97218 564734 97454
rect 564114 61774 564734 97218
rect 564114 61538 564146 61774
rect 564382 61538 564466 61774
rect 564702 61538 564734 61774
rect 564114 61454 564734 61538
rect 564114 61218 564146 61454
rect 564382 61218 564466 61454
rect 564702 61218 564734 61454
rect 560723 43174 561043 43206
rect 560723 42938 560765 43174
rect 561001 42938 561043 43174
rect 560723 42854 561043 42938
rect 560723 42618 560765 42854
rect 561001 42618 561043 42854
rect 560723 42586 561043 42618
rect 558251 39454 558571 39486
rect 558251 39218 558293 39454
rect 558529 39218 558571 39454
rect 558251 39134 558571 39218
rect 558251 38898 558293 39134
rect 558529 38898 558571 39134
rect 558251 38866 558571 38898
rect 556674 18098 556706 18334
rect 556942 18098 557026 18334
rect 557262 18098 557294 18334
rect 556674 18014 557294 18098
rect 556674 17778 556706 18014
rect 556942 17778 557026 18014
rect 557262 17778 557294 18014
rect 556674 -4186 557294 17778
rect 556674 -4422 556706 -4186
rect 556942 -4422 557026 -4186
rect 557262 -4422 557294 -4186
rect 556674 -4506 557294 -4422
rect 556674 -4742 556706 -4506
rect 556942 -4742 557026 -4506
rect 557262 -4742 557294 -4506
rect 556674 -7654 557294 -4742
rect 560394 22054 561014 30068
rect 560394 21818 560426 22054
rect 560662 21818 560746 22054
rect 560982 21818 561014 22054
rect 560394 21734 561014 21818
rect 560394 21498 560426 21734
rect 560662 21498 560746 21734
rect 560982 21498 561014 21734
rect 560394 -5146 561014 21498
rect 560394 -5382 560426 -5146
rect 560662 -5382 560746 -5146
rect 560982 -5382 561014 -5146
rect 560394 -5466 561014 -5382
rect 560394 -5702 560426 -5466
rect 560662 -5702 560746 -5466
rect 560982 -5702 561014 -5466
rect 560394 -7654 561014 -5702
rect 564114 25774 564734 61218
rect 564114 25538 564146 25774
rect 564382 25538 564466 25774
rect 564702 25538 564734 25774
rect 564114 25454 564734 25538
rect 564114 25218 564146 25454
rect 564382 25218 564466 25454
rect 564702 25218 564734 25454
rect 564114 -6106 564734 25218
rect 564114 -6342 564146 -6106
rect 564382 -6342 564466 -6106
rect 564702 -6342 564734 -6106
rect 564114 -6426 564734 -6342
rect 564114 -6662 564146 -6426
rect 564382 -6662 564466 -6426
rect 564702 -6662 564734 -6426
rect 564114 -7654 564734 -6662
rect 567834 353494 568454 388938
rect 567834 353258 567866 353494
rect 568102 353258 568186 353494
rect 568422 353258 568454 353494
rect 567834 353174 568454 353258
rect 567834 352938 567866 353174
rect 568102 352938 568186 353174
rect 568422 352938 568454 353174
rect 567834 317494 568454 352938
rect 567834 317258 567866 317494
rect 568102 317258 568186 317494
rect 568422 317258 568454 317494
rect 567834 317174 568454 317258
rect 567834 316938 567866 317174
rect 568102 316938 568186 317174
rect 568422 316938 568454 317174
rect 567834 281494 568454 316938
rect 567834 281258 567866 281494
rect 568102 281258 568186 281494
rect 568422 281258 568454 281494
rect 567834 281174 568454 281258
rect 567834 280938 567866 281174
rect 568102 280938 568186 281174
rect 568422 280938 568454 281174
rect 567834 245494 568454 280938
rect 567834 245258 567866 245494
rect 568102 245258 568186 245494
rect 568422 245258 568454 245494
rect 567834 245174 568454 245258
rect 567834 244938 567866 245174
rect 568102 244938 568186 245174
rect 568422 244938 568454 245174
rect 567834 209494 568454 244938
rect 567834 209258 567866 209494
rect 568102 209258 568186 209494
rect 568422 209258 568454 209494
rect 567834 209174 568454 209258
rect 567834 208938 567866 209174
rect 568102 208938 568186 209174
rect 568422 208938 568454 209174
rect 567834 173494 568454 208938
rect 567834 173258 567866 173494
rect 568102 173258 568186 173494
rect 568422 173258 568454 173494
rect 567834 173174 568454 173258
rect 567834 172938 567866 173174
rect 568102 172938 568186 173174
rect 568422 172938 568454 173174
rect 567834 137494 568454 172938
rect 567834 137258 567866 137494
rect 568102 137258 568186 137494
rect 568422 137258 568454 137494
rect 567834 137174 568454 137258
rect 567834 136938 567866 137174
rect 568102 136938 568186 137174
rect 568422 136938 568454 137174
rect 567834 101494 568454 136938
rect 567834 101258 567866 101494
rect 568102 101258 568186 101494
rect 568422 101258 568454 101494
rect 567834 101174 568454 101258
rect 567834 100938 567866 101174
rect 568102 100938 568186 101174
rect 568422 100938 568454 101174
rect 567834 65494 568454 100938
rect 567834 65258 567866 65494
rect 568102 65258 568186 65494
rect 568422 65258 568454 65494
rect 567834 65174 568454 65258
rect 567834 64938 567866 65174
rect 568102 64938 568186 65174
rect 568422 64938 568454 65174
rect 567834 29494 568454 64938
rect 567834 29258 567866 29494
rect 568102 29258 568186 29494
rect 568422 29258 568454 29494
rect 567834 29174 568454 29258
rect 567834 28938 567866 29174
rect 568102 28938 568186 29174
rect 568422 28938 568454 29174
rect 567834 -7066 568454 28938
rect 567834 -7302 567866 -7066
rect 568102 -7302 568186 -7066
rect 568422 -7302 568454 -7066
rect 567834 -7386 568454 -7302
rect 567834 -7622 567866 -7386
rect 568102 -7622 568186 -7386
rect 568422 -7622 568454 -7386
rect 567834 -7654 568454 -7622
rect 577794 704838 578414 711590
rect 577794 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 578414 704838
rect 577794 704518 578414 704602
rect 577794 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 578414 704518
rect 577794 687454 578414 704282
rect 577794 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 578414 687454
rect 577794 687134 578414 687218
rect 577794 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 578414 687134
rect 577794 651454 578414 686898
rect 577794 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 578414 651454
rect 577794 651134 578414 651218
rect 577794 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 578414 651134
rect 577794 615454 578414 650898
rect 577794 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 578414 615454
rect 577794 615134 578414 615218
rect 577794 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 578414 615134
rect 577794 579454 578414 614898
rect 577794 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 578414 579454
rect 577794 579134 578414 579218
rect 577794 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 578414 579134
rect 577794 543454 578414 578898
rect 577794 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 578414 543454
rect 577794 543134 578414 543218
rect 577794 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 578414 543134
rect 577794 507454 578414 542898
rect 577794 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 578414 507454
rect 577794 507134 578414 507218
rect 577794 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 578414 507134
rect 577794 471454 578414 506898
rect 577794 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 578414 471454
rect 577794 471134 578414 471218
rect 577794 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 578414 471134
rect 577794 435454 578414 470898
rect 577794 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 578414 435454
rect 577794 435134 578414 435218
rect 577794 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 578414 435134
rect 577794 399454 578414 434898
rect 577794 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 578414 399454
rect 577794 399134 578414 399218
rect 577794 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 578414 399134
rect 577794 363454 578414 398898
rect 577794 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 578414 363454
rect 577794 363134 578414 363218
rect 577794 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 578414 363134
rect 577794 327454 578414 362898
rect 577794 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 578414 327454
rect 577794 327134 578414 327218
rect 577794 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 578414 327134
rect 577794 291454 578414 326898
rect 577794 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 578414 291454
rect 577794 291134 578414 291218
rect 577794 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 578414 291134
rect 577794 255454 578414 290898
rect 577794 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 578414 255454
rect 577794 255134 578414 255218
rect 577794 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 578414 255134
rect 577794 219454 578414 254898
rect 577794 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 578414 219454
rect 577794 219134 578414 219218
rect 577794 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 578414 219134
rect 577794 183454 578414 218898
rect 577794 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 578414 183454
rect 577794 183134 578414 183218
rect 577794 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 578414 183134
rect 577794 147454 578414 182898
rect 577794 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 578414 147454
rect 577794 147134 578414 147218
rect 577794 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 578414 147134
rect 577794 111454 578414 146898
rect 577794 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 578414 111454
rect 577794 111134 578414 111218
rect 577794 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 578414 111134
rect 577794 75454 578414 110898
rect 577794 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 578414 75454
rect 577794 75134 578414 75218
rect 577794 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 578414 75134
rect 577794 39454 578414 74898
rect 577794 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 578414 39454
rect 577794 39134 578414 39218
rect 577794 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 578414 39134
rect 577794 3454 578414 38898
rect 577794 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 578414 3454
rect 577794 3134 578414 3218
rect 577794 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 578414 3134
rect 577794 -346 578414 2898
rect 577794 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 578414 -346
rect 577794 -666 578414 -582
rect 577794 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 578414 -666
rect 577794 -7654 578414 -902
rect 581514 705798 582134 711590
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 581514 705562 581546 705798
rect 581782 705562 581866 705798
rect 582102 705562 582134 705798
rect 581514 705478 582134 705562
rect 581514 705242 581546 705478
rect 581782 705242 581866 705478
rect 582102 705242 582134 705478
rect 581514 691174 582134 705242
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 581514 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 582134 691174
rect 581514 690854 582134 690938
rect 581514 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 582134 690854
rect 581514 655174 582134 690618
rect 581514 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 582134 655174
rect 581514 654854 582134 654938
rect 581514 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 582134 654854
rect 581514 619174 582134 654618
rect 581514 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 582134 619174
rect 581514 618854 582134 618938
rect 581514 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 582134 618854
rect 581514 583174 582134 618618
rect 581514 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 582134 583174
rect 581514 582854 582134 582938
rect 581514 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 582134 582854
rect 581514 547174 582134 582618
rect 581514 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 582134 547174
rect 581514 546854 582134 546938
rect 581514 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 582134 546854
rect 581514 511174 582134 546618
rect 581514 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 582134 511174
rect 581514 510854 582134 510938
rect 581514 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 582134 510854
rect 581514 475174 582134 510618
rect 581514 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 582134 475174
rect 581514 474854 582134 474938
rect 581514 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 582134 474854
rect 581514 439174 582134 474618
rect 581514 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 582134 439174
rect 581514 438854 582134 438938
rect 581514 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 582134 438854
rect 581514 403174 582134 438618
rect 581514 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 582134 403174
rect 581514 402854 582134 402938
rect 581514 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 582134 402854
rect 581514 367174 582134 402618
rect 581514 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 582134 367174
rect 581514 366854 582134 366938
rect 581514 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 582134 366854
rect 581514 331174 582134 366618
rect 581514 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 582134 331174
rect 581514 330854 582134 330938
rect 581514 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 582134 330854
rect 581514 295174 582134 330618
rect 581514 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 582134 295174
rect 581514 294854 582134 294938
rect 581514 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 582134 294854
rect 581514 259174 582134 294618
rect 581514 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 582134 259174
rect 581514 258854 582134 258938
rect 581514 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 582134 258854
rect 581514 223174 582134 258618
rect 581514 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 582134 223174
rect 581514 222854 582134 222938
rect 581514 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 582134 222854
rect 581514 187174 582134 222618
rect 581514 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 582134 187174
rect 581514 186854 582134 186938
rect 581514 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 582134 186854
rect 581514 151174 582134 186618
rect 581514 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 582134 151174
rect 581514 150854 582134 150938
rect 581514 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 582134 150854
rect 581514 115174 582134 150618
rect 581514 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 582134 115174
rect 581514 114854 582134 114938
rect 581514 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 582134 114854
rect 581514 79174 582134 114618
rect 581514 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 582134 79174
rect 581514 78854 582134 78938
rect 581514 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 582134 78854
rect 581514 43174 582134 78618
rect 581514 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 582134 43174
rect 581514 42854 582134 42938
rect 581514 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 582134 42854
rect 581514 7174 582134 42618
rect 581514 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 582134 7174
rect 581514 6854 582134 6938
rect 581514 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 582134 6854
rect 581514 -1306 582134 6618
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 687454 585930 704282
rect 585310 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 585930 687454
rect 585310 687134 585930 687218
rect 585310 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 585930 687134
rect 585310 651454 585930 686898
rect 585310 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 585930 651454
rect 585310 651134 585930 651218
rect 585310 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 585930 651134
rect 585310 615454 585930 650898
rect 585310 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 585930 615454
rect 585310 615134 585930 615218
rect 585310 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 585930 615134
rect 585310 579454 585930 614898
rect 585310 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 585930 579454
rect 585310 579134 585930 579218
rect 585310 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 585930 579134
rect 585310 543454 585930 578898
rect 585310 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 585930 543454
rect 585310 543134 585930 543218
rect 585310 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 585930 543134
rect 585310 507454 585930 542898
rect 585310 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 585930 507454
rect 585310 507134 585930 507218
rect 585310 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 585930 507134
rect 585310 471454 585930 506898
rect 585310 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 585930 471454
rect 585310 471134 585930 471218
rect 585310 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 585930 471134
rect 585310 435454 585930 470898
rect 585310 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 585930 435454
rect 585310 435134 585930 435218
rect 585310 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 585930 435134
rect 585310 399454 585930 434898
rect 585310 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 585930 399454
rect 585310 399134 585930 399218
rect 585310 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 585930 399134
rect 585310 363454 585930 398898
rect 585310 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 585930 363454
rect 585310 363134 585930 363218
rect 585310 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 585930 363134
rect 585310 327454 585930 362898
rect 585310 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 585930 327454
rect 585310 327134 585930 327218
rect 585310 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 585930 327134
rect 585310 291454 585930 326898
rect 585310 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 585930 291454
rect 585310 291134 585930 291218
rect 585310 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 585930 291134
rect 585310 255454 585930 290898
rect 585310 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 585930 255454
rect 585310 255134 585930 255218
rect 585310 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 585930 255134
rect 585310 219454 585930 254898
rect 585310 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 585930 219454
rect 585310 219134 585930 219218
rect 585310 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 585930 219134
rect 585310 183454 585930 218898
rect 585310 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 585930 183454
rect 585310 183134 585930 183218
rect 585310 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 585930 183134
rect 585310 147454 585930 182898
rect 585310 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 585930 147454
rect 585310 147134 585930 147218
rect 585310 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 585930 147134
rect 585310 111454 585930 146898
rect 585310 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 585930 111454
rect 585310 111134 585930 111218
rect 585310 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 585930 111134
rect 585310 75454 585930 110898
rect 585310 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 585930 75454
rect 585310 75134 585930 75218
rect 585310 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 585930 75134
rect 585310 39454 585930 74898
rect 585310 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 585930 39454
rect 585310 39134 585930 39218
rect 585310 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 585930 39134
rect 585310 3454 585930 38898
rect 585310 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 585930 3454
rect 585310 3134 585930 3218
rect 585310 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 585930 3134
rect 585310 -346 585930 2898
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 691174 586890 705242
rect 586270 690938 586302 691174
rect 586538 690938 586622 691174
rect 586858 690938 586890 691174
rect 586270 690854 586890 690938
rect 586270 690618 586302 690854
rect 586538 690618 586622 690854
rect 586858 690618 586890 690854
rect 586270 655174 586890 690618
rect 586270 654938 586302 655174
rect 586538 654938 586622 655174
rect 586858 654938 586890 655174
rect 586270 654854 586890 654938
rect 586270 654618 586302 654854
rect 586538 654618 586622 654854
rect 586858 654618 586890 654854
rect 586270 619174 586890 654618
rect 586270 618938 586302 619174
rect 586538 618938 586622 619174
rect 586858 618938 586890 619174
rect 586270 618854 586890 618938
rect 586270 618618 586302 618854
rect 586538 618618 586622 618854
rect 586858 618618 586890 618854
rect 586270 583174 586890 618618
rect 586270 582938 586302 583174
rect 586538 582938 586622 583174
rect 586858 582938 586890 583174
rect 586270 582854 586890 582938
rect 586270 582618 586302 582854
rect 586538 582618 586622 582854
rect 586858 582618 586890 582854
rect 586270 547174 586890 582618
rect 586270 546938 586302 547174
rect 586538 546938 586622 547174
rect 586858 546938 586890 547174
rect 586270 546854 586890 546938
rect 586270 546618 586302 546854
rect 586538 546618 586622 546854
rect 586858 546618 586890 546854
rect 586270 511174 586890 546618
rect 586270 510938 586302 511174
rect 586538 510938 586622 511174
rect 586858 510938 586890 511174
rect 586270 510854 586890 510938
rect 586270 510618 586302 510854
rect 586538 510618 586622 510854
rect 586858 510618 586890 510854
rect 586270 475174 586890 510618
rect 586270 474938 586302 475174
rect 586538 474938 586622 475174
rect 586858 474938 586890 475174
rect 586270 474854 586890 474938
rect 586270 474618 586302 474854
rect 586538 474618 586622 474854
rect 586858 474618 586890 474854
rect 586270 439174 586890 474618
rect 586270 438938 586302 439174
rect 586538 438938 586622 439174
rect 586858 438938 586890 439174
rect 586270 438854 586890 438938
rect 586270 438618 586302 438854
rect 586538 438618 586622 438854
rect 586858 438618 586890 438854
rect 586270 403174 586890 438618
rect 586270 402938 586302 403174
rect 586538 402938 586622 403174
rect 586858 402938 586890 403174
rect 586270 402854 586890 402938
rect 586270 402618 586302 402854
rect 586538 402618 586622 402854
rect 586858 402618 586890 402854
rect 586270 367174 586890 402618
rect 586270 366938 586302 367174
rect 586538 366938 586622 367174
rect 586858 366938 586890 367174
rect 586270 366854 586890 366938
rect 586270 366618 586302 366854
rect 586538 366618 586622 366854
rect 586858 366618 586890 366854
rect 586270 331174 586890 366618
rect 586270 330938 586302 331174
rect 586538 330938 586622 331174
rect 586858 330938 586890 331174
rect 586270 330854 586890 330938
rect 586270 330618 586302 330854
rect 586538 330618 586622 330854
rect 586858 330618 586890 330854
rect 586270 295174 586890 330618
rect 586270 294938 586302 295174
rect 586538 294938 586622 295174
rect 586858 294938 586890 295174
rect 586270 294854 586890 294938
rect 586270 294618 586302 294854
rect 586538 294618 586622 294854
rect 586858 294618 586890 294854
rect 586270 259174 586890 294618
rect 586270 258938 586302 259174
rect 586538 258938 586622 259174
rect 586858 258938 586890 259174
rect 586270 258854 586890 258938
rect 586270 258618 586302 258854
rect 586538 258618 586622 258854
rect 586858 258618 586890 258854
rect 586270 223174 586890 258618
rect 586270 222938 586302 223174
rect 586538 222938 586622 223174
rect 586858 222938 586890 223174
rect 586270 222854 586890 222938
rect 586270 222618 586302 222854
rect 586538 222618 586622 222854
rect 586858 222618 586890 222854
rect 586270 187174 586890 222618
rect 586270 186938 586302 187174
rect 586538 186938 586622 187174
rect 586858 186938 586890 187174
rect 586270 186854 586890 186938
rect 586270 186618 586302 186854
rect 586538 186618 586622 186854
rect 586858 186618 586890 186854
rect 586270 151174 586890 186618
rect 586270 150938 586302 151174
rect 586538 150938 586622 151174
rect 586858 150938 586890 151174
rect 586270 150854 586890 150938
rect 586270 150618 586302 150854
rect 586538 150618 586622 150854
rect 586858 150618 586890 150854
rect 586270 115174 586890 150618
rect 586270 114938 586302 115174
rect 586538 114938 586622 115174
rect 586858 114938 586890 115174
rect 586270 114854 586890 114938
rect 586270 114618 586302 114854
rect 586538 114618 586622 114854
rect 586858 114618 586890 114854
rect 586270 79174 586890 114618
rect 586270 78938 586302 79174
rect 586538 78938 586622 79174
rect 586858 78938 586890 79174
rect 586270 78854 586890 78938
rect 586270 78618 586302 78854
rect 586538 78618 586622 78854
rect 586858 78618 586890 78854
rect 586270 43174 586890 78618
rect 586270 42938 586302 43174
rect 586538 42938 586622 43174
rect 586858 42938 586890 43174
rect 586270 42854 586890 42938
rect 586270 42618 586302 42854
rect 586538 42618 586622 42854
rect 586858 42618 586890 42854
rect 586270 7174 586890 42618
rect 586270 6938 586302 7174
rect 586538 6938 586622 7174
rect 586858 6938 586890 7174
rect 586270 6854 586890 6938
rect 586270 6618 586302 6854
rect 586538 6618 586622 6854
rect 586858 6618 586890 6854
rect 581514 -1542 581546 -1306
rect 581782 -1542 581866 -1306
rect 582102 -1542 582134 -1306
rect 581514 -1626 582134 -1542
rect 581514 -1862 581546 -1626
rect 581782 -1862 581866 -1626
rect 582102 -1862 582134 -1626
rect 581514 -7654 582134 -1862
rect 586270 -1306 586890 6618
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 694894 587850 706202
rect 587230 694658 587262 694894
rect 587498 694658 587582 694894
rect 587818 694658 587850 694894
rect 587230 694574 587850 694658
rect 587230 694338 587262 694574
rect 587498 694338 587582 694574
rect 587818 694338 587850 694574
rect 587230 658894 587850 694338
rect 587230 658658 587262 658894
rect 587498 658658 587582 658894
rect 587818 658658 587850 658894
rect 587230 658574 587850 658658
rect 587230 658338 587262 658574
rect 587498 658338 587582 658574
rect 587818 658338 587850 658574
rect 587230 622894 587850 658338
rect 587230 622658 587262 622894
rect 587498 622658 587582 622894
rect 587818 622658 587850 622894
rect 587230 622574 587850 622658
rect 587230 622338 587262 622574
rect 587498 622338 587582 622574
rect 587818 622338 587850 622574
rect 587230 586894 587850 622338
rect 587230 586658 587262 586894
rect 587498 586658 587582 586894
rect 587818 586658 587850 586894
rect 587230 586574 587850 586658
rect 587230 586338 587262 586574
rect 587498 586338 587582 586574
rect 587818 586338 587850 586574
rect 587230 550894 587850 586338
rect 587230 550658 587262 550894
rect 587498 550658 587582 550894
rect 587818 550658 587850 550894
rect 587230 550574 587850 550658
rect 587230 550338 587262 550574
rect 587498 550338 587582 550574
rect 587818 550338 587850 550574
rect 587230 514894 587850 550338
rect 587230 514658 587262 514894
rect 587498 514658 587582 514894
rect 587818 514658 587850 514894
rect 587230 514574 587850 514658
rect 587230 514338 587262 514574
rect 587498 514338 587582 514574
rect 587818 514338 587850 514574
rect 587230 478894 587850 514338
rect 587230 478658 587262 478894
rect 587498 478658 587582 478894
rect 587818 478658 587850 478894
rect 587230 478574 587850 478658
rect 587230 478338 587262 478574
rect 587498 478338 587582 478574
rect 587818 478338 587850 478574
rect 587230 442894 587850 478338
rect 587230 442658 587262 442894
rect 587498 442658 587582 442894
rect 587818 442658 587850 442894
rect 587230 442574 587850 442658
rect 587230 442338 587262 442574
rect 587498 442338 587582 442574
rect 587818 442338 587850 442574
rect 587230 406894 587850 442338
rect 587230 406658 587262 406894
rect 587498 406658 587582 406894
rect 587818 406658 587850 406894
rect 587230 406574 587850 406658
rect 587230 406338 587262 406574
rect 587498 406338 587582 406574
rect 587818 406338 587850 406574
rect 587230 370894 587850 406338
rect 587230 370658 587262 370894
rect 587498 370658 587582 370894
rect 587818 370658 587850 370894
rect 587230 370574 587850 370658
rect 587230 370338 587262 370574
rect 587498 370338 587582 370574
rect 587818 370338 587850 370574
rect 587230 334894 587850 370338
rect 587230 334658 587262 334894
rect 587498 334658 587582 334894
rect 587818 334658 587850 334894
rect 587230 334574 587850 334658
rect 587230 334338 587262 334574
rect 587498 334338 587582 334574
rect 587818 334338 587850 334574
rect 587230 298894 587850 334338
rect 587230 298658 587262 298894
rect 587498 298658 587582 298894
rect 587818 298658 587850 298894
rect 587230 298574 587850 298658
rect 587230 298338 587262 298574
rect 587498 298338 587582 298574
rect 587818 298338 587850 298574
rect 587230 262894 587850 298338
rect 587230 262658 587262 262894
rect 587498 262658 587582 262894
rect 587818 262658 587850 262894
rect 587230 262574 587850 262658
rect 587230 262338 587262 262574
rect 587498 262338 587582 262574
rect 587818 262338 587850 262574
rect 587230 226894 587850 262338
rect 587230 226658 587262 226894
rect 587498 226658 587582 226894
rect 587818 226658 587850 226894
rect 587230 226574 587850 226658
rect 587230 226338 587262 226574
rect 587498 226338 587582 226574
rect 587818 226338 587850 226574
rect 587230 190894 587850 226338
rect 587230 190658 587262 190894
rect 587498 190658 587582 190894
rect 587818 190658 587850 190894
rect 587230 190574 587850 190658
rect 587230 190338 587262 190574
rect 587498 190338 587582 190574
rect 587818 190338 587850 190574
rect 587230 154894 587850 190338
rect 587230 154658 587262 154894
rect 587498 154658 587582 154894
rect 587818 154658 587850 154894
rect 587230 154574 587850 154658
rect 587230 154338 587262 154574
rect 587498 154338 587582 154574
rect 587818 154338 587850 154574
rect 587230 118894 587850 154338
rect 587230 118658 587262 118894
rect 587498 118658 587582 118894
rect 587818 118658 587850 118894
rect 587230 118574 587850 118658
rect 587230 118338 587262 118574
rect 587498 118338 587582 118574
rect 587818 118338 587850 118574
rect 587230 82894 587850 118338
rect 587230 82658 587262 82894
rect 587498 82658 587582 82894
rect 587818 82658 587850 82894
rect 587230 82574 587850 82658
rect 587230 82338 587262 82574
rect 587498 82338 587582 82574
rect 587818 82338 587850 82574
rect 587230 46894 587850 82338
rect 587230 46658 587262 46894
rect 587498 46658 587582 46894
rect 587818 46658 587850 46894
rect 587230 46574 587850 46658
rect 587230 46338 587262 46574
rect 587498 46338 587582 46574
rect 587818 46338 587850 46574
rect 587230 10894 587850 46338
rect 587230 10658 587262 10894
rect 587498 10658 587582 10894
rect 587818 10658 587850 10894
rect 587230 10574 587850 10658
rect 587230 10338 587262 10574
rect 587498 10338 587582 10574
rect 587818 10338 587850 10574
rect 587230 -2266 587850 10338
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 698614 588810 707162
rect 588190 698378 588222 698614
rect 588458 698378 588542 698614
rect 588778 698378 588810 698614
rect 588190 698294 588810 698378
rect 588190 698058 588222 698294
rect 588458 698058 588542 698294
rect 588778 698058 588810 698294
rect 588190 662614 588810 698058
rect 588190 662378 588222 662614
rect 588458 662378 588542 662614
rect 588778 662378 588810 662614
rect 588190 662294 588810 662378
rect 588190 662058 588222 662294
rect 588458 662058 588542 662294
rect 588778 662058 588810 662294
rect 588190 626614 588810 662058
rect 588190 626378 588222 626614
rect 588458 626378 588542 626614
rect 588778 626378 588810 626614
rect 588190 626294 588810 626378
rect 588190 626058 588222 626294
rect 588458 626058 588542 626294
rect 588778 626058 588810 626294
rect 588190 590614 588810 626058
rect 588190 590378 588222 590614
rect 588458 590378 588542 590614
rect 588778 590378 588810 590614
rect 588190 590294 588810 590378
rect 588190 590058 588222 590294
rect 588458 590058 588542 590294
rect 588778 590058 588810 590294
rect 588190 554614 588810 590058
rect 588190 554378 588222 554614
rect 588458 554378 588542 554614
rect 588778 554378 588810 554614
rect 588190 554294 588810 554378
rect 588190 554058 588222 554294
rect 588458 554058 588542 554294
rect 588778 554058 588810 554294
rect 588190 518614 588810 554058
rect 588190 518378 588222 518614
rect 588458 518378 588542 518614
rect 588778 518378 588810 518614
rect 588190 518294 588810 518378
rect 588190 518058 588222 518294
rect 588458 518058 588542 518294
rect 588778 518058 588810 518294
rect 588190 482614 588810 518058
rect 588190 482378 588222 482614
rect 588458 482378 588542 482614
rect 588778 482378 588810 482614
rect 588190 482294 588810 482378
rect 588190 482058 588222 482294
rect 588458 482058 588542 482294
rect 588778 482058 588810 482294
rect 588190 446614 588810 482058
rect 588190 446378 588222 446614
rect 588458 446378 588542 446614
rect 588778 446378 588810 446614
rect 588190 446294 588810 446378
rect 588190 446058 588222 446294
rect 588458 446058 588542 446294
rect 588778 446058 588810 446294
rect 588190 410614 588810 446058
rect 588190 410378 588222 410614
rect 588458 410378 588542 410614
rect 588778 410378 588810 410614
rect 588190 410294 588810 410378
rect 588190 410058 588222 410294
rect 588458 410058 588542 410294
rect 588778 410058 588810 410294
rect 588190 374614 588810 410058
rect 588190 374378 588222 374614
rect 588458 374378 588542 374614
rect 588778 374378 588810 374614
rect 588190 374294 588810 374378
rect 588190 374058 588222 374294
rect 588458 374058 588542 374294
rect 588778 374058 588810 374294
rect 588190 338614 588810 374058
rect 588190 338378 588222 338614
rect 588458 338378 588542 338614
rect 588778 338378 588810 338614
rect 588190 338294 588810 338378
rect 588190 338058 588222 338294
rect 588458 338058 588542 338294
rect 588778 338058 588810 338294
rect 588190 302614 588810 338058
rect 588190 302378 588222 302614
rect 588458 302378 588542 302614
rect 588778 302378 588810 302614
rect 588190 302294 588810 302378
rect 588190 302058 588222 302294
rect 588458 302058 588542 302294
rect 588778 302058 588810 302294
rect 588190 266614 588810 302058
rect 588190 266378 588222 266614
rect 588458 266378 588542 266614
rect 588778 266378 588810 266614
rect 588190 266294 588810 266378
rect 588190 266058 588222 266294
rect 588458 266058 588542 266294
rect 588778 266058 588810 266294
rect 588190 230614 588810 266058
rect 588190 230378 588222 230614
rect 588458 230378 588542 230614
rect 588778 230378 588810 230614
rect 588190 230294 588810 230378
rect 588190 230058 588222 230294
rect 588458 230058 588542 230294
rect 588778 230058 588810 230294
rect 588190 194614 588810 230058
rect 588190 194378 588222 194614
rect 588458 194378 588542 194614
rect 588778 194378 588810 194614
rect 588190 194294 588810 194378
rect 588190 194058 588222 194294
rect 588458 194058 588542 194294
rect 588778 194058 588810 194294
rect 588190 158614 588810 194058
rect 588190 158378 588222 158614
rect 588458 158378 588542 158614
rect 588778 158378 588810 158614
rect 588190 158294 588810 158378
rect 588190 158058 588222 158294
rect 588458 158058 588542 158294
rect 588778 158058 588810 158294
rect 588190 122614 588810 158058
rect 588190 122378 588222 122614
rect 588458 122378 588542 122614
rect 588778 122378 588810 122614
rect 588190 122294 588810 122378
rect 588190 122058 588222 122294
rect 588458 122058 588542 122294
rect 588778 122058 588810 122294
rect 588190 86614 588810 122058
rect 588190 86378 588222 86614
rect 588458 86378 588542 86614
rect 588778 86378 588810 86614
rect 588190 86294 588810 86378
rect 588190 86058 588222 86294
rect 588458 86058 588542 86294
rect 588778 86058 588810 86294
rect 588190 50614 588810 86058
rect 588190 50378 588222 50614
rect 588458 50378 588542 50614
rect 588778 50378 588810 50614
rect 588190 50294 588810 50378
rect 588190 50058 588222 50294
rect 588458 50058 588542 50294
rect 588778 50058 588810 50294
rect 588190 14614 588810 50058
rect 588190 14378 588222 14614
rect 588458 14378 588542 14614
rect 588778 14378 588810 14614
rect 588190 14294 588810 14378
rect 588190 14058 588222 14294
rect 588458 14058 588542 14294
rect 588778 14058 588810 14294
rect 588190 -3226 588810 14058
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 666334 589770 708122
rect 589150 666098 589182 666334
rect 589418 666098 589502 666334
rect 589738 666098 589770 666334
rect 589150 666014 589770 666098
rect 589150 665778 589182 666014
rect 589418 665778 589502 666014
rect 589738 665778 589770 666014
rect 589150 630334 589770 665778
rect 589150 630098 589182 630334
rect 589418 630098 589502 630334
rect 589738 630098 589770 630334
rect 589150 630014 589770 630098
rect 589150 629778 589182 630014
rect 589418 629778 589502 630014
rect 589738 629778 589770 630014
rect 589150 594334 589770 629778
rect 589150 594098 589182 594334
rect 589418 594098 589502 594334
rect 589738 594098 589770 594334
rect 589150 594014 589770 594098
rect 589150 593778 589182 594014
rect 589418 593778 589502 594014
rect 589738 593778 589770 594014
rect 589150 558334 589770 593778
rect 589150 558098 589182 558334
rect 589418 558098 589502 558334
rect 589738 558098 589770 558334
rect 589150 558014 589770 558098
rect 589150 557778 589182 558014
rect 589418 557778 589502 558014
rect 589738 557778 589770 558014
rect 589150 522334 589770 557778
rect 589150 522098 589182 522334
rect 589418 522098 589502 522334
rect 589738 522098 589770 522334
rect 589150 522014 589770 522098
rect 589150 521778 589182 522014
rect 589418 521778 589502 522014
rect 589738 521778 589770 522014
rect 589150 486334 589770 521778
rect 589150 486098 589182 486334
rect 589418 486098 589502 486334
rect 589738 486098 589770 486334
rect 589150 486014 589770 486098
rect 589150 485778 589182 486014
rect 589418 485778 589502 486014
rect 589738 485778 589770 486014
rect 589150 450334 589770 485778
rect 589150 450098 589182 450334
rect 589418 450098 589502 450334
rect 589738 450098 589770 450334
rect 589150 450014 589770 450098
rect 589150 449778 589182 450014
rect 589418 449778 589502 450014
rect 589738 449778 589770 450014
rect 589150 414334 589770 449778
rect 589150 414098 589182 414334
rect 589418 414098 589502 414334
rect 589738 414098 589770 414334
rect 589150 414014 589770 414098
rect 589150 413778 589182 414014
rect 589418 413778 589502 414014
rect 589738 413778 589770 414014
rect 589150 378334 589770 413778
rect 589150 378098 589182 378334
rect 589418 378098 589502 378334
rect 589738 378098 589770 378334
rect 589150 378014 589770 378098
rect 589150 377778 589182 378014
rect 589418 377778 589502 378014
rect 589738 377778 589770 378014
rect 589150 342334 589770 377778
rect 589150 342098 589182 342334
rect 589418 342098 589502 342334
rect 589738 342098 589770 342334
rect 589150 342014 589770 342098
rect 589150 341778 589182 342014
rect 589418 341778 589502 342014
rect 589738 341778 589770 342014
rect 589150 306334 589770 341778
rect 589150 306098 589182 306334
rect 589418 306098 589502 306334
rect 589738 306098 589770 306334
rect 589150 306014 589770 306098
rect 589150 305778 589182 306014
rect 589418 305778 589502 306014
rect 589738 305778 589770 306014
rect 589150 270334 589770 305778
rect 589150 270098 589182 270334
rect 589418 270098 589502 270334
rect 589738 270098 589770 270334
rect 589150 270014 589770 270098
rect 589150 269778 589182 270014
rect 589418 269778 589502 270014
rect 589738 269778 589770 270014
rect 589150 234334 589770 269778
rect 589150 234098 589182 234334
rect 589418 234098 589502 234334
rect 589738 234098 589770 234334
rect 589150 234014 589770 234098
rect 589150 233778 589182 234014
rect 589418 233778 589502 234014
rect 589738 233778 589770 234014
rect 589150 198334 589770 233778
rect 589150 198098 589182 198334
rect 589418 198098 589502 198334
rect 589738 198098 589770 198334
rect 589150 198014 589770 198098
rect 589150 197778 589182 198014
rect 589418 197778 589502 198014
rect 589738 197778 589770 198014
rect 589150 162334 589770 197778
rect 589150 162098 589182 162334
rect 589418 162098 589502 162334
rect 589738 162098 589770 162334
rect 589150 162014 589770 162098
rect 589150 161778 589182 162014
rect 589418 161778 589502 162014
rect 589738 161778 589770 162014
rect 589150 126334 589770 161778
rect 589150 126098 589182 126334
rect 589418 126098 589502 126334
rect 589738 126098 589770 126334
rect 589150 126014 589770 126098
rect 589150 125778 589182 126014
rect 589418 125778 589502 126014
rect 589738 125778 589770 126014
rect 589150 90334 589770 125778
rect 589150 90098 589182 90334
rect 589418 90098 589502 90334
rect 589738 90098 589770 90334
rect 589150 90014 589770 90098
rect 589150 89778 589182 90014
rect 589418 89778 589502 90014
rect 589738 89778 589770 90014
rect 589150 54334 589770 89778
rect 589150 54098 589182 54334
rect 589418 54098 589502 54334
rect 589738 54098 589770 54334
rect 589150 54014 589770 54098
rect 589150 53778 589182 54014
rect 589418 53778 589502 54014
rect 589738 53778 589770 54014
rect 589150 18334 589770 53778
rect 589150 18098 589182 18334
rect 589418 18098 589502 18334
rect 589738 18098 589770 18334
rect 589150 18014 589770 18098
rect 589150 17778 589182 18014
rect 589418 17778 589502 18014
rect 589738 17778 589770 18014
rect 589150 -4186 589770 17778
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 670054 590730 709082
rect 590110 669818 590142 670054
rect 590378 669818 590462 670054
rect 590698 669818 590730 670054
rect 590110 669734 590730 669818
rect 590110 669498 590142 669734
rect 590378 669498 590462 669734
rect 590698 669498 590730 669734
rect 590110 634054 590730 669498
rect 590110 633818 590142 634054
rect 590378 633818 590462 634054
rect 590698 633818 590730 634054
rect 590110 633734 590730 633818
rect 590110 633498 590142 633734
rect 590378 633498 590462 633734
rect 590698 633498 590730 633734
rect 590110 598054 590730 633498
rect 590110 597818 590142 598054
rect 590378 597818 590462 598054
rect 590698 597818 590730 598054
rect 590110 597734 590730 597818
rect 590110 597498 590142 597734
rect 590378 597498 590462 597734
rect 590698 597498 590730 597734
rect 590110 562054 590730 597498
rect 590110 561818 590142 562054
rect 590378 561818 590462 562054
rect 590698 561818 590730 562054
rect 590110 561734 590730 561818
rect 590110 561498 590142 561734
rect 590378 561498 590462 561734
rect 590698 561498 590730 561734
rect 590110 526054 590730 561498
rect 590110 525818 590142 526054
rect 590378 525818 590462 526054
rect 590698 525818 590730 526054
rect 590110 525734 590730 525818
rect 590110 525498 590142 525734
rect 590378 525498 590462 525734
rect 590698 525498 590730 525734
rect 590110 490054 590730 525498
rect 590110 489818 590142 490054
rect 590378 489818 590462 490054
rect 590698 489818 590730 490054
rect 590110 489734 590730 489818
rect 590110 489498 590142 489734
rect 590378 489498 590462 489734
rect 590698 489498 590730 489734
rect 590110 454054 590730 489498
rect 590110 453818 590142 454054
rect 590378 453818 590462 454054
rect 590698 453818 590730 454054
rect 590110 453734 590730 453818
rect 590110 453498 590142 453734
rect 590378 453498 590462 453734
rect 590698 453498 590730 453734
rect 590110 418054 590730 453498
rect 590110 417818 590142 418054
rect 590378 417818 590462 418054
rect 590698 417818 590730 418054
rect 590110 417734 590730 417818
rect 590110 417498 590142 417734
rect 590378 417498 590462 417734
rect 590698 417498 590730 417734
rect 590110 382054 590730 417498
rect 590110 381818 590142 382054
rect 590378 381818 590462 382054
rect 590698 381818 590730 382054
rect 590110 381734 590730 381818
rect 590110 381498 590142 381734
rect 590378 381498 590462 381734
rect 590698 381498 590730 381734
rect 590110 346054 590730 381498
rect 590110 345818 590142 346054
rect 590378 345818 590462 346054
rect 590698 345818 590730 346054
rect 590110 345734 590730 345818
rect 590110 345498 590142 345734
rect 590378 345498 590462 345734
rect 590698 345498 590730 345734
rect 590110 310054 590730 345498
rect 590110 309818 590142 310054
rect 590378 309818 590462 310054
rect 590698 309818 590730 310054
rect 590110 309734 590730 309818
rect 590110 309498 590142 309734
rect 590378 309498 590462 309734
rect 590698 309498 590730 309734
rect 590110 274054 590730 309498
rect 590110 273818 590142 274054
rect 590378 273818 590462 274054
rect 590698 273818 590730 274054
rect 590110 273734 590730 273818
rect 590110 273498 590142 273734
rect 590378 273498 590462 273734
rect 590698 273498 590730 273734
rect 590110 238054 590730 273498
rect 590110 237818 590142 238054
rect 590378 237818 590462 238054
rect 590698 237818 590730 238054
rect 590110 237734 590730 237818
rect 590110 237498 590142 237734
rect 590378 237498 590462 237734
rect 590698 237498 590730 237734
rect 590110 202054 590730 237498
rect 590110 201818 590142 202054
rect 590378 201818 590462 202054
rect 590698 201818 590730 202054
rect 590110 201734 590730 201818
rect 590110 201498 590142 201734
rect 590378 201498 590462 201734
rect 590698 201498 590730 201734
rect 590110 166054 590730 201498
rect 590110 165818 590142 166054
rect 590378 165818 590462 166054
rect 590698 165818 590730 166054
rect 590110 165734 590730 165818
rect 590110 165498 590142 165734
rect 590378 165498 590462 165734
rect 590698 165498 590730 165734
rect 590110 130054 590730 165498
rect 590110 129818 590142 130054
rect 590378 129818 590462 130054
rect 590698 129818 590730 130054
rect 590110 129734 590730 129818
rect 590110 129498 590142 129734
rect 590378 129498 590462 129734
rect 590698 129498 590730 129734
rect 590110 94054 590730 129498
rect 590110 93818 590142 94054
rect 590378 93818 590462 94054
rect 590698 93818 590730 94054
rect 590110 93734 590730 93818
rect 590110 93498 590142 93734
rect 590378 93498 590462 93734
rect 590698 93498 590730 93734
rect 590110 58054 590730 93498
rect 590110 57818 590142 58054
rect 590378 57818 590462 58054
rect 590698 57818 590730 58054
rect 590110 57734 590730 57818
rect 590110 57498 590142 57734
rect 590378 57498 590462 57734
rect 590698 57498 590730 57734
rect 590110 22054 590730 57498
rect 590110 21818 590142 22054
rect 590378 21818 590462 22054
rect 590698 21818 590730 22054
rect 590110 21734 590730 21818
rect 590110 21498 590142 21734
rect 590378 21498 590462 21734
rect 590698 21498 590730 21734
rect 590110 -5146 590730 21498
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 673774 591690 710042
rect 591070 673538 591102 673774
rect 591338 673538 591422 673774
rect 591658 673538 591690 673774
rect 591070 673454 591690 673538
rect 591070 673218 591102 673454
rect 591338 673218 591422 673454
rect 591658 673218 591690 673454
rect 591070 637774 591690 673218
rect 591070 637538 591102 637774
rect 591338 637538 591422 637774
rect 591658 637538 591690 637774
rect 591070 637454 591690 637538
rect 591070 637218 591102 637454
rect 591338 637218 591422 637454
rect 591658 637218 591690 637454
rect 591070 601774 591690 637218
rect 591070 601538 591102 601774
rect 591338 601538 591422 601774
rect 591658 601538 591690 601774
rect 591070 601454 591690 601538
rect 591070 601218 591102 601454
rect 591338 601218 591422 601454
rect 591658 601218 591690 601454
rect 591070 565774 591690 601218
rect 591070 565538 591102 565774
rect 591338 565538 591422 565774
rect 591658 565538 591690 565774
rect 591070 565454 591690 565538
rect 591070 565218 591102 565454
rect 591338 565218 591422 565454
rect 591658 565218 591690 565454
rect 591070 529774 591690 565218
rect 591070 529538 591102 529774
rect 591338 529538 591422 529774
rect 591658 529538 591690 529774
rect 591070 529454 591690 529538
rect 591070 529218 591102 529454
rect 591338 529218 591422 529454
rect 591658 529218 591690 529454
rect 591070 493774 591690 529218
rect 591070 493538 591102 493774
rect 591338 493538 591422 493774
rect 591658 493538 591690 493774
rect 591070 493454 591690 493538
rect 591070 493218 591102 493454
rect 591338 493218 591422 493454
rect 591658 493218 591690 493454
rect 591070 457774 591690 493218
rect 591070 457538 591102 457774
rect 591338 457538 591422 457774
rect 591658 457538 591690 457774
rect 591070 457454 591690 457538
rect 591070 457218 591102 457454
rect 591338 457218 591422 457454
rect 591658 457218 591690 457454
rect 591070 421774 591690 457218
rect 591070 421538 591102 421774
rect 591338 421538 591422 421774
rect 591658 421538 591690 421774
rect 591070 421454 591690 421538
rect 591070 421218 591102 421454
rect 591338 421218 591422 421454
rect 591658 421218 591690 421454
rect 591070 385774 591690 421218
rect 591070 385538 591102 385774
rect 591338 385538 591422 385774
rect 591658 385538 591690 385774
rect 591070 385454 591690 385538
rect 591070 385218 591102 385454
rect 591338 385218 591422 385454
rect 591658 385218 591690 385454
rect 591070 349774 591690 385218
rect 591070 349538 591102 349774
rect 591338 349538 591422 349774
rect 591658 349538 591690 349774
rect 591070 349454 591690 349538
rect 591070 349218 591102 349454
rect 591338 349218 591422 349454
rect 591658 349218 591690 349454
rect 591070 313774 591690 349218
rect 591070 313538 591102 313774
rect 591338 313538 591422 313774
rect 591658 313538 591690 313774
rect 591070 313454 591690 313538
rect 591070 313218 591102 313454
rect 591338 313218 591422 313454
rect 591658 313218 591690 313454
rect 591070 277774 591690 313218
rect 591070 277538 591102 277774
rect 591338 277538 591422 277774
rect 591658 277538 591690 277774
rect 591070 277454 591690 277538
rect 591070 277218 591102 277454
rect 591338 277218 591422 277454
rect 591658 277218 591690 277454
rect 591070 241774 591690 277218
rect 591070 241538 591102 241774
rect 591338 241538 591422 241774
rect 591658 241538 591690 241774
rect 591070 241454 591690 241538
rect 591070 241218 591102 241454
rect 591338 241218 591422 241454
rect 591658 241218 591690 241454
rect 591070 205774 591690 241218
rect 591070 205538 591102 205774
rect 591338 205538 591422 205774
rect 591658 205538 591690 205774
rect 591070 205454 591690 205538
rect 591070 205218 591102 205454
rect 591338 205218 591422 205454
rect 591658 205218 591690 205454
rect 591070 169774 591690 205218
rect 591070 169538 591102 169774
rect 591338 169538 591422 169774
rect 591658 169538 591690 169774
rect 591070 169454 591690 169538
rect 591070 169218 591102 169454
rect 591338 169218 591422 169454
rect 591658 169218 591690 169454
rect 591070 133774 591690 169218
rect 591070 133538 591102 133774
rect 591338 133538 591422 133774
rect 591658 133538 591690 133774
rect 591070 133454 591690 133538
rect 591070 133218 591102 133454
rect 591338 133218 591422 133454
rect 591658 133218 591690 133454
rect 591070 97774 591690 133218
rect 591070 97538 591102 97774
rect 591338 97538 591422 97774
rect 591658 97538 591690 97774
rect 591070 97454 591690 97538
rect 591070 97218 591102 97454
rect 591338 97218 591422 97454
rect 591658 97218 591690 97454
rect 591070 61774 591690 97218
rect 591070 61538 591102 61774
rect 591338 61538 591422 61774
rect 591658 61538 591690 61774
rect 591070 61454 591690 61538
rect 591070 61218 591102 61454
rect 591338 61218 591422 61454
rect 591658 61218 591690 61454
rect 591070 25774 591690 61218
rect 591070 25538 591102 25774
rect 591338 25538 591422 25774
rect 591658 25538 591690 25774
rect 591070 25454 591690 25538
rect 591070 25218 591102 25454
rect 591338 25218 591422 25454
rect 591658 25218 591690 25454
rect 591070 -6106 591690 25218
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 677494 592650 711002
rect 592030 677258 592062 677494
rect 592298 677258 592382 677494
rect 592618 677258 592650 677494
rect 592030 677174 592650 677258
rect 592030 676938 592062 677174
rect 592298 676938 592382 677174
rect 592618 676938 592650 677174
rect 592030 641494 592650 676938
rect 592030 641258 592062 641494
rect 592298 641258 592382 641494
rect 592618 641258 592650 641494
rect 592030 641174 592650 641258
rect 592030 640938 592062 641174
rect 592298 640938 592382 641174
rect 592618 640938 592650 641174
rect 592030 605494 592650 640938
rect 592030 605258 592062 605494
rect 592298 605258 592382 605494
rect 592618 605258 592650 605494
rect 592030 605174 592650 605258
rect 592030 604938 592062 605174
rect 592298 604938 592382 605174
rect 592618 604938 592650 605174
rect 592030 569494 592650 604938
rect 592030 569258 592062 569494
rect 592298 569258 592382 569494
rect 592618 569258 592650 569494
rect 592030 569174 592650 569258
rect 592030 568938 592062 569174
rect 592298 568938 592382 569174
rect 592618 568938 592650 569174
rect 592030 533494 592650 568938
rect 592030 533258 592062 533494
rect 592298 533258 592382 533494
rect 592618 533258 592650 533494
rect 592030 533174 592650 533258
rect 592030 532938 592062 533174
rect 592298 532938 592382 533174
rect 592618 532938 592650 533174
rect 592030 497494 592650 532938
rect 592030 497258 592062 497494
rect 592298 497258 592382 497494
rect 592618 497258 592650 497494
rect 592030 497174 592650 497258
rect 592030 496938 592062 497174
rect 592298 496938 592382 497174
rect 592618 496938 592650 497174
rect 592030 461494 592650 496938
rect 592030 461258 592062 461494
rect 592298 461258 592382 461494
rect 592618 461258 592650 461494
rect 592030 461174 592650 461258
rect 592030 460938 592062 461174
rect 592298 460938 592382 461174
rect 592618 460938 592650 461174
rect 592030 425494 592650 460938
rect 592030 425258 592062 425494
rect 592298 425258 592382 425494
rect 592618 425258 592650 425494
rect 592030 425174 592650 425258
rect 592030 424938 592062 425174
rect 592298 424938 592382 425174
rect 592618 424938 592650 425174
rect 592030 389494 592650 424938
rect 592030 389258 592062 389494
rect 592298 389258 592382 389494
rect 592618 389258 592650 389494
rect 592030 389174 592650 389258
rect 592030 388938 592062 389174
rect 592298 388938 592382 389174
rect 592618 388938 592650 389174
rect 592030 353494 592650 388938
rect 592030 353258 592062 353494
rect 592298 353258 592382 353494
rect 592618 353258 592650 353494
rect 592030 353174 592650 353258
rect 592030 352938 592062 353174
rect 592298 352938 592382 353174
rect 592618 352938 592650 353174
rect 592030 317494 592650 352938
rect 592030 317258 592062 317494
rect 592298 317258 592382 317494
rect 592618 317258 592650 317494
rect 592030 317174 592650 317258
rect 592030 316938 592062 317174
rect 592298 316938 592382 317174
rect 592618 316938 592650 317174
rect 592030 281494 592650 316938
rect 592030 281258 592062 281494
rect 592298 281258 592382 281494
rect 592618 281258 592650 281494
rect 592030 281174 592650 281258
rect 592030 280938 592062 281174
rect 592298 280938 592382 281174
rect 592618 280938 592650 281174
rect 592030 245494 592650 280938
rect 592030 245258 592062 245494
rect 592298 245258 592382 245494
rect 592618 245258 592650 245494
rect 592030 245174 592650 245258
rect 592030 244938 592062 245174
rect 592298 244938 592382 245174
rect 592618 244938 592650 245174
rect 592030 209494 592650 244938
rect 592030 209258 592062 209494
rect 592298 209258 592382 209494
rect 592618 209258 592650 209494
rect 592030 209174 592650 209258
rect 592030 208938 592062 209174
rect 592298 208938 592382 209174
rect 592618 208938 592650 209174
rect 592030 173494 592650 208938
rect 592030 173258 592062 173494
rect 592298 173258 592382 173494
rect 592618 173258 592650 173494
rect 592030 173174 592650 173258
rect 592030 172938 592062 173174
rect 592298 172938 592382 173174
rect 592618 172938 592650 173174
rect 592030 137494 592650 172938
rect 592030 137258 592062 137494
rect 592298 137258 592382 137494
rect 592618 137258 592650 137494
rect 592030 137174 592650 137258
rect 592030 136938 592062 137174
rect 592298 136938 592382 137174
rect 592618 136938 592650 137174
rect 592030 101494 592650 136938
rect 592030 101258 592062 101494
rect 592298 101258 592382 101494
rect 592618 101258 592650 101494
rect 592030 101174 592650 101258
rect 592030 100938 592062 101174
rect 592298 100938 592382 101174
rect 592618 100938 592650 101174
rect 592030 65494 592650 100938
rect 592030 65258 592062 65494
rect 592298 65258 592382 65494
rect 592618 65258 592650 65494
rect 592030 65174 592650 65258
rect 592030 64938 592062 65174
rect 592298 64938 592382 65174
rect 592618 64938 592650 65174
rect 592030 29494 592650 64938
rect 592030 29258 592062 29494
rect 592298 29258 592382 29494
rect 592618 29258 592650 29494
rect 592030 29174 592650 29258
rect 592030 28938 592062 29174
rect 592298 28938 592382 29174
rect 592618 28938 592650 29174
rect 592030 -7066 592650 28938
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -8694 677258 -8458 677494
rect -8374 677258 -8138 677494
rect -8694 676938 -8458 677174
rect -8374 676938 -8138 677174
rect -8694 641258 -8458 641494
rect -8374 641258 -8138 641494
rect -8694 640938 -8458 641174
rect -8374 640938 -8138 641174
rect -8694 605258 -8458 605494
rect -8374 605258 -8138 605494
rect -8694 604938 -8458 605174
rect -8374 604938 -8138 605174
rect -8694 569258 -8458 569494
rect -8374 569258 -8138 569494
rect -8694 568938 -8458 569174
rect -8374 568938 -8138 569174
rect -8694 533258 -8458 533494
rect -8374 533258 -8138 533494
rect -8694 532938 -8458 533174
rect -8374 532938 -8138 533174
rect -8694 497258 -8458 497494
rect -8374 497258 -8138 497494
rect -8694 496938 -8458 497174
rect -8374 496938 -8138 497174
rect -8694 461258 -8458 461494
rect -8374 461258 -8138 461494
rect -8694 460938 -8458 461174
rect -8374 460938 -8138 461174
rect -8694 425258 -8458 425494
rect -8374 425258 -8138 425494
rect -8694 424938 -8458 425174
rect -8374 424938 -8138 425174
rect -8694 389258 -8458 389494
rect -8374 389258 -8138 389494
rect -8694 388938 -8458 389174
rect -8374 388938 -8138 389174
rect -8694 353258 -8458 353494
rect -8374 353258 -8138 353494
rect -8694 352938 -8458 353174
rect -8374 352938 -8138 353174
rect -8694 317258 -8458 317494
rect -8374 317258 -8138 317494
rect -8694 316938 -8458 317174
rect -8374 316938 -8138 317174
rect -8694 281258 -8458 281494
rect -8374 281258 -8138 281494
rect -8694 280938 -8458 281174
rect -8374 280938 -8138 281174
rect -8694 245258 -8458 245494
rect -8374 245258 -8138 245494
rect -8694 244938 -8458 245174
rect -8374 244938 -8138 245174
rect -8694 209258 -8458 209494
rect -8374 209258 -8138 209494
rect -8694 208938 -8458 209174
rect -8374 208938 -8138 209174
rect -8694 173258 -8458 173494
rect -8374 173258 -8138 173494
rect -8694 172938 -8458 173174
rect -8374 172938 -8138 173174
rect -8694 137258 -8458 137494
rect -8374 137258 -8138 137494
rect -8694 136938 -8458 137174
rect -8374 136938 -8138 137174
rect -8694 101258 -8458 101494
rect -8374 101258 -8138 101494
rect -8694 100938 -8458 101174
rect -8374 100938 -8138 101174
rect -8694 65258 -8458 65494
rect -8374 65258 -8138 65494
rect -8694 64938 -8458 65174
rect -8374 64938 -8138 65174
rect -8694 29258 -8458 29494
rect -8374 29258 -8138 29494
rect -8694 28938 -8458 29174
rect -8374 28938 -8138 29174
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect -7734 673538 -7498 673774
rect -7414 673538 -7178 673774
rect -7734 673218 -7498 673454
rect -7414 673218 -7178 673454
rect -7734 637538 -7498 637774
rect -7414 637538 -7178 637774
rect -7734 637218 -7498 637454
rect -7414 637218 -7178 637454
rect -7734 601538 -7498 601774
rect -7414 601538 -7178 601774
rect -7734 601218 -7498 601454
rect -7414 601218 -7178 601454
rect -7734 565538 -7498 565774
rect -7414 565538 -7178 565774
rect -7734 565218 -7498 565454
rect -7414 565218 -7178 565454
rect -7734 529538 -7498 529774
rect -7414 529538 -7178 529774
rect -7734 529218 -7498 529454
rect -7414 529218 -7178 529454
rect -7734 493538 -7498 493774
rect -7414 493538 -7178 493774
rect -7734 493218 -7498 493454
rect -7414 493218 -7178 493454
rect -7734 457538 -7498 457774
rect -7414 457538 -7178 457774
rect -7734 457218 -7498 457454
rect -7414 457218 -7178 457454
rect -7734 421538 -7498 421774
rect -7414 421538 -7178 421774
rect -7734 421218 -7498 421454
rect -7414 421218 -7178 421454
rect -7734 385538 -7498 385774
rect -7414 385538 -7178 385774
rect -7734 385218 -7498 385454
rect -7414 385218 -7178 385454
rect -7734 349538 -7498 349774
rect -7414 349538 -7178 349774
rect -7734 349218 -7498 349454
rect -7414 349218 -7178 349454
rect -7734 313538 -7498 313774
rect -7414 313538 -7178 313774
rect -7734 313218 -7498 313454
rect -7414 313218 -7178 313454
rect -7734 277538 -7498 277774
rect -7414 277538 -7178 277774
rect -7734 277218 -7498 277454
rect -7414 277218 -7178 277454
rect -7734 241538 -7498 241774
rect -7414 241538 -7178 241774
rect -7734 241218 -7498 241454
rect -7414 241218 -7178 241454
rect -7734 205538 -7498 205774
rect -7414 205538 -7178 205774
rect -7734 205218 -7498 205454
rect -7414 205218 -7178 205454
rect -7734 169538 -7498 169774
rect -7414 169538 -7178 169774
rect -7734 169218 -7498 169454
rect -7414 169218 -7178 169454
rect -7734 133538 -7498 133774
rect -7414 133538 -7178 133774
rect -7734 133218 -7498 133454
rect -7414 133218 -7178 133454
rect -7734 97538 -7498 97774
rect -7414 97538 -7178 97774
rect -7734 97218 -7498 97454
rect -7414 97218 -7178 97454
rect -7734 61538 -7498 61774
rect -7414 61538 -7178 61774
rect -7734 61218 -7498 61454
rect -7414 61218 -7178 61454
rect -7734 25538 -7498 25774
rect -7414 25538 -7178 25774
rect -7734 25218 -7498 25454
rect -7414 25218 -7178 25454
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -6774 669818 -6538 670054
rect -6454 669818 -6218 670054
rect -6774 669498 -6538 669734
rect -6454 669498 -6218 669734
rect -6774 633818 -6538 634054
rect -6454 633818 -6218 634054
rect -6774 633498 -6538 633734
rect -6454 633498 -6218 633734
rect -6774 597818 -6538 598054
rect -6454 597818 -6218 598054
rect -6774 597498 -6538 597734
rect -6454 597498 -6218 597734
rect -6774 561818 -6538 562054
rect -6454 561818 -6218 562054
rect -6774 561498 -6538 561734
rect -6454 561498 -6218 561734
rect -6774 525818 -6538 526054
rect -6454 525818 -6218 526054
rect -6774 525498 -6538 525734
rect -6454 525498 -6218 525734
rect -6774 489818 -6538 490054
rect -6454 489818 -6218 490054
rect -6774 489498 -6538 489734
rect -6454 489498 -6218 489734
rect -6774 453818 -6538 454054
rect -6454 453818 -6218 454054
rect -6774 453498 -6538 453734
rect -6454 453498 -6218 453734
rect -6774 417818 -6538 418054
rect -6454 417818 -6218 418054
rect -6774 417498 -6538 417734
rect -6454 417498 -6218 417734
rect -6774 381818 -6538 382054
rect -6454 381818 -6218 382054
rect -6774 381498 -6538 381734
rect -6454 381498 -6218 381734
rect -6774 345818 -6538 346054
rect -6454 345818 -6218 346054
rect -6774 345498 -6538 345734
rect -6454 345498 -6218 345734
rect -6774 309818 -6538 310054
rect -6454 309818 -6218 310054
rect -6774 309498 -6538 309734
rect -6454 309498 -6218 309734
rect -6774 273818 -6538 274054
rect -6454 273818 -6218 274054
rect -6774 273498 -6538 273734
rect -6454 273498 -6218 273734
rect -6774 237818 -6538 238054
rect -6454 237818 -6218 238054
rect -6774 237498 -6538 237734
rect -6454 237498 -6218 237734
rect -6774 201818 -6538 202054
rect -6454 201818 -6218 202054
rect -6774 201498 -6538 201734
rect -6454 201498 -6218 201734
rect -6774 165818 -6538 166054
rect -6454 165818 -6218 166054
rect -6774 165498 -6538 165734
rect -6454 165498 -6218 165734
rect -6774 129818 -6538 130054
rect -6454 129818 -6218 130054
rect -6774 129498 -6538 129734
rect -6454 129498 -6218 129734
rect -6774 93818 -6538 94054
rect -6454 93818 -6218 94054
rect -6774 93498 -6538 93734
rect -6454 93498 -6218 93734
rect -6774 57818 -6538 58054
rect -6454 57818 -6218 58054
rect -6774 57498 -6538 57734
rect -6454 57498 -6218 57734
rect -6774 21818 -6538 22054
rect -6454 21818 -6218 22054
rect -6774 21498 -6538 21734
rect -6454 21498 -6218 21734
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect -5814 666098 -5578 666334
rect -5494 666098 -5258 666334
rect -5814 665778 -5578 666014
rect -5494 665778 -5258 666014
rect -5814 630098 -5578 630334
rect -5494 630098 -5258 630334
rect -5814 629778 -5578 630014
rect -5494 629778 -5258 630014
rect -5814 594098 -5578 594334
rect -5494 594098 -5258 594334
rect -5814 593778 -5578 594014
rect -5494 593778 -5258 594014
rect -5814 558098 -5578 558334
rect -5494 558098 -5258 558334
rect -5814 557778 -5578 558014
rect -5494 557778 -5258 558014
rect -5814 522098 -5578 522334
rect -5494 522098 -5258 522334
rect -5814 521778 -5578 522014
rect -5494 521778 -5258 522014
rect -5814 486098 -5578 486334
rect -5494 486098 -5258 486334
rect -5814 485778 -5578 486014
rect -5494 485778 -5258 486014
rect -5814 450098 -5578 450334
rect -5494 450098 -5258 450334
rect -5814 449778 -5578 450014
rect -5494 449778 -5258 450014
rect -5814 414098 -5578 414334
rect -5494 414098 -5258 414334
rect -5814 413778 -5578 414014
rect -5494 413778 -5258 414014
rect -5814 378098 -5578 378334
rect -5494 378098 -5258 378334
rect -5814 377778 -5578 378014
rect -5494 377778 -5258 378014
rect -5814 342098 -5578 342334
rect -5494 342098 -5258 342334
rect -5814 341778 -5578 342014
rect -5494 341778 -5258 342014
rect -5814 306098 -5578 306334
rect -5494 306098 -5258 306334
rect -5814 305778 -5578 306014
rect -5494 305778 -5258 306014
rect -5814 270098 -5578 270334
rect -5494 270098 -5258 270334
rect -5814 269778 -5578 270014
rect -5494 269778 -5258 270014
rect -5814 234098 -5578 234334
rect -5494 234098 -5258 234334
rect -5814 233778 -5578 234014
rect -5494 233778 -5258 234014
rect -5814 198098 -5578 198334
rect -5494 198098 -5258 198334
rect -5814 197778 -5578 198014
rect -5494 197778 -5258 198014
rect -5814 162098 -5578 162334
rect -5494 162098 -5258 162334
rect -5814 161778 -5578 162014
rect -5494 161778 -5258 162014
rect -5814 126098 -5578 126334
rect -5494 126098 -5258 126334
rect -5814 125778 -5578 126014
rect -5494 125778 -5258 126014
rect -5814 90098 -5578 90334
rect -5494 90098 -5258 90334
rect -5814 89778 -5578 90014
rect -5494 89778 -5258 90014
rect -5814 54098 -5578 54334
rect -5494 54098 -5258 54334
rect -5814 53778 -5578 54014
rect -5494 53778 -5258 54014
rect -5814 18098 -5578 18334
rect -5494 18098 -5258 18334
rect -5814 17778 -5578 18014
rect -5494 17778 -5258 18014
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -4854 698378 -4618 698614
rect -4534 698378 -4298 698614
rect -4854 698058 -4618 698294
rect -4534 698058 -4298 698294
rect -4854 662378 -4618 662614
rect -4534 662378 -4298 662614
rect -4854 662058 -4618 662294
rect -4534 662058 -4298 662294
rect -4854 626378 -4618 626614
rect -4534 626378 -4298 626614
rect -4854 626058 -4618 626294
rect -4534 626058 -4298 626294
rect -4854 590378 -4618 590614
rect -4534 590378 -4298 590614
rect -4854 590058 -4618 590294
rect -4534 590058 -4298 590294
rect -4854 554378 -4618 554614
rect -4534 554378 -4298 554614
rect -4854 554058 -4618 554294
rect -4534 554058 -4298 554294
rect -4854 518378 -4618 518614
rect -4534 518378 -4298 518614
rect -4854 518058 -4618 518294
rect -4534 518058 -4298 518294
rect -4854 482378 -4618 482614
rect -4534 482378 -4298 482614
rect -4854 482058 -4618 482294
rect -4534 482058 -4298 482294
rect -4854 446378 -4618 446614
rect -4534 446378 -4298 446614
rect -4854 446058 -4618 446294
rect -4534 446058 -4298 446294
rect -4854 410378 -4618 410614
rect -4534 410378 -4298 410614
rect -4854 410058 -4618 410294
rect -4534 410058 -4298 410294
rect -4854 374378 -4618 374614
rect -4534 374378 -4298 374614
rect -4854 374058 -4618 374294
rect -4534 374058 -4298 374294
rect -4854 338378 -4618 338614
rect -4534 338378 -4298 338614
rect -4854 338058 -4618 338294
rect -4534 338058 -4298 338294
rect -4854 302378 -4618 302614
rect -4534 302378 -4298 302614
rect -4854 302058 -4618 302294
rect -4534 302058 -4298 302294
rect -4854 266378 -4618 266614
rect -4534 266378 -4298 266614
rect -4854 266058 -4618 266294
rect -4534 266058 -4298 266294
rect -4854 230378 -4618 230614
rect -4534 230378 -4298 230614
rect -4854 230058 -4618 230294
rect -4534 230058 -4298 230294
rect -4854 194378 -4618 194614
rect -4534 194378 -4298 194614
rect -4854 194058 -4618 194294
rect -4534 194058 -4298 194294
rect -4854 158378 -4618 158614
rect -4534 158378 -4298 158614
rect -4854 158058 -4618 158294
rect -4534 158058 -4298 158294
rect -4854 122378 -4618 122614
rect -4534 122378 -4298 122614
rect -4854 122058 -4618 122294
rect -4534 122058 -4298 122294
rect -4854 86378 -4618 86614
rect -4534 86378 -4298 86614
rect -4854 86058 -4618 86294
rect -4534 86058 -4298 86294
rect -4854 50378 -4618 50614
rect -4534 50378 -4298 50614
rect -4854 50058 -4618 50294
rect -4534 50058 -4298 50294
rect -4854 14378 -4618 14614
rect -4534 14378 -4298 14614
rect -4854 14058 -4618 14294
rect -4534 14058 -4298 14294
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect -3894 694658 -3658 694894
rect -3574 694658 -3338 694894
rect -3894 694338 -3658 694574
rect -3574 694338 -3338 694574
rect -3894 658658 -3658 658894
rect -3574 658658 -3338 658894
rect -3894 658338 -3658 658574
rect -3574 658338 -3338 658574
rect -3894 622658 -3658 622894
rect -3574 622658 -3338 622894
rect -3894 622338 -3658 622574
rect -3574 622338 -3338 622574
rect -3894 586658 -3658 586894
rect -3574 586658 -3338 586894
rect -3894 586338 -3658 586574
rect -3574 586338 -3338 586574
rect -3894 550658 -3658 550894
rect -3574 550658 -3338 550894
rect -3894 550338 -3658 550574
rect -3574 550338 -3338 550574
rect -3894 514658 -3658 514894
rect -3574 514658 -3338 514894
rect -3894 514338 -3658 514574
rect -3574 514338 -3338 514574
rect -3894 478658 -3658 478894
rect -3574 478658 -3338 478894
rect -3894 478338 -3658 478574
rect -3574 478338 -3338 478574
rect -3894 442658 -3658 442894
rect -3574 442658 -3338 442894
rect -3894 442338 -3658 442574
rect -3574 442338 -3338 442574
rect -3894 406658 -3658 406894
rect -3574 406658 -3338 406894
rect -3894 406338 -3658 406574
rect -3574 406338 -3338 406574
rect -3894 370658 -3658 370894
rect -3574 370658 -3338 370894
rect -3894 370338 -3658 370574
rect -3574 370338 -3338 370574
rect -3894 334658 -3658 334894
rect -3574 334658 -3338 334894
rect -3894 334338 -3658 334574
rect -3574 334338 -3338 334574
rect -3894 298658 -3658 298894
rect -3574 298658 -3338 298894
rect -3894 298338 -3658 298574
rect -3574 298338 -3338 298574
rect -3894 262658 -3658 262894
rect -3574 262658 -3338 262894
rect -3894 262338 -3658 262574
rect -3574 262338 -3338 262574
rect -3894 226658 -3658 226894
rect -3574 226658 -3338 226894
rect -3894 226338 -3658 226574
rect -3574 226338 -3338 226574
rect -3894 190658 -3658 190894
rect -3574 190658 -3338 190894
rect -3894 190338 -3658 190574
rect -3574 190338 -3338 190574
rect -3894 154658 -3658 154894
rect -3574 154658 -3338 154894
rect -3894 154338 -3658 154574
rect -3574 154338 -3338 154574
rect -3894 118658 -3658 118894
rect -3574 118658 -3338 118894
rect -3894 118338 -3658 118574
rect -3574 118338 -3338 118574
rect -3894 82658 -3658 82894
rect -3574 82658 -3338 82894
rect -3894 82338 -3658 82574
rect -3574 82338 -3338 82574
rect -3894 46658 -3658 46894
rect -3574 46658 -3338 46894
rect -3894 46338 -3658 46574
rect -3574 46338 -3338 46574
rect -3894 10658 -3658 10894
rect -3574 10658 -3338 10894
rect -3894 10338 -3658 10574
rect -3574 10338 -3338 10574
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 690938 -2698 691174
rect -2614 690938 -2378 691174
rect -2934 690618 -2698 690854
rect -2614 690618 -2378 690854
rect -2934 654938 -2698 655174
rect -2614 654938 -2378 655174
rect -2934 654618 -2698 654854
rect -2614 654618 -2378 654854
rect -2934 618938 -2698 619174
rect -2614 618938 -2378 619174
rect -2934 618618 -2698 618854
rect -2614 618618 -2378 618854
rect -2934 582938 -2698 583174
rect -2614 582938 -2378 583174
rect -2934 582618 -2698 582854
rect -2614 582618 -2378 582854
rect -2934 546938 -2698 547174
rect -2614 546938 -2378 547174
rect -2934 546618 -2698 546854
rect -2614 546618 -2378 546854
rect -2934 510938 -2698 511174
rect -2614 510938 -2378 511174
rect -2934 510618 -2698 510854
rect -2614 510618 -2378 510854
rect -2934 474938 -2698 475174
rect -2614 474938 -2378 475174
rect -2934 474618 -2698 474854
rect -2614 474618 -2378 474854
rect -2934 438938 -2698 439174
rect -2614 438938 -2378 439174
rect -2934 438618 -2698 438854
rect -2614 438618 -2378 438854
rect -2934 402938 -2698 403174
rect -2614 402938 -2378 403174
rect -2934 402618 -2698 402854
rect -2614 402618 -2378 402854
rect -2934 366938 -2698 367174
rect -2614 366938 -2378 367174
rect -2934 366618 -2698 366854
rect -2614 366618 -2378 366854
rect -2934 330938 -2698 331174
rect -2614 330938 -2378 331174
rect -2934 330618 -2698 330854
rect -2614 330618 -2378 330854
rect -2934 294938 -2698 295174
rect -2614 294938 -2378 295174
rect -2934 294618 -2698 294854
rect -2614 294618 -2378 294854
rect -2934 258938 -2698 259174
rect -2614 258938 -2378 259174
rect -2934 258618 -2698 258854
rect -2614 258618 -2378 258854
rect -2934 222938 -2698 223174
rect -2614 222938 -2378 223174
rect -2934 222618 -2698 222854
rect -2614 222618 -2378 222854
rect -2934 186938 -2698 187174
rect -2614 186938 -2378 187174
rect -2934 186618 -2698 186854
rect -2614 186618 -2378 186854
rect -2934 150938 -2698 151174
rect -2614 150938 -2378 151174
rect -2934 150618 -2698 150854
rect -2614 150618 -2378 150854
rect -2934 114938 -2698 115174
rect -2614 114938 -2378 115174
rect -2934 114618 -2698 114854
rect -2614 114618 -2378 114854
rect -2934 78938 -2698 79174
rect -2614 78938 -2378 79174
rect -2934 78618 -2698 78854
rect -2614 78618 -2378 78854
rect -2934 42938 -2698 43174
rect -2614 42938 -2378 43174
rect -2934 42618 -2698 42854
rect -2614 42618 -2378 42854
rect -2934 6938 -2698 7174
rect -2614 6938 -2378 7174
rect -2934 6618 -2698 6854
rect -2614 6618 -2378 6854
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect -1974 687218 -1738 687454
rect -1654 687218 -1418 687454
rect -1974 686898 -1738 687134
rect -1654 686898 -1418 687134
rect -1974 651218 -1738 651454
rect -1654 651218 -1418 651454
rect -1974 650898 -1738 651134
rect -1654 650898 -1418 651134
rect -1974 615218 -1738 615454
rect -1654 615218 -1418 615454
rect -1974 614898 -1738 615134
rect -1654 614898 -1418 615134
rect -1974 579218 -1738 579454
rect -1654 579218 -1418 579454
rect -1974 578898 -1738 579134
rect -1654 578898 -1418 579134
rect -1974 543218 -1738 543454
rect -1654 543218 -1418 543454
rect -1974 542898 -1738 543134
rect -1654 542898 -1418 543134
rect -1974 507218 -1738 507454
rect -1654 507218 -1418 507454
rect -1974 506898 -1738 507134
rect -1654 506898 -1418 507134
rect -1974 471218 -1738 471454
rect -1654 471218 -1418 471454
rect -1974 470898 -1738 471134
rect -1654 470898 -1418 471134
rect -1974 435218 -1738 435454
rect -1654 435218 -1418 435454
rect -1974 434898 -1738 435134
rect -1654 434898 -1418 435134
rect -1974 399218 -1738 399454
rect -1654 399218 -1418 399454
rect -1974 398898 -1738 399134
rect -1654 398898 -1418 399134
rect -1974 363218 -1738 363454
rect -1654 363218 -1418 363454
rect -1974 362898 -1738 363134
rect -1654 362898 -1418 363134
rect -1974 327218 -1738 327454
rect -1654 327218 -1418 327454
rect -1974 326898 -1738 327134
rect -1654 326898 -1418 327134
rect -1974 291218 -1738 291454
rect -1654 291218 -1418 291454
rect -1974 290898 -1738 291134
rect -1654 290898 -1418 291134
rect -1974 255218 -1738 255454
rect -1654 255218 -1418 255454
rect -1974 254898 -1738 255134
rect -1654 254898 -1418 255134
rect -1974 219218 -1738 219454
rect -1654 219218 -1418 219454
rect -1974 218898 -1738 219134
rect -1654 218898 -1418 219134
rect -1974 183218 -1738 183454
rect -1654 183218 -1418 183454
rect -1974 182898 -1738 183134
rect -1654 182898 -1418 183134
rect -1974 147218 -1738 147454
rect -1654 147218 -1418 147454
rect -1974 146898 -1738 147134
rect -1654 146898 -1418 147134
rect -1974 111218 -1738 111454
rect -1654 111218 -1418 111454
rect -1974 110898 -1738 111134
rect -1654 110898 -1418 111134
rect -1974 75218 -1738 75454
rect -1654 75218 -1418 75454
rect -1974 74898 -1738 75134
rect -1654 74898 -1418 75134
rect -1974 39218 -1738 39454
rect -1654 39218 -1418 39454
rect -1974 38898 -1738 39134
rect -1654 38898 -1418 39134
rect -1974 3218 -1738 3454
rect -1654 3218 -1418 3454
rect -1974 2898 -1738 3134
rect -1654 2898 -1418 3134
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect 1826 704602 2062 704838
rect 2146 704602 2382 704838
rect 1826 704282 2062 704518
rect 2146 704282 2382 704518
rect 1826 687218 2062 687454
rect 2146 687218 2382 687454
rect 1826 686898 2062 687134
rect 2146 686898 2382 687134
rect 5546 705562 5782 705798
rect 5866 705562 6102 705798
rect 5546 705242 5782 705478
rect 5866 705242 6102 705478
rect 5546 690938 5782 691174
rect 5866 690938 6102 691174
rect 5546 690618 5782 690854
rect 5866 690618 6102 690854
rect 1826 651218 2062 651454
rect 2146 651218 2382 651454
rect 1826 650898 2062 651134
rect 2146 650898 2382 651134
rect 1826 615218 2062 615454
rect 2146 615218 2382 615454
rect 1826 614898 2062 615134
rect 2146 614898 2382 615134
rect 5546 654938 5782 655174
rect 5866 654938 6102 655174
rect 5546 654618 5782 654854
rect 5866 654618 6102 654854
rect 5546 618938 5782 619174
rect 5866 618938 6102 619174
rect 5546 618618 5782 618854
rect 5866 618618 6102 618854
rect 1826 579218 2062 579454
rect 2146 579218 2382 579454
rect 1826 578898 2062 579134
rect 2146 578898 2382 579134
rect 1826 543218 2062 543454
rect 2146 543218 2382 543454
rect 1826 542898 2062 543134
rect 2146 542898 2382 543134
rect 1826 507218 2062 507454
rect 2146 507218 2382 507454
rect 1826 506898 2062 507134
rect 2146 506898 2382 507134
rect 1826 471218 2062 471454
rect 2146 471218 2382 471454
rect 1826 470898 2062 471134
rect 2146 470898 2382 471134
rect 1826 435218 2062 435454
rect 2146 435218 2382 435454
rect 1826 434898 2062 435134
rect 2146 434898 2382 435134
rect 1826 399218 2062 399454
rect 2146 399218 2382 399454
rect 1826 398898 2062 399134
rect 2146 398898 2382 399134
rect 1826 363218 2062 363454
rect 2146 363218 2382 363454
rect 1826 362898 2062 363134
rect 2146 362898 2382 363134
rect 1826 327218 2062 327454
rect 2146 327218 2382 327454
rect 1826 326898 2062 327134
rect 2146 326898 2382 327134
rect 1826 291218 2062 291454
rect 2146 291218 2382 291454
rect 1826 290898 2062 291134
rect 2146 290898 2382 291134
rect 1826 255218 2062 255454
rect 2146 255218 2382 255454
rect 1826 254898 2062 255134
rect 2146 254898 2382 255134
rect 1826 219218 2062 219454
rect 2146 219218 2382 219454
rect 1826 218898 2062 219134
rect 2146 218898 2382 219134
rect 1826 183218 2062 183454
rect 2146 183218 2382 183454
rect 1826 182898 2062 183134
rect 2146 182898 2382 183134
rect 1826 147218 2062 147454
rect 2146 147218 2382 147454
rect 1826 146898 2062 147134
rect 2146 146898 2382 147134
rect 5546 582938 5782 583174
rect 5866 582938 6102 583174
rect 5546 582618 5782 582854
rect 5866 582618 6102 582854
rect 5546 546938 5782 547174
rect 5866 546938 6102 547174
rect 5546 546618 5782 546854
rect 5866 546618 6102 546854
rect 5546 510938 5782 511174
rect 5866 510938 6102 511174
rect 5546 510618 5782 510854
rect 5866 510618 6102 510854
rect 5546 474938 5782 475174
rect 5866 474938 6102 475174
rect 5546 474618 5782 474854
rect 5866 474618 6102 474854
rect 5546 438938 5782 439174
rect 5866 438938 6102 439174
rect 5546 438618 5782 438854
rect 5866 438618 6102 438854
rect 5546 402938 5782 403174
rect 5866 402938 6102 403174
rect 5546 402618 5782 402854
rect 5866 402618 6102 402854
rect 5546 366938 5782 367174
rect 5866 366938 6102 367174
rect 5546 366618 5782 366854
rect 5866 366618 6102 366854
rect 5546 330938 5782 331174
rect 5866 330938 6102 331174
rect 5546 330618 5782 330854
rect 5866 330618 6102 330854
rect 5546 294938 5782 295174
rect 5866 294938 6102 295174
rect 5546 294618 5782 294854
rect 5866 294618 6102 294854
rect 5546 258938 5782 259174
rect 5866 258938 6102 259174
rect 5546 258618 5782 258854
rect 5866 258618 6102 258854
rect 5546 222938 5782 223174
rect 5866 222938 6102 223174
rect 5546 222618 5782 222854
rect 5866 222618 6102 222854
rect 5546 186938 5782 187174
rect 5866 186938 6102 187174
rect 5546 186618 5782 186854
rect 5866 186618 6102 186854
rect 5546 150938 5782 151174
rect 5866 150938 6102 151174
rect 5546 150618 5782 150854
rect 5866 150618 6102 150854
rect 1826 111218 2062 111454
rect 2146 111218 2382 111454
rect 1826 110898 2062 111134
rect 2146 110898 2382 111134
rect 5546 114938 5782 115174
rect 5866 114938 6102 115174
rect 5546 114618 5782 114854
rect 5866 114618 6102 114854
rect 1826 75218 2062 75454
rect 2146 75218 2382 75454
rect 1826 74898 2062 75134
rect 2146 74898 2382 75134
rect 5546 78938 5782 79174
rect 5866 78938 6102 79174
rect 5546 78618 5782 78854
rect 5866 78618 6102 78854
rect 1826 39218 2062 39454
rect 2146 39218 2382 39454
rect 1826 38898 2062 39134
rect 2146 38898 2382 39134
rect 1826 3218 2062 3454
rect 2146 3218 2382 3454
rect 1826 2898 2062 3134
rect 2146 2898 2382 3134
rect 1826 -582 2062 -346
rect 2146 -582 2382 -346
rect 1826 -902 2062 -666
rect 2146 -902 2382 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 5546 42938 5782 43174
rect 5866 42938 6102 43174
rect 5546 42618 5782 42854
rect 5866 42618 6102 42854
rect 5546 6938 5782 7174
rect 5866 6938 6102 7174
rect 5546 6618 5782 6854
rect 5866 6618 6102 6854
rect 5546 -1542 5782 -1306
rect 5866 -1542 6102 -1306
rect 5546 -1862 5782 -1626
rect 5866 -1862 6102 -1626
rect 9266 706522 9502 706758
rect 9586 706522 9822 706758
rect 9266 706202 9502 706438
rect 9586 706202 9822 706438
rect 9266 694658 9502 694894
rect 9586 694658 9822 694894
rect 9266 694338 9502 694574
rect 9586 694338 9822 694574
rect 9266 658658 9502 658894
rect 9586 658658 9822 658894
rect 9266 658338 9502 658574
rect 9586 658338 9822 658574
rect 9266 622658 9502 622894
rect 9586 622658 9822 622894
rect 9266 622338 9502 622574
rect 9586 622338 9822 622574
rect 9266 586658 9502 586894
rect 9586 586658 9822 586894
rect 9266 586338 9502 586574
rect 9586 586338 9822 586574
rect 9266 550658 9502 550894
rect 9586 550658 9822 550894
rect 9266 550338 9502 550574
rect 9586 550338 9822 550574
rect 9266 514658 9502 514894
rect 9586 514658 9822 514894
rect 9266 514338 9502 514574
rect 9586 514338 9822 514574
rect 9266 478658 9502 478894
rect 9586 478658 9822 478894
rect 9266 478338 9502 478574
rect 9586 478338 9822 478574
rect 9266 442658 9502 442894
rect 9586 442658 9822 442894
rect 9266 442338 9502 442574
rect 9586 442338 9822 442574
rect 9266 406658 9502 406894
rect 9586 406658 9822 406894
rect 9266 406338 9502 406574
rect 9586 406338 9822 406574
rect 9266 370658 9502 370894
rect 9586 370658 9822 370894
rect 9266 370338 9502 370574
rect 9586 370338 9822 370574
rect 9266 334658 9502 334894
rect 9586 334658 9822 334894
rect 9266 334338 9502 334574
rect 9586 334338 9822 334574
rect 9266 298658 9502 298894
rect 9586 298658 9822 298894
rect 9266 298338 9502 298574
rect 9586 298338 9822 298574
rect 9266 262658 9502 262894
rect 9586 262658 9822 262894
rect 9266 262338 9502 262574
rect 9586 262338 9822 262574
rect 9266 226658 9502 226894
rect 9586 226658 9822 226894
rect 9266 226338 9502 226574
rect 9586 226338 9822 226574
rect 9266 190658 9502 190894
rect 9586 190658 9822 190894
rect 9266 190338 9502 190574
rect 9586 190338 9822 190574
rect 9266 154658 9502 154894
rect 9586 154658 9822 154894
rect 9266 154338 9502 154574
rect 9586 154338 9822 154574
rect 9266 118658 9502 118894
rect 9586 118658 9822 118894
rect 9266 118338 9502 118574
rect 9586 118338 9822 118574
rect 9266 82658 9502 82894
rect 9586 82658 9822 82894
rect 9266 82338 9502 82574
rect 9586 82338 9822 82574
rect 9266 46658 9502 46894
rect 9586 46658 9822 46894
rect 9266 46338 9502 46574
rect 9586 46338 9822 46574
rect 9266 10658 9502 10894
rect 9586 10658 9822 10894
rect 9266 10338 9502 10574
rect 9586 10338 9822 10574
rect 9266 -2502 9502 -2266
rect 9586 -2502 9822 -2266
rect 9266 -2822 9502 -2586
rect 9586 -2822 9822 -2586
rect 12986 707482 13222 707718
rect 13306 707482 13542 707718
rect 12986 707162 13222 707398
rect 13306 707162 13542 707398
rect 12986 698378 13222 698614
rect 13306 698378 13542 698614
rect 12986 698058 13222 698294
rect 13306 698058 13542 698294
rect 12986 662378 13222 662614
rect 13306 662378 13542 662614
rect 12986 662058 13222 662294
rect 13306 662058 13542 662294
rect 12986 626378 13222 626614
rect 13306 626378 13542 626614
rect 12986 626058 13222 626294
rect 13306 626058 13542 626294
rect 12986 590378 13222 590614
rect 13306 590378 13542 590614
rect 12986 590058 13222 590294
rect 13306 590058 13542 590294
rect 12986 554378 13222 554614
rect 13306 554378 13542 554614
rect 12986 554058 13222 554294
rect 13306 554058 13542 554294
rect 12986 518378 13222 518614
rect 13306 518378 13542 518614
rect 12986 518058 13222 518294
rect 13306 518058 13542 518294
rect 12986 482378 13222 482614
rect 13306 482378 13542 482614
rect 12986 482058 13222 482294
rect 13306 482058 13542 482294
rect 12986 446378 13222 446614
rect 13306 446378 13542 446614
rect 12986 446058 13222 446294
rect 13306 446058 13542 446294
rect 12986 410378 13222 410614
rect 13306 410378 13542 410614
rect 12986 410058 13222 410294
rect 13306 410058 13542 410294
rect 12986 374378 13222 374614
rect 13306 374378 13542 374614
rect 12986 374058 13222 374294
rect 13306 374058 13542 374294
rect 12986 338378 13222 338614
rect 13306 338378 13542 338614
rect 12986 338058 13222 338294
rect 13306 338058 13542 338294
rect 12986 302378 13222 302614
rect 13306 302378 13542 302614
rect 12986 302058 13222 302294
rect 13306 302058 13542 302294
rect 12986 266378 13222 266614
rect 13306 266378 13542 266614
rect 12986 266058 13222 266294
rect 13306 266058 13542 266294
rect 12986 230378 13222 230614
rect 13306 230378 13542 230614
rect 12986 230058 13222 230294
rect 13306 230058 13542 230294
rect 12986 194378 13222 194614
rect 13306 194378 13542 194614
rect 12986 194058 13222 194294
rect 13306 194058 13542 194294
rect 12986 158378 13222 158614
rect 13306 158378 13542 158614
rect 12986 158058 13222 158294
rect 13306 158058 13542 158294
rect 12986 122378 13222 122614
rect 13306 122378 13542 122614
rect 12986 122058 13222 122294
rect 13306 122058 13542 122294
rect 12986 86378 13222 86614
rect 13306 86378 13542 86614
rect 12986 86058 13222 86294
rect 13306 86058 13542 86294
rect 12986 50378 13222 50614
rect 13306 50378 13542 50614
rect 12986 50058 13222 50294
rect 13306 50058 13542 50294
rect 12986 14378 13222 14614
rect 13306 14378 13542 14614
rect 12986 14058 13222 14294
rect 13306 14058 13542 14294
rect 12986 -3462 13222 -3226
rect 13306 -3462 13542 -3226
rect 12986 -3782 13222 -3546
rect 13306 -3782 13542 -3546
rect 16706 708442 16942 708678
rect 17026 708442 17262 708678
rect 16706 708122 16942 708358
rect 17026 708122 17262 708358
rect 16706 666098 16942 666334
rect 17026 666098 17262 666334
rect 16706 665778 16942 666014
rect 17026 665778 17262 666014
rect 16706 630098 16942 630334
rect 17026 630098 17262 630334
rect 16706 629778 16942 630014
rect 17026 629778 17262 630014
rect 16706 594098 16942 594334
rect 17026 594098 17262 594334
rect 16706 593778 16942 594014
rect 17026 593778 17262 594014
rect 16706 558098 16942 558334
rect 17026 558098 17262 558334
rect 16706 557778 16942 558014
rect 17026 557778 17262 558014
rect 16706 522098 16942 522334
rect 17026 522098 17262 522334
rect 16706 521778 16942 522014
rect 17026 521778 17262 522014
rect 16706 486098 16942 486334
rect 17026 486098 17262 486334
rect 16706 485778 16942 486014
rect 17026 485778 17262 486014
rect 16706 450098 16942 450334
rect 17026 450098 17262 450334
rect 16706 449778 16942 450014
rect 17026 449778 17262 450014
rect 16706 414098 16942 414334
rect 17026 414098 17262 414334
rect 16706 413778 16942 414014
rect 17026 413778 17262 414014
rect 16706 378098 16942 378334
rect 17026 378098 17262 378334
rect 16706 377778 16942 378014
rect 17026 377778 17262 378014
rect 16706 342098 16942 342334
rect 17026 342098 17262 342334
rect 16706 341778 16942 342014
rect 17026 341778 17262 342014
rect 16706 306098 16942 306334
rect 17026 306098 17262 306334
rect 16706 305778 16942 306014
rect 17026 305778 17262 306014
rect 16706 270098 16942 270334
rect 17026 270098 17262 270334
rect 16706 269778 16942 270014
rect 17026 269778 17262 270014
rect 16706 234098 16942 234334
rect 17026 234098 17262 234334
rect 16706 233778 16942 234014
rect 17026 233778 17262 234014
rect 16706 198098 16942 198334
rect 17026 198098 17262 198334
rect 16706 197778 16942 198014
rect 17026 197778 17262 198014
rect 16706 162098 16942 162334
rect 17026 162098 17262 162334
rect 16706 161778 16942 162014
rect 17026 161778 17262 162014
rect 16706 126098 16942 126334
rect 17026 126098 17262 126334
rect 16706 125778 16942 126014
rect 17026 125778 17262 126014
rect 16706 90098 16942 90334
rect 17026 90098 17262 90334
rect 16706 89778 16942 90014
rect 17026 89778 17262 90014
rect 16706 54098 16942 54334
rect 17026 54098 17262 54334
rect 16706 53778 16942 54014
rect 17026 53778 17262 54014
rect 16706 18098 16942 18334
rect 17026 18098 17262 18334
rect 16706 17778 16942 18014
rect 17026 17778 17262 18014
rect 16706 -4422 16942 -4186
rect 17026 -4422 17262 -4186
rect 16706 -4742 16942 -4506
rect 17026 -4742 17262 -4506
rect 20426 709402 20662 709638
rect 20746 709402 20982 709638
rect 20426 709082 20662 709318
rect 20746 709082 20982 709318
rect 20426 669818 20662 670054
rect 20746 669818 20982 670054
rect 20426 669498 20662 669734
rect 20746 669498 20982 669734
rect 27866 711322 28102 711558
rect 28186 711322 28422 711558
rect 27866 711002 28102 711238
rect 28186 711002 28422 711238
rect 27866 677258 28102 677494
rect 28186 677258 28422 677494
rect 27866 676938 28102 677174
rect 28186 676938 28422 677174
rect 24250 651218 24486 651454
rect 24250 650898 24486 651134
rect 20426 633818 20662 634054
rect 20746 633818 20982 634054
rect 20426 633498 20662 633734
rect 20746 633498 20982 633734
rect 37826 704602 38062 704838
rect 38146 704602 38382 704838
rect 37826 704282 38062 704518
rect 38146 704282 38382 704518
rect 37826 687218 38062 687454
rect 38146 687218 38382 687454
rect 37826 686898 38062 687134
rect 38146 686898 38382 687134
rect 41546 705562 41782 705798
rect 41866 705562 42102 705798
rect 41546 705242 41782 705478
rect 41866 705242 42102 705478
rect 41546 690938 41782 691174
rect 41866 690938 42102 691174
rect 41546 690618 41782 690854
rect 41866 690618 42102 690854
rect 45266 706522 45502 706758
rect 45586 706522 45822 706758
rect 45266 706202 45502 706438
rect 45586 706202 45822 706438
rect 45266 694658 45502 694894
rect 45586 694658 45822 694894
rect 45266 694338 45502 694574
rect 45586 694338 45822 694574
rect 48986 707482 49222 707718
rect 49306 707482 49542 707718
rect 48986 707162 49222 707398
rect 49306 707162 49542 707398
rect 48986 698378 49222 698614
rect 49306 698378 49542 698614
rect 48986 698058 49222 698294
rect 49306 698058 49542 698294
rect 63866 711322 64102 711558
rect 64186 711322 64422 711558
rect 63866 711002 64102 711238
rect 64186 711002 64422 711238
rect 63866 677258 64102 677494
rect 64186 677258 64422 677494
rect 63866 676938 64102 677174
rect 64186 676938 64422 677174
rect 73826 704602 74062 704838
rect 74146 704602 74382 704838
rect 73826 704282 74062 704518
rect 74146 704282 74382 704518
rect 73826 687218 74062 687454
rect 74146 687218 74382 687454
rect 73826 686898 74062 687134
rect 74146 686898 74382 687134
rect 77546 705562 77782 705798
rect 77866 705562 78102 705798
rect 77546 705242 77782 705478
rect 77866 705242 78102 705478
rect 77546 690938 77782 691174
rect 77866 690938 78102 691174
rect 77546 690618 77782 690854
rect 77866 690618 78102 690854
rect 81266 706522 81502 706758
rect 81586 706522 81822 706758
rect 81266 706202 81502 706438
rect 81586 706202 81822 706438
rect 81266 694658 81502 694894
rect 81586 694658 81822 694894
rect 81266 694338 81502 694574
rect 81586 694338 81822 694574
rect 84986 707482 85222 707718
rect 85306 707482 85542 707718
rect 84986 707162 85222 707398
rect 85306 707162 85542 707398
rect 84986 698378 85222 698614
rect 85306 698378 85542 698614
rect 84986 698058 85222 698294
rect 85306 698058 85542 698294
rect 99866 711322 100102 711558
rect 100186 711322 100422 711558
rect 99866 711002 100102 711238
rect 100186 711002 100422 711238
rect 99866 677258 100102 677494
rect 100186 677258 100422 677494
rect 99866 676938 100102 677174
rect 100186 676938 100422 677174
rect 109826 704602 110062 704838
rect 110146 704602 110382 704838
rect 109826 704282 110062 704518
rect 110146 704282 110382 704518
rect 109826 687218 110062 687454
rect 110146 687218 110382 687454
rect 109826 686898 110062 687134
rect 110146 686898 110382 687134
rect 113546 705562 113782 705798
rect 113866 705562 114102 705798
rect 113546 705242 113782 705478
rect 113866 705242 114102 705478
rect 113546 690938 113782 691174
rect 113866 690938 114102 691174
rect 113546 690618 113782 690854
rect 113866 690618 114102 690854
rect 117266 706522 117502 706758
rect 117586 706522 117822 706758
rect 117266 706202 117502 706438
rect 117586 706202 117822 706438
rect 117266 694658 117502 694894
rect 117586 694658 117822 694894
rect 117266 694338 117502 694574
rect 117586 694338 117822 694574
rect 120986 707482 121222 707718
rect 121306 707482 121542 707718
rect 120986 707162 121222 707398
rect 121306 707162 121542 707398
rect 120986 698378 121222 698614
rect 121306 698378 121542 698614
rect 120986 698058 121222 698294
rect 121306 698058 121542 698294
rect 135866 711322 136102 711558
rect 136186 711322 136422 711558
rect 135866 711002 136102 711238
rect 136186 711002 136422 711238
rect 135866 677258 136102 677494
rect 136186 677258 136422 677494
rect 135866 676938 136102 677174
rect 136186 676938 136422 677174
rect 145826 704602 146062 704838
rect 146146 704602 146382 704838
rect 145826 704282 146062 704518
rect 146146 704282 146382 704518
rect 145826 687218 146062 687454
rect 146146 687218 146382 687454
rect 145826 686898 146062 687134
rect 146146 686898 146382 687134
rect 149546 705562 149782 705798
rect 149866 705562 150102 705798
rect 149546 705242 149782 705478
rect 149866 705242 150102 705478
rect 149546 690938 149782 691174
rect 149866 690938 150102 691174
rect 149546 690618 149782 690854
rect 149866 690618 150102 690854
rect 153266 706522 153502 706758
rect 153586 706522 153822 706758
rect 153266 706202 153502 706438
rect 153586 706202 153822 706438
rect 153266 694658 153502 694894
rect 153586 694658 153822 694894
rect 153266 694338 153502 694574
rect 153586 694338 153822 694574
rect 156986 707482 157222 707718
rect 157306 707482 157542 707718
rect 156986 707162 157222 707398
rect 157306 707162 157542 707398
rect 156986 698378 157222 698614
rect 157306 698378 157542 698614
rect 156986 698058 157222 698294
rect 157306 698058 157542 698294
rect 171866 711322 172102 711558
rect 172186 711322 172422 711558
rect 171866 711002 172102 711238
rect 172186 711002 172422 711238
rect 171866 677258 172102 677494
rect 172186 677258 172422 677494
rect 171866 676938 172102 677174
rect 172186 676938 172422 677174
rect 181826 704602 182062 704838
rect 182146 704602 182382 704838
rect 181826 704282 182062 704518
rect 182146 704282 182382 704518
rect 181826 687218 182062 687454
rect 182146 687218 182382 687454
rect 181826 686898 182062 687134
rect 182146 686898 182382 687134
rect 185546 705562 185782 705798
rect 185866 705562 186102 705798
rect 185546 705242 185782 705478
rect 185866 705242 186102 705478
rect 185546 690938 185782 691174
rect 185866 690938 186102 691174
rect 185546 690618 185782 690854
rect 185866 690618 186102 690854
rect 189266 706522 189502 706758
rect 189586 706522 189822 706758
rect 189266 706202 189502 706438
rect 189586 706202 189822 706438
rect 189266 694658 189502 694894
rect 189586 694658 189822 694894
rect 189266 694338 189502 694574
rect 189586 694338 189822 694574
rect 192986 707482 193222 707718
rect 193306 707482 193542 707718
rect 192986 707162 193222 707398
rect 193306 707162 193542 707398
rect 192986 698378 193222 698614
rect 193306 698378 193542 698614
rect 192986 698058 193222 698294
rect 193306 698058 193542 698294
rect 207866 711322 208102 711558
rect 208186 711322 208422 711558
rect 207866 711002 208102 711238
rect 208186 711002 208422 711238
rect 207866 677258 208102 677494
rect 208186 677258 208422 677494
rect 207866 676938 208102 677174
rect 208186 676938 208422 677174
rect 217826 704602 218062 704838
rect 218146 704602 218382 704838
rect 217826 704282 218062 704518
rect 218146 704282 218382 704518
rect 217826 687218 218062 687454
rect 218146 687218 218382 687454
rect 217826 686898 218062 687134
rect 218146 686898 218382 687134
rect 221546 705562 221782 705798
rect 221866 705562 222102 705798
rect 221546 705242 221782 705478
rect 221866 705242 222102 705478
rect 221546 690938 221782 691174
rect 221866 690938 222102 691174
rect 221546 690618 221782 690854
rect 221866 690618 222102 690854
rect 225266 706522 225502 706758
rect 225586 706522 225822 706758
rect 225266 706202 225502 706438
rect 225586 706202 225822 706438
rect 225266 694658 225502 694894
rect 225586 694658 225822 694894
rect 225266 694338 225502 694574
rect 225586 694338 225822 694574
rect 228986 707482 229222 707718
rect 229306 707482 229542 707718
rect 228986 707162 229222 707398
rect 229306 707162 229542 707398
rect 228986 698378 229222 698614
rect 229306 698378 229542 698614
rect 228986 698058 229222 698294
rect 229306 698058 229542 698294
rect 243866 711322 244102 711558
rect 244186 711322 244422 711558
rect 243866 711002 244102 711238
rect 244186 711002 244422 711238
rect 243866 677258 244102 677494
rect 244186 677258 244422 677494
rect 243866 676938 244102 677174
rect 244186 676938 244422 677174
rect 253826 704602 254062 704838
rect 254146 704602 254382 704838
rect 253826 704282 254062 704518
rect 254146 704282 254382 704518
rect 253826 687218 254062 687454
rect 254146 687218 254382 687454
rect 253826 686898 254062 687134
rect 254146 686898 254382 687134
rect 257546 705562 257782 705798
rect 257866 705562 258102 705798
rect 257546 705242 257782 705478
rect 257866 705242 258102 705478
rect 257546 690938 257782 691174
rect 257866 690938 258102 691174
rect 257546 690618 257782 690854
rect 257866 690618 258102 690854
rect 261266 706522 261502 706758
rect 261586 706522 261822 706758
rect 261266 706202 261502 706438
rect 261586 706202 261822 706438
rect 261266 694658 261502 694894
rect 261586 694658 261822 694894
rect 261266 694338 261502 694574
rect 261586 694338 261822 694574
rect 264986 707482 265222 707718
rect 265306 707482 265542 707718
rect 264986 707162 265222 707398
rect 265306 707162 265542 707398
rect 264986 698378 265222 698614
rect 265306 698378 265542 698614
rect 264986 698058 265222 698294
rect 265306 698058 265542 698294
rect 279866 711322 280102 711558
rect 280186 711322 280422 711558
rect 279866 711002 280102 711238
rect 280186 711002 280422 711238
rect 279866 677258 280102 677494
rect 280186 677258 280422 677494
rect 279866 676938 280102 677174
rect 280186 676938 280422 677174
rect 289826 704602 290062 704838
rect 290146 704602 290382 704838
rect 289826 704282 290062 704518
rect 290146 704282 290382 704518
rect 289826 687218 290062 687454
rect 290146 687218 290382 687454
rect 289826 686898 290062 687134
rect 290146 686898 290382 687134
rect 293546 705562 293782 705798
rect 293866 705562 294102 705798
rect 293546 705242 293782 705478
rect 293866 705242 294102 705478
rect 293546 690938 293782 691174
rect 293866 690938 294102 691174
rect 293546 690618 293782 690854
rect 293866 690618 294102 690854
rect 297266 706522 297502 706758
rect 297586 706522 297822 706758
rect 297266 706202 297502 706438
rect 297586 706202 297822 706438
rect 297266 694658 297502 694894
rect 297586 694658 297822 694894
rect 297266 694338 297502 694574
rect 297586 694338 297822 694574
rect 300986 707482 301222 707718
rect 301306 707482 301542 707718
rect 300986 707162 301222 707398
rect 301306 707162 301542 707398
rect 300986 698378 301222 698614
rect 301306 698378 301542 698614
rect 300986 698058 301222 698294
rect 301306 698058 301542 698294
rect 325826 704602 326062 704838
rect 326146 704602 326382 704838
rect 325826 704282 326062 704518
rect 326146 704282 326382 704518
rect 325826 687218 326062 687454
rect 326146 687218 326382 687454
rect 325826 686898 326062 687134
rect 326146 686898 326382 687134
rect 329546 705562 329782 705798
rect 329866 705562 330102 705798
rect 329546 705242 329782 705478
rect 329866 705242 330102 705478
rect 329546 690938 329782 691174
rect 329866 690938 330102 691174
rect 329546 690618 329782 690854
rect 329866 690618 330102 690854
rect 333266 706522 333502 706758
rect 333586 706522 333822 706758
rect 333266 706202 333502 706438
rect 333586 706202 333822 706438
rect 333266 694658 333502 694894
rect 333586 694658 333822 694894
rect 333266 694338 333502 694574
rect 333586 694338 333822 694574
rect 336986 707482 337222 707718
rect 337306 707482 337542 707718
rect 336986 707162 337222 707398
rect 337306 707162 337542 707398
rect 336986 698378 337222 698614
rect 337306 698378 337542 698614
rect 336986 698058 337222 698294
rect 337306 698058 337542 698294
rect 351866 711322 352102 711558
rect 352186 711322 352422 711558
rect 351866 711002 352102 711238
rect 352186 711002 352422 711238
rect 351866 677258 352102 677494
rect 352186 677258 352422 677494
rect 351866 676938 352102 677174
rect 352186 676938 352422 677174
rect 361826 704602 362062 704838
rect 362146 704602 362382 704838
rect 361826 704282 362062 704518
rect 362146 704282 362382 704518
rect 361826 687218 362062 687454
rect 362146 687218 362382 687454
rect 361826 686898 362062 687134
rect 362146 686898 362382 687134
rect 39610 654938 39846 655174
rect 39610 654618 39846 654854
rect 70330 654938 70566 655174
rect 70330 654618 70566 654854
rect 101050 654938 101286 655174
rect 101050 654618 101286 654854
rect 131770 654938 132006 655174
rect 131770 654618 132006 654854
rect 162490 654938 162726 655174
rect 162490 654618 162726 654854
rect 193210 654938 193446 655174
rect 193210 654618 193446 654854
rect 223930 654938 224166 655174
rect 223930 654618 224166 654854
rect 254650 654938 254886 655174
rect 254650 654618 254886 654854
rect 285370 654938 285606 655174
rect 285370 654618 285606 654854
rect 316090 654938 316326 655174
rect 316090 654618 316326 654854
rect 346810 654938 347046 655174
rect 346810 654618 347046 654854
rect 54970 651218 55206 651454
rect 54970 650898 55206 651134
rect 85690 651218 85926 651454
rect 85690 650898 85926 651134
rect 116410 651218 116646 651454
rect 116410 650898 116646 651134
rect 147130 651218 147366 651454
rect 147130 650898 147366 651134
rect 177850 651218 178086 651454
rect 177850 650898 178086 651134
rect 208570 651218 208806 651454
rect 208570 650898 208806 651134
rect 239290 651218 239526 651454
rect 239290 650898 239526 651134
rect 270010 651218 270246 651454
rect 270010 650898 270246 651134
rect 300730 651218 300966 651454
rect 300730 650898 300966 651134
rect 331450 651218 331686 651454
rect 331450 650898 331686 651134
rect 361826 651218 362062 651454
rect 362146 651218 362382 651454
rect 361826 650898 362062 651134
rect 362146 650898 362382 651134
rect 27866 641258 28102 641494
rect 28186 641258 28422 641494
rect 27866 640938 28102 641174
rect 28186 640938 28422 641174
rect 24250 615218 24486 615454
rect 24250 614898 24486 615134
rect 20426 597818 20662 598054
rect 20746 597818 20982 598054
rect 20426 597498 20662 597734
rect 20746 597498 20982 597734
rect 39610 618938 39846 619174
rect 39610 618618 39846 618854
rect 70330 618938 70566 619174
rect 70330 618618 70566 618854
rect 101050 618938 101286 619174
rect 101050 618618 101286 618854
rect 131770 618938 132006 619174
rect 131770 618618 132006 618854
rect 162490 618938 162726 619174
rect 162490 618618 162726 618854
rect 193210 618938 193446 619174
rect 193210 618618 193446 618854
rect 223930 618938 224166 619174
rect 223930 618618 224166 618854
rect 254650 618938 254886 619174
rect 254650 618618 254886 618854
rect 285370 618938 285606 619174
rect 285370 618618 285606 618854
rect 316090 618938 316326 619174
rect 316090 618618 316326 618854
rect 346810 618938 347046 619174
rect 346810 618618 347046 618854
rect 54970 615218 55206 615454
rect 54970 614898 55206 615134
rect 85690 615218 85926 615454
rect 85690 614898 85926 615134
rect 116410 615218 116646 615454
rect 116410 614898 116646 615134
rect 147130 615218 147366 615454
rect 147130 614898 147366 615134
rect 177850 615218 178086 615454
rect 177850 614898 178086 615134
rect 208570 615218 208806 615454
rect 208570 614898 208806 615134
rect 239290 615218 239526 615454
rect 239290 614898 239526 615134
rect 270010 615218 270246 615454
rect 270010 614898 270246 615134
rect 300730 615218 300966 615454
rect 300730 614898 300966 615134
rect 331450 615218 331686 615454
rect 331450 614898 331686 615134
rect 361826 615218 362062 615454
rect 362146 615218 362382 615454
rect 361826 614898 362062 615134
rect 362146 614898 362382 615134
rect 27866 605258 28102 605494
rect 28186 605258 28422 605494
rect 27866 604938 28102 605174
rect 28186 604938 28422 605174
rect 24250 579218 24486 579454
rect 24250 578898 24486 579134
rect 20426 561818 20662 562054
rect 20746 561818 20982 562054
rect 20426 561498 20662 561734
rect 20746 561498 20982 561734
rect 39610 582938 39846 583174
rect 39610 582618 39846 582854
rect 70330 582938 70566 583174
rect 70330 582618 70566 582854
rect 101050 582938 101286 583174
rect 101050 582618 101286 582854
rect 131770 582938 132006 583174
rect 131770 582618 132006 582854
rect 162490 582938 162726 583174
rect 162490 582618 162726 582854
rect 193210 582938 193446 583174
rect 193210 582618 193446 582854
rect 223930 582938 224166 583174
rect 223930 582618 224166 582854
rect 254650 582938 254886 583174
rect 254650 582618 254886 582854
rect 285370 582938 285606 583174
rect 285370 582618 285606 582854
rect 316090 582938 316326 583174
rect 316090 582618 316326 582854
rect 346810 582938 347046 583174
rect 346810 582618 347046 582854
rect 54970 579218 55206 579454
rect 54970 578898 55206 579134
rect 85690 579218 85926 579454
rect 85690 578898 85926 579134
rect 116410 579218 116646 579454
rect 116410 578898 116646 579134
rect 147130 579218 147366 579454
rect 147130 578898 147366 579134
rect 177850 579218 178086 579454
rect 177850 578898 178086 579134
rect 208570 579218 208806 579454
rect 208570 578898 208806 579134
rect 239290 579218 239526 579454
rect 239290 578898 239526 579134
rect 270010 579218 270246 579454
rect 270010 578898 270246 579134
rect 300730 579218 300966 579454
rect 300730 578898 300966 579134
rect 331450 579218 331686 579454
rect 331450 578898 331686 579134
rect 361826 579218 362062 579454
rect 362146 579218 362382 579454
rect 361826 578898 362062 579134
rect 362146 578898 362382 579134
rect 27866 569258 28102 569494
rect 28186 569258 28422 569494
rect 27866 568938 28102 569174
rect 28186 568938 28422 569174
rect 24250 543218 24486 543454
rect 24250 542898 24486 543134
rect 20426 525818 20662 526054
rect 20746 525818 20982 526054
rect 20426 525498 20662 525734
rect 20746 525498 20982 525734
rect 39610 546938 39846 547174
rect 39610 546618 39846 546854
rect 70330 546938 70566 547174
rect 70330 546618 70566 546854
rect 101050 546938 101286 547174
rect 101050 546618 101286 546854
rect 131770 546938 132006 547174
rect 131770 546618 132006 546854
rect 162490 546938 162726 547174
rect 162490 546618 162726 546854
rect 193210 546938 193446 547174
rect 193210 546618 193446 546854
rect 223930 546938 224166 547174
rect 223930 546618 224166 546854
rect 254650 546938 254886 547174
rect 254650 546618 254886 546854
rect 285370 546938 285606 547174
rect 285370 546618 285606 546854
rect 316090 546938 316326 547174
rect 316090 546618 316326 546854
rect 346810 546938 347046 547174
rect 346810 546618 347046 546854
rect 54970 543218 55206 543454
rect 54970 542898 55206 543134
rect 85690 543218 85926 543454
rect 85690 542898 85926 543134
rect 116410 543218 116646 543454
rect 116410 542898 116646 543134
rect 147130 543218 147366 543454
rect 147130 542898 147366 543134
rect 177850 543218 178086 543454
rect 177850 542898 178086 543134
rect 208570 543218 208806 543454
rect 208570 542898 208806 543134
rect 239290 543218 239526 543454
rect 239290 542898 239526 543134
rect 270010 543218 270246 543454
rect 270010 542898 270246 543134
rect 300730 543218 300966 543454
rect 300730 542898 300966 543134
rect 331450 543218 331686 543454
rect 331450 542898 331686 543134
rect 361826 543218 362062 543454
rect 362146 543218 362382 543454
rect 361826 542898 362062 543134
rect 362146 542898 362382 543134
rect 27866 533258 28102 533494
rect 28186 533258 28422 533494
rect 27866 532938 28102 533174
rect 28186 532938 28422 533174
rect 24250 507218 24486 507454
rect 24250 506898 24486 507134
rect 20426 489818 20662 490054
rect 20746 489818 20982 490054
rect 20426 489498 20662 489734
rect 20746 489498 20982 489734
rect 39610 510938 39846 511174
rect 39610 510618 39846 510854
rect 70330 510938 70566 511174
rect 70330 510618 70566 510854
rect 101050 510938 101286 511174
rect 101050 510618 101286 510854
rect 131770 510938 132006 511174
rect 131770 510618 132006 510854
rect 162490 510938 162726 511174
rect 162490 510618 162726 510854
rect 193210 510938 193446 511174
rect 193210 510618 193446 510854
rect 223930 510938 224166 511174
rect 223930 510618 224166 510854
rect 254650 510938 254886 511174
rect 254650 510618 254886 510854
rect 285370 510938 285606 511174
rect 285370 510618 285606 510854
rect 316090 510938 316326 511174
rect 316090 510618 316326 510854
rect 346810 510938 347046 511174
rect 346810 510618 347046 510854
rect 54970 507218 55206 507454
rect 54970 506898 55206 507134
rect 85690 507218 85926 507454
rect 85690 506898 85926 507134
rect 116410 507218 116646 507454
rect 116410 506898 116646 507134
rect 147130 507218 147366 507454
rect 147130 506898 147366 507134
rect 177850 507218 178086 507454
rect 177850 506898 178086 507134
rect 208570 507218 208806 507454
rect 208570 506898 208806 507134
rect 239290 507218 239526 507454
rect 239290 506898 239526 507134
rect 270010 507218 270246 507454
rect 270010 506898 270246 507134
rect 300730 507218 300966 507454
rect 300730 506898 300966 507134
rect 331450 507218 331686 507454
rect 331450 506898 331686 507134
rect 361826 507218 362062 507454
rect 362146 507218 362382 507454
rect 361826 506898 362062 507134
rect 362146 506898 362382 507134
rect 27866 497258 28102 497494
rect 28186 497258 28422 497494
rect 27866 496938 28102 497174
rect 28186 496938 28422 497174
rect 24250 471218 24486 471454
rect 24250 470898 24486 471134
rect 20426 453818 20662 454054
rect 20746 453818 20982 454054
rect 20426 453498 20662 453734
rect 20746 453498 20982 453734
rect 39610 474938 39846 475174
rect 39610 474618 39846 474854
rect 70330 474938 70566 475174
rect 70330 474618 70566 474854
rect 101050 474938 101286 475174
rect 101050 474618 101286 474854
rect 131770 474938 132006 475174
rect 131770 474618 132006 474854
rect 162490 474938 162726 475174
rect 162490 474618 162726 474854
rect 193210 474938 193446 475174
rect 193210 474618 193446 474854
rect 223930 474938 224166 475174
rect 223930 474618 224166 474854
rect 254650 474938 254886 475174
rect 254650 474618 254886 474854
rect 285370 474938 285606 475174
rect 285370 474618 285606 474854
rect 316090 474938 316326 475174
rect 316090 474618 316326 474854
rect 346810 474938 347046 475174
rect 346810 474618 347046 474854
rect 54970 471218 55206 471454
rect 54970 470898 55206 471134
rect 85690 471218 85926 471454
rect 85690 470898 85926 471134
rect 116410 471218 116646 471454
rect 116410 470898 116646 471134
rect 147130 471218 147366 471454
rect 147130 470898 147366 471134
rect 177850 471218 178086 471454
rect 177850 470898 178086 471134
rect 208570 471218 208806 471454
rect 208570 470898 208806 471134
rect 239290 471218 239526 471454
rect 239290 470898 239526 471134
rect 270010 471218 270246 471454
rect 270010 470898 270246 471134
rect 300730 471218 300966 471454
rect 300730 470898 300966 471134
rect 331450 471218 331686 471454
rect 331450 470898 331686 471134
rect 361826 471218 362062 471454
rect 362146 471218 362382 471454
rect 361826 470898 362062 471134
rect 362146 470898 362382 471134
rect 27866 461258 28102 461494
rect 28186 461258 28422 461494
rect 27866 460938 28102 461174
rect 28186 460938 28422 461174
rect 24250 435218 24486 435454
rect 24250 434898 24486 435134
rect 20426 417818 20662 418054
rect 20746 417818 20982 418054
rect 20426 417498 20662 417734
rect 20746 417498 20982 417734
rect 39610 438938 39846 439174
rect 39610 438618 39846 438854
rect 70330 438938 70566 439174
rect 70330 438618 70566 438854
rect 101050 438938 101286 439174
rect 101050 438618 101286 438854
rect 131770 438938 132006 439174
rect 131770 438618 132006 438854
rect 162490 438938 162726 439174
rect 162490 438618 162726 438854
rect 193210 438938 193446 439174
rect 193210 438618 193446 438854
rect 223930 438938 224166 439174
rect 223930 438618 224166 438854
rect 254650 438938 254886 439174
rect 254650 438618 254886 438854
rect 285370 438938 285606 439174
rect 285370 438618 285606 438854
rect 316090 438938 316326 439174
rect 316090 438618 316326 438854
rect 346810 438938 347046 439174
rect 346810 438618 347046 438854
rect 54970 435218 55206 435454
rect 54970 434898 55206 435134
rect 85690 435218 85926 435454
rect 85690 434898 85926 435134
rect 116410 435218 116646 435454
rect 116410 434898 116646 435134
rect 147130 435218 147366 435454
rect 147130 434898 147366 435134
rect 177850 435218 178086 435454
rect 177850 434898 178086 435134
rect 208570 435218 208806 435454
rect 208570 434898 208806 435134
rect 239290 435218 239526 435454
rect 239290 434898 239526 435134
rect 270010 435218 270246 435454
rect 270010 434898 270246 435134
rect 300730 435218 300966 435454
rect 300730 434898 300966 435134
rect 331450 435218 331686 435454
rect 331450 434898 331686 435134
rect 361826 435218 362062 435454
rect 362146 435218 362382 435454
rect 361826 434898 362062 435134
rect 362146 434898 362382 435134
rect 27866 425258 28102 425494
rect 28186 425258 28422 425494
rect 27866 424938 28102 425174
rect 28186 424938 28422 425174
rect 24250 399218 24486 399454
rect 24250 398898 24486 399134
rect 20426 381818 20662 382054
rect 20746 381818 20982 382054
rect 20426 381498 20662 381734
rect 20746 381498 20982 381734
rect 39610 402938 39846 403174
rect 39610 402618 39846 402854
rect 70330 402938 70566 403174
rect 70330 402618 70566 402854
rect 101050 402938 101286 403174
rect 101050 402618 101286 402854
rect 131770 402938 132006 403174
rect 131770 402618 132006 402854
rect 162490 402938 162726 403174
rect 162490 402618 162726 402854
rect 193210 402938 193446 403174
rect 193210 402618 193446 402854
rect 223930 402938 224166 403174
rect 223930 402618 224166 402854
rect 254650 402938 254886 403174
rect 254650 402618 254886 402854
rect 285370 402938 285606 403174
rect 285370 402618 285606 402854
rect 316090 402938 316326 403174
rect 316090 402618 316326 402854
rect 346810 402938 347046 403174
rect 346810 402618 347046 402854
rect 54970 399218 55206 399454
rect 54970 398898 55206 399134
rect 85690 399218 85926 399454
rect 85690 398898 85926 399134
rect 116410 399218 116646 399454
rect 116410 398898 116646 399134
rect 147130 399218 147366 399454
rect 147130 398898 147366 399134
rect 177850 399218 178086 399454
rect 177850 398898 178086 399134
rect 208570 399218 208806 399454
rect 208570 398898 208806 399134
rect 239290 399218 239526 399454
rect 239290 398898 239526 399134
rect 270010 399218 270246 399454
rect 270010 398898 270246 399134
rect 300730 399218 300966 399454
rect 300730 398898 300966 399134
rect 331450 399218 331686 399454
rect 331450 398898 331686 399134
rect 361826 399218 362062 399454
rect 362146 399218 362382 399454
rect 361826 398898 362062 399134
rect 362146 398898 362382 399134
rect 27866 389258 28102 389494
rect 28186 389258 28422 389494
rect 27866 388938 28102 389174
rect 28186 388938 28422 389174
rect 24250 363218 24486 363454
rect 24250 362898 24486 363134
rect 20426 345818 20662 346054
rect 20746 345818 20982 346054
rect 20426 345498 20662 345734
rect 20746 345498 20982 345734
rect 39610 366938 39846 367174
rect 39610 366618 39846 366854
rect 70330 366938 70566 367174
rect 70330 366618 70566 366854
rect 101050 366938 101286 367174
rect 101050 366618 101286 366854
rect 131770 366938 132006 367174
rect 131770 366618 132006 366854
rect 162490 366938 162726 367174
rect 162490 366618 162726 366854
rect 193210 366938 193446 367174
rect 193210 366618 193446 366854
rect 223930 366938 224166 367174
rect 223930 366618 224166 366854
rect 254650 366938 254886 367174
rect 254650 366618 254886 366854
rect 285370 366938 285606 367174
rect 285370 366618 285606 366854
rect 316090 366938 316326 367174
rect 316090 366618 316326 366854
rect 346810 366938 347046 367174
rect 346810 366618 347046 366854
rect 54970 363218 55206 363454
rect 54970 362898 55206 363134
rect 85690 363218 85926 363454
rect 85690 362898 85926 363134
rect 116410 363218 116646 363454
rect 116410 362898 116646 363134
rect 147130 363218 147366 363454
rect 147130 362898 147366 363134
rect 177850 363218 178086 363454
rect 177850 362898 178086 363134
rect 208570 363218 208806 363454
rect 208570 362898 208806 363134
rect 239290 363218 239526 363454
rect 239290 362898 239526 363134
rect 270010 363218 270246 363454
rect 270010 362898 270246 363134
rect 300730 363218 300966 363454
rect 300730 362898 300966 363134
rect 331450 363218 331686 363454
rect 331450 362898 331686 363134
rect 361826 363218 362062 363454
rect 362146 363218 362382 363454
rect 361826 362898 362062 363134
rect 362146 362898 362382 363134
rect 27866 353258 28102 353494
rect 28186 353258 28422 353494
rect 27866 352938 28102 353174
rect 28186 352938 28422 353174
rect 24250 327218 24486 327454
rect 24250 326898 24486 327134
rect 20426 309818 20662 310054
rect 20746 309818 20982 310054
rect 20426 309498 20662 309734
rect 20746 309498 20982 309734
rect 39610 330938 39846 331174
rect 39610 330618 39846 330854
rect 70330 330938 70566 331174
rect 70330 330618 70566 330854
rect 101050 330938 101286 331174
rect 101050 330618 101286 330854
rect 131770 330938 132006 331174
rect 131770 330618 132006 330854
rect 162490 330938 162726 331174
rect 162490 330618 162726 330854
rect 193210 330938 193446 331174
rect 193210 330618 193446 330854
rect 223930 330938 224166 331174
rect 223930 330618 224166 330854
rect 254650 330938 254886 331174
rect 254650 330618 254886 330854
rect 285370 330938 285606 331174
rect 285370 330618 285606 330854
rect 316090 330938 316326 331174
rect 316090 330618 316326 330854
rect 346810 330938 347046 331174
rect 346810 330618 347046 330854
rect 54970 327218 55206 327454
rect 54970 326898 55206 327134
rect 85690 327218 85926 327454
rect 85690 326898 85926 327134
rect 116410 327218 116646 327454
rect 116410 326898 116646 327134
rect 147130 327218 147366 327454
rect 147130 326898 147366 327134
rect 177850 327218 178086 327454
rect 177850 326898 178086 327134
rect 208570 327218 208806 327454
rect 208570 326898 208806 327134
rect 239290 327218 239526 327454
rect 239290 326898 239526 327134
rect 270010 327218 270246 327454
rect 270010 326898 270246 327134
rect 300730 327218 300966 327454
rect 300730 326898 300966 327134
rect 331450 327218 331686 327454
rect 331450 326898 331686 327134
rect 361826 327218 362062 327454
rect 362146 327218 362382 327454
rect 361826 326898 362062 327134
rect 362146 326898 362382 327134
rect 27866 317258 28102 317494
rect 28186 317258 28422 317494
rect 27866 316938 28102 317174
rect 28186 316938 28422 317174
rect 24250 291218 24486 291454
rect 24250 290898 24486 291134
rect 20426 273818 20662 274054
rect 20746 273818 20982 274054
rect 20426 273498 20662 273734
rect 20746 273498 20982 273734
rect 39610 294938 39846 295174
rect 39610 294618 39846 294854
rect 70330 294938 70566 295174
rect 70330 294618 70566 294854
rect 101050 294938 101286 295174
rect 101050 294618 101286 294854
rect 131770 294938 132006 295174
rect 131770 294618 132006 294854
rect 162490 294938 162726 295174
rect 162490 294618 162726 294854
rect 193210 294938 193446 295174
rect 193210 294618 193446 294854
rect 223930 294938 224166 295174
rect 223930 294618 224166 294854
rect 254650 294938 254886 295174
rect 254650 294618 254886 294854
rect 285370 294938 285606 295174
rect 285370 294618 285606 294854
rect 316090 294938 316326 295174
rect 316090 294618 316326 294854
rect 346810 294938 347046 295174
rect 346810 294618 347046 294854
rect 54970 291218 55206 291454
rect 54970 290898 55206 291134
rect 85690 291218 85926 291454
rect 85690 290898 85926 291134
rect 116410 291218 116646 291454
rect 116410 290898 116646 291134
rect 147130 291218 147366 291454
rect 147130 290898 147366 291134
rect 177850 291218 178086 291454
rect 177850 290898 178086 291134
rect 208570 291218 208806 291454
rect 208570 290898 208806 291134
rect 239290 291218 239526 291454
rect 239290 290898 239526 291134
rect 270010 291218 270246 291454
rect 270010 290898 270246 291134
rect 300730 291218 300966 291454
rect 300730 290898 300966 291134
rect 331450 291218 331686 291454
rect 331450 290898 331686 291134
rect 361826 291218 362062 291454
rect 362146 291218 362382 291454
rect 361826 290898 362062 291134
rect 362146 290898 362382 291134
rect 27866 281258 28102 281494
rect 28186 281258 28422 281494
rect 27866 280938 28102 281174
rect 28186 280938 28422 281174
rect 24250 255218 24486 255454
rect 24250 254898 24486 255134
rect 20426 237818 20662 238054
rect 20746 237818 20982 238054
rect 20426 237498 20662 237734
rect 20746 237498 20982 237734
rect 39610 258938 39846 259174
rect 39610 258618 39846 258854
rect 70330 258938 70566 259174
rect 70330 258618 70566 258854
rect 101050 258938 101286 259174
rect 101050 258618 101286 258854
rect 131770 258938 132006 259174
rect 131770 258618 132006 258854
rect 162490 258938 162726 259174
rect 162490 258618 162726 258854
rect 193210 258938 193446 259174
rect 193210 258618 193446 258854
rect 223930 258938 224166 259174
rect 223930 258618 224166 258854
rect 254650 258938 254886 259174
rect 254650 258618 254886 258854
rect 285370 258938 285606 259174
rect 285370 258618 285606 258854
rect 316090 258938 316326 259174
rect 316090 258618 316326 258854
rect 346810 258938 347046 259174
rect 346810 258618 347046 258854
rect 54970 255218 55206 255454
rect 54970 254898 55206 255134
rect 85690 255218 85926 255454
rect 85690 254898 85926 255134
rect 116410 255218 116646 255454
rect 116410 254898 116646 255134
rect 147130 255218 147366 255454
rect 147130 254898 147366 255134
rect 177850 255218 178086 255454
rect 177850 254898 178086 255134
rect 208570 255218 208806 255454
rect 208570 254898 208806 255134
rect 239290 255218 239526 255454
rect 239290 254898 239526 255134
rect 270010 255218 270246 255454
rect 270010 254898 270246 255134
rect 300730 255218 300966 255454
rect 300730 254898 300966 255134
rect 331450 255218 331686 255454
rect 331450 254898 331686 255134
rect 361826 255218 362062 255454
rect 362146 255218 362382 255454
rect 361826 254898 362062 255134
rect 362146 254898 362382 255134
rect 27866 245258 28102 245494
rect 28186 245258 28422 245494
rect 27866 244938 28102 245174
rect 28186 244938 28422 245174
rect 24250 219218 24486 219454
rect 24250 218898 24486 219134
rect 20426 201818 20662 202054
rect 20746 201818 20982 202054
rect 20426 201498 20662 201734
rect 20746 201498 20982 201734
rect 39610 222938 39846 223174
rect 39610 222618 39846 222854
rect 70330 222938 70566 223174
rect 70330 222618 70566 222854
rect 101050 222938 101286 223174
rect 101050 222618 101286 222854
rect 131770 222938 132006 223174
rect 131770 222618 132006 222854
rect 162490 222938 162726 223174
rect 162490 222618 162726 222854
rect 193210 222938 193446 223174
rect 193210 222618 193446 222854
rect 223930 222938 224166 223174
rect 223930 222618 224166 222854
rect 254650 222938 254886 223174
rect 254650 222618 254886 222854
rect 285370 222938 285606 223174
rect 285370 222618 285606 222854
rect 316090 222938 316326 223174
rect 316090 222618 316326 222854
rect 346810 222938 347046 223174
rect 346810 222618 347046 222854
rect 54970 219218 55206 219454
rect 54970 218898 55206 219134
rect 85690 219218 85926 219454
rect 85690 218898 85926 219134
rect 116410 219218 116646 219454
rect 116410 218898 116646 219134
rect 147130 219218 147366 219454
rect 147130 218898 147366 219134
rect 177850 219218 178086 219454
rect 177850 218898 178086 219134
rect 208570 219218 208806 219454
rect 208570 218898 208806 219134
rect 239290 219218 239526 219454
rect 239290 218898 239526 219134
rect 270010 219218 270246 219454
rect 270010 218898 270246 219134
rect 300730 219218 300966 219454
rect 300730 218898 300966 219134
rect 331450 219218 331686 219454
rect 331450 218898 331686 219134
rect 361826 219218 362062 219454
rect 362146 219218 362382 219454
rect 361826 218898 362062 219134
rect 362146 218898 362382 219134
rect 27866 209258 28102 209494
rect 28186 209258 28422 209494
rect 27866 208938 28102 209174
rect 28186 208938 28422 209174
rect 24250 183218 24486 183454
rect 24250 182898 24486 183134
rect 20426 165818 20662 166054
rect 20746 165818 20982 166054
rect 20426 165498 20662 165734
rect 20746 165498 20982 165734
rect 39610 186938 39846 187174
rect 39610 186618 39846 186854
rect 70330 186938 70566 187174
rect 70330 186618 70566 186854
rect 101050 186938 101286 187174
rect 101050 186618 101286 186854
rect 131770 186938 132006 187174
rect 131770 186618 132006 186854
rect 162490 186938 162726 187174
rect 162490 186618 162726 186854
rect 193210 186938 193446 187174
rect 193210 186618 193446 186854
rect 223930 186938 224166 187174
rect 223930 186618 224166 186854
rect 254650 186938 254886 187174
rect 254650 186618 254886 186854
rect 285370 186938 285606 187174
rect 285370 186618 285606 186854
rect 316090 186938 316326 187174
rect 316090 186618 316326 186854
rect 346810 186938 347046 187174
rect 346810 186618 347046 186854
rect 54970 183218 55206 183454
rect 54970 182898 55206 183134
rect 85690 183218 85926 183454
rect 85690 182898 85926 183134
rect 116410 183218 116646 183454
rect 116410 182898 116646 183134
rect 147130 183218 147366 183454
rect 147130 182898 147366 183134
rect 177850 183218 178086 183454
rect 177850 182898 178086 183134
rect 208570 183218 208806 183454
rect 208570 182898 208806 183134
rect 239290 183218 239526 183454
rect 239290 182898 239526 183134
rect 270010 183218 270246 183454
rect 270010 182898 270246 183134
rect 300730 183218 300966 183454
rect 300730 182898 300966 183134
rect 331450 183218 331686 183454
rect 331450 182898 331686 183134
rect 361826 183218 362062 183454
rect 362146 183218 362382 183454
rect 361826 182898 362062 183134
rect 362146 182898 362382 183134
rect 27866 173258 28102 173494
rect 28186 173258 28422 173494
rect 27866 172938 28102 173174
rect 28186 172938 28422 173174
rect 24250 147218 24486 147454
rect 24250 146898 24486 147134
rect 20426 129818 20662 130054
rect 20746 129818 20982 130054
rect 20426 129498 20662 129734
rect 20746 129498 20982 129734
rect 39610 150938 39846 151174
rect 39610 150618 39846 150854
rect 70330 150938 70566 151174
rect 70330 150618 70566 150854
rect 101050 150938 101286 151174
rect 101050 150618 101286 150854
rect 131770 150938 132006 151174
rect 131770 150618 132006 150854
rect 162490 150938 162726 151174
rect 162490 150618 162726 150854
rect 193210 150938 193446 151174
rect 193210 150618 193446 150854
rect 223930 150938 224166 151174
rect 223930 150618 224166 150854
rect 254650 150938 254886 151174
rect 254650 150618 254886 150854
rect 285370 150938 285606 151174
rect 285370 150618 285606 150854
rect 316090 150938 316326 151174
rect 316090 150618 316326 150854
rect 346810 150938 347046 151174
rect 346810 150618 347046 150854
rect 54970 147218 55206 147454
rect 54970 146898 55206 147134
rect 85690 147218 85926 147454
rect 85690 146898 85926 147134
rect 116410 147218 116646 147454
rect 116410 146898 116646 147134
rect 147130 147218 147366 147454
rect 147130 146898 147366 147134
rect 177850 147218 178086 147454
rect 177850 146898 178086 147134
rect 208570 147218 208806 147454
rect 208570 146898 208806 147134
rect 239290 147218 239526 147454
rect 239290 146898 239526 147134
rect 270010 147218 270246 147454
rect 270010 146898 270246 147134
rect 300730 147218 300966 147454
rect 300730 146898 300966 147134
rect 331450 147218 331686 147454
rect 331450 146898 331686 147134
rect 361826 147218 362062 147454
rect 362146 147218 362382 147454
rect 361826 146898 362062 147134
rect 362146 146898 362382 147134
rect 27866 137258 28102 137494
rect 28186 137258 28422 137494
rect 27866 136938 28102 137174
rect 28186 136938 28422 137174
rect 24250 111218 24486 111454
rect 24250 110898 24486 111134
rect 20426 93818 20662 94054
rect 20746 93818 20982 94054
rect 20426 93498 20662 93734
rect 20746 93498 20982 93734
rect 39610 114938 39846 115174
rect 39610 114618 39846 114854
rect 70330 114938 70566 115174
rect 70330 114618 70566 114854
rect 101050 114938 101286 115174
rect 101050 114618 101286 114854
rect 131770 114938 132006 115174
rect 131770 114618 132006 114854
rect 162490 114938 162726 115174
rect 162490 114618 162726 114854
rect 193210 114938 193446 115174
rect 193210 114618 193446 114854
rect 223930 114938 224166 115174
rect 223930 114618 224166 114854
rect 254650 114938 254886 115174
rect 254650 114618 254886 114854
rect 285370 114938 285606 115174
rect 285370 114618 285606 114854
rect 316090 114938 316326 115174
rect 316090 114618 316326 114854
rect 346810 114938 347046 115174
rect 346810 114618 347046 114854
rect 54970 111218 55206 111454
rect 54970 110898 55206 111134
rect 85690 111218 85926 111454
rect 85690 110898 85926 111134
rect 116410 111218 116646 111454
rect 116410 110898 116646 111134
rect 147130 111218 147366 111454
rect 147130 110898 147366 111134
rect 177850 111218 178086 111454
rect 177850 110898 178086 111134
rect 208570 111218 208806 111454
rect 208570 110898 208806 111134
rect 239290 111218 239526 111454
rect 239290 110898 239526 111134
rect 270010 111218 270246 111454
rect 270010 110898 270246 111134
rect 300730 111218 300966 111454
rect 300730 110898 300966 111134
rect 331450 111218 331686 111454
rect 331450 110898 331686 111134
rect 361826 111218 362062 111454
rect 362146 111218 362382 111454
rect 361826 110898 362062 111134
rect 362146 110898 362382 111134
rect 27866 101258 28102 101494
rect 28186 101258 28422 101494
rect 27866 100938 28102 101174
rect 28186 100938 28422 101174
rect 24250 75218 24486 75454
rect 24250 74898 24486 75134
rect 20426 57818 20662 58054
rect 20746 57818 20982 58054
rect 20426 57498 20662 57734
rect 20746 57498 20982 57734
rect 39610 78938 39846 79174
rect 39610 78618 39846 78854
rect 70330 78938 70566 79174
rect 70330 78618 70566 78854
rect 101050 78938 101286 79174
rect 101050 78618 101286 78854
rect 131770 78938 132006 79174
rect 131770 78618 132006 78854
rect 162490 78938 162726 79174
rect 162490 78618 162726 78854
rect 193210 78938 193446 79174
rect 193210 78618 193446 78854
rect 223930 78938 224166 79174
rect 223930 78618 224166 78854
rect 254650 78938 254886 79174
rect 254650 78618 254886 78854
rect 285370 78938 285606 79174
rect 285370 78618 285606 78854
rect 316090 78938 316326 79174
rect 316090 78618 316326 78854
rect 346810 78938 347046 79174
rect 346810 78618 347046 78854
rect 54970 75218 55206 75454
rect 54970 74898 55206 75134
rect 85690 75218 85926 75454
rect 85690 74898 85926 75134
rect 116410 75218 116646 75454
rect 116410 74898 116646 75134
rect 147130 75218 147366 75454
rect 147130 74898 147366 75134
rect 177850 75218 178086 75454
rect 177850 74898 178086 75134
rect 208570 75218 208806 75454
rect 208570 74898 208806 75134
rect 239290 75218 239526 75454
rect 239290 74898 239526 75134
rect 270010 75218 270246 75454
rect 270010 74898 270246 75134
rect 300730 75218 300966 75454
rect 300730 74898 300966 75134
rect 331450 75218 331686 75454
rect 331450 74898 331686 75134
rect 361826 75218 362062 75454
rect 362146 75218 362382 75454
rect 361826 74898 362062 75134
rect 362146 74898 362382 75134
rect 27866 65258 28102 65494
rect 28186 65258 28422 65494
rect 27866 64938 28102 65174
rect 28186 64938 28422 65174
rect 20426 21818 20662 22054
rect 20746 21818 20982 22054
rect 20426 21498 20662 21734
rect 20746 21498 20982 21734
rect 20426 -5382 20662 -5146
rect 20746 -5382 20982 -5146
rect 20426 -5702 20662 -5466
rect 20746 -5702 20982 -5466
rect 24146 25538 24382 25774
rect 24466 25538 24702 25774
rect 24146 25218 24382 25454
rect 24466 25218 24702 25454
rect 24146 -6342 24382 -6106
rect 24466 -6342 24702 -6106
rect 24146 -6662 24382 -6426
rect 24466 -6662 24702 -6426
rect 27866 29258 28102 29494
rect 28186 29258 28422 29494
rect 27866 28938 28102 29174
rect 28186 28938 28422 29174
rect 27866 -7302 28102 -7066
rect 28186 -7302 28422 -7066
rect 27866 -7622 28102 -7386
rect 28186 -7622 28422 -7386
rect 37826 39218 38062 39454
rect 38146 39218 38382 39454
rect 37826 38898 38062 39134
rect 38146 38898 38382 39134
rect 37826 3218 38062 3454
rect 38146 3218 38382 3454
rect 37826 2898 38062 3134
rect 38146 2898 38382 3134
rect 37826 -582 38062 -346
rect 38146 -582 38382 -346
rect 37826 -902 38062 -666
rect 38146 -902 38382 -666
rect 41546 42938 41782 43174
rect 41866 42938 42102 43174
rect 41546 42618 41782 42854
rect 41866 42618 42102 42854
rect 41546 6938 41782 7174
rect 41866 6938 42102 7174
rect 41546 6618 41782 6854
rect 41866 6618 42102 6854
rect 41546 -1542 41782 -1306
rect 41866 -1542 42102 -1306
rect 41546 -1862 41782 -1626
rect 41866 -1862 42102 -1626
rect 45266 46658 45502 46894
rect 45586 46658 45822 46894
rect 45266 46338 45502 46574
rect 45586 46338 45822 46574
rect 45266 10658 45502 10894
rect 45586 10658 45822 10894
rect 45266 10338 45502 10574
rect 45586 10338 45822 10574
rect 45266 -2502 45502 -2266
rect 45586 -2502 45822 -2266
rect 45266 -2822 45502 -2586
rect 45586 -2822 45822 -2586
rect 48986 14378 49222 14614
rect 49306 14378 49542 14614
rect 48986 14058 49222 14294
rect 49306 14058 49542 14294
rect 48986 -3462 49222 -3226
rect 49306 -3462 49542 -3226
rect 48986 -3782 49222 -3546
rect 49306 -3782 49542 -3546
rect 52706 18098 52942 18334
rect 53026 18098 53262 18334
rect 52706 17778 52942 18014
rect 53026 17778 53262 18014
rect 52706 -4422 52942 -4186
rect 53026 -4422 53262 -4186
rect 52706 -4742 52942 -4506
rect 53026 -4742 53262 -4506
rect 56426 21818 56662 22054
rect 56746 21818 56982 22054
rect 56426 21498 56662 21734
rect 56746 21498 56982 21734
rect 56426 -5382 56662 -5146
rect 56746 -5382 56982 -5146
rect 56426 -5702 56662 -5466
rect 56746 -5702 56982 -5466
rect 60146 25538 60382 25774
rect 60466 25538 60702 25774
rect 60146 25218 60382 25454
rect 60466 25218 60702 25454
rect 60146 -6342 60382 -6106
rect 60466 -6342 60702 -6106
rect 60146 -6662 60382 -6426
rect 60466 -6662 60702 -6426
rect 63866 29258 64102 29494
rect 64186 29258 64422 29494
rect 63866 28938 64102 29174
rect 64186 28938 64422 29174
rect 63866 -7302 64102 -7066
rect 64186 -7302 64422 -7066
rect 63866 -7622 64102 -7386
rect 64186 -7622 64422 -7386
rect 73826 39218 74062 39454
rect 74146 39218 74382 39454
rect 73826 38898 74062 39134
rect 74146 38898 74382 39134
rect 73826 3218 74062 3454
rect 74146 3218 74382 3454
rect 73826 2898 74062 3134
rect 74146 2898 74382 3134
rect 73826 -582 74062 -346
rect 74146 -582 74382 -346
rect 73826 -902 74062 -666
rect 74146 -902 74382 -666
rect 77546 42938 77782 43174
rect 77866 42938 78102 43174
rect 77546 42618 77782 42854
rect 77866 42618 78102 42854
rect 77546 6938 77782 7174
rect 77866 6938 78102 7174
rect 77546 6618 77782 6854
rect 77866 6618 78102 6854
rect 77546 -1542 77782 -1306
rect 77866 -1542 78102 -1306
rect 77546 -1862 77782 -1626
rect 77866 -1862 78102 -1626
rect 81266 46658 81502 46894
rect 81586 46658 81822 46894
rect 81266 46338 81502 46574
rect 81586 46338 81822 46574
rect 81266 10658 81502 10894
rect 81586 10658 81822 10894
rect 81266 10338 81502 10574
rect 81586 10338 81822 10574
rect 81266 -2502 81502 -2266
rect 81586 -2502 81822 -2266
rect 81266 -2822 81502 -2586
rect 81586 -2822 81822 -2586
rect 84986 14378 85222 14614
rect 85306 14378 85542 14614
rect 84986 14058 85222 14294
rect 85306 14058 85542 14294
rect 84986 -3462 85222 -3226
rect 85306 -3462 85542 -3226
rect 84986 -3782 85222 -3546
rect 85306 -3782 85542 -3546
rect 88706 18098 88942 18334
rect 89026 18098 89262 18334
rect 88706 17778 88942 18014
rect 89026 17778 89262 18014
rect 88706 -4422 88942 -4186
rect 89026 -4422 89262 -4186
rect 88706 -4742 88942 -4506
rect 89026 -4742 89262 -4506
rect 92426 21818 92662 22054
rect 92746 21818 92982 22054
rect 92426 21498 92662 21734
rect 92746 21498 92982 21734
rect 92426 -5382 92662 -5146
rect 92746 -5382 92982 -5146
rect 92426 -5702 92662 -5466
rect 92746 -5702 92982 -5466
rect 96146 25538 96382 25774
rect 96466 25538 96702 25774
rect 96146 25218 96382 25454
rect 96466 25218 96702 25454
rect 96146 -6342 96382 -6106
rect 96466 -6342 96702 -6106
rect 96146 -6662 96382 -6426
rect 96466 -6662 96702 -6426
rect 99866 29258 100102 29494
rect 100186 29258 100422 29494
rect 99866 28938 100102 29174
rect 100186 28938 100422 29174
rect 99866 -7302 100102 -7066
rect 100186 -7302 100422 -7066
rect 99866 -7622 100102 -7386
rect 100186 -7622 100422 -7386
rect 109826 39218 110062 39454
rect 110146 39218 110382 39454
rect 109826 38898 110062 39134
rect 110146 38898 110382 39134
rect 109826 3218 110062 3454
rect 110146 3218 110382 3454
rect 109826 2898 110062 3134
rect 110146 2898 110382 3134
rect 109826 -582 110062 -346
rect 110146 -582 110382 -346
rect 109826 -902 110062 -666
rect 110146 -902 110382 -666
rect 113546 42938 113782 43174
rect 113866 42938 114102 43174
rect 113546 42618 113782 42854
rect 113866 42618 114102 42854
rect 113546 6938 113782 7174
rect 113866 6938 114102 7174
rect 113546 6618 113782 6854
rect 113866 6618 114102 6854
rect 113546 -1542 113782 -1306
rect 113866 -1542 114102 -1306
rect 113546 -1862 113782 -1626
rect 113866 -1862 114102 -1626
rect 117266 46658 117502 46894
rect 117586 46658 117822 46894
rect 117266 46338 117502 46574
rect 117586 46338 117822 46574
rect 117266 10658 117502 10894
rect 117586 10658 117822 10894
rect 117266 10338 117502 10574
rect 117586 10338 117822 10574
rect 117266 -2502 117502 -2266
rect 117586 -2502 117822 -2266
rect 117266 -2822 117502 -2586
rect 117586 -2822 117822 -2586
rect 120986 14378 121222 14614
rect 121306 14378 121542 14614
rect 120986 14058 121222 14294
rect 121306 14058 121542 14294
rect 120986 -3462 121222 -3226
rect 121306 -3462 121542 -3226
rect 120986 -3782 121222 -3546
rect 121306 -3782 121542 -3546
rect 124706 18098 124942 18334
rect 125026 18098 125262 18334
rect 124706 17778 124942 18014
rect 125026 17778 125262 18014
rect 124706 -4422 124942 -4186
rect 125026 -4422 125262 -4186
rect 124706 -4742 124942 -4506
rect 125026 -4742 125262 -4506
rect 128426 21818 128662 22054
rect 128746 21818 128982 22054
rect 128426 21498 128662 21734
rect 128746 21498 128982 21734
rect 128426 -5382 128662 -5146
rect 128746 -5382 128982 -5146
rect 128426 -5702 128662 -5466
rect 128746 -5702 128982 -5466
rect 132146 25538 132382 25774
rect 132466 25538 132702 25774
rect 132146 25218 132382 25454
rect 132466 25218 132702 25454
rect 132146 -6342 132382 -6106
rect 132466 -6342 132702 -6106
rect 132146 -6662 132382 -6426
rect 132466 -6662 132702 -6426
rect 135866 29258 136102 29494
rect 136186 29258 136422 29494
rect 135866 28938 136102 29174
rect 136186 28938 136422 29174
rect 135866 -7302 136102 -7066
rect 136186 -7302 136422 -7066
rect 135866 -7622 136102 -7386
rect 136186 -7622 136422 -7386
rect 145826 39218 146062 39454
rect 146146 39218 146382 39454
rect 145826 38898 146062 39134
rect 146146 38898 146382 39134
rect 145826 3218 146062 3454
rect 146146 3218 146382 3454
rect 145826 2898 146062 3134
rect 146146 2898 146382 3134
rect 145826 -582 146062 -346
rect 146146 -582 146382 -346
rect 145826 -902 146062 -666
rect 146146 -902 146382 -666
rect 149546 42938 149782 43174
rect 149866 42938 150102 43174
rect 149546 42618 149782 42854
rect 149866 42618 150102 42854
rect 149546 6938 149782 7174
rect 149866 6938 150102 7174
rect 149546 6618 149782 6854
rect 149866 6618 150102 6854
rect 149546 -1542 149782 -1306
rect 149866 -1542 150102 -1306
rect 149546 -1862 149782 -1626
rect 149866 -1862 150102 -1626
rect 153266 46658 153502 46894
rect 153586 46658 153822 46894
rect 153266 46338 153502 46574
rect 153586 46338 153822 46574
rect 153266 10658 153502 10894
rect 153586 10658 153822 10894
rect 153266 10338 153502 10574
rect 153586 10338 153822 10574
rect 153266 -2502 153502 -2266
rect 153586 -2502 153822 -2266
rect 153266 -2822 153502 -2586
rect 153586 -2822 153822 -2586
rect 156986 14378 157222 14614
rect 157306 14378 157542 14614
rect 156986 14058 157222 14294
rect 157306 14058 157542 14294
rect 156986 -3462 157222 -3226
rect 157306 -3462 157542 -3226
rect 156986 -3782 157222 -3546
rect 157306 -3782 157542 -3546
rect 160706 18098 160942 18334
rect 161026 18098 161262 18334
rect 160706 17778 160942 18014
rect 161026 17778 161262 18014
rect 160706 -4422 160942 -4186
rect 161026 -4422 161262 -4186
rect 160706 -4742 160942 -4506
rect 161026 -4742 161262 -4506
rect 164426 21818 164662 22054
rect 164746 21818 164982 22054
rect 164426 21498 164662 21734
rect 164746 21498 164982 21734
rect 164426 -5382 164662 -5146
rect 164746 -5382 164982 -5146
rect 164426 -5702 164662 -5466
rect 164746 -5702 164982 -5466
rect 168146 25538 168382 25774
rect 168466 25538 168702 25774
rect 168146 25218 168382 25454
rect 168466 25218 168702 25454
rect 168146 -6342 168382 -6106
rect 168466 -6342 168702 -6106
rect 168146 -6662 168382 -6426
rect 168466 -6662 168702 -6426
rect 171866 29258 172102 29494
rect 172186 29258 172422 29494
rect 171866 28938 172102 29174
rect 172186 28938 172422 29174
rect 171866 -7302 172102 -7066
rect 172186 -7302 172422 -7066
rect 171866 -7622 172102 -7386
rect 172186 -7622 172422 -7386
rect 181826 39218 182062 39454
rect 182146 39218 182382 39454
rect 181826 38898 182062 39134
rect 182146 38898 182382 39134
rect 181826 3218 182062 3454
rect 182146 3218 182382 3454
rect 181826 2898 182062 3134
rect 182146 2898 182382 3134
rect 181826 -582 182062 -346
rect 182146 -582 182382 -346
rect 181826 -902 182062 -666
rect 182146 -902 182382 -666
rect 185546 42938 185782 43174
rect 185866 42938 186102 43174
rect 185546 42618 185782 42854
rect 185866 42618 186102 42854
rect 185546 6938 185782 7174
rect 185866 6938 186102 7174
rect 185546 6618 185782 6854
rect 185866 6618 186102 6854
rect 185546 -1542 185782 -1306
rect 185866 -1542 186102 -1306
rect 185546 -1862 185782 -1626
rect 185866 -1862 186102 -1626
rect 189266 46658 189502 46894
rect 189586 46658 189822 46894
rect 189266 46338 189502 46574
rect 189586 46338 189822 46574
rect 189266 10658 189502 10894
rect 189586 10658 189822 10894
rect 189266 10338 189502 10574
rect 189586 10338 189822 10574
rect 189266 -2502 189502 -2266
rect 189586 -2502 189822 -2266
rect 189266 -2822 189502 -2586
rect 189586 -2822 189822 -2586
rect 192986 14378 193222 14614
rect 193306 14378 193542 14614
rect 192986 14058 193222 14294
rect 193306 14058 193542 14294
rect 192986 -3462 193222 -3226
rect 193306 -3462 193542 -3226
rect 192986 -3782 193222 -3546
rect 193306 -3782 193542 -3546
rect 196706 18098 196942 18334
rect 197026 18098 197262 18334
rect 196706 17778 196942 18014
rect 197026 17778 197262 18014
rect 196706 -4422 196942 -4186
rect 197026 -4422 197262 -4186
rect 196706 -4742 196942 -4506
rect 197026 -4742 197262 -4506
rect 200426 21818 200662 22054
rect 200746 21818 200982 22054
rect 200426 21498 200662 21734
rect 200746 21498 200982 21734
rect 200426 -5382 200662 -5146
rect 200746 -5382 200982 -5146
rect 200426 -5702 200662 -5466
rect 200746 -5702 200982 -5466
rect 204146 25538 204382 25774
rect 204466 25538 204702 25774
rect 204146 25218 204382 25454
rect 204466 25218 204702 25454
rect 204146 -6342 204382 -6106
rect 204466 -6342 204702 -6106
rect 204146 -6662 204382 -6426
rect 204466 -6662 204702 -6426
rect 207866 29258 208102 29494
rect 208186 29258 208422 29494
rect 207866 28938 208102 29174
rect 208186 28938 208422 29174
rect 207866 -7302 208102 -7066
rect 208186 -7302 208422 -7066
rect 207866 -7622 208102 -7386
rect 208186 -7622 208422 -7386
rect 217826 39218 218062 39454
rect 218146 39218 218382 39454
rect 217826 38898 218062 39134
rect 218146 38898 218382 39134
rect 217826 3218 218062 3454
rect 218146 3218 218382 3454
rect 217826 2898 218062 3134
rect 218146 2898 218382 3134
rect 217826 -582 218062 -346
rect 218146 -582 218382 -346
rect 217826 -902 218062 -666
rect 218146 -902 218382 -666
rect 221546 42938 221782 43174
rect 221866 42938 222102 43174
rect 221546 42618 221782 42854
rect 221866 42618 222102 42854
rect 221546 6938 221782 7174
rect 221866 6938 222102 7174
rect 221546 6618 221782 6854
rect 221866 6618 222102 6854
rect 221546 -1542 221782 -1306
rect 221866 -1542 222102 -1306
rect 221546 -1862 221782 -1626
rect 221866 -1862 222102 -1626
rect 225266 46658 225502 46894
rect 225586 46658 225822 46894
rect 225266 46338 225502 46574
rect 225586 46338 225822 46574
rect 225266 10658 225502 10894
rect 225586 10658 225822 10894
rect 225266 10338 225502 10574
rect 225586 10338 225822 10574
rect 225266 -2502 225502 -2266
rect 225586 -2502 225822 -2266
rect 225266 -2822 225502 -2586
rect 225586 -2822 225822 -2586
rect 228986 14378 229222 14614
rect 229306 14378 229542 14614
rect 228986 14058 229222 14294
rect 229306 14058 229542 14294
rect 228986 -3462 229222 -3226
rect 229306 -3462 229542 -3226
rect 228986 -3782 229222 -3546
rect 229306 -3782 229542 -3546
rect 232706 18098 232942 18334
rect 233026 18098 233262 18334
rect 232706 17778 232942 18014
rect 233026 17778 233262 18014
rect 232706 -4422 232942 -4186
rect 233026 -4422 233262 -4186
rect 232706 -4742 232942 -4506
rect 233026 -4742 233262 -4506
rect 236426 21818 236662 22054
rect 236746 21818 236982 22054
rect 236426 21498 236662 21734
rect 236746 21498 236982 21734
rect 236426 -5382 236662 -5146
rect 236746 -5382 236982 -5146
rect 236426 -5702 236662 -5466
rect 236746 -5702 236982 -5466
rect 240146 25538 240382 25774
rect 240466 25538 240702 25774
rect 240146 25218 240382 25454
rect 240466 25218 240702 25454
rect 240146 -6342 240382 -6106
rect 240466 -6342 240702 -6106
rect 240146 -6662 240382 -6426
rect 240466 -6662 240702 -6426
rect 243866 29258 244102 29494
rect 244186 29258 244422 29494
rect 243866 28938 244102 29174
rect 244186 28938 244422 29174
rect 243866 -7302 244102 -7066
rect 244186 -7302 244422 -7066
rect 243866 -7622 244102 -7386
rect 244186 -7622 244422 -7386
rect 253826 39218 254062 39454
rect 254146 39218 254382 39454
rect 253826 38898 254062 39134
rect 254146 38898 254382 39134
rect 253826 3218 254062 3454
rect 254146 3218 254382 3454
rect 253826 2898 254062 3134
rect 254146 2898 254382 3134
rect 253826 -582 254062 -346
rect 254146 -582 254382 -346
rect 253826 -902 254062 -666
rect 254146 -902 254382 -666
rect 257546 42938 257782 43174
rect 257866 42938 258102 43174
rect 257546 42618 257782 42854
rect 257866 42618 258102 42854
rect 257546 6938 257782 7174
rect 257866 6938 258102 7174
rect 257546 6618 257782 6854
rect 257866 6618 258102 6854
rect 257546 -1542 257782 -1306
rect 257866 -1542 258102 -1306
rect 257546 -1862 257782 -1626
rect 257866 -1862 258102 -1626
rect 261266 46658 261502 46894
rect 261586 46658 261822 46894
rect 261266 46338 261502 46574
rect 261586 46338 261822 46574
rect 261266 10658 261502 10894
rect 261586 10658 261822 10894
rect 261266 10338 261502 10574
rect 261586 10338 261822 10574
rect 261266 -2502 261502 -2266
rect 261586 -2502 261822 -2266
rect 261266 -2822 261502 -2586
rect 261586 -2822 261822 -2586
rect 264986 14378 265222 14614
rect 265306 14378 265542 14614
rect 264986 14058 265222 14294
rect 265306 14058 265542 14294
rect 264986 -3462 265222 -3226
rect 265306 -3462 265542 -3226
rect 264986 -3782 265222 -3546
rect 265306 -3782 265542 -3546
rect 268706 18098 268942 18334
rect 269026 18098 269262 18334
rect 268706 17778 268942 18014
rect 269026 17778 269262 18014
rect 268706 -4422 268942 -4186
rect 269026 -4422 269262 -4186
rect 268706 -4742 268942 -4506
rect 269026 -4742 269262 -4506
rect 272426 21818 272662 22054
rect 272746 21818 272982 22054
rect 272426 21498 272662 21734
rect 272746 21498 272982 21734
rect 272426 -5382 272662 -5146
rect 272746 -5382 272982 -5146
rect 272426 -5702 272662 -5466
rect 272746 -5702 272982 -5466
rect 276146 25538 276382 25774
rect 276466 25538 276702 25774
rect 276146 25218 276382 25454
rect 276466 25218 276702 25454
rect 276146 -6342 276382 -6106
rect 276466 -6342 276702 -6106
rect 276146 -6662 276382 -6426
rect 276466 -6662 276702 -6426
rect 279866 29258 280102 29494
rect 280186 29258 280422 29494
rect 279866 28938 280102 29174
rect 280186 28938 280422 29174
rect 279866 -7302 280102 -7066
rect 280186 -7302 280422 -7066
rect 279866 -7622 280102 -7386
rect 280186 -7622 280422 -7386
rect 289826 39218 290062 39454
rect 290146 39218 290382 39454
rect 289826 38898 290062 39134
rect 290146 38898 290382 39134
rect 289826 3218 290062 3454
rect 290146 3218 290382 3454
rect 289826 2898 290062 3134
rect 290146 2898 290382 3134
rect 289826 -582 290062 -346
rect 290146 -582 290382 -346
rect 289826 -902 290062 -666
rect 290146 -902 290382 -666
rect 293546 42938 293782 43174
rect 293866 42938 294102 43174
rect 293546 42618 293782 42854
rect 293866 42618 294102 42854
rect 293546 6938 293782 7174
rect 293866 6938 294102 7174
rect 293546 6618 293782 6854
rect 293866 6618 294102 6854
rect 293546 -1542 293782 -1306
rect 293866 -1542 294102 -1306
rect 293546 -1862 293782 -1626
rect 293866 -1862 294102 -1626
rect 297266 46658 297502 46894
rect 297586 46658 297822 46894
rect 297266 46338 297502 46574
rect 297586 46338 297822 46574
rect 297266 10658 297502 10894
rect 297586 10658 297822 10894
rect 297266 10338 297502 10574
rect 297586 10338 297822 10574
rect 297266 -2502 297502 -2266
rect 297586 -2502 297822 -2266
rect 297266 -2822 297502 -2586
rect 297586 -2822 297822 -2586
rect 300986 14378 301222 14614
rect 301306 14378 301542 14614
rect 300986 14058 301222 14294
rect 301306 14058 301542 14294
rect 300986 -3462 301222 -3226
rect 301306 -3462 301542 -3226
rect 300986 -3782 301222 -3546
rect 301306 -3782 301542 -3546
rect 304706 18098 304942 18334
rect 305026 18098 305262 18334
rect 304706 17778 304942 18014
rect 305026 17778 305262 18014
rect 304706 -4422 304942 -4186
rect 305026 -4422 305262 -4186
rect 304706 -4742 304942 -4506
rect 305026 -4742 305262 -4506
rect 308426 21818 308662 22054
rect 308746 21818 308982 22054
rect 308426 21498 308662 21734
rect 308746 21498 308982 21734
rect 308426 -5382 308662 -5146
rect 308746 -5382 308982 -5146
rect 308426 -5702 308662 -5466
rect 308746 -5702 308982 -5466
rect 312146 25538 312382 25774
rect 312466 25538 312702 25774
rect 312146 25218 312382 25454
rect 312466 25218 312702 25454
rect 312146 -6342 312382 -6106
rect 312466 -6342 312702 -6106
rect 312146 -6662 312382 -6426
rect 312466 -6662 312702 -6426
rect 315866 29258 316102 29494
rect 316186 29258 316422 29494
rect 315866 28938 316102 29174
rect 316186 28938 316422 29174
rect 315866 -7302 316102 -7066
rect 316186 -7302 316422 -7066
rect 315866 -7622 316102 -7386
rect 316186 -7622 316422 -7386
rect 325826 39218 326062 39454
rect 326146 39218 326382 39454
rect 325826 38898 326062 39134
rect 326146 38898 326382 39134
rect 325826 3218 326062 3454
rect 326146 3218 326382 3454
rect 325826 2898 326062 3134
rect 326146 2898 326382 3134
rect 325826 -582 326062 -346
rect 326146 -582 326382 -346
rect 325826 -902 326062 -666
rect 326146 -902 326382 -666
rect 329546 42938 329782 43174
rect 329866 42938 330102 43174
rect 329546 42618 329782 42854
rect 329866 42618 330102 42854
rect 329546 6938 329782 7174
rect 329866 6938 330102 7174
rect 329546 6618 329782 6854
rect 329866 6618 330102 6854
rect 329546 -1542 329782 -1306
rect 329866 -1542 330102 -1306
rect 329546 -1862 329782 -1626
rect 329866 -1862 330102 -1626
rect 333266 46658 333502 46894
rect 333586 46658 333822 46894
rect 333266 46338 333502 46574
rect 333586 46338 333822 46574
rect 333266 10658 333502 10894
rect 333586 10658 333822 10894
rect 333266 10338 333502 10574
rect 333586 10338 333822 10574
rect 333266 -2502 333502 -2266
rect 333586 -2502 333822 -2266
rect 333266 -2822 333502 -2586
rect 333586 -2822 333822 -2586
rect 336986 14378 337222 14614
rect 337306 14378 337542 14614
rect 336986 14058 337222 14294
rect 337306 14058 337542 14294
rect 336986 -3462 337222 -3226
rect 337306 -3462 337542 -3226
rect 336986 -3782 337222 -3546
rect 337306 -3782 337542 -3546
rect 340706 18098 340942 18334
rect 341026 18098 341262 18334
rect 340706 17778 340942 18014
rect 341026 17778 341262 18014
rect 340706 -4422 340942 -4186
rect 341026 -4422 341262 -4186
rect 340706 -4742 340942 -4506
rect 341026 -4742 341262 -4506
rect 344426 21818 344662 22054
rect 344746 21818 344982 22054
rect 344426 21498 344662 21734
rect 344746 21498 344982 21734
rect 344426 -5382 344662 -5146
rect 344746 -5382 344982 -5146
rect 344426 -5702 344662 -5466
rect 344746 -5702 344982 -5466
rect 348146 25538 348382 25774
rect 348466 25538 348702 25774
rect 348146 25218 348382 25454
rect 348466 25218 348702 25454
rect 348146 -6342 348382 -6106
rect 348466 -6342 348702 -6106
rect 348146 -6662 348382 -6426
rect 348466 -6662 348702 -6426
rect 351866 29258 352102 29494
rect 352186 29258 352422 29494
rect 351866 28938 352102 29174
rect 352186 28938 352422 29174
rect 351866 -7302 352102 -7066
rect 352186 -7302 352422 -7066
rect 351866 -7622 352102 -7386
rect 352186 -7622 352422 -7386
rect 361826 39218 362062 39454
rect 362146 39218 362382 39454
rect 361826 38898 362062 39134
rect 362146 38898 362382 39134
rect 361826 3218 362062 3454
rect 362146 3218 362382 3454
rect 361826 2898 362062 3134
rect 362146 2898 362382 3134
rect 361826 -582 362062 -346
rect 362146 -582 362382 -346
rect 361826 -902 362062 -666
rect 362146 -902 362382 -666
rect 365546 705562 365782 705798
rect 365866 705562 366102 705798
rect 365546 705242 365782 705478
rect 365866 705242 366102 705478
rect 365546 690938 365782 691174
rect 365866 690938 366102 691174
rect 365546 690618 365782 690854
rect 365866 690618 366102 690854
rect 365546 654938 365782 655174
rect 365866 654938 366102 655174
rect 365546 654618 365782 654854
rect 365866 654618 366102 654854
rect 365546 618938 365782 619174
rect 365866 618938 366102 619174
rect 365546 618618 365782 618854
rect 365866 618618 366102 618854
rect 365546 582938 365782 583174
rect 365866 582938 366102 583174
rect 365546 582618 365782 582854
rect 365866 582618 366102 582854
rect 365546 546938 365782 547174
rect 365866 546938 366102 547174
rect 365546 546618 365782 546854
rect 365866 546618 366102 546854
rect 365546 510938 365782 511174
rect 365866 510938 366102 511174
rect 365546 510618 365782 510854
rect 365866 510618 366102 510854
rect 365546 474938 365782 475174
rect 365866 474938 366102 475174
rect 365546 474618 365782 474854
rect 365866 474618 366102 474854
rect 365546 438938 365782 439174
rect 365866 438938 366102 439174
rect 365546 438618 365782 438854
rect 365866 438618 366102 438854
rect 365546 402938 365782 403174
rect 365866 402938 366102 403174
rect 365546 402618 365782 402854
rect 365866 402618 366102 402854
rect 365546 366938 365782 367174
rect 365866 366938 366102 367174
rect 365546 366618 365782 366854
rect 365866 366618 366102 366854
rect 365546 330938 365782 331174
rect 365866 330938 366102 331174
rect 365546 330618 365782 330854
rect 365866 330618 366102 330854
rect 365546 294938 365782 295174
rect 365866 294938 366102 295174
rect 365546 294618 365782 294854
rect 365866 294618 366102 294854
rect 365546 258938 365782 259174
rect 365866 258938 366102 259174
rect 365546 258618 365782 258854
rect 365866 258618 366102 258854
rect 365546 222938 365782 223174
rect 365866 222938 366102 223174
rect 365546 222618 365782 222854
rect 365866 222618 366102 222854
rect 365546 186938 365782 187174
rect 365866 186938 366102 187174
rect 365546 186618 365782 186854
rect 365866 186618 366102 186854
rect 365546 150938 365782 151174
rect 365866 150938 366102 151174
rect 365546 150618 365782 150854
rect 365866 150618 366102 150854
rect 365546 114938 365782 115174
rect 365866 114938 366102 115174
rect 365546 114618 365782 114854
rect 365866 114618 366102 114854
rect 365546 78938 365782 79174
rect 365866 78938 366102 79174
rect 365546 78618 365782 78854
rect 365866 78618 366102 78854
rect 365546 42938 365782 43174
rect 365866 42938 366102 43174
rect 365546 42618 365782 42854
rect 365866 42618 366102 42854
rect 365546 6938 365782 7174
rect 365866 6938 366102 7174
rect 365546 6618 365782 6854
rect 365866 6618 366102 6854
rect 365546 -1542 365782 -1306
rect 365866 -1542 366102 -1306
rect 365546 -1862 365782 -1626
rect 365866 -1862 366102 -1626
rect 369266 706522 369502 706758
rect 369586 706522 369822 706758
rect 369266 706202 369502 706438
rect 369586 706202 369822 706438
rect 369266 694658 369502 694894
rect 369586 694658 369822 694894
rect 369266 694338 369502 694574
rect 369586 694338 369822 694574
rect 369266 658658 369502 658894
rect 369586 658658 369822 658894
rect 369266 658338 369502 658574
rect 369586 658338 369822 658574
rect 369266 622658 369502 622894
rect 369586 622658 369822 622894
rect 369266 622338 369502 622574
rect 369586 622338 369822 622574
rect 369266 586658 369502 586894
rect 369586 586658 369822 586894
rect 369266 586338 369502 586574
rect 369586 586338 369822 586574
rect 369266 550658 369502 550894
rect 369586 550658 369822 550894
rect 369266 550338 369502 550574
rect 369586 550338 369822 550574
rect 369266 514658 369502 514894
rect 369586 514658 369822 514894
rect 369266 514338 369502 514574
rect 369586 514338 369822 514574
rect 369266 478658 369502 478894
rect 369586 478658 369822 478894
rect 369266 478338 369502 478574
rect 369586 478338 369822 478574
rect 369266 442658 369502 442894
rect 369586 442658 369822 442894
rect 369266 442338 369502 442574
rect 369586 442338 369822 442574
rect 369266 406658 369502 406894
rect 369586 406658 369822 406894
rect 369266 406338 369502 406574
rect 369586 406338 369822 406574
rect 369266 370658 369502 370894
rect 369586 370658 369822 370894
rect 369266 370338 369502 370574
rect 369586 370338 369822 370574
rect 369266 334658 369502 334894
rect 369586 334658 369822 334894
rect 369266 334338 369502 334574
rect 369586 334338 369822 334574
rect 369266 298658 369502 298894
rect 369586 298658 369822 298894
rect 369266 298338 369502 298574
rect 369586 298338 369822 298574
rect 369266 262658 369502 262894
rect 369586 262658 369822 262894
rect 369266 262338 369502 262574
rect 369586 262338 369822 262574
rect 369266 226658 369502 226894
rect 369586 226658 369822 226894
rect 369266 226338 369502 226574
rect 369586 226338 369822 226574
rect 369266 190658 369502 190894
rect 369586 190658 369822 190894
rect 369266 190338 369502 190574
rect 369586 190338 369822 190574
rect 369266 154658 369502 154894
rect 369586 154658 369822 154894
rect 369266 154338 369502 154574
rect 369586 154338 369822 154574
rect 369266 118658 369502 118894
rect 369586 118658 369822 118894
rect 369266 118338 369502 118574
rect 369586 118338 369822 118574
rect 369266 82658 369502 82894
rect 369586 82658 369822 82894
rect 369266 82338 369502 82574
rect 369586 82338 369822 82574
rect 369266 46658 369502 46894
rect 369586 46658 369822 46894
rect 369266 46338 369502 46574
rect 369586 46338 369822 46574
rect 369266 10658 369502 10894
rect 369586 10658 369822 10894
rect 369266 10338 369502 10574
rect 369586 10338 369822 10574
rect 369266 -2502 369502 -2266
rect 369586 -2502 369822 -2266
rect 369266 -2822 369502 -2586
rect 369586 -2822 369822 -2586
rect 372986 707482 373222 707718
rect 373306 707482 373542 707718
rect 372986 707162 373222 707398
rect 373306 707162 373542 707398
rect 372986 698378 373222 698614
rect 373306 698378 373542 698614
rect 372986 698058 373222 698294
rect 373306 698058 373542 698294
rect 372986 662378 373222 662614
rect 373306 662378 373542 662614
rect 372986 662058 373222 662294
rect 373306 662058 373542 662294
rect 372986 626378 373222 626614
rect 373306 626378 373542 626614
rect 372986 626058 373222 626294
rect 373306 626058 373542 626294
rect 372986 590378 373222 590614
rect 373306 590378 373542 590614
rect 372986 590058 373222 590294
rect 373306 590058 373542 590294
rect 372986 554378 373222 554614
rect 373306 554378 373542 554614
rect 372986 554058 373222 554294
rect 373306 554058 373542 554294
rect 372986 518378 373222 518614
rect 373306 518378 373542 518614
rect 372986 518058 373222 518294
rect 373306 518058 373542 518294
rect 372986 482378 373222 482614
rect 373306 482378 373542 482614
rect 372986 482058 373222 482294
rect 373306 482058 373542 482294
rect 372986 446378 373222 446614
rect 373306 446378 373542 446614
rect 372986 446058 373222 446294
rect 373306 446058 373542 446294
rect 372986 410378 373222 410614
rect 373306 410378 373542 410614
rect 372986 410058 373222 410294
rect 373306 410058 373542 410294
rect 372986 374378 373222 374614
rect 373306 374378 373542 374614
rect 372986 374058 373222 374294
rect 373306 374058 373542 374294
rect 372986 338378 373222 338614
rect 373306 338378 373542 338614
rect 372986 338058 373222 338294
rect 373306 338058 373542 338294
rect 372986 302378 373222 302614
rect 373306 302378 373542 302614
rect 372986 302058 373222 302294
rect 373306 302058 373542 302294
rect 372986 266378 373222 266614
rect 373306 266378 373542 266614
rect 372986 266058 373222 266294
rect 373306 266058 373542 266294
rect 372986 230378 373222 230614
rect 373306 230378 373542 230614
rect 372986 230058 373222 230294
rect 373306 230058 373542 230294
rect 372986 194378 373222 194614
rect 373306 194378 373542 194614
rect 372986 194058 373222 194294
rect 373306 194058 373542 194294
rect 372986 158378 373222 158614
rect 373306 158378 373542 158614
rect 372986 158058 373222 158294
rect 373306 158058 373542 158294
rect 372986 122378 373222 122614
rect 373306 122378 373542 122614
rect 372986 122058 373222 122294
rect 373306 122058 373542 122294
rect 372986 86378 373222 86614
rect 373306 86378 373542 86614
rect 372986 86058 373222 86294
rect 373306 86058 373542 86294
rect 372986 50378 373222 50614
rect 373306 50378 373542 50614
rect 372986 50058 373222 50294
rect 373306 50058 373542 50294
rect 372986 14378 373222 14614
rect 373306 14378 373542 14614
rect 372986 14058 373222 14294
rect 373306 14058 373542 14294
rect 372986 -3462 373222 -3226
rect 373306 -3462 373542 -3226
rect 372986 -3782 373222 -3546
rect 373306 -3782 373542 -3546
rect 376706 708442 376942 708678
rect 377026 708442 377262 708678
rect 376706 708122 376942 708358
rect 377026 708122 377262 708358
rect 376706 666098 376942 666334
rect 377026 666098 377262 666334
rect 376706 665778 376942 666014
rect 377026 665778 377262 666014
rect 376706 630098 376942 630334
rect 377026 630098 377262 630334
rect 376706 629778 376942 630014
rect 377026 629778 377262 630014
rect 376706 594098 376942 594334
rect 377026 594098 377262 594334
rect 376706 593778 376942 594014
rect 377026 593778 377262 594014
rect 376706 558098 376942 558334
rect 377026 558098 377262 558334
rect 376706 557778 376942 558014
rect 377026 557778 377262 558014
rect 376706 522098 376942 522334
rect 377026 522098 377262 522334
rect 376706 521778 376942 522014
rect 377026 521778 377262 522014
rect 376706 486098 376942 486334
rect 377026 486098 377262 486334
rect 376706 485778 376942 486014
rect 377026 485778 377262 486014
rect 376706 450098 376942 450334
rect 377026 450098 377262 450334
rect 376706 449778 376942 450014
rect 377026 449778 377262 450014
rect 376706 414098 376942 414334
rect 377026 414098 377262 414334
rect 376706 413778 376942 414014
rect 377026 413778 377262 414014
rect 376706 378098 376942 378334
rect 377026 378098 377262 378334
rect 376706 377778 376942 378014
rect 377026 377778 377262 378014
rect 376706 342098 376942 342334
rect 377026 342098 377262 342334
rect 376706 341778 376942 342014
rect 377026 341778 377262 342014
rect 376706 306098 376942 306334
rect 377026 306098 377262 306334
rect 376706 305778 376942 306014
rect 377026 305778 377262 306014
rect 376706 270098 376942 270334
rect 377026 270098 377262 270334
rect 376706 269778 376942 270014
rect 377026 269778 377262 270014
rect 376706 234098 376942 234334
rect 377026 234098 377262 234334
rect 376706 233778 376942 234014
rect 377026 233778 377262 234014
rect 376706 198098 376942 198334
rect 377026 198098 377262 198334
rect 376706 197778 376942 198014
rect 377026 197778 377262 198014
rect 376706 162098 376942 162334
rect 377026 162098 377262 162334
rect 376706 161778 376942 162014
rect 377026 161778 377262 162014
rect 376706 126098 376942 126334
rect 377026 126098 377262 126334
rect 376706 125778 376942 126014
rect 377026 125778 377262 126014
rect 376706 90098 376942 90334
rect 377026 90098 377262 90334
rect 376706 89778 376942 90014
rect 377026 89778 377262 90014
rect 376706 54098 376942 54334
rect 377026 54098 377262 54334
rect 376706 53778 376942 54014
rect 377026 53778 377262 54014
rect 376706 18098 376942 18334
rect 377026 18098 377262 18334
rect 376706 17778 376942 18014
rect 377026 17778 377262 18014
rect 376706 -4422 376942 -4186
rect 377026 -4422 377262 -4186
rect 376706 -4742 376942 -4506
rect 377026 -4742 377262 -4506
rect 380426 709402 380662 709638
rect 380746 709402 380982 709638
rect 380426 709082 380662 709318
rect 380746 709082 380982 709318
rect 380426 669818 380662 670054
rect 380746 669818 380982 670054
rect 380426 669498 380662 669734
rect 380746 669498 380982 669734
rect 380426 633818 380662 634054
rect 380746 633818 380982 634054
rect 380426 633498 380662 633734
rect 380746 633498 380982 633734
rect 380426 597818 380662 598054
rect 380746 597818 380982 598054
rect 380426 597498 380662 597734
rect 380746 597498 380982 597734
rect 380426 561818 380662 562054
rect 380746 561818 380982 562054
rect 380426 561498 380662 561734
rect 380746 561498 380982 561734
rect 380426 525818 380662 526054
rect 380746 525818 380982 526054
rect 380426 525498 380662 525734
rect 380746 525498 380982 525734
rect 380426 489818 380662 490054
rect 380746 489818 380982 490054
rect 380426 489498 380662 489734
rect 380746 489498 380982 489734
rect 380426 453818 380662 454054
rect 380746 453818 380982 454054
rect 380426 453498 380662 453734
rect 380746 453498 380982 453734
rect 380426 417818 380662 418054
rect 380746 417818 380982 418054
rect 380426 417498 380662 417734
rect 380746 417498 380982 417734
rect 380426 381818 380662 382054
rect 380746 381818 380982 382054
rect 380426 381498 380662 381734
rect 380746 381498 380982 381734
rect 380426 345818 380662 346054
rect 380746 345818 380982 346054
rect 380426 345498 380662 345734
rect 380746 345498 380982 345734
rect 380426 309818 380662 310054
rect 380746 309818 380982 310054
rect 380426 309498 380662 309734
rect 380746 309498 380982 309734
rect 380426 273818 380662 274054
rect 380746 273818 380982 274054
rect 380426 273498 380662 273734
rect 380746 273498 380982 273734
rect 380426 237818 380662 238054
rect 380746 237818 380982 238054
rect 380426 237498 380662 237734
rect 380746 237498 380982 237734
rect 380426 201818 380662 202054
rect 380746 201818 380982 202054
rect 380426 201498 380662 201734
rect 380746 201498 380982 201734
rect 380426 165818 380662 166054
rect 380746 165818 380982 166054
rect 380426 165498 380662 165734
rect 380746 165498 380982 165734
rect 380426 129818 380662 130054
rect 380746 129818 380982 130054
rect 380426 129498 380662 129734
rect 380746 129498 380982 129734
rect 380426 93818 380662 94054
rect 380746 93818 380982 94054
rect 380426 93498 380662 93734
rect 380746 93498 380982 93734
rect 380426 57818 380662 58054
rect 380746 57818 380982 58054
rect 380426 57498 380662 57734
rect 380746 57498 380982 57734
rect 380426 21818 380662 22054
rect 380746 21818 380982 22054
rect 380426 21498 380662 21734
rect 380746 21498 380982 21734
rect 380426 -5382 380662 -5146
rect 380746 -5382 380982 -5146
rect 380426 -5702 380662 -5466
rect 380746 -5702 380982 -5466
rect 384146 710362 384382 710598
rect 384466 710362 384702 710598
rect 384146 710042 384382 710278
rect 384466 710042 384702 710278
rect 384146 673538 384382 673774
rect 384466 673538 384702 673774
rect 384146 673218 384382 673454
rect 384466 673218 384702 673454
rect 384146 637538 384382 637774
rect 384466 637538 384702 637774
rect 384146 637218 384382 637454
rect 384466 637218 384702 637454
rect 384146 601538 384382 601774
rect 384466 601538 384702 601774
rect 384146 601218 384382 601454
rect 384466 601218 384702 601454
rect 384146 565538 384382 565774
rect 384466 565538 384702 565774
rect 384146 565218 384382 565454
rect 384466 565218 384702 565454
rect 384146 529538 384382 529774
rect 384466 529538 384702 529774
rect 384146 529218 384382 529454
rect 384466 529218 384702 529454
rect 384146 493538 384382 493774
rect 384466 493538 384702 493774
rect 384146 493218 384382 493454
rect 384466 493218 384702 493454
rect 384146 457538 384382 457774
rect 384466 457538 384702 457774
rect 384146 457218 384382 457454
rect 384466 457218 384702 457454
rect 384146 421538 384382 421774
rect 384466 421538 384702 421774
rect 384146 421218 384382 421454
rect 384466 421218 384702 421454
rect 384146 385538 384382 385774
rect 384466 385538 384702 385774
rect 384146 385218 384382 385454
rect 384466 385218 384702 385454
rect 384146 349538 384382 349774
rect 384466 349538 384702 349774
rect 384146 349218 384382 349454
rect 384466 349218 384702 349454
rect 384146 313538 384382 313774
rect 384466 313538 384702 313774
rect 384146 313218 384382 313454
rect 384466 313218 384702 313454
rect 384146 277538 384382 277774
rect 384466 277538 384702 277774
rect 384146 277218 384382 277454
rect 384466 277218 384702 277454
rect 384146 241538 384382 241774
rect 384466 241538 384702 241774
rect 384146 241218 384382 241454
rect 384466 241218 384702 241454
rect 384146 205538 384382 205774
rect 384466 205538 384702 205774
rect 384146 205218 384382 205454
rect 384466 205218 384702 205454
rect 384146 169538 384382 169774
rect 384466 169538 384702 169774
rect 384146 169218 384382 169454
rect 384466 169218 384702 169454
rect 384146 133538 384382 133774
rect 384466 133538 384702 133774
rect 384146 133218 384382 133454
rect 384466 133218 384702 133454
rect 384146 97538 384382 97774
rect 384466 97538 384702 97774
rect 384146 97218 384382 97454
rect 384466 97218 384702 97454
rect 387866 711322 388102 711558
rect 388186 711322 388422 711558
rect 387866 711002 388102 711238
rect 388186 711002 388422 711238
rect 387866 677258 388102 677494
rect 388186 677258 388422 677494
rect 387866 676938 388102 677174
rect 388186 676938 388422 677174
rect 387866 641258 388102 641494
rect 388186 641258 388422 641494
rect 387866 640938 388102 641174
rect 388186 640938 388422 641174
rect 387866 605258 388102 605494
rect 388186 605258 388422 605494
rect 387866 604938 388102 605174
rect 388186 604938 388422 605174
rect 387866 569258 388102 569494
rect 388186 569258 388422 569494
rect 387866 568938 388102 569174
rect 388186 568938 388422 569174
rect 387866 533258 388102 533494
rect 388186 533258 388422 533494
rect 387866 532938 388102 533174
rect 388186 532938 388422 533174
rect 387866 497258 388102 497494
rect 388186 497258 388422 497494
rect 387866 496938 388102 497174
rect 388186 496938 388422 497174
rect 387866 461258 388102 461494
rect 388186 461258 388422 461494
rect 387866 460938 388102 461174
rect 388186 460938 388422 461174
rect 387866 425258 388102 425494
rect 388186 425258 388422 425494
rect 387866 424938 388102 425174
rect 388186 424938 388422 425174
rect 387866 389258 388102 389494
rect 388186 389258 388422 389494
rect 387866 388938 388102 389174
rect 388186 388938 388422 389174
rect 387866 353258 388102 353494
rect 388186 353258 388422 353494
rect 387866 352938 388102 353174
rect 388186 352938 388422 353174
rect 387866 317258 388102 317494
rect 388186 317258 388422 317494
rect 387866 316938 388102 317174
rect 388186 316938 388422 317174
rect 387866 281258 388102 281494
rect 388186 281258 388422 281494
rect 387866 280938 388102 281174
rect 388186 280938 388422 281174
rect 387866 245258 388102 245494
rect 388186 245258 388422 245494
rect 387866 244938 388102 245174
rect 388186 244938 388422 245174
rect 387866 209258 388102 209494
rect 388186 209258 388422 209494
rect 387866 208938 388102 209174
rect 388186 208938 388422 209174
rect 387866 173258 388102 173494
rect 388186 173258 388422 173494
rect 387866 172938 388102 173174
rect 388186 172938 388422 173174
rect 387866 137258 388102 137494
rect 388186 137258 388422 137494
rect 387866 136938 388102 137174
rect 388186 136938 388422 137174
rect 387866 101258 388102 101494
rect 388186 101258 388422 101494
rect 387866 100938 388102 101174
rect 388186 100938 388422 101174
rect 397826 704602 398062 704838
rect 398146 704602 398382 704838
rect 397826 704282 398062 704518
rect 398146 704282 398382 704518
rect 397826 687218 398062 687454
rect 398146 687218 398382 687454
rect 397826 686898 398062 687134
rect 398146 686898 398382 687134
rect 397826 651218 398062 651454
rect 398146 651218 398382 651454
rect 397826 650898 398062 651134
rect 398146 650898 398382 651134
rect 397826 615218 398062 615454
rect 398146 615218 398382 615454
rect 397826 614898 398062 615134
rect 398146 614898 398382 615134
rect 397826 579218 398062 579454
rect 398146 579218 398382 579454
rect 397826 578898 398062 579134
rect 398146 578898 398382 579134
rect 397826 543218 398062 543454
rect 398146 543218 398382 543454
rect 397826 542898 398062 543134
rect 398146 542898 398382 543134
rect 397826 507218 398062 507454
rect 398146 507218 398382 507454
rect 397826 506898 398062 507134
rect 398146 506898 398382 507134
rect 397826 471218 398062 471454
rect 398146 471218 398382 471454
rect 397826 470898 398062 471134
rect 398146 470898 398382 471134
rect 397826 435218 398062 435454
rect 398146 435218 398382 435454
rect 397826 434898 398062 435134
rect 398146 434898 398382 435134
rect 397826 399218 398062 399454
rect 398146 399218 398382 399454
rect 397826 398898 398062 399134
rect 398146 398898 398382 399134
rect 397826 363218 398062 363454
rect 398146 363218 398382 363454
rect 397826 362898 398062 363134
rect 398146 362898 398382 363134
rect 397826 327218 398062 327454
rect 398146 327218 398382 327454
rect 397826 326898 398062 327134
rect 398146 326898 398382 327134
rect 397826 291218 398062 291454
rect 398146 291218 398382 291454
rect 397826 290898 398062 291134
rect 398146 290898 398382 291134
rect 397826 255218 398062 255454
rect 398146 255218 398382 255454
rect 397826 254898 398062 255134
rect 398146 254898 398382 255134
rect 397826 219218 398062 219454
rect 398146 219218 398382 219454
rect 397826 218898 398062 219134
rect 398146 218898 398382 219134
rect 397826 183218 398062 183454
rect 398146 183218 398382 183454
rect 397826 182898 398062 183134
rect 398146 182898 398382 183134
rect 397826 147218 398062 147454
rect 398146 147218 398382 147454
rect 397826 146898 398062 147134
rect 398146 146898 398382 147134
rect 397826 111218 398062 111454
rect 398146 111218 398382 111454
rect 397826 110898 398062 111134
rect 398146 110898 398382 111134
rect 401546 705562 401782 705798
rect 401866 705562 402102 705798
rect 401546 705242 401782 705478
rect 401866 705242 402102 705478
rect 401546 690938 401782 691174
rect 401866 690938 402102 691174
rect 401546 690618 401782 690854
rect 401866 690618 402102 690854
rect 401546 654938 401782 655174
rect 401866 654938 402102 655174
rect 401546 654618 401782 654854
rect 401866 654618 402102 654854
rect 401546 618938 401782 619174
rect 401866 618938 402102 619174
rect 401546 618618 401782 618854
rect 401866 618618 402102 618854
rect 401546 582938 401782 583174
rect 401866 582938 402102 583174
rect 401546 582618 401782 582854
rect 401866 582618 402102 582854
rect 401546 546938 401782 547174
rect 401866 546938 402102 547174
rect 401546 546618 401782 546854
rect 401866 546618 402102 546854
rect 401546 510938 401782 511174
rect 401866 510938 402102 511174
rect 401546 510618 401782 510854
rect 401866 510618 402102 510854
rect 401546 474938 401782 475174
rect 401866 474938 402102 475174
rect 401546 474618 401782 474854
rect 401866 474618 402102 474854
rect 401546 438938 401782 439174
rect 401866 438938 402102 439174
rect 401546 438618 401782 438854
rect 401866 438618 402102 438854
rect 401546 402938 401782 403174
rect 401866 402938 402102 403174
rect 401546 402618 401782 402854
rect 401866 402618 402102 402854
rect 401546 366938 401782 367174
rect 401866 366938 402102 367174
rect 401546 366618 401782 366854
rect 401866 366618 402102 366854
rect 401546 330938 401782 331174
rect 401866 330938 402102 331174
rect 401546 330618 401782 330854
rect 401866 330618 402102 330854
rect 405266 706522 405502 706758
rect 405586 706522 405822 706758
rect 405266 706202 405502 706438
rect 405586 706202 405822 706438
rect 405266 694658 405502 694894
rect 405586 694658 405822 694894
rect 405266 694338 405502 694574
rect 405586 694338 405822 694574
rect 405266 658658 405502 658894
rect 405586 658658 405822 658894
rect 405266 658338 405502 658574
rect 405586 658338 405822 658574
rect 405266 622658 405502 622894
rect 405586 622658 405822 622894
rect 405266 622338 405502 622574
rect 405586 622338 405822 622574
rect 405266 586658 405502 586894
rect 405586 586658 405822 586894
rect 405266 586338 405502 586574
rect 405586 586338 405822 586574
rect 405266 550658 405502 550894
rect 405586 550658 405822 550894
rect 405266 550338 405502 550574
rect 405586 550338 405822 550574
rect 405266 514658 405502 514894
rect 405586 514658 405822 514894
rect 405266 514338 405502 514574
rect 405586 514338 405822 514574
rect 405266 478658 405502 478894
rect 405586 478658 405822 478894
rect 405266 478338 405502 478574
rect 405586 478338 405822 478574
rect 405266 442658 405502 442894
rect 405586 442658 405822 442894
rect 405266 442338 405502 442574
rect 405586 442338 405822 442574
rect 405266 406658 405502 406894
rect 405586 406658 405822 406894
rect 405266 406338 405502 406574
rect 405586 406338 405822 406574
rect 405266 370658 405502 370894
rect 405586 370658 405822 370894
rect 405266 370338 405502 370574
rect 405586 370338 405822 370574
rect 405266 334658 405502 334894
rect 405586 334658 405822 334894
rect 405266 334338 405502 334574
rect 405586 334338 405822 334574
rect 404459 327218 404695 327454
rect 404459 326898 404695 327134
rect 401546 294938 401782 295174
rect 401866 294938 402102 295174
rect 401546 294618 401782 294854
rect 401866 294618 402102 294854
rect 401546 258938 401782 259174
rect 401866 258938 402102 259174
rect 401546 258618 401782 258854
rect 401866 258618 402102 258854
rect 401546 222938 401782 223174
rect 401866 222938 402102 223174
rect 401546 222618 401782 222854
rect 401866 222618 402102 222854
rect 401546 186938 401782 187174
rect 401866 186938 402102 187174
rect 401546 186618 401782 186854
rect 401866 186618 402102 186854
rect 401546 150938 401782 151174
rect 401866 150938 402102 151174
rect 401546 150618 401782 150854
rect 401866 150618 402102 150854
rect 401546 114938 401782 115174
rect 401866 114938 402102 115174
rect 401546 114618 401782 114854
rect 401866 114618 402102 114854
rect 408986 707482 409222 707718
rect 409306 707482 409542 707718
rect 408986 707162 409222 707398
rect 409306 707162 409542 707398
rect 408986 698378 409222 698614
rect 409306 698378 409542 698614
rect 408986 698058 409222 698294
rect 409306 698058 409542 698294
rect 408986 662378 409222 662614
rect 409306 662378 409542 662614
rect 408986 662058 409222 662294
rect 409306 662058 409542 662294
rect 408986 626378 409222 626614
rect 409306 626378 409542 626614
rect 408986 626058 409222 626294
rect 409306 626058 409542 626294
rect 408986 590378 409222 590614
rect 409306 590378 409542 590614
rect 408986 590058 409222 590294
rect 409306 590058 409542 590294
rect 408986 554378 409222 554614
rect 409306 554378 409542 554614
rect 408986 554058 409222 554294
rect 409306 554058 409542 554294
rect 408986 518378 409222 518614
rect 409306 518378 409542 518614
rect 408986 518058 409222 518294
rect 409306 518058 409542 518294
rect 408986 482378 409222 482614
rect 409306 482378 409542 482614
rect 408986 482058 409222 482294
rect 409306 482058 409542 482294
rect 408986 446378 409222 446614
rect 409306 446378 409542 446614
rect 408986 446058 409222 446294
rect 409306 446058 409542 446294
rect 408986 410378 409222 410614
rect 409306 410378 409542 410614
rect 408986 410058 409222 410294
rect 409306 410058 409542 410294
rect 408986 374378 409222 374614
rect 409306 374378 409542 374614
rect 408986 374058 409222 374294
rect 409306 374058 409542 374294
rect 408986 338378 409222 338614
rect 409306 338378 409542 338614
rect 408986 338058 409222 338294
rect 409306 338058 409542 338294
rect 407932 330938 408168 331174
rect 407932 330618 408168 330854
rect 405266 298658 405502 298894
rect 405586 298658 405822 298894
rect 405266 298338 405502 298574
rect 405586 298338 405822 298574
rect 405266 262658 405502 262894
rect 405586 262658 405822 262894
rect 405266 262338 405502 262574
rect 405586 262338 405822 262574
rect 405266 226658 405502 226894
rect 405586 226658 405822 226894
rect 405266 226338 405502 226574
rect 405586 226338 405822 226574
rect 405266 190658 405502 190894
rect 405586 190658 405822 190894
rect 405266 190338 405502 190574
rect 405586 190338 405822 190574
rect 405266 154658 405502 154894
rect 405586 154658 405822 154894
rect 405266 154338 405502 154574
rect 405586 154338 405822 154574
rect 405266 118658 405502 118894
rect 405586 118658 405822 118894
rect 405266 118338 405502 118574
rect 405586 118338 405822 118574
rect 412706 708442 412942 708678
rect 413026 708442 413262 708678
rect 412706 708122 412942 708358
rect 413026 708122 413262 708358
rect 412706 666098 412942 666334
rect 413026 666098 413262 666334
rect 412706 665778 412942 666014
rect 413026 665778 413262 666014
rect 412706 630098 412942 630334
rect 413026 630098 413262 630334
rect 412706 629778 412942 630014
rect 413026 629778 413262 630014
rect 412706 594098 412942 594334
rect 413026 594098 413262 594334
rect 412706 593778 412942 594014
rect 413026 593778 413262 594014
rect 412706 558098 412942 558334
rect 413026 558098 413262 558334
rect 412706 557778 412942 558014
rect 413026 557778 413262 558014
rect 412706 522098 412942 522334
rect 413026 522098 413262 522334
rect 412706 521778 412942 522014
rect 413026 521778 413262 522014
rect 412706 486098 412942 486334
rect 413026 486098 413262 486334
rect 412706 485778 412942 486014
rect 413026 485778 413262 486014
rect 412706 450098 412942 450334
rect 413026 450098 413262 450334
rect 412706 449778 412942 450014
rect 413026 449778 413262 450014
rect 412706 414098 412942 414334
rect 413026 414098 413262 414334
rect 412706 413778 412942 414014
rect 413026 413778 413262 414014
rect 412706 378098 412942 378334
rect 413026 378098 413262 378334
rect 412706 377778 412942 378014
rect 413026 377778 413262 378014
rect 412706 342098 412942 342334
rect 413026 342098 413262 342334
rect 412706 341778 412942 342014
rect 413026 341778 413262 342014
rect 411405 327218 411641 327454
rect 411405 326898 411641 327134
rect 408986 302378 409222 302614
rect 409306 302378 409542 302614
rect 408986 302058 409222 302294
rect 409306 302058 409542 302294
rect 408986 266378 409222 266614
rect 409306 266378 409542 266614
rect 408986 266058 409222 266294
rect 409306 266058 409542 266294
rect 408986 230378 409222 230614
rect 409306 230378 409542 230614
rect 408986 230058 409222 230294
rect 409306 230058 409542 230294
rect 408986 194378 409222 194614
rect 409306 194378 409542 194614
rect 408986 194058 409222 194294
rect 409306 194058 409542 194294
rect 408986 158378 409222 158614
rect 409306 158378 409542 158614
rect 408986 158058 409222 158294
rect 409306 158058 409542 158294
rect 408986 122378 409222 122614
rect 409306 122378 409542 122614
rect 408986 122058 409222 122294
rect 409306 122058 409542 122294
rect 416426 709402 416662 709638
rect 416746 709402 416982 709638
rect 416426 709082 416662 709318
rect 416746 709082 416982 709318
rect 416426 669818 416662 670054
rect 416746 669818 416982 670054
rect 416426 669498 416662 669734
rect 416746 669498 416982 669734
rect 416426 633818 416662 634054
rect 416746 633818 416982 634054
rect 416426 633498 416662 633734
rect 416746 633498 416982 633734
rect 416426 597818 416662 598054
rect 416746 597818 416982 598054
rect 416426 597498 416662 597734
rect 416746 597498 416982 597734
rect 416426 561818 416662 562054
rect 416746 561818 416982 562054
rect 416426 561498 416662 561734
rect 416746 561498 416982 561734
rect 416426 525818 416662 526054
rect 416746 525818 416982 526054
rect 416426 525498 416662 525734
rect 416746 525498 416982 525734
rect 416426 489818 416662 490054
rect 416746 489818 416982 490054
rect 416426 489498 416662 489734
rect 416746 489498 416982 489734
rect 416426 453818 416662 454054
rect 416746 453818 416982 454054
rect 416426 453498 416662 453734
rect 416746 453498 416982 453734
rect 416426 417818 416662 418054
rect 416746 417818 416982 418054
rect 416426 417498 416662 417734
rect 416746 417498 416982 417734
rect 416426 381818 416662 382054
rect 416746 381818 416982 382054
rect 416426 381498 416662 381734
rect 416746 381498 416982 381734
rect 416426 345818 416662 346054
rect 416746 345818 416982 346054
rect 416426 345498 416662 345734
rect 416746 345498 416982 345734
rect 414878 330938 415114 331174
rect 414878 330618 415114 330854
rect 412706 306098 412942 306334
rect 413026 306098 413262 306334
rect 412706 305778 412942 306014
rect 413026 305778 413262 306014
rect 412706 270098 412942 270334
rect 413026 270098 413262 270334
rect 412706 269778 412942 270014
rect 413026 269778 413262 270014
rect 412706 234098 412942 234334
rect 413026 234098 413262 234334
rect 412706 233778 412942 234014
rect 413026 233778 413262 234014
rect 412706 198098 412942 198334
rect 413026 198098 413262 198334
rect 412706 197778 412942 198014
rect 413026 197778 413262 198014
rect 412706 162098 412942 162334
rect 413026 162098 413262 162334
rect 412706 161778 412942 162014
rect 413026 161778 413262 162014
rect 420146 710362 420382 710598
rect 420466 710362 420702 710598
rect 420146 710042 420382 710278
rect 420466 710042 420702 710278
rect 420146 673538 420382 673774
rect 420466 673538 420702 673774
rect 420146 673218 420382 673454
rect 420466 673218 420702 673454
rect 420146 637538 420382 637774
rect 420466 637538 420702 637774
rect 420146 637218 420382 637454
rect 420466 637218 420702 637454
rect 420146 601538 420382 601774
rect 420466 601538 420702 601774
rect 420146 601218 420382 601454
rect 420466 601218 420702 601454
rect 420146 565538 420382 565774
rect 420466 565538 420702 565774
rect 420146 565218 420382 565454
rect 420466 565218 420702 565454
rect 420146 529538 420382 529774
rect 420466 529538 420702 529774
rect 420146 529218 420382 529454
rect 420466 529218 420702 529454
rect 420146 493538 420382 493774
rect 420466 493538 420702 493774
rect 420146 493218 420382 493454
rect 420466 493218 420702 493454
rect 420146 457538 420382 457774
rect 420466 457538 420702 457774
rect 420146 457218 420382 457454
rect 420466 457218 420702 457454
rect 423866 711322 424102 711558
rect 424186 711322 424422 711558
rect 423866 711002 424102 711238
rect 424186 711002 424422 711238
rect 423866 677258 424102 677494
rect 424186 677258 424422 677494
rect 423866 676938 424102 677174
rect 424186 676938 424422 677174
rect 423866 641258 424102 641494
rect 424186 641258 424422 641494
rect 423866 640938 424102 641174
rect 424186 640938 424422 641174
rect 423866 605258 424102 605494
rect 424186 605258 424422 605494
rect 423866 604938 424102 605174
rect 424186 604938 424422 605174
rect 423866 569258 424102 569494
rect 424186 569258 424422 569494
rect 423866 568938 424102 569174
rect 424186 568938 424422 569174
rect 423866 533258 424102 533494
rect 424186 533258 424422 533494
rect 423866 532938 424102 533174
rect 424186 532938 424422 533174
rect 423866 497258 424102 497494
rect 424186 497258 424422 497494
rect 423866 496938 424102 497174
rect 424186 496938 424422 497174
rect 423866 461258 424102 461494
rect 424186 461258 424422 461494
rect 423866 460938 424102 461174
rect 424186 460938 424422 461174
rect 433826 704602 434062 704838
rect 434146 704602 434382 704838
rect 433826 704282 434062 704518
rect 434146 704282 434382 704518
rect 433826 687218 434062 687454
rect 434146 687218 434382 687454
rect 433826 686898 434062 687134
rect 434146 686898 434382 687134
rect 433826 651218 434062 651454
rect 434146 651218 434382 651454
rect 433826 650898 434062 651134
rect 434146 650898 434382 651134
rect 433826 615218 434062 615454
rect 434146 615218 434382 615454
rect 433826 614898 434062 615134
rect 434146 614898 434382 615134
rect 433826 579218 434062 579454
rect 434146 579218 434382 579454
rect 433826 578898 434062 579134
rect 434146 578898 434382 579134
rect 433826 543218 434062 543454
rect 434146 543218 434382 543454
rect 433826 542898 434062 543134
rect 434146 542898 434382 543134
rect 433826 507218 434062 507454
rect 434146 507218 434382 507454
rect 433826 506898 434062 507134
rect 434146 506898 434382 507134
rect 433826 471218 434062 471454
rect 434146 471218 434382 471454
rect 433826 470898 434062 471134
rect 434146 470898 434382 471134
rect 437546 705562 437782 705798
rect 437866 705562 438102 705798
rect 437546 705242 437782 705478
rect 437866 705242 438102 705478
rect 437546 690938 437782 691174
rect 437866 690938 438102 691174
rect 437546 690618 437782 690854
rect 437866 690618 438102 690854
rect 437546 654938 437782 655174
rect 437866 654938 438102 655174
rect 437546 654618 437782 654854
rect 437866 654618 438102 654854
rect 437546 618938 437782 619174
rect 437866 618938 438102 619174
rect 437546 618618 437782 618854
rect 437866 618618 438102 618854
rect 437546 582938 437782 583174
rect 437866 582938 438102 583174
rect 437546 582618 437782 582854
rect 437866 582618 438102 582854
rect 437546 546938 437782 547174
rect 437866 546938 438102 547174
rect 437546 546618 437782 546854
rect 437866 546618 438102 546854
rect 437546 510938 437782 511174
rect 437866 510938 438102 511174
rect 437546 510618 437782 510854
rect 437866 510618 438102 510854
rect 437546 474938 437782 475174
rect 437866 474938 438102 475174
rect 437546 474618 437782 474854
rect 437866 474618 438102 474854
rect 441266 706522 441502 706758
rect 441586 706522 441822 706758
rect 441266 706202 441502 706438
rect 441586 706202 441822 706438
rect 441266 694658 441502 694894
rect 441586 694658 441822 694894
rect 441266 694338 441502 694574
rect 441586 694338 441822 694574
rect 444986 707482 445222 707718
rect 445306 707482 445542 707718
rect 444986 707162 445222 707398
rect 445306 707162 445542 707398
rect 448706 708442 448942 708678
rect 449026 708442 449262 708678
rect 448706 708122 448942 708358
rect 449026 708122 449262 708358
rect 444986 698378 445222 698614
rect 445306 698378 445542 698614
rect 444986 698058 445222 698294
rect 445306 698058 445542 698294
rect 441266 658658 441502 658894
rect 441586 658658 441822 658894
rect 441266 658338 441502 658574
rect 441586 658338 441822 658574
rect 441266 622658 441502 622894
rect 441586 622658 441822 622894
rect 441266 622338 441502 622574
rect 441586 622338 441822 622574
rect 441266 586658 441502 586894
rect 441586 586658 441822 586894
rect 441266 586338 441502 586574
rect 441586 586338 441822 586574
rect 441266 550658 441502 550894
rect 441586 550658 441822 550894
rect 441266 550338 441502 550574
rect 441586 550338 441822 550574
rect 441266 514658 441502 514894
rect 441586 514658 441822 514894
rect 441266 514338 441502 514574
rect 441586 514338 441822 514574
rect 441266 478658 441502 478894
rect 441586 478658 441822 478894
rect 441266 478338 441502 478574
rect 441586 478338 441822 478574
rect 426666 438938 426902 439174
rect 426666 438618 426902 438854
rect 432347 438938 432583 439174
rect 432347 438618 432583 438854
rect 438028 438938 438264 439174
rect 438028 438618 438264 438854
rect 443709 438938 443945 439174
rect 443709 438618 443945 438854
rect 423826 435218 424062 435454
rect 423826 434898 424062 435134
rect 429507 435218 429743 435454
rect 429507 434898 429743 435134
rect 435188 435218 435424 435454
rect 435188 434898 435424 435134
rect 440869 435218 441105 435454
rect 440869 434898 441105 435134
rect 420146 421538 420382 421774
rect 420466 421538 420702 421774
rect 420146 421218 420382 421454
rect 420466 421218 420702 421454
rect 420146 385538 420382 385774
rect 420466 385538 420702 385774
rect 420146 385218 420382 385454
rect 420466 385218 420702 385454
rect 420146 349538 420382 349774
rect 420466 349538 420702 349774
rect 420146 349218 420382 349454
rect 420466 349218 420702 349454
rect 418351 327218 418587 327454
rect 418351 326898 418587 327134
rect 416426 309818 416662 310054
rect 416746 309818 416982 310054
rect 416426 309498 416662 309734
rect 416746 309498 416982 309734
rect 416426 273818 416662 274054
rect 416746 273818 416982 274054
rect 416426 273498 416662 273734
rect 416746 273498 416982 273734
rect 416426 237818 416662 238054
rect 416746 237818 416982 238054
rect 416426 237498 416662 237734
rect 416746 237498 416982 237734
rect 416426 201818 416662 202054
rect 416746 201818 416982 202054
rect 416426 201498 416662 201734
rect 416746 201498 416982 201734
rect 416426 165818 416662 166054
rect 416746 165818 416982 166054
rect 416426 165498 416662 165734
rect 416746 165498 416982 165734
rect 423866 389258 424102 389494
rect 424186 389258 424422 389494
rect 423866 388938 424102 389174
rect 424186 388938 424422 389174
rect 423866 353258 424102 353494
rect 424186 353258 424422 353494
rect 423866 352938 424102 353174
rect 424186 352938 424422 353174
rect 420146 313538 420382 313774
rect 420466 313538 420702 313774
rect 420146 313218 420382 313454
rect 420466 313218 420702 313454
rect 420146 277538 420382 277774
rect 420466 277538 420702 277774
rect 420146 277218 420382 277454
rect 420466 277218 420702 277454
rect 420146 241538 420382 241774
rect 420466 241538 420702 241774
rect 420146 241218 420382 241454
rect 420466 241218 420702 241454
rect 420146 205538 420382 205774
rect 420466 205538 420702 205774
rect 420146 205218 420382 205454
rect 420466 205218 420702 205454
rect 420146 169538 420382 169774
rect 420466 169538 420702 169774
rect 420146 169218 420382 169454
rect 420466 169218 420702 169454
rect 421824 330938 422060 331174
rect 421824 330618 422060 330854
rect 433826 399218 434062 399454
rect 434146 399218 434382 399454
rect 433826 398898 434062 399134
rect 434146 398898 434382 399134
rect 433826 363218 434062 363454
rect 434146 363218 434382 363454
rect 433826 362898 434062 363134
rect 434146 362898 434382 363134
rect 425297 327218 425533 327454
rect 425297 326898 425533 327134
rect 423866 317258 424102 317494
rect 424186 317258 424422 317494
rect 423866 316938 424102 317174
rect 424186 316938 424422 317174
rect 423866 281258 424102 281494
rect 424186 281258 424422 281494
rect 423866 280938 424102 281174
rect 424186 280938 424422 281174
rect 423866 245258 424102 245494
rect 424186 245258 424422 245494
rect 423866 244938 424102 245174
rect 424186 244938 424422 245174
rect 423866 209258 424102 209494
rect 424186 209258 424422 209494
rect 423866 208938 424102 209174
rect 424186 208938 424422 209174
rect 423866 173258 424102 173494
rect 424186 173258 424422 173494
rect 423866 172938 424102 173174
rect 424186 172938 424422 173174
rect 428770 330938 429006 331174
rect 428770 330618 429006 330854
rect 433826 327218 434062 327454
rect 434146 327218 434382 327454
rect 433826 326898 434062 327134
rect 434146 326898 434382 327134
rect 433826 291218 434062 291454
rect 434146 291218 434382 291454
rect 433826 290898 434062 291134
rect 434146 290898 434382 291134
rect 433826 255218 434062 255454
rect 434146 255218 434382 255454
rect 433826 254898 434062 255134
rect 434146 254898 434382 255134
rect 433826 219218 434062 219454
rect 434146 219218 434382 219454
rect 433826 218898 434062 219134
rect 434146 218898 434382 219134
rect 433826 183218 434062 183454
rect 434146 183218 434382 183454
rect 433826 182898 434062 183134
rect 434146 182898 434382 183134
rect 437546 402938 437782 403174
rect 437866 402938 438102 403174
rect 437546 402618 437782 402854
rect 437866 402618 438102 402854
rect 437546 366938 437782 367174
rect 437866 366938 438102 367174
rect 437546 366618 437782 366854
rect 437866 366618 438102 366854
rect 437546 330938 437782 331174
rect 437866 330938 438102 331174
rect 437546 330618 437782 330854
rect 437866 330618 438102 330854
rect 437546 294938 437782 295174
rect 437866 294938 438102 295174
rect 437546 294618 437782 294854
rect 437866 294618 438102 294854
rect 437546 258938 437782 259174
rect 437866 258938 438102 259174
rect 437546 258618 437782 258854
rect 437866 258618 438102 258854
rect 437546 222938 437782 223174
rect 437866 222938 438102 223174
rect 437546 222618 437782 222854
rect 437866 222618 438102 222854
rect 437546 186938 437782 187174
rect 437866 186938 438102 187174
rect 437546 186618 437782 186854
rect 437866 186618 438102 186854
rect 441266 406658 441502 406894
rect 441586 406658 441822 406894
rect 441266 406338 441502 406574
rect 441586 406338 441822 406574
rect 441266 370658 441502 370894
rect 441586 370658 441822 370894
rect 441266 370338 441502 370574
rect 441586 370338 441822 370574
rect 441266 334658 441502 334894
rect 441586 334658 441822 334894
rect 441266 334338 441502 334574
rect 441586 334338 441822 334574
rect 444986 662378 445222 662614
rect 445306 662378 445542 662614
rect 444986 662058 445222 662294
rect 445306 662058 445542 662294
rect 444986 626378 445222 626614
rect 445306 626378 445542 626614
rect 444986 626058 445222 626294
rect 445306 626058 445542 626294
rect 444986 590378 445222 590614
rect 445306 590378 445542 590614
rect 444986 590058 445222 590294
rect 445306 590058 445542 590294
rect 444986 554378 445222 554614
rect 445306 554378 445542 554614
rect 444986 554058 445222 554294
rect 445306 554058 445542 554294
rect 444986 518378 445222 518614
rect 445306 518378 445542 518614
rect 444986 518058 445222 518294
rect 445306 518058 445542 518294
rect 444986 482378 445222 482614
rect 445306 482378 445542 482614
rect 444986 482058 445222 482294
rect 445306 482058 445542 482294
rect 444986 446378 445222 446614
rect 445306 446378 445542 446614
rect 444986 446058 445222 446294
rect 445306 446058 445542 446294
rect 444986 410378 445222 410614
rect 445306 410378 445542 410614
rect 444986 410058 445222 410294
rect 445306 410058 445542 410294
rect 444986 374378 445222 374614
rect 445306 374378 445542 374614
rect 444986 374058 445222 374294
rect 445306 374058 445542 374294
rect 444986 338378 445222 338614
rect 445306 338378 445542 338614
rect 444986 338058 445222 338294
rect 445306 338058 445542 338294
rect 441266 298658 441502 298894
rect 441586 298658 441822 298894
rect 441266 298338 441502 298574
rect 441586 298338 441822 298574
rect 441266 262658 441502 262894
rect 441586 262658 441822 262894
rect 441266 262338 441502 262574
rect 441586 262338 441822 262574
rect 441266 226658 441502 226894
rect 441586 226658 441822 226894
rect 441266 226338 441502 226574
rect 441586 226338 441822 226574
rect 441266 190658 441502 190894
rect 441586 190658 441822 190894
rect 441266 190338 441502 190574
rect 441586 190338 441822 190574
rect 452426 709402 452662 709638
rect 452746 709402 452982 709638
rect 452426 709082 452662 709318
rect 452746 709082 452982 709318
rect 448706 666098 448942 666334
rect 449026 666098 449262 666334
rect 448706 665778 448942 666014
rect 449026 665778 449262 666014
rect 448706 630098 448942 630334
rect 449026 630098 449262 630334
rect 448706 629778 448942 630014
rect 449026 629778 449262 630014
rect 448706 594098 448942 594334
rect 449026 594098 449262 594334
rect 448706 593778 448942 594014
rect 449026 593778 449262 594014
rect 448706 558098 448942 558334
rect 449026 558098 449262 558334
rect 448706 557778 448942 558014
rect 449026 557778 449262 558014
rect 448706 522098 448942 522334
rect 449026 522098 449262 522334
rect 448706 521778 448942 522014
rect 449026 521778 449262 522014
rect 448706 486098 448942 486334
rect 449026 486098 449262 486334
rect 448706 485778 448942 486014
rect 449026 485778 449262 486014
rect 448706 450098 448942 450334
rect 449026 450098 449262 450334
rect 448706 449778 448942 450014
rect 449026 449778 449262 450014
rect 448706 414098 448942 414334
rect 449026 414098 449262 414334
rect 448706 413778 448942 414014
rect 449026 413778 449262 414014
rect 448706 378098 448942 378334
rect 449026 378098 449262 378334
rect 448706 377778 448942 378014
rect 449026 377778 449262 378014
rect 448706 342098 448942 342334
rect 449026 342098 449262 342334
rect 448706 341778 448942 342014
rect 449026 341778 449262 342014
rect 444986 302378 445222 302614
rect 445306 302378 445542 302614
rect 444986 302058 445222 302294
rect 445306 302058 445542 302294
rect 444986 266378 445222 266614
rect 445306 266378 445542 266614
rect 444986 266058 445222 266294
rect 445306 266058 445542 266294
rect 444986 230378 445222 230614
rect 445306 230378 445542 230614
rect 444986 230058 445222 230294
rect 445306 230058 445542 230294
rect 444986 194378 445222 194614
rect 445306 194378 445542 194614
rect 444986 194058 445222 194294
rect 445306 194058 445542 194294
rect 452426 669818 452662 670054
rect 452746 669818 452982 670054
rect 452426 669498 452662 669734
rect 452746 669498 452982 669734
rect 452426 633818 452662 634054
rect 452746 633818 452982 634054
rect 452426 633498 452662 633734
rect 452746 633498 452982 633734
rect 452426 597818 452662 598054
rect 452746 597818 452982 598054
rect 452426 597498 452662 597734
rect 452746 597498 452982 597734
rect 452426 561818 452662 562054
rect 452746 561818 452982 562054
rect 452426 561498 452662 561734
rect 452746 561498 452982 561734
rect 452426 525818 452662 526054
rect 452746 525818 452982 526054
rect 452426 525498 452662 525734
rect 452746 525498 452982 525734
rect 456146 710362 456382 710598
rect 456466 710362 456702 710598
rect 456146 710042 456382 710278
rect 456466 710042 456702 710278
rect 456146 673538 456382 673774
rect 456466 673538 456702 673774
rect 456146 673218 456382 673454
rect 456466 673218 456702 673454
rect 459866 711322 460102 711558
rect 460186 711322 460422 711558
rect 459866 711002 460102 711238
rect 460186 711002 460422 711238
rect 459866 677258 460102 677494
rect 460186 677258 460422 677494
rect 459866 676938 460102 677174
rect 460186 676938 460422 677174
rect 469826 704602 470062 704838
rect 470146 704602 470382 704838
rect 469826 704282 470062 704518
rect 470146 704282 470382 704518
rect 469826 687218 470062 687454
rect 470146 687218 470382 687454
rect 469826 686898 470062 687134
rect 470146 686898 470382 687134
rect 473546 705562 473782 705798
rect 473866 705562 474102 705798
rect 473546 705242 473782 705478
rect 473866 705242 474102 705478
rect 473546 690938 473782 691174
rect 473866 690938 474102 691174
rect 473546 690618 473782 690854
rect 473866 690618 474102 690854
rect 477266 706522 477502 706758
rect 477586 706522 477822 706758
rect 477266 706202 477502 706438
rect 477586 706202 477822 706438
rect 477266 694658 477502 694894
rect 477586 694658 477822 694894
rect 477266 694338 477502 694574
rect 477586 694338 477822 694574
rect 480986 707482 481222 707718
rect 481306 707482 481542 707718
rect 480986 707162 481222 707398
rect 481306 707162 481542 707398
rect 480986 698378 481222 698614
rect 481306 698378 481542 698614
rect 480986 698058 481222 698294
rect 481306 698058 481542 698294
rect 488426 709402 488662 709638
rect 488746 709402 488982 709638
rect 488426 709082 488662 709318
rect 488746 709082 488982 709318
rect 488426 669818 488662 670054
rect 488746 669818 488982 670054
rect 488426 669498 488662 669734
rect 488746 669498 488982 669734
rect 492146 710362 492382 710598
rect 492466 710362 492702 710598
rect 492146 710042 492382 710278
rect 492466 710042 492702 710278
rect 492146 673538 492382 673774
rect 492466 673538 492702 673774
rect 492146 673218 492382 673454
rect 492466 673218 492702 673454
rect 495866 711322 496102 711558
rect 496186 711322 496422 711558
rect 495866 711002 496102 711238
rect 496186 711002 496422 711238
rect 495866 677258 496102 677494
rect 496186 677258 496422 677494
rect 495866 676938 496102 677174
rect 496186 676938 496422 677174
rect 505826 704602 506062 704838
rect 506146 704602 506382 704838
rect 505826 704282 506062 704518
rect 506146 704282 506382 704518
rect 505826 687218 506062 687454
rect 506146 687218 506382 687454
rect 505826 686898 506062 687134
rect 506146 686898 506382 687134
rect 509546 705562 509782 705798
rect 509866 705562 510102 705798
rect 509546 705242 509782 705478
rect 509866 705242 510102 705478
rect 509546 690938 509782 691174
rect 509866 690938 510102 691174
rect 509546 690618 509782 690854
rect 509866 690618 510102 690854
rect 513266 706522 513502 706758
rect 513586 706522 513822 706758
rect 513266 706202 513502 706438
rect 513586 706202 513822 706438
rect 513266 694658 513502 694894
rect 513586 694658 513822 694894
rect 513266 694338 513502 694574
rect 513586 694338 513822 694574
rect 516986 707482 517222 707718
rect 517306 707482 517542 707718
rect 516986 707162 517222 707398
rect 517306 707162 517542 707398
rect 516986 698378 517222 698614
rect 517306 698378 517542 698614
rect 516986 698058 517222 698294
rect 517306 698058 517542 698294
rect 520706 708442 520942 708678
rect 521026 708442 521262 708678
rect 520706 708122 520942 708358
rect 521026 708122 521262 708358
rect 520706 666098 520942 666334
rect 521026 666098 521262 666334
rect 520706 665778 520942 666014
rect 521026 665778 521262 666014
rect 456146 637538 456382 637774
rect 456466 637538 456702 637774
rect 456146 637218 456382 637454
rect 456466 637218 456702 637454
rect 456146 601538 456382 601774
rect 456466 601538 456702 601774
rect 456146 601218 456382 601454
rect 456466 601218 456702 601454
rect 456146 565538 456382 565774
rect 456466 565538 456702 565774
rect 456146 565218 456382 565454
rect 456466 565218 456702 565454
rect 456146 529538 456382 529774
rect 456466 529538 456702 529774
rect 456146 529218 456382 529454
rect 456466 529218 456702 529454
rect 479610 654938 479846 655174
rect 479610 654618 479846 654854
rect 510330 654938 510566 655174
rect 510330 654618 510566 654854
rect 464250 651218 464486 651454
rect 464250 650898 464486 651134
rect 494970 651218 495206 651454
rect 494970 650898 495206 651134
rect 520706 630098 520942 630334
rect 521026 630098 521262 630334
rect 520706 629778 520942 630014
rect 521026 629778 521262 630014
rect 479610 618938 479846 619174
rect 479610 618618 479846 618854
rect 510330 618938 510566 619174
rect 510330 618618 510566 618854
rect 464250 615218 464486 615454
rect 464250 614898 464486 615134
rect 494970 615218 495206 615454
rect 494970 614898 495206 615134
rect 459866 569258 460102 569494
rect 460186 569258 460422 569494
rect 459866 568938 460102 569174
rect 460186 568938 460422 569174
rect 459866 533258 460102 533494
rect 460186 533258 460422 533494
rect 459866 532938 460102 533174
rect 460186 532938 460422 533174
rect 469826 579218 470062 579454
rect 470146 579218 470382 579454
rect 469826 578898 470062 579134
rect 470146 578898 470382 579134
rect 469826 543218 470062 543454
rect 470146 543218 470382 543454
rect 469826 542898 470062 543134
rect 470146 542898 470382 543134
rect 453424 510938 453660 511174
rect 453424 510618 453660 510854
rect 455862 510938 456098 511174
rect 455862 510618 456098 510854
rect 458300 510938 458536 511174
rect 458300 510618 458536 510854
rect 460738 510938 460974 511174
rect 460738 510618 460974 510854
rect 452205 507218 452441 507454
rect 452205 506898 452441 507134
rect 454643 507218 454879 507454
rect 454643 506898 454879 507134
rect 457081 507218 457317 507454
rect 457081 506898 457317 507134
rect 459519 507218 459755 507454
rect 459519 506898 459755 507134
rect 469826 507218 470062 507454
rect 470146 507218 470382 507454
rect 469826 506898 470062 507134
rect 470146 506898 470382 507134
rect 452426 489818 452662 490054
rect 452746 489818 452982 490054
rect 452426 489498 452662 489734
rect 452746 489498 452982 489734
rect 452426 453818 452662 454054
rect 452746 453818 452982 454054
rect 452426 453498 452662 453734
rect 452746 453498 452982 453734
rect 452426 417818 452662 418054
rect 452746 417818 452982 418054
rect 452426 417498 452662 417734
rect 452746 417498 452982 417734
rect 452426 381818 452662 382054
rect 452746 381818 452982 382054
rect 452426 381498 452662 381734
rect 452746 381498 452982 381734
rect 456146 493538 456382 493774
rect 456466 493538 456702 493774
rect 456146 493218 456382 493454
rect 456466 493218 456702 493454
rect 456146 457538 456382 457774
rect 456466 457538 456702 457774
rect 456146 457218 456382 457454
rect 456466 457218 456702 457454
rect 456146 421538 456382 421774
rect 456466 421538 456702 421774
rect 456146 421218 456382 421454
rect 456466 421218 456702 421454
rect 456146 385538 456382 385774
rect 456466 385538 456702 385774
rect 456146 385218 456382 385454
rect 456466 385218 456702 385454
rect 454250 363218 454486 363454
rect 454250 362898 454486 363134
rect 452426 345818 452662 346054
rect 452746 345818 452982 346054
rect 452426 345498 452662 345734
rect 452746 345498 452982 345734
rect 448706 306098 448942 306334
rect 449026 306098 449262 306334
rect 448706 305778 448942 306014
rect 449026 305778 449262 306014
rect 448706 270098 448942 270334
rect 449026 270098 449262 270334
rect 448706 269778 448942 270014
rect 449026 269778 449262 270014
rect 448706 234098 448942 234334
rect 449026 234098 449262 234334
rect 448706 233778 448942 234014
rect 449026 233778 449262 234014
rect 448706 198098 448942 198334
rect 449026 198098 449262 198334
rect 448706 197778 448942 198014
rect 449026 197778 449262 198014
rect 448706 162098 448942 162334
rect 449026 162098 449262 162334
rect 448706 161778 448942 162014
rect 449026 161778 449262 162014
rect 429610 150938 429846 151174
rect 429610 150618 429846 150854
rect 414250 147218 414486 147454
rect 414250 146898 414486 147134
rect 444970 147218 445206 147454
rect 444970 146898 445206 147134
rect 412706 126098 412942 126334
rect 413026 126098 413262 126334
rect 412706 125778 412942 126014
rect 413026 125778 413262 126014
rect 416426 93818 416662 94054
rect 416746 93818 416982 94054
rect 416426 93498 416662 93734
rect 416746 93498 416982 93734
rect 420146 97538 420382 97774
rect 420466 97538 420702 97774
rect 420146 97218 420382 97454
rect 420466 97218 420702 97454
rect 423866 101258 424102 101494
rect 424186 101258 424422 101494
rect 423866 100938 424102 101174
rect 424186 100938 424422 101174
rect 448706 126098 448942 126334
rect 449026 126098 449262 126334
rect 448706 125778 448942 126014
rect 449026 125778 449262 126014
rect 456146 349538 456382 349774
rect 456466 349538 456702 349774
rect 456146 349218 456382 349454
rect 456466 349218 456702 349454
rect 454250 327218 454486 327454
rect 454250 326898 454486 327134
rect 452426 309818 452662 310054
rect 452746 309818 452982 310054
rect 452426 309498 452662 309734
rect 452746 309498 452982 309734
rect 452426 273818 452662 274054
rect 452746 273818 452982 274054
rect 452426 273498 452662 273734
rect 452746 273498 452982 273734
rect 452426 237818 452662 238054
rect 452746 237818 452982 238054
rect 452426 237498 452662 237734
rect 452746 237498 452982 237734
rect 452426 201818 452662 202054
rect 452746 201818 452982 202054
rect 452426 201498 452662 201734
rect 452746 201498 452982 201734
rect 452426 165818 452662 166054
rect 452746 165818 452982 166054
rect 452426 165498 452662 165734
rect 452746 165498 452982 165734
rect 452426 129818 452662 130054
rect 452746 129818 452982 130054
rect 452426 129498 452662 129734
rect 452746 129498 452982 129734
rect 452426 93818 452662 94054
rect 452746 93818 452982 94054
rect 452426 93498 452662 93734
rect 452746 93498 452982 93734
rect 456146 313538 456382 313774
rect 456466 313538 456702 313774
rect 456146 313218 456382 313454
rect 456466 313218 456702 313454
rect 456146 277538 456382 277774
rect 456466 277538 456702 277774
rect 456146 277218 456382 277454
rect 456466 277218 456702 277454
rect 456146 241538 456382 241774
rect 456466 241538 456702 241774
rect 456146 241218 456382 241454
rect 456466 241218 456702 241454
rect 456146 205538 456382 205774
rect 456466 205538 456702 205774
rect 456146 205218 456382 205454
rect 456466 205218 456702 205454
rect 456146 169538 456382 169774
rect 456466 169538 456702 169774
rect 456146 169218 456382 169454
rect 456466 169218 456702 169454
rect 456146 133538 456382 133774
rect 456466 133538 456702 133774
rect 456146 133218 456382 133454
rect 456466 133218 456702 133454
rect 456146 97538 456382 97774
rect 456466 97538 456702 97774
rect 456146 97218 456382 97454
rect 456466 97218 456702 97454
rect 459866 497258 460102 497494
rect 460186 497258 460422 497494
rect 459866 496938 460102 497174
rect 460186 496938 460422 497174
rect 459866 461258 460102 461494
rect 460186 461258 460422 461494
rect 459866 460938 460102 461174
rect 460186 460938 460422 461174
rect 459866 425258 460102 425494
rect 460186 425258 460422 425494
rect 459866 424938 460102 425174
rect 460186 424938 460422 425174
rect 459866 389258 460102 389494
rect 460186 389258 460422 389494
rect 459866 388938 460102 389174
rect 460186 388938 460422 389174
rect 469826 471218 470062 471454
rect 470146 471218 470382 471454
rect 469826 470898 470062 471134
rect 470146 470898 470382 471134
rect 469826 435218 470062 435454
rect 470146 435218 470382 435454
rect 469826 434898 470062 435134
rect 470146 434898 470382 435134
rect 469826 399218 470062 399454
rect 470146 399218 470382 399454
rect 469826 398898 470062 399134
rect 470146 398898 470382 399134
rect 473546 582938 473782 583174
rect 473866 582938 474102 583174
rect 473546 582618 473782 582854
rect 473866 582618 474102 582854
rect 473546 546938 473782 547174
rect 473866 546938 474102 547174
rect 473546 546618 473782 546854
rect 473866 546618 474102 546854
rect 473546 510938 473782 511174
rect 473866 510938 474102 511174
rect 473546 510618 473782 510854
rect 473866 510618 474102 510854
rect 473546 474938 473782 475174
rect 473866 474938 474102 475174
rect 473546 474618 473782 474854
rect 473866 474618 474102 474854
rect 473458 435218 473694 435454
rect 473458 434898 473694 435134
rect 475930 438938 476166 439174
rect 475930 438618 476166 438854
rect 477266 586658 477502 586894
rect 477586 586658 477822 586894
rect 477266 586338 477502 586574
rect 477586 586338 477822 586574
rect 477266 550658 477502 550894
rect 477586 550658 477822 550894
rect 477266 550338 477502 550574
rect 477586 550338 477822 550574
rect 477266 514658 477502 514894
rect 477586 514658 477822 514894
rect 477266 514338 477502 514574
rect 477586 514338 477822 514574
rect 477266 478658 477502 478894
rect 477586 478658 477822 478894
rect 477266 478338 477502 478574
rect 477586 478338 477822 478574
rect 477266 442658 477502 442894
rect 477586 442658 477822 442894
rect 477266 442338 477502 442574
rect 477586 442338 477822 442574
rect 478403 435218 478639 435454
rect 478403 434898 478639 435134
rect 477266 406658 477502 406894
rect 477586 406658 477822 406894
rect 477266 406338 477502 406574
rect 477586 406338 477822 406574
rect 480986 590378 481222 590614
rect 481306 590378 481542 590614
rect 480986 590058 481222 590294
rect 481306 590058 481542 590294
rect 480986 554378 481222 554614
rect 481306 554378 481542 554614
rect 480986 554058 481222 554294
rect 481306 554058 481542 554294
rect 480986 518378 481222 518614
rect 481306 518378 481542 518614
rect 480986 518058 481222 518294
rect 481306 518058 481542 518294
rect 484706 594098 484942 594334
rect 485026 594098 485262 594334
rect 484706 593778 484942 594014
rect 485026 593778 485262 594014
rect 484706 558098 484942 558334
rect 485026 558098 485262 558334
rect 484706 557778 484942 558014
rect 485026 557778 485262 558014
rect 484706 522098 484942 522334
rect 485026 522098 485262 522334
rect 484706 521778 484942 522014
rect 485026 521778 485262 522014
rect 488426 597818 488662 598054
rect 488746 597818 488982 598054
rect 488426 597498 488662 597734
rect 488746 597498 488982 597734
rect 488426 561818 488662 562054
rect 488746 561818 488982 562054
rect 488426 561498 488662 561734
rect 488746 561498 488982 561734
rect 488426 525818 488662 526054
rect 488746 525818 488982 526054
rect 488426 525498 488662 525734
rect 488746 525498 488982 525734
rect 492146 565538 492382 565774
rect 492466 565538 492702 565774
rect 492146 565218 492382 565454
rect 492466 565218 492702 565454
rect 492146 529538 492382 529774
rect 492466 529538 492702 529774
rect 492146 529218 492382 529454
rect 492466 529218 492702 529454
rect 482205 507218 482441 507454
rect 482205 506898 482441 507134
rect 480986 482378 481222 482614
rect 481306 482378 481542 482614
rect 480986 482058 481222 482294
rect 481306 482058 481542 482294
rect 483424 510938 483660 511174
rect 483424 510618 483660 510854
rect 485862 510938 486098 511174
rect 485862 510618 486098 510854
rect 488300 510938 488536 511174
rect 488300 510618 488536 510854
rect 490738 510938 490974 511174
rect 490738 510618 490974 510854
rect 484643 507218 484879 507454
rect 484643 506898 484879 507134
rect 487081 507218 487317 507454
rect 487081 506898 487317 507134
rect 489519 507218 489755 507454
rect 489519 506898 489755 507134
rect 484706 486098 484942 486334
rect 485026 486098 485262 486334
rect 484706 485778 484942 486014
rect 485026 485778 485262 486014
rect 488426 489818 488662 490054
rect 488746 489818 488982 490054
rect 488426 489498 488662 489734
rect 488746 489498 488982 489734
rect 488426 453771 488662 454007
rect 488746 453771 488982 454007
rect 484706 450098 484942 450334
rect 485026 450098 485262 450334
rect 484706 449778 484942 450014
rect 485026 449778 485262 450014
rect 480875 438938 481111 439174
rect 480875 438618 481111 438854
rect 483348 435218 483584 435454
rect 483348 434898 483584 435134
rect 485820 438938 486056 439174
rect 485820 438618 486056 438854
rect 488293 435218 488529 435454
rect 488293 434898 488529 435134
rect 484706 414098 484942 414334
rect 485026 414098 485262 414334
rect 484706 413778 484942 414014
rect 485026 413778 485262 414014
rect 492146 493538 492382 493774
rect 492466 493538 492702 493774
rect 492146 493218 492382 493454
rect 492466 493218 492702 493454
rect 492146 457538 492382 457774
rect 492466 457538 492702 457774
rect 492146 457218 492382 457454
rect 492466 457218 492702 457454
rect 490765 438938 491001 439174
rect 490765 438618 491001 438854
rect 492146 421538 492382 421774
rect 492466 421538 492702 421774
rect 492146 421218 492382 421454
rect 492466 421218 492702 421454
rect 492146 385538 492382 385774
rect 492466 385538 492702 385774
rect 492146 385218 492382 385454
rect 492466 385218 492702 385454
rect 495866 569258 496102 569494
rect 496186 569258 496422 569494
rect 495866 568938 496102 569174
rect 496186 568938 496422 569174
rect 495866 533258 496102 533494
rect 496186 533258 496422 533494
rect 495866 532938 496102 533174
rect 496186 532938 496422 533174
rect 495866 497258 496102 497494
rect 496186 497258 496422 497494
rect 495866 496938 496102 497174
rect 496186 496938 496422 497174
rect 495866 461258 496102 461494
rect 496186 461258 496422 461494
rect 495866 460938 496102 461174
rect 496186 460938 496422 461174
rect 495866 425258 496102 425494
rect 496186 425258 496422 425494
rect 495866 424938 496102 425174
rect 496186 424938 496422 425174
rect 495866 389258 496102 389494
rect 496186 389258 496422 389494
rect 495866 388938 496102 389174
rect 496186 388938 496422 389174
rect 505826 579218 506062 579454
rect 506146 579218 506382 579454
rect 505826 578898 506062 579134
rect 506146 578898 506382 579134
rect 505826 543218 506062 543454
rect 506146 543218 506382 543454
rect 505826 542898 506062 543134
rect 506146 542898 506382 543134
rect 505826 507218 506062 507454
rect 506146 507218 506382 507454
rect 505826 506898 506062 507134
rect 506146 506898 506382 507134
rect 505826 471218 506062 471454
rect 506146 471218 506382 471454
rect 505826 470898 506062 471134
rect 506146 470898 506382 471134
rect 505826 435218 506062 435454
rect 506146 435218 506382 435454
rect 505826 434898 506062 435134
rect 506146 434898 506382 435134
rect 505826 399218 506062 399454
rect 506146 399218 506382 399454
rect 505826 398898 506062 399134
rect 506146 398898 506382 399134
rect 469610 366938 469846 367174
rect 469610 366618 469846 366854
rect 500330 366938 500566 367174
rect 500330 366618 500566 366854
rect 484970 363218 485206 363454
rect 484970 362898 485206 363134
rect 505826 363218 506062 363454
rect 506146 363218 506382 363454
rect 505826 362898 506062 363134
rect 506146 362898 506382 363134
rect 459866 353258 460102 353494
rect 460186 353258 460422 353494
rect 459866 352938 460102 353174
rect 460186 352938 460422 353174
rect 469610 330938 469846 331174
rect 469610 330618 469846 330854
rect 500330 330938 500566 331174
rect 500330 330618 500566 330854
rect 484970 327218 485206 327454
rect 484970 326898 485206 327134
rect 505826 327218 506062 327454
rect 506146 327218 506382 327454
rect 505826 326898 506062 327134
rect 506146 326898 506382 327134
rect 459866 317258 460102 317494
rect 460186 317258 460422 317494
rect 459866 316938 460102 317174
rect 460186 316938 460422 317174
rect 459866 281258 460102 281494
rect 460186 281258 460422 281494
rect 459866 280938 460102 281174
rect 460186 280938 460422 281174
rect 459866 245258 460102 245494
rect 460186 245258 460422 245494
rect 459866 244938 460102 245174
rect 460186 244938 460422 245174
rect 459866 209258 460102 209494
rect 460186 209258 460422 209494
rect 459866 208938 460102 209174
rect 460186 208938 460422 209174
rect 459866 173258 460102 173494
rect 460186 173258 460422 173494
rect 459866 172938 460102 173174
rect 460186 172938 460422 173174
rect 459866 137258 460102 137494
rect 460186 137258 460422 137494
rect 459866 136938 460102 137174
rect 460186 136938 460422 137174
rect 459866 101258 460102 101494
rect 460186 101258 460422 101494
rect 459866 100938 460102 101174
rect 460186 100938 460422 101174
rect 405610 78938 405846 79174
rect 405610 78618 405846 78854
rect 436330 78938 436566 79174
rect 436330 78618 436566 78854
rect 390250 75218 390486 75454
rect 390250 74898 390486 75134
rect 420970 75218 421206 75454
rect 420970 74898 421206 75134
rect 451690 75218 451926 75454
rect 451690 74898 451926 75134
rect 384146 61538 384382 61774
rect 384466 61538 384702 61774
rect 384146 61218 384382 61454
rect 384466 61218 384702 61454
rect 459866 65258 460102 65494
rect 460186 65258 460422 65494
rect 459866 64938 460102 65174
rect 460186 64938 460422 65174
rect 405610 42938 405846 43174
rect 405610 42618 405846 42854
rect 436330 42938 436566 43174
rect 436330 42618 436566 42854
rect 390250 39218 390486 39454
rect 390250 38898 390486 39134
rect 420970 39218 421206 39454
rect 420970 38898 421206 39134
rect 451690 39218 451926 39454
rect 451690 38898 451926 39134
rect 384146 25538 384382 25774
rect 384466 25538 384702 25774
rect 384146 25218 384382 25454
rect 384466 25218 384702 25454
rect 384146 -6342 384382 -6106
rect 384466 -6342 384702 -6106
rect 384146 -6662 384382 -6426
rect 384466 -6662 384702 -6426
rect 387866 29258 388102 29494
rect 388186 29258 388422 29494
rect 387866 28938 388102 29174
rect 388186 28938 388422 29174
rect 387866 -7302 388102 -7066
rect 388186 -7302 388422 -7066
rect 387866 -7622 388102 -7386
rect 388186 -7622 388422 -7386
rect 397826 3218 398062 3454
rect 398146 3218 398382 3454
rect 397826 2898 398062 3134
rect 398146 2898 398382 3134
rect 397826 -582 398062 -346
rect 398146 -582 398382 -346
rect 397826 -902 398062 -666
rect 398146 -902 398382 -666
rect 401546 6938 401782 7174
rect 401866 6938 402102 7174
rect 401546 6618 401782 6854
rect 401866 6618 402102 6854
rect 401546 -1542 401782 -1306
rect 401866 -1542 402102 -1306
rect 401546 -1862 401782 -1626
rect 401866 -1862 402102 -1626
rect 405266 10658 405502 10894
rect 405586 10658 405822 10894
rect 405266 10338 405502 10574
rect 405586 10338 405822 10574
rect 405266 -2502 405502 -2266
rect 405586 -2502 405822 -2266
rect 405266 -2822 405502 -2586
rect 405586 -2822 405822 -2586
rect 408986 14378 409222 14614
rect 409306 14378 409542 14614
rect 408986 14058 409222 14294
rect 409306 14058 409542 14294
rect 408986 -3462 409222 -3226
rect 409306 -3462 409542 -3226
rect 408986 -3782 409222 -3546
rect 409306 -3782 409542 -3546
rect 412706 18098 412942 18334
rect 413026 18098 413262 18334
rect 412706 17778 412942 18014
rect 413026 17778 413262 18014
rect 412706 -4422 412942 -4186
rect 413026 -4422 413262 -4186
rect 412706 -4742 412942 -4506
rect 413026 -4742 413262 -4506
rect 416426 21818 416662 22054
rect 416746 21818 416982 22054
rect 416426 21498 416662 21734
rect 416746 21498 416982 21734
rect 416426 -5382 416662 -5146
rect 416746 -5382 416982 -5146
rect 416426 -5702 416662 -5466
rect 416746 -5702 416982 -5466
rect 420146 25538 420382 25774
rect 420466 25538 420702 25774
rect 420146 25218 420382 25454
rect 420466 25218 420702 25454
rect 420146 -6342 420382 -6106
rect 420466 -6342 420702 -6106
rect 420146 -6662 420382 -6426
rect 420466 -6662 420702 -6426
rect 423866 29258 424102 29494
rect 424186 29258 424422 29494
rect 423866 28938 424102 29174
rect 424186 28938 424422 29174
rect 423866 -7302 424102 -7066
rect 424186 -7302 424422 -7066
rect 423866 -7622 424102 -7386
rect 424186 -7622 424422 -7386
rect 433826 3218 434062 3454
rect 434146 3218 434382 3454
rect 433826 2898 434062 3134
rect 434146 2898 434382 3134
rect 433826 -582 434062 -346
rect 434146 -582 434382 -346
rect 433826 -902 434062 -666
rect 434146 -902 434382 -666
rect 437546 6938 437782 7174
rect 437866 6938 438102 7174
rect 437546 6618 437782 6854
rect 437866 6618 438102 6854
rect 437546 -1542 437782 -1306
rect 437866 -1542 438102 -1306
rect 437546 -1862 437782 -1626
rect 437866 -1862 438102 -1626
rect 441266 10658 441502 10894
rect 441586 10658 441822 10894
rect 441266 10338 441502 10574
rect 441586 10338 441822 10574
rect 441266 -2502 441502 -2266
rect 441586 -2502 441822 -2266
rect 441266 -2822 441502 -2586
rect 441586 -2822 441822 -2586
rect 444986 14378 445222 14614
rect 445306 14378 445542 14614
rect 444986 14058 445222 14294
rect 445306 14058 445542 14294
rect 444986 -3462 445222 -3226
rect 445306 -3462 445542 -3226
rect 444986 -3782 445222 -3546
rect 445306 -3782 445542 -3546
rect 448706 18098 448942 18334
rect 449026 18098 449262 18334
rect 448706 17778 448942 18014
rect 449026 17778 449262 18014
rect 448706 -4422 448942 -4186
rect 449026 -4422 449262 -4186
rect 448706 -4742 448942 -4506
rect 449026 -4742 449262 -4506
rect 452426 21818 452662 22054
rect 452746 21818 452982 22054
rect 452426 21498 452662 21734
rect 452746 21498 452982 21734
rect 452426 -5382 452662 -5146
rect 452746 -5382 452982 -5146
rect 452426 -5702 452662 -5466
rect 452746 -5702 452982 -5466
rect 456146 25538 456382 25774
rect 456466 25538 456702 25774
rect 456146 25218 456382 25454
rect 456466 25218 456702 25454
rect 456146 -6342 456382 -6106
rect 456466 -6342 456702 -6106
rect 456146 -6662 456382 -6426
rect 456466 -6662 456702 -6426
rect 459866 29258 460102 29494
rect 460186 29258 460422 29494
rect 459866 28938 460102 29174
rect 460186 28938 460422 29174
rect 477266 298658 477502 298894
rect 477586 298658 477822 298894
rect 477266 298338 477502 298574
rect 477586 298338 477822 298574
rect 477266 262658 477502 262894
rect 477586 262658 477822 262894
rect 477266 262338 477502 262574
rect 477586 262338 477822 262574
rect 480986 302378 481222 302614
rect 481306 302378 481542 302614
rect 480986 302058 481222 302294
rect 481306 302058 481542 302294
rect 480986 266378 481222 266614
rect 481306 266378 481542 266614
rect 480986 266058 481222 266294
rect 481306 266058 481542 266294
rect 484706 306098 484942 306334
rect 485026 306098 485262 306334
rect 484706 305778 484942 306014
rect 485026 305778 485262 306014
rect 484706 270098 484942 270334
rect 485026 270098 485262 270334
rect 484706 269778 484942 270014
rect 485026 269778 485262 270014
rect 488426 309818 488662 310054
rect 488746 309818 488982 310054
rect 488426 309498 488662 309734
rect 488746 309498 488982 309734
rect 488426 273818 488662 274054
rect 488746 273818 488982 274054
rect 488426 273498 488662 273734
rect 488746 273498 488982 273734
rect 492146 313538 492382 313774
rect 492466 313538 492702 313774
rect 492146 313218 492382 313454
rect 492466 313218 492702 313454
rect 492146 277538 492382 277774
rect 492466 277538 492702 277774
rect 492146 277218 492382 277454
rect 492466 277218 492702 277454
rect 495866 317258 496102 317494
rect 496186 317258 496422 317494
rect 495866 316938 496102 317174
rect 496186 316938 496422 317174
rect 495866 281258 496102 281494
rect 496186 281258 496422 281494
rect 495866 280938 496102 281174
rect 496186 280938 496422 281174
rect 509546 582938 509782 583174
rect 509866 582938 510102 583174
rect 509546 582618 509782 582854
rect 509866 582618 510102 582854
rect 509546 546938 509782 547174
rect 509866 546938 510102 547174
rect 509546 546618 509782 546854
rect 509866 546618 510102 546854
rect 509546 510938 509782 511174
rect 509866 510938 510102 511174
rect 509546 510618 509782 510854
rect 509866 510618 510102 510854
rect 509546 474938 509782 475174
rect 509866 474938 510102 475174
rect 509546 474618 509782 474854
rect 509866 474618 510102 474854
rect 509546 438938 509782 439174
rect 509866 438938 510102 439174
rect 509546 438618 509782 438854
rect 509866 438618 510102 438854
rect 509546 402938 509782 403174
rect 509866 402938 510102 403174
rect 509546 402618 509782 402854
rect 509866 402618 510102 402854
rect 509546 366938 509782 367174
rect 509866 366938 510102 367174
rect 509546 366618 509782 366854
rect 509866 366618 510102 366854
rect 513266 586658 513502 586894
rect 513586 586658 513822 586894
rect 513266 586338 513502 586574
rect 513586 586338 513822 586574
rect 513266 550658 513502 550894
rect 513586 550658 513822 550894
rect 513266 550338 513502 550574
rect 513586 550338 513822 550574
rect 513266 514658 513502 514894
rect 513586 514658 513822 514894
rect 513266 514338 513502 514574
rect 513586 514338 513822 514574
rect 513266 478658 513502 478894
rect 513586 478658 513822 478894
rect 513266 478338 513502 478574
rect 513586 478338 513822 478574
rect 513266 442658 513502 442894
rect 513586 442658 513822 442894
rect 513266 442338 513502 442574
rect 513586 442338 513822 442574
rect 513266 406658 513502 406894
rect 513586 406658 513822 406894
rect 513266 406338 513502 406574
rect 513586 406338 513822 406574
rect 513266 370658 513502 370894
rect 513586 370658 513822 370894
rect 513266 370338 513502 370574
rect 513586 370338 513822 370574
rect 509546 330938 509782 331174
rect 509866 330938 510102 331174
rect 509546 330618 509782 330854
rect 509866 330618 510102 330854
rect 505826 291218 506062 291454
rect 506146 291218 506382 291454
rect 505826 290898 506062 291134
rect 506146 290898 506382 291134
rect 513266 334658 513502 334894
rect 513586 334658 513822 334894
rect 513266 334338 513502 334574
rect 513586 334338 513822 334574
rect 516986 590378 517222 590614
rect 517306 590378 517542 590614
rect 516986 590058 517222 590294
rect 517306 590058 517542 590294
rect 516986 554378 517222 554614
rect 517306 554378 517542 554614
rect 516986 554058 517222 554294
rect 517306 554058 517542 554294
rect 516986 518378 517222 518614
rect 517306 518378 517542 518614
rect 516986 518058 517222 518294
rect 517306 518058 517542 518294
rect 516986 482378 517222 482614
rect 517306 482378 517542 482614
rect 516986 482058 517222 482294
rect 517306 482058 517542 482294
rect 516986 446378 517222 446614
rect 517306 446378 517542 446614
rect 516986 446058 517222 446294
rect 517306 446058 517542 446294
rect 516986 410378 517222 410614
rect 517306 410378 517542 410614
rect 516986 410058 517222 410294
rect 517306 410058 517542 410294
rect 516986 374378 517222 374614
rect 517306 374378 517542 374614
rect 516986 374058 517222 374294
rect 517306 374058 517542 374294
rect 516986 338378 517222 338614
rect 517306 338378 517542 338614
rect 516986 338058 517222 338294
rect 517306 338058 517542 338294
rect 513266 298658 513502 298894
rect 513586 298658 513822 298894
rect 513266 298338 513502 298574
rect 513586 298338 513822 298574
rect 509546 294938 509782 295174
rect 509866 294938 510102 295174
rect 509546 294618 509782 294854
rect 509866 294618 510102 294854
rect 520706 594098 520942 594334
rect 521026 594098 521262 594334
rect 520706 593778 520942 594014
rect 521026 593778 521262 594014
rect 520706 558098 520942 558334
rect 521026 558098 521262 558334
rect 520706 557778 520942 558014
rect 521026 557778 521262 558014
rect 520706 522098 520942 522334
rect 521026 522098 521262 522334
rect 520706 521778 520942 522014
rect 521026 521778 521262 522014
rect 520706 486098 520942 486334
rect 521026 486098 521262 486334
rect 520706 485778 520942 486014
rect 521026 485778 521262 486014
rect 520706 450098 520942 450334
rect 521026 450098 521262 450334
rect 520706 449778 520942 450014
rect 521026 449778 521262 450014
rect 520706 414098 520942 414334
rect 521026 414098 521262 414334
rect 520706 413778 520942 414014
rect 521026 413778 521262 414014
rect 520706 378098 520942 378334
rect 521026 378098 521262 378334
rect 520706 377778 520942 378014
rect 521026 377778 521262 378014
rect 520706 342098 520942 342334
rect 521026 342098 521262 342334
rect 520706 341778 520942 342014
rect 521026 341778 521262 342014
rect 516986 302378 517222 302614
rect 517306 302378 517542 302614
rect 516986 302058 517222 302294
rect 517306 302058 517542 302294
rect 513266 262658 513502 262894
rect 513586 262658 513822 262894
rect 513266 262338 513502 262574
rect 513586 262338 513822 262574
rect 520706 306098 520942 306334
rect 521026 306098 521262 306334
rect 520706 305778 520942 306014
rect 521026 305778 521262 306014
rect 516986 266378 517222 266614
rect 517306 266378 517542 266614
rect 516986 266058 517222 266294
rect 517306 266058 517542 266294
rect 520706 270098 520942 270334
rect 521026 270098 521262 270334
rect 520706 269778 520942 270014
rect 521026 269778 521262 270014
rect 524426 709402 524662 709638
rect 524746 709402 524982 709638
rect 524426 709082 524662 709318
rect 524746 709082 524982 709318
rect 528146 710362 528382 710598
rect 528466 710362 528702 710598
rect 528146 710042 528382 710278
rect 528466 710042 528702 710278
rect 524426 669818 524662 670054
rect 524746 669818 524982 670054
rect 524426 669498 524662 669734
rect 524746 669498 524982 669734
rect 525690 651218 525926 651454
rect 525690 650898 525926 651134
rect 524426 633818 524662 634054
rect 524746 633818 524982 634054
rect 524426 633498 524662 633734
rect 524746 633498 524982 633734
rect 525690 615218 525926 615454
rect 525690 614898 525926 615134
rect 524426 597818 524662 598054
rect 524746 597818 524982 598054
rect 524426 597498 524662 597734
rect 524746 597498 524982 597734
rect 524426 561818 524662 562054
rect 524746 561818 524982 562054
rect 524426 561498 524662 561734
rect 524746 561498 524982 561734
rect 524426 525818 524662 526054
rect 524746 525818 524982 526054
rect 524426 525498 524662 525734
rect 524746 525498 524982 525734
rect 531866 711322 532102 711558
rect 532186 711322 532422 711558
rect 531866 711002 532102 711238
rect 532186 711002 532422 711238
rect 528146 673538 528382 673774
rect 528466 673538 528702 673774
rect 528146 673218 528382 673454
rect 528466 673218 528702 673454
rect 528146 637538 528382 637774
rect 528466 637538 528702 637774
rect 528146 637218 528382 637454
rect 528466 637218 528702 637454
rect 528146 601538 528382 601774
rect 528466 601538 528702 601774
rect 528146 601218 528382 601454
rect 528466 601218 528702 601454
rect 528146 565538 528382 565774
rect 528466 565538 528702 565774
rect 528146 565218 528382 565454
rect 528466 565218 528702 565454
rect 528146 529538 528382 529774
rect 528466 529538 528702 529774
rect 528146 529218 528382 529454
rect 528466 529218 528702 529454
rect 524426 489818 524662 490054
rect 524746 489818 524982 490054
rect 524426 489498 524662 489734
rect 524746 489498 524982 489734
rect 524426 453818 524662 454054
rect 524746 453818 524982 454054
rect 524426 453498 524662 453734
rect 524746 453498 524982 453734
rect 528146 493538 528382 493774
rect 528466 493538 528702 493774
rect 528146 493218 528382 493454
rect 528466 493218 528702 493454
rect 528146 457538 528382 457774
rect 528466 457538 528702 457774
rect 528146 457218 528382 457454
rect 528466 457218 528702 457454
rect 525206 435218 525442 435454
rect 525206 434898 525442 435134
rect 524426 417818 524662 418054
rect 524746 417818 524982 418054
rect 524426 417498 524662 417734
rect 524746 417498 524982 417734
rect 524426 381818 524662 382054
rect 524746 381818 524982 382054
rect 524426 381498 524662 381734
rect 524746 381498 524982 381734
rect 524426 345818 524662 346054
rect 524746 345818 524982 346054
rect 524426 345498 524662 345734
rect 524746 345498 524982 345734
rect 524426 309818 524662 310054
rect 524746 309818 524982 310054
rect 524426 309498 524662 309734
rect 524746 309498 524982 309734
rect 524426 273818 524662 274054
rect 524746 273818 524982 274054
rect 524426 273498 524662 273734
rect 524746 273498 524982 273734
rect 529426 438938 529662 439174
rect 529426 438618 529662 438854
rect 528146 421538 528382 421774
rect 528466 421538 528702 421774
rect 528146 421218 528382 421454
rect 528466 421218 528702 421454
rect 528146 385538 528382 385774
rect 528466 385538 528702 385774
rect 528146 385218 528382 385454
rect 528466 385218 528702 385454
rect 528146 349538 528382 349774
rect 528466 349538 528702 349774
rect 528146 349218 528382 349454
rect 528466 349218 528702 349454
rect 531866 677258 532102 677494
rect 532186 677258 532422 677494
rect 531866 676938 532102 677174
rect 532186 676938 532422 677174
rect 531866 641258 532102 641494
rect 532186 641258 532422 641494
rect 531866 640938 532102 641174
rect 532186 640938 532422 641174
rect 531866 605258 532102 605494
rect 532186 605258 532422 605494
rect 531866 604938 532102 605174
rect 532186 604938 532422 605174
rect 531866 569258 532102 569494
rect 532186 569258 532422 569494
rect 531866 568938 532102 569174
rect 532186 568938 532422 569174
rect 531866 533258 532102 533494
rect 532186 533258 532422 533494
rect 531866 532938 532102 533174
rect 532186 532938 532422 533174
rect 531866 497258 532102 497494
rect 532186 497258 532422 497494
rect 531866 496938 532102 497174
rect 532186 496938 532422 497174
rect 531866 461258 532102 461494
rect 532186 461258 532422 461494
rect 531866 460938 532102 461174
rect 532186 460938 532422 461174
rect 541826 704602 542062 704838
rect 542146 704602 542382 704838
rect 541826 704282 542062 704518
rect 542146 704282 542382 704518
rect 541826 687218 542062 687454
rect 542146 687218 542382 687454
rect 541826 686898 542062 687134
rect 542146 686898 542382 687134
rect 541826 651218 542062 651454
rect 542146 651218 542382 651454
rect 541826 650898 542062 651134
rect 542146 650898 542382 651134
rect 541826 615218 542062 615454
rect 542146 615218 542382 615454
rect 541826 614898 542062 615134
rect 542146 614898 542382 615134
rect 541826 579218 542062 579454
rect 542146 579218 542382 579454
rect 541826 578898 542062 579134
rect 542146 578898 542382 579134
rect 541826 543218 542062 543454
rect 542146 543218 542382 543454
rect 541826 542898 542062 543134
rect 542146 542898 542382 543134
rect 541826 507218 542062 507454
rect 542146 507218 542382 507454
rect 541826 506898 542062 507134
rect 542146 506898 542382 507134
rect 541826 471218 542062 471454
rect 542146 471218 542382 471454
rect 541826 470898 542062 471134
rect 542146 470898 542382 471134
rect 545546 705562 545782 705798
rect 545866 705562 546102 705798
rect 545546 705242 545782 705478
rect 545866 705242 546102 705478
rect 545546 690938 545782 691174
rect 545866 690938 546102 691174
rect 545546 690618 545782 690854
rect 545866 690618 546102 690854
rect 545546 654938 545782 655174
rect 545866 654938 546102 655174
rect 545546 654618 545782 654854
rect 545866 654618 546102 654854
rect 545546 618938 545782 619174
rect 545866 618938 546102 619174
rect 545546 618618 545782 618854
rect 545866 618618 546102 618854
rect 545546 582938 545782 583174
rect 545866 582938 546102 583174
rect 545546 582618 545782 582854
rect 545866 582618 546102 582854
rect 545546 546938 545782 547174
rect 545866 546938 546102 547174
rect 545546 546618 545782 546854
rect 545866 546618 546102 546854
rect 545546 510938 545782 511174
rect 545866 510938 546102 511174
rect 545546 510618 545782 510854
rect 545866 510618 546102 510854
rect 545546 474938 545782 475174
rect 545866 474938 546102 475174
rect 545546 474618 545782 474854
rect 545866 474618 546102 474854
rect 537867 438938 538103 439174
rect 537867 438618 538103 438854
rect 549266 706522 549502 706758
rect 549586 706522 549822 706758
rect 549266 706202 549502 706438
rect 549586 706202 549822 706438
rect 549266 694658 549502 694894
rect 549586 694658 549822 694894
rect 549266 694338 549502 694574
rect 549586 694338 549822 694574
rect 549266 658658 549502 658894
rect 549586 658658 549822 658894
rect 549266 658338 549502 658574
rect 549586 658338 549822 658574
rect 549266 622658 549502 622894
rect 549586 622658 549822 622894
rect 549266 622338 549502 622574
rect 549586 622338 549822 622574
rect 549266 586658 549502 586894
rect 549586 586658 549822 586894
rect 549266 586338 549502 586574
rect 549586 586338 549822 586574
rect 549266 550658 549502 550894
rect 549586 550658 549822 550894
rect 549266 550338 549502 550574
rect 549586 550338 549822 550574
rect 549266 514658 549502 514894
rect 549586 514658 549822 514894
rect 549266 514338 549502 514574
rect 549586 514338 549822 514574
rect 549266 478658 549502 478894
rect 549586 478658 549822 478894
rect 549266 478338 549502 478574
rect 549586 478338 549822 478574
rect 549266 442658 549502 442894
rect 549586 442658 549822 442894
rect 549266 442338 549502 442574
rect 549586 442338 549822 442574
rect 545546 438938 545782 439174
rect 545866 438938 546102 439174
rect 545546 438618 545782 438854
rect 545866 438618 546102 438854
rect 533647 435218 533883 435454
rect 533647 434898 533883 435134
rect 542088 435218 542324 435454
rect 542088 434898 542324 435134
rect 531866 425258 532102 425494
rect 532186 425258 532422 425494
rect 531866 424938 532102 425174
rect 532186 424938 532422 425174
rect 531866 389258 532102 389494
rect 532186 389258 532422 389494
rect 531866 388938 532102 389174
rect 532186 388938 532422 389174
rect 531866 353258 532102 353494
rect 532186 353258 532422 353494
rect 531866 352938 532102 353174
rect 532186 352938 532422 353174
rect 528146 313538 528382 313774
rect 528466 313538 528702 313774
rect 528146 313218 528382 313454
rect 528466 313218 528702 313454
rect 528146 277538 528382 277774
rect 528466 277538 528702 277774
rect 528146 277218 528382 277454
rect 528466 277218 528702 277454
rect 531866 317258 532102 317494
rect 532186 317258 532422 317494
rect 531866 316938 532102 317174
rect 532186 316938 532422 317174
rect 541826 399218 542062 399454
rect 542146 399218 542382 399454
rect 541826 398898 542062 399134
rect 542146 398898 542382 399134
rect 541826 363218 542062 363454
rect 542146 363218 542382 363454
rect 541826 362898 542062 363134
rect 542146 362898 542382 363134
rect 541826 327218 542062 327454
rect 542146 327218 542382 327454
rect 541826 326898 542062 327134
rect 542146 326898 542382 327134
rect 531866 281258 532102 281494
rect 532186 281258 532422 281494
rect 531866 280938 532102 281174
rect 532186 280938 532422 281174
rect 479610 258938 479846 259174
rect 479610 258618 479846 258854
rect 510330 258938 510566 259174
rect 510330 258618 510566 258854
rect 464250 255218 464486 255454
rect 464250 254898 464486 255134
rect 494970 255218 495206 255454
rect 494970 254898 495206 255134
rect 525690 255218 525926 255454
rect 525690 254898 525926 255134
rect 531866 245258 532102 245494
rect 532186 245258 532422 245494
rect 531866 244938 532102 245174
rect 532186 244938 532422 245174
rect 479610 222938 479846 223174
rect 479610 222618 479846 222854
rect 510330 222938 510566 223174
rect 510330 222618 510566 222854
rect 464250 219218 464486 219454
rect 464250 218898 464486 219134
rect 494970 219218 495206 219454
rect 494970 218898 495206 219134
rect 525690 219218 525926 219454
rect 525690 218898 525926 219134
rect 531866 209258 532102 209494
rect 532186 209258 532422 209494
rect 531866 208938 532102 209174
rect 532186 208938 532422 209174
rect 469826 183218 470062 183454
rect 470146 183218 470382 183454
rect 469826 182898 470062 183134
rect 470146 182898 470382 183134
rect 469826 147218 470062 147454
rect 470146 147218 470382 147454
rect 469826 146898 470062 147134
rect 470146 146898 470382 147134
rect 469826 111218 470062 111454
rect 470146 111218 470382 111454
rect 469826 110898 470062 111134
rect 470146 110898 470382 111134
rect 469826 75218 470062 75454
rect 470146 75218 470382 75454
rect 469826 74898 470062 75134
rect 470146 74898 470382 75134
rect 469826 39218 470062 39454
rect 470146 39218 470382 39454
rect 469826 38898 470062 39134
rect 470146 38898 470382 39134
rect 459866 -7302 460102 -7066
rect 460186 -7302 460422 -7066
rect 459866 -7622 460102 -7386
rect 460186 -7622 460422 -7386
rect 469826 3218 470062 3454
rect 470146 3218 470382 3454
rect 469826 2898 470062 3134
rect 470146 2898 470382 3134
rect 469826 -582 470062 -346
rect 470146 -582 470382 -346
rect 469826 -902 470062 -666
rect 470146 -902 470382 -666
rect 473546 186938 473782 187174
rect 473866 186938 474102 187174
rect 473546 186618 473782 186854
rect 473866 186618 474102 186854
rect 473546 150938 473782 151174
rect 473866 150938 474102 151174
rect 473546 150618 473782 150854
rect 473866 150618 474102 150854
rect 473546 114938 473782 115174
rect 473866 114938 474102 115174
rect 473546 114618 473782 114854
rect 473866 114618 474102 114854
rect 473546 78938 473782 79174
rect 473866 78938 474102 79174
rect 473546 78618 473782 78854
rect 473866 78618 474102 78854
rect 473546 42938 473782 43174
rect 473866 42938 474102 43174
rect 473546 42618 473782 42854
rect 473866 42618 474102 42854
rect 473546 6938 473782 7174
rect 473866 6938 474102 7174
rect 473546 6618 473782 6854
rect 473866 6618 474102 6854
rect 473546 -1542 473782 -1306
rect 473866 -1542 474102 -1306
rect 473546 -1862 473782 -1626
rect 473866 -1862 474102 -1626
rect 477266 190658 477502 190894
rect 477586 190658 477822 190894
rect 477266 190338 477502 190574
rect 477586 190338 477822 190574
rect 477266 154658 477502 154894
rect 477586 154658 477822 154894
rect 477266 154338 477502 154574
rect 477586 154338 477822 154574
rect 477266 118658 477502 118894
rect 477586 118658 477822 118894
rect 477266 118338 477502 118574
rect 477586 118338 477822 118574
rect 477266 82658 477502 82894
rect 477586 82658 477822 82894
rect 477266 82338 477502 82574
rect 477586 82338 477822 82574
rect 477266 46658 477502 46894
rect 477586 46658 477822 46894
rect 477266 46338 477502 46574
rect 477586 46338 477822 46574
rect 477266 10658 477502 10894
rect 477586 10658 477822 10894
rect 477266 10338 477502 10574
rect 477586 10338 477822 10574
rect 477266 -2502 477502 -2266
rect 477586 -2502 477822 -2266
rect 477266 -2822 477502 -2586
rect 477586 -2822 477822 -2586
rect 480986 194378 481222 194614
rect 481306 194378 481542 194614
rect 480986 194058 481222 194294
rect 481306 194058 481542 194294
rect 480986 158378 481222 158614
rect 481306 158378 481542 158614
rect 480986 158058 481222 158294
rect 481306 158058 481542 158294
rect 480986 122378 481222 122614
rect 481306 122378 481542 122614
rect 480986 122058 481222 122294
rect 481306 122058 481542 122294
rect 484706 198098 484942 198334
rect 485026 198098 485262 198334
rect 484706 197778 484942 198014
rect 485026 197778 485262 198014
rect 484706 162098 484942 162334
rect 485026 162098 485262 162334
rect 484706 161778 484942 162014
rect 485026 161778 485262 162014
rect 488426 165818 488662 166054
rect 488746 165818 488982 166054
rect 488426 165498 488662 165734
rect 488746 165498 488982 165734
rect 505826 183218 506062 183454
rect 506146 183218 506382 183454
rect 505826 182898 506062 183134
rect 506146 182898 506382 183134
rect 505826 147218 506062 147454
rect 506146 147218 506382 147454
rect 505826 146898 506062 147134
rect 506146 146898 506382 147134
rect 509546 186938 509782 187174
rect 509866 186938 510102 187174
rect 509546 186618 509782 186854
rect 509866 186618 510102 186854
rect 509546 150938 509782 151174
rect 509866 150938 510102 151174
rect 509546 150618 509782 150854
rect 509866 150618 510102 150854
rect 513266 190658 513502 190894
rect 513586 190658 513822 190894
rect 513266 190338 513502 190574
rect 513586 190338 513822 190574
rect 513266 154658 513502 154894
rect 513586 154658 513822 154894
rect 513266 154338 513502 154574
rect 513586 154338 513822 154574
rect 516986 194378 517222 194614
rect 517306 194378 517542 194614
rect 516986 194058 517222 194294
rect 517306 194058 517542 194294
rect 516986 158378 517222 158614
rect 517306 158378 517542 158614
rect 516986 158058 517222 158294
rect 517306 158058 517542 158294
rect 520706 198098 520942 198334
rect 521026 198098 521262 198334
rect 520706 197778 520942 198014
rect 521026 197778 521262 198014
rect 520706 162098 520942 162334
rect 521026 162098 521262 162334
rect 520706 161778 520942 162014
rect 521026 161778 521262 162014
rect 524426 165818 524662 166054
rect 524746 165818 524982 166054
rect 524426 165498 524662 165734
rect 524746 165498 524982 165734
rect 531866 173258 532102 173494
rect 532186 173258 532422 173494
rect 531866 172938 532102 173174
rect 532186 172938 532422 173174
rect 541826 291218 542062 291454
rect 542146 291218 542382 291454
rect 541826 290898 542062 291134
rect 542146 290898 542382 291134
rect 541826 255218 542062 255454
rect 542146 255218 542382 255454
rect 541826 254898 542062 255134
rect 542146 254898 542382 255134
rect 541826 219218 542062 219454
rect 542146 219218 542382 219454
rect 541826 218898 542062 219134
rect 542146 218898 542382 219134
rect 541826 183218 542062 183454
rect 542146 183218 542382 183454
rect 541826 182898 542062 183134
rect 542146 182898 542382 183134
rect 541826 147218 542062 147454
rect 542146 147218 542382 147454
rect 541826 146898 542062 147134
rect 542146 146898 542382 147134
rect 484706 126098 484942 126334
rect 485026 126098 485262 126334
rect 484706 125778 484942 126014
rect 485026 125778 485262 126014
rect 484250 111218 484486 111454
rect 484250 110898 484486 111134
rect 480986 86378 481222 86614
rect 481306 86378 481542 86614
rect 480986 86058 481222 86294
rect 481306 86058 481542 86294
rect 480986 50378 481222 50614
rect 481306 50378 481542 50614
rect 480986 50058 481222 50294
rect 481306 50058 481542 50294
rect 480986 14378 481222 14614
rect 481306 14378 481542 14614
rect 480986 14058 481222 14294
rect 481306 14058 481542 14294
rect 480986 -3462 481222 -3226
rect 481306 -3462 481542 -3226
rect 480986 -3782 481222 -3546
rect 481306 -3782 481542 -3546
rect 499610 114938 499846 115174
rect 499610 114618 499846 114854
rect 530330 114938 530566 115174
rect 530330 114618 530566 114854
rect 514970 111218 515206 111454
rect 514970 110898 515206 111134
rect 541826 111218 542062 111454
rect 542146 111218 542382 111454
rect 541826 110898 542062 111134
rect 542146 110898 542382 111134
rect 484706 90098 484942 90334
rect 485026 90098 485262 90334
rect 484706 89778 484942 90014
rect 485026 89778 485262 90014
rect 484706 54098 484942 54334
rect 485026 54098 485262 54334
rect 484706 53778 484942 54014
rect 485026 53778 485262 54014
rect 484706 18098 484942 18334
rect 485026 18098 485262 18334
rect 484706 17778 484942 18014
rect 485026 17778 485262 18014
rect 484706 -4422 484942 -4186
rect 485026 -4422 485262 -4186
rect 484706 -4742 484942 -4506
rect 485026 -4742 485262 -4506
rect 488426 57818 488662 58054
rect 488746 57818 488982 58054
rect 488426 57498 488662 57734
rect 488746 57498 488982 57734
rect 488426 21818 488662 22054
rect 488746 21818 488982 22054
rect 488426 21498 488662 21734
rect 488746 21498 488982 21734
rect 488426 -5382 488662 -5146
rect 488746 -5382 488982 -5146
rect 488426 -5702 488662 -5466
rect 488746 -5702 488982 -5466
rect 492146 61538 492382 61774
rect 492466 61538 492702 61774
rect 492146 61218 492382 61454
rect 492466 61218 492702 61454
rect 492146 25538 492382 25774
rect 492466 25538 492702 25774
rect 492146 25218 492382 25454
rect 492466 25218 492702 25454
rect 492146 -6342 492382 -6106
rect 492466 -6342 492702 -6106
rect 492146 -6662 492382 -6426
rect 492466 -6662 492702 -6426
rect 495866 65258 496102 65494
rect 496186 65258 496422 65494
rect 495866 64938 496102 65174
rect 496186 64938 496422 65174
rect 495866 29258 496102 29494
rect 496186 29258 496422 29494
rect 495866 28938 496102 29174
rect 496186 28938 496422 29174
rect 495866 -7302 496102 -7066
rect 496186 -7302 496422 -7066
rect 495866 -7622 496102 -7386
rect 496186 -7622 496422 -7386
rect 505826 75218 506062 75454
rect 506146 75218 506382 75454
rect 505826 74898 506062 75134
rect 506146 74898 506382 75134
rect 505826 39218 506062 39454
rect 506146 39218 506382 39454
rect 505826 38898 506062 39134
rect 506146 38898 506382 39134
rect 505826 3218 506062 3454
rect 506146 3218 506382 3454
rect 505826 2898 506062 3134
rect 506146 2898 506382 3134
rect 505826 -582 506062 -346
rect 506146 -582 506382 -346
rect 505826 -902 506062 -666
rect 506146 -902 506382 -666
rect 509546 78938 509782 79174
rect 509866 78938 510102 79174
rect 509546 78618 509782 78854
rect 509866 78618 510102 78854
rect 509546 42938 509782 43174
rect 509866 42938 510102 43174
rect 509546 42618 509782 42854
rect 509866 42618 510102 42854
rect 509546 6938 509782 7174
rect 509866 6938 510102 7174
rect 509546 6618 509782 6854
rect 509866 6618 510102 6854
rect 509546 -1542 509782 -1306
rect 509866 -1542 510102 -1306
rect 509546 -1862 509782 -1626
rect 509866 -1862 510102 -1626
rect 513266 46658 513502 46894
rect 513586 46658 513822 46894
rect 513266 46338 513502 46574
rect 513586 46338 513822 46574
rect 513266 10658 513502 10894
rect 513586 10658 513822 10894
rect 513266 10338 513502 10574
rect 513586 10338 513822 10574
rect 513266 -2502 513502 -2266
rect 513586 -2502 513822 -2266
rect 513266 -2822 513502 -2586
rect 513586 -2822 513822 -2586
rect 516986 50378 517222 50614
rect 517306 50378 517542 50614
rect 516986 50058 517222 50294
rect 517306 50058 517542 50294
rect 516986 14378 517222 14614
rect 517306 14378 517542 14614
rect 516986 14058 517222 14294
rect 517306 14058 517542 14294
rect 516986 -3462 517222 -3226
rect 517306 -3462 517542 -3226
rect 516986 -3782 517222 -3546
rect 517306 -3782 517542 -3546
rect 520706 54098 520942 54334
rect 521026 54098 521262 54334
rect 520706 53778 520942 54014
rect 521026 53778 521262 54014
rect 520706 18098 520942 18334
rect 521026 18098 521262 18334
rect 520706 17778 520942 18014
rect 521026 17778 521262 18014
rect 520706 -4422 520942 -4186
rect 521026 -4422 521262 -4186
rect 520706 -4742 520942 -4506
rect 521026 -4742 521262 -4506
rect 524426 57818 524662 58054
rect 524746 57818 524982 58054
rect 524426 57498 524662 57734
rect 524746 57498 524982 57734
rect 524426 21818 524662 22054
rect 524746 21818 524982 22054
rect 524426 21498 524662 21734
rect 524746 21498 524982 21734
rect 524426 -5382 524662 -5146
rect 524746 -5382 524982 -5146
rect 524426 -5702 524662 -5466
rect 524746 -5702 524982 -5466
rect 528146 61538 528382 61774
rect 528466 61538 528702 61774
rect 528146 61218 528382 61454
rect 528466 61218 528702 61454
rect 528146 25538 528382 25774
rect 528466 25538 528702 25774
rect 528146 25218 528382 25454
rect 528466 25218 528702 25454
rect 528146 -6342 528382 -6106
rect 528466 -6342 528702 -6106
rect 528146 -6662 528382 -6426
rect 528466 -6662 528702 -6426
rect 531866 65258 532102 65494
rect 532186 65258 532422 65494
rect 531866 64938 532102 65174
rect 532186 64938 532422 65174
rect 531866 29258 532102 29494
rect 532186 29258 532422 29494
rect 531866 28938 532102 29174
rect 532186 28938 532422 29174
rect 531866 -7302 532102 -7066
rect 532186 -7302 532422 -7066
rect 531866 -7622 532102 -7386
rect 532186 -7622 532422 -7386
rect 541826 75218 542062 75454
rect 542146 75218 542382 75454
rect 541826 74898 542062 75134
rect 542146 74898 542382 75134
rect 546308 438938 546544 439174
rect 546308 438618 546544 438854
rect 545546 402938 545782 403174
rect 545866 402938 546102 403174
rect 545546 402618 545782 402854
rect 545866 402618 546102 402854
rect 545546 366938 545782 367174
rect 545866 366938 546102 367174
rect 545546 366618 545782 366854
rect 545866 366618 546102 366854
rect 545546 330938 545782 331174
rect 545866 330938 546102 331174
rect 545546 330618 545782 330854
rect 545866 330618 546102 330854
rect 545546 294938 545782 295174
rect 545866 294938 546102 295174
rect 545546 294618 545782 294854
rect 545866 294618 546102 294854
rect 545546 258938 545782 259174
rect 545866 258938 546102 259174
rect 545546 258618 545782 258854
rect 545866 258618 546102 258854
rect 545546 222938 545782 223174
rect 545866 222938 546102 223174
rect 545546 222618 545782 222854
rect 545866 222618 546102 222854
rect 545546 186938 545782 187174
rect 545866 186938 546102 187174
rect 545546 186618 545782 186854
rect 545866 186618 546102 186854
rect 545546 150938 545782 151174
rect 545866 150938 546102 151174
rect 545546 150618 545782 150854
rect 545866 150618 546102 150854
rect 545546 114938 545782 115174
rect 545866 114938 546102 115174
rect 545546 114618 545782 114854
rect 545866 114618 546102 114854
rect 545546 78938 545782 79174
rect 545866 78938 546102 79174
rect 545546 78618 545782 78854
rect 545866 78618 546102 78854
rect 552986 707482 553222 707718
rect 553306 707482 553542 707718
rect 552986 707162 553222 707398
rect 553306 707162 553542 707398
rect 552986 698378 553222 698614
rect 553306 698378 553542 698614
rect 552986 698058 553222 698294
rect 553306 698058 553542 698294
rect 552986 662378 553222 662614
rect 553306 662378 553542 662614
rect 552986 662058 553222 662294
rect 553306 662058 553542 662294
rect 552986 626378 553222 626614
rect 553306 626378 553542 626614
rect 552986 626058 553222 626294
rect 553306 626058 553542 626294
rect 552986 590378 553222 590614
rect 553306 590378 553542 590614
rect 552986 590058 553222 590294
rect 553306 590058 553542 590294
rect 552986 554378 553222 554614
rect 553306 554378 553542 554614
rect 552986 554058 553222 554294
rect 553306 554058 553542 554294
rect 552986 518378 553222 518614
rect 553306 518378 553542 518614
rect 552986 518058 553222 518294
rect 553306 518058 553542 518294
rect 552986 482378 553222 482614
rect 553306 482378 553542 482614
rect 552986 482058 553222 482294
rect 553306 482058 553542 482294
rect 552986 446378 553222 446614
rect 553306 446378 553542 446614
rect 552986 446058 553222 446294
rect 553306 446058 553542 446294
rect 550529 435218 550765 435454
rect 550529 434898 550765 435134
rect 549266 406658 549502 406894
rect 549586 406658 549822 406894
rect 549266 406338 549502 406574
rect 549586 406338 549822 406574
rect 556706 708442 556942 708678
rect 557026 708442 557262 708678
rect 556706 708122 556942 708358
rect 557026 708122 557262 708358
rect 560426 709402 560662 709638
rect 560746 709402 560982 709638
rect 560426 709082 560662 709318
rect 560746 709082 560982 709318
rect 556706 666098 556942 666334
rect 557026 666098 557262 666334
rect 556706 665778 556942 666014
rect 557026 665778 557262 666014
rect 556706 630098 556942 630334
rect 557026 630098 557262 630334
rect 556706 629778 556942 630014
rect 557026 629778 557262 630014
rect 556706 594098 556942 594334
rect 557026 594098 557262 594334
rect 556706 593778 556942 594014
rect 557026 593778 557262 594014
rect 556706 558098 556942 558334
rect 557026 558098 557262 558334
rect 556706 557778 556942 558014
rect 557026 557778 557262 558014
rect 556706 522098 556942 522334
rect 557026 522098 557262 522334
rect 556706 521778 556942 522014
rect 557026 521778 557262 522014
rect 556706 486098 556942 486334
rect 557026 486098 557262 486334
rect 556706 485778 556942 486014
rect 557026 485778 557262 486014
rect 556706 450098 556942 450334
rect 557026 450098 557262 450334
rect 556706 449778 556942 450014
rect 557026 449778 557262 450014
rect 554749 438938 554985 439174
rect 554749 438618 554985 438854
rect 552986 410378 553222 410614
rect 553306 410378 553542 410614
rect 552986 410058 553222 410294
rect 553306 410058 553542 410294
rect 556706 414098 556942 414334
rect 557026 414098 557262 414334
rect 556706 413778 556942 414014
rect 557026 413778 557262 414014
rect 556706 378007 556942 378243
rect 557026 378007 557262 378243
rect 549266 370658 549502 370894
rect 549586 370658 549822 370894
rect 549266 370338 549502 370574
rect 549586 370338 549822 370574
rect 554918 366938 555154 367174
rect 554918 366618 555154 366854
rect 552952 363218 553188 363454
rect 552952 362898 553188 363134
rect 556885 363218 557121 363454
rect 556885 362898 557121 363134
rect 549266 334658 549502 334894
rect 549586 334658 549822 334894
rect 549266 334338 549502 334574
rect 549586 334338 549822 334574
rect 549266 298658 549502 298894
rect 549586 298658 549822 298894
rect 549266 298338 549502 298574
rect 549586 298338 549822 298574
rect 549266 262658 549502 262894
rect 549586 262658 549822 262894
rect 549266 262338 549502 262574
rect 549586 262338 549822 262574
rect 549266 226658 549502 226894
rect 549586 226658 549822 226894
rect 549266 226338 549502 226574
rect 549586 226338 549822 226574
rect 549266 190658 549502 190894
rect 549586 190658 549822 190894
rect 549266 190338 549502 190574
rect 549586 190338 549822 190574
rect 549266 154658 549502 154894
rect 549586 154658 549822 154894
rect 549266 154338 549502 154574
rect 549586 154338 549822 154574
rect 549266 118658 549502 118894
rect 549586 118658 549822 118894
rect 549266 118338 549502 118574
rect 549586 118338 549822 118574
rect 549266 82658 549502 82894
rect 549586 82658 549822 82894
rect 549266 82338 549502 82574
rect 549586 82338 549822 82574
rect 552986 338378 553222 338614
rect 553306 338378 553542 338614
rect 552986 338058 553222 338294
rect 553306 338058 553542 338294
rect 552986 302378 553222 302614
rect 553306 302378 553542 302614
rect 552986 302058 553222 302294
rect 553306 302058 553542 302294
rect 552986 266378 553222 266614
rect 553306 266378 553542 266614
rect 552986 266058 553222 266294
rect 553306 266058 553542 266294
rect 552986 230378 553222 230614
rect 553306 230378 553542 230614
rect 552986 230058 553222 230294
rect 553306 230058 553542 230294
rect 552986 194378 553222 194614
rect 553306 194378 553542 194614
rect 552986 194058 553222 194294
rect 553306 194058 553542 194294
rect 552986 158378 553222 158614
rect 553306 158378 553542 158614
rect 552986 158058 553222 158294
rect 553306 158058 553542 158294
rect 552986 122378 553222 122614
rect 553306 122378 553542 122614
rect 552986 122058 553222 122294
rect 553306 122058 553542 122294
rect 552986 86378 553222 86614
rect 553306 86378 553542 86614
rect 552986 86058 553222 86294
rect 553306 86058 553542 86294
rect 556706 342098 556942 342334
rect 557026 342098 557262 342334
rect 556706 341778 556942 342014
rect 557026 341778 557262 342014
rect 560426 669818 560662 670054
rect 560746 669818 560982 670054
rect 560426 669498 560662 669734
rect 560746 669498 560982 669734
rect 560426 633818 560662 634054
rect 560746 633818 560982 634054
rect 560426 633498 560662 633734
rect 560746 633498 560982 633734
rect 560426 597818 560662 598054
rect 560746 597818 560982 598054
rect 560426 597498 560662 597734
rect 560746 597498 560982 597734
rect 560426 561818 560662 562054
rect 560746 561818 560982 562054
rect 560426 561498 560662 561734
rect 560746 561498 560982 561734
rect 560426 525818 560662 526054
rect 560746 525818 560982 526054
rect 560426 525498 560662 525734
rect 560746 525498 560982 525734
rect 560426 489818 560662 490054
rect 560746 489818 560982 490054
rect 560426 489498 560662 489734
rect 560746 489498 560982 489734
rect 560426 453818 560662 454054
rect 560746 453818 560982 454054
rect 560426 453498 560662 453734
rect 560746 453498 560982 453734
rect 560426 417818 560662 418054
rect 560746 417818 560982 418054
rect 560426 417498 560662 417734
rect 560746 417498 560982 417734
rect 560426 381818 560662 382054
rect 560746 381818 560982 382054
rect 560426 381498 560662 381734
rect 560746 381498 560982 381734
rect 564146 710362 564382 710598
rect 564466 710362 564702 710598
rect 564146 710042 564382 710278
rect 564466 710042 564702 710278
rect 564146 673538 564382 673774
rect 564466 673538 564702 673774
rect 564146 673218 564382 673454
rect 564466 673218 564702 673454
rect 564146 637538 564382 637774
rect 564466 637538 564702 637774
rect 564146 637218 564382 637454
rect 564466 637218 564702 637454
rect 564146 601538 564382 601774
rect 564466 601538 564702 601774
rect 564146 601218 564382 601454
rect 564466 601218 564702 601454
rect 564146 565538 564382 565774
rect 564466 565538 564702 565774
rect 564146 565218 564382 565454
rect 564466 565218 564702 565454
rect 564146 529538 564382 529774
rect 564466 529538 564702 529774
rect 564146 529218 564382 529454
rect 564466 529218 564702 529454
rect 564146 493538 564382 493774
rect 564466 493538 564702 493774
rect 564146 493218 564382 493454
rect 564466 493218 564702 493454
rect 564146 457538 564382 457774
rect 564466 457538 564702 457774
rect 564146 457218 564382 457454
rect 564466 457218 564702 457454
rect 564146 421538 564382 421774
rect 564466 421538 564702 421774
rect 564146 421218 564382 421454
rect 564466 421218 564702 421454
rect 564146 385538 564382 385774
rect 564466 385538 564702 385774
rect 564146 385218 564382 385454
rect 564466 385218 564702 385454
rect 567866 711322 568102 711558
rect 568186 711322 568422 711558
rect 567866 711002 568102 711238
rect 568186 711002 568422 711238
rect 567866 677258 568102 677494
rect 568186 677258 568422 677494
rect 567866 676938 568102 677174
rect 568186 676938 568422 677174
rect 567866 641258 568102 641494
rect 568186 641258 568422 641494
rect 567866 640938 568102 641174
rect 568186 640938 568422 641174
rect 567866 605258 568102 605494
rect 568186 605258 568422 605494
rect 567866 604938 568102 605174
rect 568186 604938 568422 605174
rect 567866 569258 568102 569494
rect 568186 569258 568422 569494
rect 567866 568938 568102 569174
rect 568186 568938 568422 569174
rect 567866 533258 568102 533494
rect 568186 533258 568422 533494
rect 567866 532938 568102 533174
rect 568186 532938 568422 533174
rect 567866 497258 568102 497494
rect 568186 497258 568422 497494
rect 567866 496938 568102 497174
rect 568186 496938 568422 497174
rect 567866 461258 568102 461494
rect 568186 461258 568422 461494
rect 567866 460938 568102 461174
rect 568186 460938 568422 461174
rect 567866 425258 568102 425494
rect 568186 425258 568422 425494
rect 567866 424938 568102 425174
rect 568186 424938 568422 425174
rect 567866 389258 568102 389494
rect 568186 389258 568422 389494
rect 567866 388938 568102 389174
rect 568186 388938 568422 389174
rect 558851 366938 559087 367174
rect 558851 366618 559087 366854
rect 562784 366938 563020 367174
rect 562784 366618 563020 366854
rect 566717 366938 566953 367174
rect 566717 366618 566953 366854
rect 560818 363218 561054 363454
rect 560818 362898 561054 363134
rect 564751 363218 564987 363454
rect 564751 362898 564987 363134
rect 560426 345818 560662 346054
rect 560746 345818 560982 346054
rect 560426 345498 560662 345734
rect 560746 345498 560982 345734
rect 556706 306098 556942 306334
rect 557026 306098 557262 306334
rect 556706 305778 556942 306014
rect 557026 305778 557262 306014
rect 556706 270098 556942 270334
rect 557026 270098 557262 270334
rect 556706 269778 556942 270014
rect 557026 269778 557262 270014
rect 556706 234098 556942 234334
rect 557026 234098 557262 234334
rect 556706 233778 556942 234014
rect 557026 233778 557262 234014
rect 556706 198098 556942 198334
rect 557026 198098 557262 198334
rect 556706 197778 556942 198014
rect 557026 197778 557262 198014
rect 556706 162098 556942 162334
rect 557026 162098 557262 162334
rect 556706 161778 556942 162014
rect 557026 161778 557262 162014
rect 556706 126098 556942 126334
rect 557026 126098 557262 126334
rect 556706 125778 556942 126014
rect 557026 125778 557262 126014
rect 556706 90098 556942 90334
rect 557026 90098 557262 90334
rect 556706 89778 556942 90014
rect 557026 89778 557262 90014
rect 556706 54098 556942 54334
rect 557026 54098 557262 54334
rect 556706 53778 556942 54014
rect 557026 53778 557262 54014
rect 549266 46658 549502 46894
rect 549586 46658 549822 46894
rect 549266 46338 549502 46574
rect 549586 46338 549822 46574
rect 545930 42938 546166 43174
rect 545930 42618 546166 42854
rect 541826 39218 542062 39454
rect 542146 39218 542382 39454
rect 541826 38898 542062 39134
rect 542146 38898 542382 39134
rect 543458 39218 543694 39454
rect 543458 38898 543694 39134
rect 548403 39218 548639 39454
rect 548403 38898 548639 39134
rect 541826 3218 542062 3454
rect 542146 3218 542382 3454
rect 541826 2898 542062 3134
rect 542146 2898 542382 3134
rect 541826 -582 542062 -346
rect 542146 -582 542382 -346
rect 541826 -902 542062 -666
rect 542146 -902 542382 -666
rect 545546 6938 545782 7174
rect 545866 6938 546102 7174
rect 545546 6618 545782 6854
rect 545866 6618 546102 6854
rect 545546 -1542 545782 -1306
rect 545866 -1542 546102 -1306
rect 545546 -1862 545782 -1626
rect 545866 -1862 546102 -1626
rect 550875 42938 551111 43174
rect 550875 42618 551111 42854
rect 555820 42938 556056 43174
rect 555820 42618 556056 42854
rect 553348 39218 553584 39454
rect 553348 38898 553584 39134
rect 549266 10658 549502 10894
rect 549586 10658 549822 10894
rect 549266 10338 549502 10574
rect 549586 10338 549822 10574
rect 549266 -2502 549502 -2266
rect 549586 -2502 549822 -2266
rect 549266 -2822 549502 -2586
rect 549586 -2822 549822 -2586
rect 552986 14378 553222 14614
rect 553306 14378 553542 14614
rect 552986 14058 553222 14294
rect 553306 14058 553542 14294
rect 552986 -3462 553222 -3226
rect 553306 -3462 553542 -3226
rect 552986 -3782 553222 -3546
rect 553306 -3782 553542 -3546
rect 560426 309818 560662 310054
rect 560746 309818 560982 310054
rect 560426 309498 560662 309734
rect 560746 309498 560982 309734
rect 560426 273818 560662 274054
rect 560746 273818 560982 274054
rect 560426 273498 560662 273734
rect 560746 273498 560982 273734
rect 560426 237818 560662 238054
rect 560746 237818 560982 238054
rect 560426 237498 560662 237734
rect 560746 237498 560982 237734
rect 560426 201818 560662 202054
rect 560746 201818 560982 202054
rect 560426 201498 560662 201734
rect 560746 201498 560982 201734
rect 560426 165818 560662 166054
rect 560746 165818 560982 166054
rect 560426 165498 560662 165734
rect 560746 165498 560982 165734
rect 560426 129818 560662 130054
rect 560746 129818 560982 130054
rect 560426 129498 560662 129734
rect 560746 129498 560982 129734
rect 560426 93818 560662 94054
rect 560746 93818 560982 94054
rect 560426 93498 560662 93734
rect 560746 93498 560982 93734
rect 560426 57818 560662 58054
rect 560746 57818 560982 58054
rect 560426 57498 560662 57734
rect 560746 57498 560982 57734
rect 564146 349538 564382 349774
rect 564466 349538 564702 349774
rect 564146 349218 564382 349454
rect 564466 349218 564702 349454
rect 564146 313538 564382 313774
rect 564466 313538 564702 313774
rect 564146 313218 564382 313454
rect 564466 313218 564702 313454
rect 564146 277538 564382 277774
rect 564466 277538 564702 277774
rect 564146 277218 564382 277454
rect 564466 277218 564702 277454
rect 564146 241538 564382 241774
rect 564466 241538 564702 241774
rect 564146 241218 564382 241454
rect 564466 241218 564702 241454
rect 564146 205538 564382 205774
rect 564466 205538 564702 205774
rect 564146 205218 564382 205454
rect 564466 205218 564702 205454
rect 564146 169538 564382 169774
rect 564466 169538 564702 169774
rect 564146 169218 564382 169454
rect 564466 169218 564702 169454
rect 564146 133538 564382 133774
rect 564466 133538 564702 133774
rect 564146 133218 564382 133454
rect 564466 133218 564702 133454
rect 564146 97538 564382 97774
rect 564466 97538 564702 97774
rect 564146 97218 564382 97454
rect 564466 97218 564702 97454
rect 564146 61538 564382 61774
rect 564466 61538 564702 61774
rect 564146 61218 564382 61454
rect 564466 61218 564702 61454
rect 560765 42938 561001 43174
rect 560765 42618 561001 42854
rect 558293 39218 558529 39454
rect 558293 38898 558529 39134
rect 556706 18098 556942 18334
rect 557026 18098 557262 18334
rect 556706 17778 556942 18014
rect 557026 17778 557262 18014
rect 556706 -4422 556942 -4186
rect 557026 -4422 557262 -4186
rect 556706 -4742 556942 -4506
rect 557026 -4742 557262 -4506
rect 560426 21818 560662 22054
rect 560746 21818 560982 22054
rect 560426 21498 560662 21734
rect 560746 21498 560982 21734
rect 560426 -5382 560662 -5146
rect 560746 -5382 560982 -5146
rect 560426 -5702 560662 -5466
rect 560746 -5702 560982 -5466
rect 564146 25538 564382 25774
rect 564466 25538 564702 25774
rect 564146 25218 564382 25454
rect 564466 25218 564702 25454
rect 564146 -6342 564382 -6106
rect 564466 -6342 564702 -6106
rect 564146 -6662 564382 -6426
rect 564466 -6662 564702 -6426
rect 567866 353258 568102 353494
rect 568186 353258 568422 353494
rect 567866 352938 568102 353174
rect 568186 352938 568422 353174
rect 567866 317258 568102 317494
rect 568186 317258 568422 317494
rect 567866 316938 568102 317174
rect 568186 316938 568422 317174
rect 567866 281258 568102 281494
rect 568186 281258 568422 281494
rect 567866 280938 568102 281174
rect 568186 280938 568422 281174
rect 567866 245258 568102 245494
rect 568186 245258 568422 245494
rect 567866 244938 568102 245174
rect 568186 244938 568422 245174
rect 567866 209258 568102 209494
rect 568186 209258 568422 209494
rect 567866 208938 568102 209174
rect 568186 208938 568422 209174
rect 567866 173258 568102 173494
rect 568186 173258 568422 173494
rect 567866 172938 568102 173174
rect 568186 172938 568422 173174
rect 567866 137258 568102 137494
rect 568186 137258 568422 137494
rect 567866 136938 568102 137174
rect 568186 136938 568422 137174
rect 567866 101258 568102 101494
rect 568186 101258 568422 101494
rect 567866 100938 568102 101174
rect 568186 100938 568422 101174
rect 567866 65258 568102 65494
rect 568186 65258 568422 65494
rect 567866 64938 568102 65174
rect 568186 64938 568422 65174
rect 567866 29258 568102 29494
rect 568186 29258 568422 29494
rect 567866 28938 568102 29174
rect 568186 28938 568422 29174
rect 567866 -7302 568102 -7066
rect 568186 -7302 568422 -7066
rect 567866 -7622 568102 -7386
rect 568186 -7622 568422 -7386
rect 577826 704602 578062 704838
rect 578146 704602 578382 704838
rect 577826 704282 578062 704518
rect 578146 704282 578382 704518
rect 577826 687218 578062 687454
rect 578146 687218 578382 687454
rect 577826 686898 578062 687134
rect 578146 686898 578382 687134
rect 577826 651218 578062 651454
rect 578146 651218 578382 651454
rect 577826 650898 578062 651134
rect 578146 650898 578382 651134
rect 577826 615218 578062 615454
rect 578146 615218 578382 615454
rect 577826 614898 578062 615134
rect 578146 614898 578382 615134
rect 577826 579218 578062 579454
rect 578146 579218 578382 579454
rect 577826 578898 578062 579134
rect 578146 578898 578382 579134
rect 577826 543218 578062 543454
rect 578146 543218 578382 543454
rect 577826 542898 578062 543134
rect 578146 542898 578382 543134
rect 577826 507218 578062 507454
rect 578146 507218 578382 507454
rect 577826 506898 578062 507134
rect 578146 506898 578382 507134
rect 577826 471218 578062 471454
rect 578146 471218 578382 471454
rect 577826 470898 578062 471134
rect 578146 470898 578382 471134
rect 577826 435218 578062 435454
rect 578146 435218 578382 435454
rect 577826 434898 578062 435134
rect 578146 434898 578382 435134
rect 577826 399218 578062 399454
rect 578146 399218 578382 399454
rect 577826 398898 578062 399134
rect 578146 398898 578382 399134
rect 577826 363218 578062 363454
rect 578146 363218 578382 363454
rect 577826 362898 578062 363134
rect 578146 362898 578382 363134
rect 577826 327218 578062 327454
rect 578146 327218 578382 327454
rect 577826 326898 578062 327134
rect 578146 326898 578382 327134
rect 577826 291218 578062 291454
rect 578146 291218 578382 291454
rect 577826 290898 578062 291134
rect 578146 290898 578382 291134
rect 577826 255218 578062 255454
rect 578146 255218 578382 255454
rect 577826 254898 578062 255134
rect 578146 254898 578382 255134
rect 577826 219218 578062 219454
rect 578146 219218 578382 219454
rect 577826 218898 578062 219134
rect 578146 218898 578382 219134
rect 577826 183218 578062 183454
rect 578146 183218 578382 183454
rect 577826 182898 578062 183134
rect 578146 182898 578382 183134
rect 577826 147218 578062 147454
rect 578146 147218 578382 147454
rect 577826 146898 578062 147134
rect 578146 146898 578382 147134
rect 577826 111218 578062 111454
rect 578146 111218 578382 111454
rect 577826 110898 578062 111134
rect 578146 110898 578382 111134
rect 577826 75218 578062 75454
rect 578146 75218 578382 75454
rect 577826 74898 578062 75134
rect 578146 74898 578382 75134
rect 577826 39218 578062 39454
rect 578146 39218 578382 39454
rect 577826 38898 578062 39134
rect 578146 38898 578382 39134
rect 577826 3218 578062 3454
rect 578146 3218 578382 3454
rect 577826 2898 578062 3134
rect 578146 2898 578382 3134
rect 577826 -582 578062 -346
rect 578146 -582 578382 -346
rect 577826 -902 578062 -666
rect 578146 -902 578382 -666
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 581546 705562 581782 705798
rect 581866 705562 582102 705798
rect 581546 705242 581782 705478
rect 581866 705242 582102 705478
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 581546 690938 581782 691174
rect 581866 690938 582102 691174
rect 581546 690618 581782 690854
rect 581866 690618 582102 690854
rect 581546 654938 581782 655174
rect 581866 654938 582102 655174
rect 581546 654618 581782 654854
rect 581866 654618 582102 654854
rect 581546 618938 581782 619174
rect 581866 618938 582102 619174
rect 581546 618618 581782 618854
rect 581866 618618 582102 618854
rect 581546 582938 581782 583174
rect 581866 582938 582102 583174
rect 581546 582618 581782 582854
rect 581866 582618 582102 582854
rect 581546 546938 581782 547174
rect 581866 546938 582102 547174
rect 581546 546618 581782 546854
rect 581866 546618 582102 546854
rect 581546 510938 581782 511174
rect 581866 510938 582102 511174
rect 581546 510618 581782 510854
rect 581866 510618 582102 510854
rect 581546 474938 581782 475174
rect 581866 474938 582102 475174
rect 581546 474618 581782 474854
rect 581866 474618 582102 474854
rect 581546 438938 581782 439174
rect 581866 438938 582102 439174
rect 581546 438618 581782 438854
rect 581866 438618 582102 438854
rect 581546 402938 581782 403174
rect 581866 402938 582102 403174
rect 581546 402618 581782 402854
rect 581866 402618 582102 402854
rect 581546 366938 581782 367174
rect 581866 366938 582102 367174
rect 581546 366618 581782 366854
rect 581866 366618 582102 366854
rect 581546 330938 581782 331174
rect 581866 330938 582102 331174
rect 581546 330618 581782 330854
rect 581866 330618 582102 330854
rect 581546 294938 581782 295174
rect 581866 294938 582102 295174
rect 581546 294618 581782 294854
rect 581866 294618 582102 294854
rect 581546 258938 581782 259174
rect 581866 258938 582102 259174
rect 581546 258618 581782 258854
rect 581866 258618 582102 258854
rect 581546 222938 581782 223174
rect 581866 222938 582102 223174
rect 581546 222618 581782 222854
rect 581866 222618 582102 222854
rect 581546 186938 581782 187174
rect 581866 186938 582102 187174
rect 581546 186618 581782 186854
rect 581866 186618 582102 186854
rect 581546 150938 581782 151174
rect 581866 150938 582102 151174
rect 581546 150618 581782 150854
rect 581866 150618 582102 150854
rect 581546 114938 581782 115174
rect 581866 114938 582102 115174
rect 581546 114618 581782 114854
rect 581866 114618 582102 114854
rect 581546 78938 581782 79174
rect 581866 78938 582102 79174
rect 581546 78618 581782 78854
rect 581866 78618 582102 78854
rect 581546 42938 581782 43174
rect 581866 42938 582102 43174
rect 581546 42618 581782 42854
rect 581866 42618 582102 42854
rect 581546 6938 581782 7174
rect 581866 6938 582102 7174
rect 581546 6618 581782 6854
rect 581866 6618 582102 6854
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 687218 585578 687454
rect 585662 687218 585898 687454
rect 585342 686898 585578 687134
rect 585662 686898 585898 687134
rect 585342 651218 585578 651454
rect 585662 651218 585898 651454
rect 585342 650898 585578 651134
rect 585662 650898 585898 651134
rect 585342 615218 585578 615454
rect 585662 615218 585898 615454
rect 585342 614898 585578 615134
rect 585662 614898 585898 615134
rect 585342 579218 585578 579454
rect 585662 579218 585898 579454
rect 585342 578898 585578 579134
rect 585662 578898 585898 579134
rect 585342 543218 585578 543454
rect 585662 543218 585898 543454
rect 585342 542898 585578 543134
rect 585662 542898 585898 543134
rect 585342 507218 585578 507454
rect 585662 507218 585898 507454
rect 585342 506898 585578 507134
rect 585662 506898 585898 507134
rect 585342 471218 585578 471454
rect 585662 471218 585898 471454
rect 585342 470898 585578 471134
rect 585662 470898 585898 471134
rect 585342 435218 585578 435454
rect 585662 435218 585898 435454
rect 585342 434898 585578 435134
rect 585662 434898 585898 435134
rect 585342 399218 585578 399454
rect 585662 399218 585898 399454
rect 585342 398898 585578 399134
rect 585662 398898 585898 399134
rect 585342 363218 585578 363454
rect 585662 363218 585898 363454
rect 585342 362898 585578 363134
rect 585662 362898 585898 363134
rect 585342 327218 585578 327454
rect 585662 327218 585898 327454
rect 585342 326898 585578 327134
rect 585662 326898 585898 327134
rect 585342 291218 585578 291454
rect 585662 291218 585898 291454
rect 585342 290898 585578 291134
rect 585662 290898 585898 291134
rect 585342 255218 585578 255454
rect 585662 255218 585898 255454
rect 585342 254898 585578 255134
rect 585662 254898 585898 255134
rect 585342 219218 585578 219454
rect 585662 219218 585898 219454
rect 585342 218898 585578 219134
rect 585662 218898 585898 219134
rect 585342 183218 585578 183454
rect 585662 183218 585898 183454
rect 585342 182898 585578 183134
rect 585662 182898 585898 183134
rect 585342 147218 585578 147454
rect 585662 147218 585898 147454
rect 585342 146898 585578 147134
rect 585662 146898 585898 147134
rect 585342 111218 585578 111454
rect 585662 111218 585898 111454
rect 585342 110898 585578 111134
rect 585662 110898 585898 111134
rect 585342 75218 585578 75454
rect 585662 75218 585898 75454
rect 585342 74898 585578 75134
rect 585662 74898 585898 75134
rect 585342 39218 585578 39454
rect 585662 39218 585898 39454
rect 585342 38898 585578 39134
rect 585662 38898 585898 39134
rect 585342 3218 585578 3454
rect 585662 3218 585898 3454
rect 585342 2898 585578 3134
rect 585662 2898 585898 3134
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 690938 586538 691174
rect 586622 690938 586858 691174
rect 586302 690618 586538 690854
rect 586622 690618 586858 690854
rect 586302 654938 586538 655174
rect 586622 654938 586858 655174
rect 586302 654618 586538 654854
rect 586622 654618 586858 654854
rect 586302 618938 586538 619174
rect 586622 618938 586858 619174
rect 586302 618618 586538 618854
rect 586622 618618 586858 618854
rect 586302 582938 586538 583174
rect 586622 582938 586858 583174
rect 586302 582618 586538 582854
rect 586622 582618 586858 582854
rect 586302 546938 586538 547174
rect 586622 546938 586858 547174
rect 586302 546618 586538 546854
rect 586622 546618 586858 546854
rect 586302 510938 586538 511174
rect 586622 510938 586858 511174
rect 586302 510618 586538 510854
rect 586622 510618 586858 510854
rect 586302 474938 586538 475174
rect 586622 474938 586858 475174
rect 586302 474618 586538 474854
rect 586622 474618 586858 474854
rect 586302 438938 586538 439174
rect 586622 438938 586858 439174
rect 586302 438618 586538 438854
rect 586622 438618 586858 438854
rect 586302 402938 586538 403174
rect 586622 402938 586858 403174
rect 586302 402618 586538 402854
rect 586622 402618 586858 402854
rect 586302 366938 586538 367174
rect 586622 366938 586858 367174
rect 586302 366618 586538 366854
rect 586622 366618 586858 366854
rect 586302 330938 586538 331174
rect 586622 330938 586858 331174
rect 586302 330618 586538 330854
rect 586622 330618 586858 330854
rect 586302 294938 586538 295174
rect 586622 294938 586858 295174
rect 586302 294618 586538 294854
rect 586622 294618 586858 294854
rect 586302 258938 586538 259174
rect 586622 258938 586858 259174
rect 586302 258618 586538 258854
rect 586622 258618 586858 258854
rect 586302 222938 586538 223174
rect 586622 222938 586858 223174
rect 586302 222618 586538 222854
rect 586622 222618 586858 222854
rect 586302 186938 586538 187174
rect 586622 186938 586858 187174
rect 586302 186618 586538 186854
rect 586622 186618 586858 186854
rect 586302 150938 586538 151174
rect 586622 150938 586858 151174
rect 586302 150618 586538 150854
rect 586622 150618 586858 150854
rect 586302 114938 586538 115174
rect 586622 114938 586858 115174
rect 586302 114618 586538 114854
rect 586622 114618 586858 114854
rect 586302 78938 586538 79174
rect 586622 78938 586858 79174
rect 586302 78618 586538 78854
rect 586622 78618 586858 78854
rect 586302 42938 586538 43174
rect 586622 42938 586858 43174
rect 586302 42618 586538 42854
rect 586622 42618 586858 42854
rect 586302 6938 586538 7174
rect 586622 6938 586858 7174
rect 586302 6618 586538 6854
rect 586622 6618 586858 6854
rect 581546 -1542 581782 -1306
rect 581866 -1542 582102 -1306
rect 581546 -1862 581782 -1626
rect 581866 -1862 582102 -1626
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 694658 587498 694894
rect 587582 694658 587818 694894
rect 587262 694338 587498 694574
rect 587582 694338 587818 694574
rect 587262 658658 587498 658894
rect 587582 658658 587818 658894
rect 587262 658338 587498 658574
rect 587582 658338 587818 658574
rect 587262 622658 587498 622894
rect 587582 622658 587818 622894
rect 587262 622338 587498 622574
rect 587582 622338 587818 622574
rect 587262 586658 587498 586894
rect 587582 586658 587818 586894
rect 587262 586338 587498 586574
rect 587582 586338 587818 586574
rect 587262 550658 587498 550894
rect 587582 550658 587818 550894
rect 587262 550338 587498 550574
rect 587582 550338 587818 550574
rect 587262 514658 587498 514894
rect 587582 514658 587818 514894
rect 587262 514338 587498 514574
rect 587582 514338 587818 514574
rect 587262 478658 587498 478894
rect 587582 478658 587818 478894
rect 587262 478338 587498 478574
rect 587582 478338 587818 478574
rect 587262 442658 587498 442894
rect 587582 442658 587818 442894
rect 587262 442338 587498 442574
rect 587582 442338 587818 442574
rect 587262 406658 587498 406894
rect 587582 406658 587818 406894
rect 587262 406338 587498 406574
rect 587582 406338 587818 406574
rect 587262 370658 587498 370894
rect 587582 370658 587818 370894
rect 587262 370338 587498 370574
rect 587582 370338 587818 370574
rect 587262 334658 587498 334894
rect 587582 334658 587818 334894
rect 587262 334338 587498 334574
rect 587582 334338 587818 334574
rect 587262 298658 587498 298894
rect 587582 298658 587818 298894
rect 587262 298338 587498 298574
rect 587582 298338 587818 298574
rect 587262 262658 587498 262894
rect 587582 262658 587818 262894
rect 587262 262338 587498 262574
rect 587582 262338 587818 262574
rect 587262 226658 587498 226894
rect 587582 226658 587818 226894
rect 587262 226338 587498 226574
rect 587582 226338 587818 226574
rect 587262 190658 587498 190894
rect 587582 190658 587818 190894
rect 587262 190338 587498 190574
rect 587582 190338 587818 190574
rect 587262 154658 587498 154894
rect 587582 154658 587818 154894
rect 587262 154338 587498 154574
rect 587582 154338 587818 154574
rect 587262 118658 587498 118894
rect 587582 118658 587818 118894
rect 587262 118338 587498 118574
rect 587582 118338 587818 118574
rect 587262 82658 587498 82894
rect 587582 82658 587818 82894
rect 587262 82338 587498 82574
rect 587582 82338 587818 82574
rect 587262 46658 587498 46894
rect 587582 46658 587818 46894
rect 587262 46338 587498 46574
rect 587582 46338 587818 46574
rect 587262 10658 587498 10894
rect 587582 10658 587818 10894
rect 587262 10338 587498 10574
rect 587582 10338 587818 10574
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 698378 588458 698614
rect 588542 698378 588778 698614
rect 588222 698058 588458 698294
rect 588542 698058 588778 698294
rect 588222 662378 588458 662614
rect 588542 662378 588778 662614
rect 588222 662058 588458 662294
rect 588542 662058 588778 662294
rect 588222 626378 588458 626614
rect 588542 626378 588778 626614
rect 588222 626058 588458 626294
rect 588542 626058 588778 626294
rect 588222 590378 588458 590614
rect 588542 590378 588778 590614
rect 588222 590058 588458 590294
rect 588542 590058 588778 590294
rect 588222 554378 588458 554614
rect 588542 554378 588778 554614
rect 588222 554058 588458 554294
rect 588542 554058 588778 554294
rect 588222 518378 588458 518614
rect 588542 518378 588778 518614
rect 588222 518058 588458 518294
rect 588542 518058 588778 518294
rect 588222 482378 588458 482614
rect 588542 482378 588778 482614
rect 588222 482058 588458 482294
rect 588542 482058 588778 482294
rect 588222 446378 588458 446614
rect 588542 446378 588778 446614
rect 588222 446058 588458 446294
rect 588542 446058 588778 446294
rect 588222 410378 588458 410614
rect 588542 410378 588778 410614
rect 588222 410058 588458 410294
rect 588542 410058 588778 410294
rect 588222 374378 588458 374614
rect 588542 374378 588778 374614
rect 588222 374058 588458 374294
rect 588542 374058 588778 374294
rect 588222 338378 588458 338614
rect 588542 338378 588778 338614
rect 588222 338058 588458 338294
rect 588542 338058 588778 338294
rect 588222 302378 588458 302614
rect 588542 302378 588778 302614
rect 588222 302058 588458 302294
rect 588542 302058 588778 302294
rect 588222 266378 588458 266614
rect 588542 266378 588778 266614
rect 588222 266058 588458 266294
rect 588542 266058 588778 266294
rect 588222 230378 588458 230614
rect 588542 230378 588778 230614
rect 588222 230058 588458 230294
rect 588542 230058 588778 230294
rect 588222 194378 588458 194614
rect 588542 194378 588778 194614
rect 588222 194058 588458 194294
rect 588542 194058 588778 194294
rect 588222 158378 588458 158614
rect 588542 158378 588778 158614
rect 588222 158058 588458 158294
rect 588542 158058 588778 158294
rect 588222 122378 588458 122614
rect 588542 122378 588778 122614
rect 588222 122058 588458 122294
rect 588542 122058 588778 122294
rect 588222 86378 588458 86614
rect 588542 86378 588778 86614
rect 588222 86058 588458 86294
rect 588542 86058 588778 86294
rect 588222 50378 588458 50614
rect 588542 50378 588778 50614
rect 588222 50058 588458 50294
rect 588542 50058 588778 50294
rect 588222 14378 588458 14614
rect 588542 14378 588778 14614
rect 588222 14058 588458 14294
rect 588542 14058 588778 14294
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 666098 589418 666334
rect 589502 666098 589738 666334
rect 589182 665778 589418 666014
rect 589502 665778 589738 666014
rect 589182 630098 589418 630334
rect 589502 630098 589738 630334
rect 589182 629778 589418 630014
rect 589502 629778 589738 630014
rect 589182 594098 589418 594334
rect 589502 594098 589738 594334
rect 589182 593778 589418 594014
rect 589502 593778 589738 594014
rect 589182 558098 589418 558334
rect 589502 558098 589738 558334
rect 589182 557778 589418 558014
rect 589502 557778 589738 558014
rect 589182 522098 589418 522334
rect 589502 522098 589738 522334
rect 589182 521778 589418 522014
rect 589502 521778 589738 522014
rect 589182 486098 589418 486334
rect 589502 486098 589738 486334
rect 589182 485778 589418 486014
rect 589502 485778 589738 486014
rect 589182 450098 589418 450334
rect 589502 450098 589738 450334
rect 589182 449778 589418 450014
rect 589502 449778 589738 450014
rect 589182 414098 589418 414334
rect 589502 414098 589738 414334
rect 589182 413778 589418 414014
rect 589502 413778 589738 414014
rect 589182 378098 589418 378334
rect 589502 378098 589738 378334
rect 589182 377778 589418 378014
rect 589502 377778 589738 378014
rect 589182 342098 589418 342334
rect 589502 342098 589738 342334
rect 589182 341778 589418 342014
rect 589502 341778 589738 342014
rect 589182 306098 589418 306334
rect 589502 306098 589738 306334
rect 589182 305778 589418 306014
rect 589502 305778 589738 306014
rect 589182 270098 589418 270334
rect 589502 270098 589738 270334
rect 589182 269778 589418 270014
rect 589502 269778 589738 270014
rect 589182 234098 589418 234334
rect 589502 234098 589738 234334
rect 589182 233778 589418 234014
rect 589502 233778 589738 234014
rect 589182 198098 589418 198334
rect 589502 198098 589738 198334
rect 589182 197778 589418 198014
rect 589502 197778 589738 198014
rect 589182 162098 589418 162334
rect 589502 162098 589738 162334
rect 589182 161778 589418 162014
rect 589502 161778 589738 162014
rect 589182 126098 589418 126334
rect 589502 126098 589738 126334
rect 589182 125778 589418 126014
rect 589502 125778 589738 126014
rect 589182 90098 589418 90334
rect 589502 90098 589738 90334
rect 589182 89778 589418 90014
rect 589502 89778 589738 90014
rect 589182 54098 589418 54334
rect 589502 54098 589738 54334
rect 589182 53778 589418 54014
rect 589502 53778 589738 54014
rect 589182 18098 589418 18334
rect 589502 18098 589738 18334
rect 589182 17778 589418 18014
rect 589502 17778 589738 18014
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 669818 590378 670054
rect 590462 669818 590698 670054
rect 590142 669498 590378 669734
rect 590462 669498 590698 669734
rect 590142 633818 590378 634054
rect 590462 633818 590698 634054
rect 590142 633498 590378 633734
rect 590462 633498 590698 633734
rect 590142 597818 590378 598054
rect 590462 597818 590698 598054
rect 590142 597498 590378 597734
rect 590462 597498 590698 597734
rect 590142 561818 590378 562054
rect 590462 561818 590698 562054
rect 590142 561498 590378 561734
rect 590462 561498 590698 561734
rect 590142 525818 590378 526054
rect 590462 525818 590698 526054
rect 590142 525498 590378 525734
rect 590462 525498 590698 525734
rect 590142 489818 590378 490054
rect 590462 489818 590698 490054
rect 590142 489498 590378 489734
rect 590462 489498 590698 489734
rect 590142 453818 590378 454054
rect 590462 453818 590698 454054
rect 590142 453498 590378 453734
rect 590462 453498 590698 453734
rect 590142 417818 590378 418054
rect 590462 417818 590698 418054
rect 590142 417498 590378 417734
rect 590462 417498 590698 417734
rect 590142 381818 590378 382054
rect 590462 381818 590698 382054
rect 590142 381498 590378 381734
rect 590462 381498 590698 381734
rect 590142 345818 590378 346054
rect 590462 345818 590698 346054
rect 590142 345498 590378 345734
rect 590462 345498 590698 345734
rect 590142 309818 590378 310054
rect 590462 309818 590698 310054
rect 590142 309498 590378 309734
rect 590462 309498 590698 309734
rect 590142 273818 590378 274054
rect 590462 273818 590698 274054
rect 590142 273498 590378 273734
rect 590462 273498 590698 273734
rect 590142 237818 590378 238054
rect 590462 237818 590698 238054
rect 590142 237498 590378 237734
rect 590462 237498 590698 237734
rect 590142 201818 590378 202054
rect 590462 201818 590698 202054
rect 590142 201498 590378 201734
rect 590462 201498 590698 201734
rect 590142 165818 590378 166054
rect 590462 165818 590698 166054
rect 590142 165498 590378 165734
rect 590462 165498 590698 165734
rect 590142 129818 590378 130054
rect 590462 129818 590698 130054
rect 590142 129498 590378 129734
rect 590462 129498 590698 129734
rect 590142 93818 590378 94054
rect 590462 93818 590698 94054
rect 590142 93498 590378 93734
rect 590462 93498 590698 93734
rect 590142 57818 590378 58054
rect 590462 57818 590698 58054
rect 590142 57498 590378 57734
rect 590462 57498 590698 57734
rect 590142 21818 590378 22054
rect 590462 21818 590698 22054
rect 590142 21498 590378 21734
rect 590462 21498 590698 21734
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 673538 591338 673774
rect 591422 673538 591658 673774
rect 591102 673218 591338 673454
rect 591422 673218 591658 673454
rect 591102 637538 591338 637774
rect 591422 637538 591658 637774
rect 591102 637218 591338 637454
rect 591422 637218 591658 637454
rect 591102 601538 591338 601774
rect 591422 601538 591658 601774
rect 591102 601218 591338 601454
rect 591422 601218 591658 601454
rect 591102 565538 591338 565774
rect 591422 565538 591658 565774
rect 591102 565218 591338 565454
rect 591422 565218 591658 565454
rect 591102 529538 591338 529774
rect 591422 529538 591658 529774
rect 591102 529218 591338 529454
rect 591422 529218 591658 529454
rect 591102 493538 591338 493774
rect 591422 493538 591658 493774
rect 591102 493218 591338 493454
rect 591422 493218 591658 493454
rect 591102 457538 591338 457774
rect 591422 457538 591658 457774
rect 591102 457218 591338 457454
rect 591422 457218 591658 457454
rect 591102 421538 591338 421774
rect 591422 421538 591658 421774
rect 591102 421218 591338 421454
rect 591422 421218 591658 421454
rect 591102 385538 591338 385774
rect 591422 385538 591658 385774
rect 591102 385218 591338 385454
rect 591422 385218 591658 385454
rect 591102 349538 591338 349774
rect 591422 349538 591658 349774
rect 591102 349218 591338 349454
rect 591422 349218 591658 349454
rect 591102 313538 591338 313774
rect 591422 313538 591658 313774
rect 591102 313218 591338 313454
rect 591422 313218 591658 313454
rect 591102 277538 591338 277774
rect 591422 277538 591658 277774
rect 591102 277218 591338 277454
rect 591422 277218 591658 277454
rect 591102 241538 591338 241774
rect 591422 241538 591658 241774
rect 591102 241218 591338 241454
rect 591422 241218 591658 241454
rect 591102 205538 591338 205774
rect 591422 205538 591658 205774
rect 591102 205218 591338 205454
rect 591422 205218 591658 205454
rect 591102 169538 591338 169774
rect 591422 169538 591658 169774
rect 591102 169218 591338 169454
rect 591422 169218 591658 169454
rect 591102 133538 591338 133774
rect 591422 133538 591658 133774
rect 591102 133218 591338 133454
rect 591422 133218 591658 133454
rect 591102 97538 591338 97774
rect 591422 97538 591658 97774
rect 591102 97218 591338 97454
rect 591422 97218 591658 97454
rect 591102 61538 591338 61774
rect 591422 61538 591658 61774
rect 591102 61218 591338 61454
rect 591422 61218 591658 61454
rect 591102 25538 591338 25774
rect 591422 25538 591658 25774
rect 591102 25218 591338 25454
rect 591422 25218 591658 25454
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 677258 592298 677494
rect 592382 677258 592618 677494
rect 592062 676938 592298 677174
rect 592382 676938 592618 677174
rect 592062 641258 592298 641494
rect 592382 641258 592618 641494
rect 592062 640938 592298 641174
rect 592382 640938 592618 641174
rect 592062 605258 592298 605494
rect 592382 605258 592618 605494
rect 592062 604938 592298 605174
rect 592382 604938 592618 605174
rect 592062 569258 592298 569494
rect 592382 569258 592618 569494
rect 592062 568938 592298 569174
rect 592382 568938 592618 569174
rect 592062 533258 592298 533494
rect 592382 533258 592618 533494
rect 592062 532938 592298 533174
rect 592382 532938 592618 533174
rect 592062 497258 592298 497494
rect 592382 497258 592618 497494
rect 592062 496938 592298 497174
rect 592382 496938 592618 497174
rect 592062 461258 592298 461494
rect 592382 461258 592618 461494
rect 592062 460938 592298 461174
rect 592382 460938 592618 461174
rect 592062 425258 592298 425494
rect 592382 425258 592618 425494
rect 592062 424938 592298 425174
rect 592382 424938 592618 425174
rect 592062 389258 592298 389494
rect 592382 389258 592618 389494
rect 592062 388938 592298 389174
rect 592382 388938 592618 389174
rect 592062 353258 592298 353494
rect 592382 353258 592618 353494
rect 592062 352938 592298 353174
rect 592382 352938 592618 353174
rect 592062 317258 592298 317494
rect 592382 317258 592618 317494
rect 592062 316938 592298 317174
rect 592382 316938 592618 317174
rect 592062 281258 592298 281494
rect 592382 281258 592618 281494
rect 592062 280938 592298 281174
rect 592382 280938 592618 281174
rect 592062 245258 592298 245494
rect 592382 245258 592618 245494
rect 592062 244938 592298 245174
rect 592382 244938 592618 245174
rect 592062 209258 592298 209494
rect 592382 209258 592618 209494
rect 592062 208938 592298 209174
rect 592382 208938 592618 209174
rect 592062 173258 592298 173494
rect 592382 173258 592618 173494
rect 592062 172938 592298 173174
rect 592382 172938 592618 173174
rect 592062 137258 592298 137494
rect 592382 137258 592618 137494
rect 592062 136938 592298 137174
rect 592382 136938 592618 137174
rect 592062 101258 592298 101494
rect 592382 101258 592618 101494
rect 592062 100938 592298 101174
rect 592382 100938 592618 101174
rect 592062 65258 592298 65494
rect 592382 65258 592618 65494
rect 592062 64938 592298 65174
rect 592382 64938 592618 65174
rect 592062 29258 592298 29494
rect 592382 29258 592618 29494
rect 592062 28938 592298 29174
rect 592382 28938 592618 29174
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 27866 711558
rect 28102 711322 28186 711558
rect 28422 711322 63866 711558
rect 64102 711322 64186 711558
rect 64422 711322 99866 711558
rect 100102 711322 100186 711558
rect 100422 711322 135866 711558
rect 136102 711322 136186 711558
rect 136422 711322 171866 711558
rect 172102 711322 172186 711558
rect 172422 711322 207866 711558
rect 208102 711322 208186 711558
rect 208422 711322 243866 711558
rect 244102 711322 244186 711558
rect 244422 711322 279866 711558
rect 280102 711322 280186 711558
rect 280422 711322 351866 711558
rect 352102 711322 352186 711558
rect 352422 711322 387866 711558
rect 388102 711322 388186 711558
rect 388422 711322 423866 711558
rect 424102 711322 424186 711558
rect 424422 711322 459866 711558
rect 460102 711322 460186 711558
rect 460422 711322 495866 711558
rect 496102 711322 496186 711558
rect 496422 711322 531866 711558
rect 532102 711322 532186 711558
rect 532422 711322 567866 711558
rect 568102 711322 568186 711558
rect 568422 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 27866 711238
rect 28102 711002 28186 711238
rect 28422 711002 63866 711238
rect 64102 711002 64186 711238
rect 64422 711002 99866 711238
rect 100102 711002 100186 711238
rect 100422 711002 135866 711238
rect 136102 711002 136186 711238
rect 136422 711002 171866 711238
rect 172102 711002 172186 711238
rect 172422 711002 207866 711238
rect 208102 711002 208186 711238
rect 208422 711002 243866 711238
rect 244102 711002 244186 711238
rect 244422 711002 279866 711238
rect 280102 711002 280186 711238
rect 280422 711002 351866 711238
rect 352102 711002 352186 711238
rect 352422 711002 387866 711238
rect 388102 711002 388186 711238
rect 388422 711002 423866 711238
rect 424102 711002 424186 711238
rect 424422 711002 459866 711238
rect 460102 711002 460186 711238
rect 460422 711002 495866 711238
rect 496102 711002 496186 711238
rect 496422 711002 531866 711238
rect 532102 711002 532186 711238
rect 532422 711002 567866 711238
rect 568102 711002 568186 711238
rect 568422 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 384146 710598
rect 384382 710362 384466 710598
rect 384702 710362 420146 710598
rect 420382 710362 420466 710598
rect 420702 710362 456146 710598
rect 456382 710362 456466 710598
rect 456702 710362 492146 710598
rect 492382 710362 492466 710598
rect 492702 710362 528146 710598
rect 528382 710362 528466 710598
rect 528702 710362 564146 710598
rect 564382 710362 564466 710598
rect 564702 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 384146 710278
rect 384382 710042 384466 710278
rect 384702 710042 420146 710278
rect 420382 710042 420466 710278
rect 420702 710042 456146 710278
rect 456382 710042 456466 710278
rect 456702 710042 492146 710278
rect 492382 710042 492466 710278
rect 492702 710042 528146 710278
rect 528382 710042 528466 710278
rect 528702 710042 564146 710278
rect 564382 710042 564466 710278
rect 564702 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 20426 709638
rect 20662 709402 20746 709638
rect 20982 709402 380426 709638
rect 380662 709402 380746 709638
rect 380982 709402 416426 709638
rect 416662 709402 416746 709638
rect 416982 709402 452426 709638
rect 452662 709402 452746 709638
rect 452982 709402 488426 709638
rect 488662 709402 488746 709638
rect 488982 709402 524426 709638
rect 524662 709402 524746 709638
rect 524982 709402 560426 709638
rect 560662 709402 560746 709638
rect 560982 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 20426 709318
rect 20662 709082 20746 709318
rect 20982 709082 380426 709318
rect 380662 709082 380746 709318
rect 380982 709082 416426 709318
rect 416662 709082 416746 709318
rect 416982 709082 452426 709318
rect 452662 709082 452746 709318
rect 452982 709082 488426 709318
rect 488662 709082 488746 709318
rect 488982 709082 524426 709318
rect 524662 709082 524746 709318
rect 524982 709082 560426 709318
rect 560662 709082 560746 709318
rect 560982 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 16706 708678
rect 16942 708442 17026 708678
rect 17262 708442 376706 708678
rect 376942 708442 377026 708678
rect 377262 708442 412706 708678
rect 412942 708442 413026 708678
rect 413262 708442 448706 708678
rect 448942 708442 449026 708678
rect 449262 708442 520706 708678
rect 520942 708442 521026 708678
rect 521262 708442 556706 708678
rect 556942 708442 557026 708678
rect 557262 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 16706 708358
rect 16942 708122 17026 708358
rect 17262 708122 376706 708358
rect 376942 708122 377026 708358
rect 377262 708122 412706 708358
rect 412942 708122 413026 708358
rect 413262 708122 448706 708358
rect 448942 708122 449026 708358
rect 449262 708122 520706 708358
rect 520942 708122 521026 708358
rect 521262 708122 556706 708358
rect 556942 708122 557026 708358
rect 557262 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 12986 707718
rect 13222 707482 13306 707718
rect 13542 707482 48986 707718
rect 49222 707482 49306 707718
rect 49542 707482 84986 707718
rect 85222 707482 85306 707718
rect 85542 707482 120986 707718
rect 121222 707482 121306 707718
rect 121542 707482 156986 707718
rect 157222 707482 157306 707718
rect 157542 707482 192986 707718
rect 193222 707482 193306 707718
rect 193542 707482 228986 707718
rect 229222 707482 229306 707718
rect 229542 707482 264986 707718
rect 265222 707482 265306 707718
rect 265542 707482 300986 707718
rect 301222 707482 301306 707718
rect 301542 707482 336986 707718
rect 337222 707482 337306 707718
rect 337542 707482 372986 707718
rect 373222 707482 373306 707718
rect 373542 707482 408986 707718
rect 409222 707482 409306 707718
rect 409542 707482 444986 707718
rect 445222 707482 445306 707718
rect 445542 707482 480986 707718
rect 481222 707482 481306 707718
rect 481542 707482 516986 707718
rect 517222 707482 517306 707718
rect 517542 707482 552986 707718
rect 553222 707482 553306 707718
rect 553542 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 12986 707398
rect 13222 707162 13306 707398
rect 13542 707162 48986 707398
rect 49222 707162 49306 707398
rect 49542 707162 84986 707398
rect 85222 707162 85306 707398
rect 85542 707162 120986 707398
rect 121222 707162 121306 707398
rect 121542 707162 156986 707398
rect 157222 707162 157306 707398
rect 157542 707162 192986 707398
rect 193222 707162 193306 707398
rect 193542 707162 228986 707398
rect 229222 707162 229306 707398
rect 229542 707162 264986 707398
rect 265222 707162 265306 707398
rect 265542 707162 300986 707398
rect 301222 707162 301306 707398
rect 301542 707162 336986 707398
rect 337222 707162 337306 707398
rect 337542 707162 372986 707398
rect 373222 707162 373306 707398
rect 373542 707162 408986 707398
rect 409222 707162 409306 707398
rect 409542 707162 444986 707398
rect 445222 707162 445306 707398
rect 445542 707162 480986 707398
rect 481222 707162 481306 707398
rect 481542 707162 516986 707398
rect 517222 707162 517306 707398
rect 517542 707162 552986 707398
rect 553222 707162 553306 707398
rect 553542 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 9266 706758
rect 9502 706522 9586 706758
rect 9822 706522 45266 706758
rect 45502 706522 45586 706758
rect 45822 706522 81266 706758
rect 81502 706522 81586 706758
rect 81822 706522 117266 706758
rect 117502 706522 117586 706758
rect 117822 706522 153266 706758
rect 153502 706522 153586 706758
rect 153822 706522 189266 706758
rect 189502 706522 189586 706758
rect 189822 706522 225266 706758
rect 225502 706522 225586 706758
rect 225822 706522 261266 706758
rect 261502 706522 261586 706758
rect 261822 706522 297266 706758
rect 297502 706522 297586 706758
rect 297822 706522 333266 706758
rect 333502 706522 333586 706758
rect 333822 706522 369266 706758
rect 369502 706522 369586 706758
rect 369822 706522 405266 706758
rect 405502 706522 405586 706758
rect 405822 706522 441266 706758
rect 441502 706522 441586 706758
rect 441822 706522 477266 706758
rect 477502 706522 477586 706758
rect 477822 706522 513266 706758
rect 513502 706522 513586 706758
rect 513822 706522 549266 706758
rect 549502 706522 549586 706758
rect 549822 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 9266 706438
rect 9502 706202 9586 706438
rect 9822 706202 45266 706438
rect 45502 706202 45586 706438
rect 45822 706202 81266 706438
rect 81502 706202 81586 706438
rect 81822 706202 117266 706438
rect 117502 706202 117586 706438
rect 117822 706202 153266 706438
rect 153502 706202 153586 706438
rect 153822 706202 189266 706438
rect 189502 706202 189586 706438
rect 189822 706202 225266 706438
rect 225502 706202 225586 706438
rect 225822 706202 261266 706438
rect 261502 706202 261586 706438
rect 261822 706202 297266 706438
rect 297502 706202 297586 706438
rect 297822 706202 333266 706438
rect 333502 706202 333586 706438
rect 333822 706202 369266 706438
rect 369502 706202 369586 706438
rect 369822 706202 405266 706438
rect 405502 706202 405586 706438
rect 405822 706202 441266 706438
rect 441502 706202 441586 706438
rect 441822 706202 477266 706438
rect 477502 706202 477586 706438
rect 477822 706202 513266 706438
rect 513502 706202 513586 706438
rect 513822 706202 549266 706438
rect 549502 706202 549586 706438
rect 549822 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 5546 705798
rect 5782 705562 5866 705798
rect 6102 705562 41546 705798
rect 41782 705562 41866 705798
rect 42102 705562 77546 705798
rect 77782 705562 77866 705798
rect 78102 705562 113546 705798
rect 113782 705562 113866 705798
rect 114102 705562 149546 705798
rect 149782 705562 149866 705798
rect 150102 705562 185546 705798
rect 185782 705562 185866 705798
rect 186102 705562 221546 705798
rect 221782 705562 221866 705798
rect 222102 705562 257546 705798
rect 257782 705562 257866 705798
rect 258102 705562 293546 705798
rect 293782 705562 293866 705798
rect 294102 705562 329546 705798
rect 329782 705562 329866 705798
rect 330102 705562 365546 705798
rect 365782 705562 365866 705798
rect 366102 705562 401546 705798
rect 401782 705562 401866 705798
rect 402102 705562 437546 705798
rect 437782 705562 437866 705798
rect 438102 705562 473546 705798
rect 473782 705562 473866 705798
rect 474102 705562 509546 705798
rect 509782 705562 509866 705798
rect 510102 705562 545546 705798
rect 545782 705562 545866 705798
rect 546102 705562 581546 705798
rect 581782 705562 581866 705798
rect 582102 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 5546 705478
rect 5782 705242 5866 705478
rect 6102 705242 41546 705478
rect 41782 705242 41866 705478
rect 42102 705242 77546 705478
rect 77782 705242 77866 705478
rect 78102 705242 113546 705478
rect 113782 705242 113866 705478
rect 114102 705242 149546 705478
rect 149782 705242 149866 705478
rect 150102 705242 185546 705478
rect 185782 705242 185866 705478
rect 186102 705242 221546 705478
rect 221782 705242 221866 705478
rect 222102 705242 257546 705478
rect 257782 705242 257866 705478
rect 258102 705242 293546 705478
rect 293782 705242 293866 705478
rect 294102 705242 329546 705478
rect 329782 705242 329866 705478
rect 330102 705242 365546 705478
rect 365782 705242 365866 705478
rect 366102 705242 401546 705478
rect 401782 705242 401866 705478
rect 402102 705242 437546 705478
rect 437782 705242 437866 705478
rect 438102 705242 473546 705478
rect 473782 705242 473866 705478
rect 474102 705242 509546 705478
rect 509782 705242 509866 705478
rect 510102 705242 545546 705478
rect 545782 705242 545866 705478
rect 546102 705242 581546 705478
rect 581782 705242 581866 705478
rect 582102 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 698614 592650 698646
rect -8726 698378 -4854 698614
rect -4618 698378 -4534 698614
rect -4298 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 588222 698614
rect 588458 698378 588542 698614
rect 588778 698378 592650 698614
rect -8726 698294 592650 698378
rect -8726 698058 -4854 698294
rect -4618 698058 -4534 698294
rect -4298 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 588222 698294
rect 588458 698058 588542 698294
rect 588778 698058 592650 698294
rect -8726 698026 592650 698058
rect -8726 694894 592650 694926
rect -8726 694658 -3894 694894
rect -3658 694658 -3574 694894
rect -3338 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 587262 694894
rect 587498 694658 587582 694894
rect 587818 694658 592650 694894
rect -8726 694574 592650 694658
rect -8726 694338 -3894 694574
rect -3658 694338 -3574 694574
rect -3338 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 587262 694574
rect 587498 694338 587582 694574
rect 587818 694338 592650 694574
rect -8726 694306 592650 694338
rect -8726 691174 592650 691206
rect -8726 690938 -2934 691174
rect -2698 690938 -2614 691174
rect -2378 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 586302 691174
rect 586538 690938 586622 691174
rect 586858 690938 592650 691174
rect -8726 690854 592650 690938
rect -8726 690618 -2934 690854
rect -2698 690618 -2614 690854
rect -2378 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 586302 690854
rect 586538 690618 586622 690854
rect 586858 690618 592650 690854
rect -8726 690586 592650 690618
rect -8726 687454 592650 687486
rect -8726 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 592650 687454
rect -8726 687134 592650 687218
rect -8726 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 592650 687134
rect -8726 686866 592650 686898
rect -8726 677494 592650 677526
rect -8726 677258 -8694 677494
rect -8458 677258 -8374 677494
rect -8138 677258 27866 677494
rect 28102 677258 28186 677494
rect 28422 677258 63866 677494
rect 64102 677258 64186 677494
rect 64422 677258 99866 677494
rect 100102 677258 100186 677494
rect 100422 677258 135866 677494
rect 136102 677258 136186 677494
rect 136422 677258 171866 677494
rect 172102 677258 172186 677494
rect 172422 677258 207866 677494
rect 208102 677258 208186 677494
rect 208422 677258 243866 677494
rect 244102 677258 244186 677494
rect 244422 677258 279866 677494
rect 280102 677258 280186 677494
rect 280422 677258 351866 677494
rect 352102 677258 352186 677494
rect 352422 677258 387866 677494
rect 388102 677258 388186 677494
rect 388422 677258 423866 677494
rect 424102 677258 424186 677494
rect 424422 677258 459866 677494
rect 460102 677258 460186 677494
rect 460422 677258 495866 677494
rect 496102 677258 496186 677494
rect 496422 677258 531866 677494
rect 532102 677258 532186 677494
rect 532422 677258 567866 677494
rect 568102 677258 568186 677494
rect 568422 677258 592062 677494
rect 592298 677258 592382 677494
rect 592618 677258 592650 677494
rect -8726 677174 592650 677258
rect -8726 676938 -8694 677174
rect -8458 676938 -8374 677174
rect -8138 676938 27866 677174
rect 28102 676938 28186 677174
rect 28422 676938 63866 677174
rect 64102 676938 64186 677174
rect 64422 676938 99866 677174
rect 100102 676938 100186 677174
rect 100422 676938 135866 677174
rect 136102 676938 136186 677174
rect 136422 676938 171866 677174
rect 172102 676938 172186 677174
rect 172422 676938 207866 677174
rect 208102 676938 208186 677174
rect 208422 676938 243866 677174
rect 244102 676938 244186 677174
rect 244422 676938 279866 677174
rect 280102 676938 280186 677174
rect 280422 676938 351866 677174
rect 352102 676938 352186 677174
rect 352422 676938 387866 677174
rect 388102 676938 388186 677174
rect 388422 676938 423866 677174
rect 424102 676938 424186 677174
rect 424422 676938 459866 677174
rect 460102 676938 460186 677174
rect 460422 676938 495866 677174
rect 496102 676938 496186 677174
rect 496422 676938 531866 677174
rect 532102 676938 532186 677174
rect 532422 676938 567866 677174
rect 568102 676938 568186 677174
rect 568422 676938 592062 677174
rect 592298 676938 592382 677174
rect 592618 676938 592650 677174
rect -8726 676906 592650 676938
rect -8726 673774 592650 673806
rect -8726 673538 -7734 673774
rect -7498 673538 -7414 673774
rect -7178 673538 384146 673774
rect 384382 673538 384466 673774
rect 384702 673538 420146 673774
rect 420382 673538 420466 673774
rect 420702 673538 456146 673774
rect 456382 673538 456466 673774
rect 456702 673538 492146 673774
rect 492382 673538 492466 673774
rect 492702 673538 528146 673774
rect 528382 673538 528466 673774
rect 528702 673538 564146 673774
rect 564382 673538 564466 673774
rect 564702 673538 591102 673774
rect 591338 673538 591422 673774
rect 591658 673538 592650 673774
rect -8726 673454 592650 673538
rect -8726 673218 -7734 673454
rect -7498 673218 -7414 673454
rect -7178 673218 384146 673454
rect 384382 673218 384466 673454
rect 384702 673218 420146 673454
rect 420382 673218 420466 673454
rect 420702 673218 456146 673454
rect 456382 673218 456466 673454
rect 456702 673218 492146 673454
rect 492382 673218 492466 673454
rect 492702 673218 528146 673454
rect 528382 673218 528466 673454
rect 528702 673218 564146 673454
rect 564382 673218 564466 673454
rect 564702 673218 591102 673454
rect 591338 673218 591422 673454
rect 591658 673218 592650 673454
rect -8726 673186 592650 673218
rect -8726 670054 592650 670086
rect -8726 669818 -6774 670054
rect -6538 669818 -6454 670054
rect -6218 669818 20426 670054
rect 20662 669818 20746 670054
rect 20982 669818 380426 670054
rect 380662 669818 380746 670054
rect 380982 669818 416426 670054
rect 416662 669818 416746 670054
rect 416982 669818 452426 670054
rect 452662 669818 452746 670054
rect 452982 669818 488426 670054
rect 488662 669818 488746 670054
rect 488982 669818 524426 670054
rect 524662 669818 524746 670054
rect 524982 669818 560426 670054
rect 560662 669818 560746 670054
rect 560982 669818 590142 670054
rect 590378 669818 590462 670054
rect 590698 669818 592650 670054
rect -8726 669734 592650 669818
rect -8726 669498 -6774 669734
rect -6538 669498 -6454 669734
rect -6218 669498 20426 669734
rect 20662 669498 20746 669734
rect 20982 669498 380426 669734
rect 380662 669498 380746 669734
rect 380982 669498 416426 669734
rect 416662 669498 416746 669734
rect 416982 669498 452426 669734
rect 452662 669498 452746 669734
rect 452982 669498 488426 669734
rect 488662 669498 488746 669734
rect 488982 669498 524426 669734
rect 524662 669498 524746 669734
rect 524982 669498 560426 669734
rect 560662 669498 560746 669734
rect 560982 669498 590142 669734
rect 590378 669498 590462 669734
rect 590698 669498 592650 669734
rect -8726 669466 592650 669498
rect -8726 666334 592650 666366
rect -8726 666098 -5814 666334
rect -5578 666098 -5494 666334
rect -5258 666098 16706 666334
rect 16942 666098 17026 666334
rect 17262 666098 376706 666334
rect 376942 666098 377026 666334
rect 377262 666098 412706 666334
rect 412942 666098 413026 666334
rect 413262 666098 448706 666334
rect 448942 666098 449026 666334
rect 449262 666098 520706 666334
rect 520942 666098 521026 666334
rect 521262 666098 556706 666334
rect 556942 666098 557026 666334
rect 557262 666098 589182 666334
rect 589418 666098 589502 666334
rect 589738 666098 592650 666334
rect -8726 666014 592650 666098
rect -8726 665778 -5814 666014
rect -5578 665778 -5494 666014
rect -5258 665778 16706 666014
rect 16942 665778 17026 666014
rect 17262 665778 376706 666014
rect 376942 665778 377026 666014
rect 377262 665778 412706 666014
rect 412942 665778 413026 666014
rect 413262 665778 448706 666014
rect 448942 665778 449026 666014
rect 449262 665778 520706 666014
rect 520942 665778 521026 666014
rect 521262 665778 556706 666014
rect 556942 665778 557026 666014
rect 557262 665778 589182 666014
rect 589418 665778 589502 666014
rect 589738 665778 592650 666014
rect -8726 665746 592650 665778
rect -8726 662614 592650 662646
rect -8726 662378 -4854 662614
rect -4618 662378 -4534 662614
rect -4298 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 588222 662614
rect 588458 662378 588542 662614
rect 588778 662378 592650 662614
rect -8726 662294 592650 662378
rect -8726 662058 -4854 662294
rect -4618 662058 -4534 662294
rect -4298 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 588222 662294
rect 588458 662058 588542 662294
rect 588778 662058 592650 662294
rect -8726 662026 592650 662058
rect -8726 658894 592650 658926
rect -8726 658658 -3894 658894
rect -3658 658658 -3574 658894
rect -3338 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 587262 658894
rect 587498 658658 587582 658894
rect 587818 658658 592650 658894
rect -8726 658574 592650 658658
rect -8726 658338 -3894 658574
rect -3658 658338 -3574 658574
rect -3338 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 587262 658574
rect 587498 658338 587582 658574
rect 587818 658338 592650 658574
rect -8726 658306 592650 658338
rect -8726 655174 592650 655206
rect -8726 654938 -2934 655174
rect -2698 654938 -2614 655174
rect -2378 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 39610 655174
rect 39846 654938 70330 655174
rect 70566 654938 101050 655174
rect 101286 654938 131770 655174
rect 132006 654938 162490 655174
rect 162726 654938 193210 655174
rect 193446 654938 223930 655174
rect 224166 654938 254650 655174
rect 254886 654938 285370 655174
rect 285606 654938 316090 655174
rect 316326 654938 346810 655174
rect 347046 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 479610 655174
rect 479846 654938 510330 655174
rect 510566 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 586302 655174
rect 586538 654938 586622 655174
rect 586858 654938 592650 655174
rect -8726 654854 592650 654938
rect -8726 654618 -2934 654854
rect -2698 654618 -2614 654854
rect -2378 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 39610 654854
rect 39846 654618 70330 654854
rect 70566 654618 101050 654854
rect 101286 654618 131770 654854
rect 132006 654618 162490 654854
rect 162726 654618 193210 654854
rect 193446 654618 223930 654854
rect 224166 654618 254650 654854
rect 254886 654618 285370 654854
rect 285606 654618 316090 654854
rect 316326 654618 346810 654854
rect 347046 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 479610 654854
rect 479846 654618 510330 654854
rect 510566 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 586302 654854
rect 586538 654618 586622 654854
rect 586858 654618 592650 654854
rect -8726 654586 592650 654618
rect -8726 651454 592650 651486
rect -8726 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 24250 651454
rect 24486 651218 54970 651454
rect 55206 651218 85690 651454
rect 85926 651218 116410 651454
rect 116646 651218 147130 651454
rect 147366 651218 177850 651454
rect 178086 651218 208570 651454
rect 208806 651218 239290 651454
rect 239526 651218 270010 651454
rect 270246 651218 300730 651454
rect 300966 651218 331450 651454
rect 331686 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 464250 651454
rect 464486 651218 494970 651454
rect 495206 651218 525690 651454
rect 525926 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 592650 651454
rect -8726 651134 592650 651218
rect -8726 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 24250 651134
rect 24486 650898 54970 651134
rect 55206 650898 85690 651134
rect 85926 650898 116410 651134
rect 116646 650898 147130 651134
rect 147366 650898 177850 651134
rect 178086 650898 208570 651134
rect 208806 650898 239290 651134
rect 239526 650898 270010 651134
rect 270246 650898 300730 651134
rect 300966 650898 331450 651134
rect 331686 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 464250 651134
rect 464486 650898 494970 651134
rect 495206 650898 525690 651134
rect 525926 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 592650 651134
rect -8726 650866 592650 650898
rect -8726 641494 592650 641526
rect -8726 641258 -8694 641494
rect -8458 641258 -8374 641494
rect -8138 641258 27866 641494
rect 28102 641258 28186 641494
rect 28422 641258 387866 641494
rect 388102 641258 388186 641494
rect 388422 641258 423866 641494
rect 424102 641258 424186 641494
rect 424422 641258 531866 641494
rect 532102 641258 532186 641494
rect 532422 641258 567866 641494
rect 568102 641258 568186 641494
rect 568422 641258 592062 641494
rect 592298 641258 592382 641494
rect 592618 641258 592650 641494
rect -8726 641174 592650 641258
rect -8726 640938 -8694 641174
rect -8458 640938 -8374 641174
rect -8138 640938 27866 641174
rect 28102 640938 28186 641174
rect 28422 640938 387866 641174
rect 388102 640938 388186 641174
rect 388422 640938 423866 641174
rect 424102 640938 424186 641174
rect 424422 640938 531866 641174
rect 532102 640938 532186 641174
rect 532422 640938 567866 641174
rect 568102 640938 568186 641174
rect 568422 640938 592062 641174
rect 592298 640938 592382 641174
rect 592618 640938 592650 641174
rect -8726 640906 592650 640938
rect -8726 637774 592650 637806
rect -8726 637538 -7734 637774
rect -7498 637538 -7414 637774
rect -7178 637538 384146 637774
rect 384382 637538 384466 637774
rect 384702 637538 420146 637774
rect 420382 637538 420466 637774
rect 420702 637538 456146 637774
rect 456382 637538 456466 637774
rect 456702 637538 528146 637774
rect 528382 637538 528466 637774
rect 528702 637538 564146 637774
rect 564382 637538 564466 637774
rect 564702 637538 591102 637774
rect 591338 637538 591422 637774
rect 591658 637538 592650 637774
rect -8726 637454 592650 637538
rect -8726 637218 -7734 637454
rect -7498 637218 -7414 637454
rect -7178 637218 384146 637454
rect 384382 637218 384466 637454
rect 384702 637218 420146 637454
rect 420382 637218 420466 637454
rect 420702 637218 456146 637454
rect 456382 637218 456466 637454
rect 456702 637218 528146 637454
rect 528382 637218 528466 637454
rect 528702 637218 564146 637454
rect 564382 637218 564466 637454
rect 564702 637218 591102 637454
rect 591338 637218 591422 637454
rect 591658 637218 592650 637454
rect -8726 637186 592650 637218
rect -8726 634054 592650 634086
rect -8726 633818 -6774 634054
rect -6538 633818 -6454 634054
rect -6218 633818 20426 634054
rect 20662 633818 20746 634054
rect 20982 633818 380426 634054
rect 380662 633818 380746 634054
rect 380982 633818 416426 634054
rect 416662 633818 416746 634054
rect 416982 633818 452426 634054
rect 452662 633818 452746 634054
rect 452982 633818 524426 634054
rect 524662 633818 524746 634054
rect 524982 633818 560426 634054
rect 560662 633818 560746 634054
rect 560982 633818 590142 634054
rect 590378 633818 590462 634054
rect 590698 633818 592650 634054
rect -8726 633734 592650 633818
rect -8726 633498 -6774 633734
rect -6538 633498 -6454 633734
rect -6218 633498 20426 633734
rect 20662 633498 20746 633734
rect 20982 633498 380426 633734
rect 380662 633498 380746 633734
rect 380982 633498 416426 633734
rect 416662 633498 416746 633734
rect 416982 633498 452426 633734
rect 452662 633498 452746 633734
rect 452982 633498 524426 633734
rect 524662 633498 524746 633734
rect 524982 633498 560426 633734
rect 560662 633498 560746 633734
rect 560982 633498 590142 633734
rect 590378 633498 590462 633734
rect 590698 633498 592650 633734
rect -8726 633466 592650 633498
rect -8726 630334 592650 630366
rect -8726 630098 -5814 630334
rect -5578 630098 -5494 630334
rect -5258 630098 16706 630334
rect 16942 630098 17026 630334
rect 17262 630098 376706 630334
rect 376942 630098 377026 630334
rect 377262 630098 412706 630334
rect 412942 630098 413026 630334
rect 413262 630098 448706 630334
rect 448942 630098 449026 630334
rect 449262 630098 520706 630334
rect 520942 630098 521026 630334
rect 521262 630098 556706 630334
rect 556942 630098 557026 630334
rect 557262 630098 589182 630334
rect 589418 630098 589502 630334
rect 589738 630098 592650 630334
rect -8726 630014 592650 630098
rect -8726 629778 -5814 630014
rect -5578 629778 -5494 630014
rect -5258 629778 16706 630014
rect 16942 629778 17026 630014
rect 17262 629778 376706 630014
rect 376942 629778 377026 630014
rect 377262 629778 412706 630014
rect 412942 629778 413026 630014
rect 413262 629778 448706 630014
rect 448942 629778 449026 630014
rect 449262 629778 520706 630014
rect 520942 629778 521026 630014
rect 521262 629778 556706 630014
rect 556942 629778 557026 630014
rect 557262 629778 589182 630014
rect 589418 629778 589502 630014
rect 589738 629778 592650 630014
rect -8726 629746 592650 629778
rect -8726 626614 592650 626646
rect -8726 626378 -4854 626614
rect -4618 626378 -4534 626614
rect -4298 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 372986 626614
rect 373222 626378 373306 626614
rect 373542 626378 408986 626614
rect 409222 626378 409306 626614
rect 409542 626378 444986 626614
rect 445222 626378 445306 626614
rect 445542 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 588222 626614
rect 588458 626378 588542 626614
rect 588778 626378 592650 626614
rect -8726 626294 592650 626378
rect -8726 626058 -4854 626294
rect -4618 626058 -4534 626294
rect -4298 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 372986 626294
rect 373222 626058 373306 626294
rect 373542 626058 408986 626294
rect 409222 626058 409306 626294
rect 409542 626058 444986 626294
rect 445222 626058 445306 626294
rect 445542 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 588222 626294
rect 588458 626058 588542 626294
rect 588778 626058 592650 626294
rect -8726 626026 592650 626058
rect -8726 622894 592650 622926
rect -8726 622658 -3894 622894
rect -3658 622658 -3574 622894
rect -3338 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 369266 622894
rect 369502 622658 369586 622894
rect 369822 622658 405266 622894
rect 405502 622658 405586 622894
rect 405822 622658 441266 622894
rect 441502 622658 441586 622894
rect 441822 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 587262 622894
rect 587498 622658 587582 622894
rect 587818 622658 592650 622894
rect -8726 622574 592650 622658
rect -8726 622338 -3894 622574
rect -3658 622338 -3574 622574
rect -3338 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 369266 622574
rect 369502 622338 369586 622574
rect 369822 622338 405266 622574
rect 405502 622338 405586 622574
rect 405822 622338 441266 622574
rect 441502 622338 441586 622574
rect 441822 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 587262 622574
rect 587498 622338 587582 622574
rect 587818 622338 592650 622574
rect -8726 622306 592650 622338
rect -8726 619174 592650 619206
rect -8726 618938 -2934 619174
rect -2698 618938 -2614 619174
rect -2378 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 39610 619174
rect 39846 618938 70330 619174
rect 70566 618938 101050 619174
rect 101286 618938 131770 619174
rect 132006 618938 162490 619174
rect 162726 618938 193210 619174
rect 193446 618938 223930 619174
rect 224166 618938 254650 619174
rect 254886 618938 285370 619174
rect 285606 618938 316090 619174
rect 316326 618938 346810 619174
rect 347046 618938 365546 619174
rect 365782 618938 365866 619174
rect 366102 618938 401546 619174
rect 401782 618938 401866 619174
rect 402102 618938 437546 619174
rect 437782 618938 437866 619174
rect 438102 618938 479610 619174
rect 479846 618938 510330 619174
rect 510566 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 586302 619174
rect 586538 618938 586622 619174
rect 586858 618938 592650 619174
rect -8726 618854 592650 618938
rect -8726 618618 -2934 618854
rect -2698 618618 -2614 618854
rect -2378 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 39610 618854
rect 39846 618618 70330 618854
rect 70566 618618 101050 618854
rect 101286 618618 131770 618854
rect 132006 618618 162490 618854
rect 162726 618618 193210 618854
rect 193446 618618 223930 618854
rect 224166 618618 254650 618854
rect 254886 618618 285370 618854
rect 285606 618618 316090 618854
rect 316326 618618 346810 618854
rect 347046 618618 365546 618854
rect 365782 618618 365866 618854
rect 366102 618618 401546 618854
rect 401782 618618 401866 618854
rect 402102 618618 437546 618854
rect 437782 618618 437866 618854
rect 438102 618618 479610 618854
rect 479846 618618 510330 618854
rect 510566 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 586302 618854
rect 586538 618618 586622 618854
rect 586858 618618 592650 618854
rect -8726 618586 592650 618618
rect -8726 615454 592650 615486
rect -8726 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 24250 615454
rect 24486 615218 54970 615454
rect 55206 615218 85690 615454
rect 85926 615218 116410 615454
rect 116646 615218 147130 615454
rect 147366 615218 177850 615454
rect 178086 615218 208570 615454
rect 208806 615218 239290 615454
rect 239526 615218 270010 615454
rect 270246 615218 300730 615454
rect 300966 615218 331450 615454
rect 331686 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 464250 615454
rect 464486 615218 494970 615454
rect 495206 615218 525690 615454
rect 525926 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 592650 615454
rect -8726 615134 592650 615218
rect -8726 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 24250 615134
rect 24486 614898 54970 615134
rect 55206 614898 85690 615134
rect 85926 614898 116410 615134
rect 116646 614898 147130 615134
rect 147366 614898 177850 615134
rect 178086 614898 208570 615134
rect 208806 614898 239290 615134
rect 239526 614898 270010 615134
rect 270246 614898 300730 615134
rect 300966 614898 331450 615134
rect 331686 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 464250 615134
rect 464486 614898 494970 615134
rect 495206 614898 525690 615134
rect 525926 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 592650 615134
rect -8726 614866 592650 614898
rect -8726 605494 592650 605526
rect -8726 605258 -8694 605494
rect -8458 605258 -8374 605494
rect -8138 605258 27866 605494
rect 28102 605258 28186 605494
rect 28422 605258 387866 605494
rect 388102 605258 388186 605494
rect 388422 605258 423866 605494
rect 424102 605258 424186 605494
rect 424422 605258 531866 605494
rect 532102 605258 532186 605494
rect 532422 605258 567866 605494
rect 568102 605258 568186 605494
rect 568422 605258 592062 605494
rect 592298 605258 592382 605494
rect 592618 605258 592650 605494
rect -8726 605174 592650 605258
rect -8726 604938 -8694 605174
rect -8458 604938 -8374 605174
rect -8138 604938 27866 605174
rect 28102 604938 28186 605174
rect 28422 604938 387866 605174
rect 388102 604938 388186 605174
rect 388422 604938 423866 605174
rect 424102 604938 424186 605174
rect 424422 604938 531866 605174
rect 532102 604938 532186 605174
rect 532422 604938 567866 605174
rect 568102 604938 568186 605174
rect 568422 604938 592062 605174
rect 592298 604938 592382 605174
rect 592618 604938 592650 605174
rect -8726 604906 592650 604938
rect -8726 601774 592650 601806
rect -8726 601538 -7734 601774
rect -7498 601538 -7414 601774
rect -7178 601538 384146 601774
rect 384382 601538 384466 601774
rect 384702 601538 420146 601774
rect 420382 601538 420466 601774
rect 420702 601538 456146 601774
rect 456382 601538 456466 601774
rect 456702 601538 528146 601774
rect 528382 601538 528466 601774
rect 528702 601538 564146 601774
rect 564382 601538 564466 601774
rect 564702 601538 591102 601774
rect 591338 601538 591422 601774
rect 591658 601538 592650 601774
rect -8726 601454 592650 601538
rect -8726 601218 -7734 601454
rect -7498 601218 -7414 601454
rect -7178 601218 384146 601454
rect 384382 601218 384466 601454
rect 384702 601218 420146 601454
rect 420382 601218 420466 601454
rect 420702 601218 456146 601454
rect 456382 601218 456466 601454
rect 456702 601218 528146 601454
rect 528382 601218 528466 601454
rect 528702 601218 564146 601454
rect 564382 601218 564466 601454
rect 564702 601218 591102 601454
rect 591338 601218 591422 601454
rect 591658 601218 592650 601454
rect -8726 601186 592650 601218
rect -8726 598054 592650 598086
rect -8726 597818 -6774 598054
rect -6538 597818 -6454 598054
rect -6218 597818 20426 598054
rect 20662 597818 20746 598054
rect 20982 597818 380426 598054
rect 380662 597818 380746 598054
rect 380982 597818 416426 598054
rect 416662 597818 416746 598054
rect 416982 597818 452426 598054
rect 452662 597818 452746 598054
rect 452982 597818 488426 598054
rect 488662 597818 488746 598054
rect 488982 597818 524426 598054
rect 524662 597818 524746 598054
rect 524982 597818 560426 598054
rect 560662 597818 560746 598054
rect 560982 597818 590142 598054
rect 590378 597818 590462 598054
rect 590698 597818 592650 598054
rect -8726 597734 592650 597818
rect -8726 597498 -6774 597734
rect -6538 597498 -6454 597734
rect -6218 597498 20426 597734
rect 20662 597498 20746 597734
rect 20982 597498 380426 597734
rect 380662 597498 380746 597734
rect 380982 597498 416426 597734
rect 416662 597498 416746 597734
rect 416982 597498 452426 597734
rect 452662 597498 452746 597734
rect 452982 597498 488426 597734
rect 488662 597498 488746 597734
rect 488982 597498 524426 597734
rect 524662 597498 524746 597734
rect 524982 597498 560426 597734
rect 560662 597498 560746 597734
rect 560982 597498 590142 597734
rect 590378 597498 590462 597734
rect 590698 597498 592650 597734
rect -8726 597466 592650 597498
rect -8726 594334 592650 594366
rect -8726 594098 -5814 594334
rect -5578 594098 -5494 594334
rect -5258 594098 16706 594334
rect 16942 594098 17026 594334
rect 17262 594098 376706 594334
rect 376942 594098 377026 594334
rect 377262 594098 412706 594334
rect 412942 594098 413026 594334
rect 413262 594098 448706 594334
rect 448942 594098 449026 594334
rect 449262 594098 484706 594334
rect 484942 594098 485026 594334
rect 485262 594098 520706 594334
rect 520942 594098 521026 594334
rect 521262 594098 556706 594334
rect 556942 594098 557026 594334
rect 557262 594098 589182 594334
rect 589418 594098 589502 594334
rect 589738 594098 592650 594334
rect -8726 594014 592650 594098
rect -8726 593778 -5814 594014
rect -5578 593778 -5494 594014
rect -5258 593778 16706 594014
rect 16942 593778 17026 594014
rect 17262 593778 376706 594014
rect 376942 593778 377026 594014
rect 377262 593778 412706 594014
rect 412942 593778 413026 594014
rect 413262 593778 448706 594014
rect 448942 593778 449026 594014
rect 449262 593778 484706 594014
rect 484942 593778 485026 594014
rect 485262 593778 520706 594014
rect 520942 593778 521026 594014
rect 521262 593778 556706 594014
rect 556942 593778 557026 594014
rect 557262 593778 589182 594014
rect 589418 593778 589502 594014
rect 589738 593778 592650 594014
rect -8726 593746 592650 593778
rect -8726 590614 592650 590646
rect -8726 590378 -4854 590614
rect -4618 590378 -4534 590614
rect -4298 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 372986 590614
rect 373222 590378 373306 590614
rect 373542 590378 408986 590614
rect 409222 590378 409306 590614
rect 409542 590378 444986 590614
rect 445222 590378 445306 590614
rect 445542 590378 480986 590614
rect 481222 590378 481306 590614
rect 481542 590378 516986 590614
rect 517222 590378 517306 590614
rect 517542 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 588222 590614
rect 588458 590378 588542 590614
rect 588778 590378 592650 590614
rect -8726 590294 592650 590378
rect -8726 590058 -4854 590294
rect -4618 590058 -4534 590294
rect -4298 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 372986 590294
rect 373222 590058 373306 590294
rect 373542 590058 408986 590294
rect 409222 590058 409306 590294
rect 409542 590058 444986 590294
rect 445222 590058 445306 590294
rect 445542 590058 480986 590294
rect 481222 590058 481306 590294
rect 481542 590058 516986 590294
rect 517222 590058 517306 590294
rect 517542 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 588222 590294
rect 588458 590058 588542 590294
rect 588778 590058 592650 590294
rect -8726 590026 592650 590058
rect -8726 586894 592650 586926
rect -8726 586658 -3894 586894
rect -3658 586658 -3574 586894
rect -3338 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 369266 586894
rect 369502 586658 369586 586894
rect 369822 586658 405266 586894
rect 405502 586658 405586 586894
rect 405822 586658 441266 586894
rect 441502 586658 441586 586894
rect 441822 586658 477266 586894
rect 477502 586658 477586 586894
rect 477822 586658 513266 586894
rect 513502 586658 513586 586894
rect 513822 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 587262 586894
rect 587498 586658 587582 586894
rect 587818 586658 592650 586894
rect -8726 586574 592650 586658
rect -8726 586338 -3894 586574
rect -3658 586338 -3574 586574
rect -3338 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 369266 586574
rect 369502 586338 369586 586574
rect 369822 586338 405266 586574
rect 405502 586338 405586 586574
rect 405822 586338 441266 586574
rect 441502 586338 441586 586574
rect 441822 586338 477266 586574
rect 477502 586338 477586 586574
rect 477822 586338 513266 586574
rect 513502 586338 513586 586574
rect 513822 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 587262 586574
rect 587498 586338 587582 586574
rect 587818 586338 592650 586574
rect -8726 586306 592650 586338
rect -8726 583174 592650 583206
rect -8726 582938 -2934 583174
rect -2698 582938 -2614 583174
rect -2378 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 39610 583174
rect 39846 582938 70330 583174
rect 70566 582938 101050 583174
rect 101286 582938 131770 583174
rect 132006 582938 162490 583174
rect 162726 582938 193210 583174
rect 193446 582938 223930 583174
rect 224166 582938 254650 583174
rect 254886 582938 285370 583174
rect 285606 582938 316090 583174
rect 316326 582938 346810 583174
rect 347046 582938 365546 583174
rect 365782 582938 365866 583174
rect 366102 582938 401546 583174
rect 401782 582938 401866 583174
rect 402102 582938 437546 583174
rect 437782 582938 437866 583174
rect 438102 582938 473546 583174
rect 473782 582938 473866 583174
rect 474102 582938 509546 583174
rect 509782 582938 509866 583174
rect 510102 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 586302 583174
rect 586538 582938 586622 583174
rect 586858 582938 592650 583174
rect -8726 582854 592650 582938
rect -8726 582618 -2934 582854
rect -2698 582618 -2614 582854
rect -2378 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 39610 582854
rect 39846 582618 70330 582854
rect 70566 582618 101050 582854
rect 101286 582618 131770 582854
rect 132006 582618 162490 582854
rect 162726 582618 193210 582854
rect 193446 582618 223930 582854
rect 224166 582618 254650 582854
rect 254886 582618 285370 582854
rect 285606 582618 316090 582854
rect 316326 582618 346810 582854
rect 347046 582618 365546 582854
rect 365782 582618 365866 582854
rect 366102 582618 401546 582854
rect 401782 582618 401866 582854
rect 402102 582618 437546 582854
rect 437782 582618 437866 582854
rect 438102 582618 473546 582854
rect 473782 582618 473866 582854
rect 474102 582618 509546 582854
rect 509782 582618 509866 582854
rect 510102 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 586302 582854
rect 586538 582618 586622 582854
rect 586858 582618 592650 582854
rect -8726 582586 592650 582618
rect -8726 579454 592650 579486
rect -8726 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 24250 579454
rect 24486 579218 54970 579454
rect 55206 579218 85690 579454
rect 85926 579218 116410 579454
rect 116646 579218 147130 579454
rect 147366 579218 177850 579454
rect 178086 579218 208570 579454
rect 208806 579218 239290 579454
rect 239526 579218 270010 579454
rect 270246 579218 300730 579454
rect 300966 579218 331450 579454
rect 331686 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 592650 579454
rect -8726 579134 592650 579218
rect -8726 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 24250 579134
rect 24486 578898 54970 579134
rect 55206 578898 85690 579134
rect 85926 578898 116410 579134
rect 116646 578898 147130 579134
rect 147366 578898 177850 579134
rect 178086 578898 208570 579134
rect 208806 578898 239290 579134
rect 239526 578898 270010 579134
rect 270246 578898 300730 579134
rect 300966 578898 331450 579134
rect 331686 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 592650 579134
rect -8726 578866 592650 578898
rect -8726 569494 592650 569526
rect -8726 569258 -8694 569494
rect -8458 569258 -8374 569494
rect -8138 569258 27866 569494
rect 28102 569258 28186 569494
rect 28422 569258 387866 569494
rect 388102 569258 388186 569494
rect 388422 569258 423866 569494
rect 424102 569258 424186 569494
rect 424422 569258 459866 569494
rect 460102 569258 460186 569494
rect 460422 569258 495866 569494
rect 496102 569258 496186 569494
rect 496422 569258 531866 569494
rect 532102 569258 532186 569494
rect 532422 569258 567866 569494
rect 568102 569258 568186 569494
rect 568422 569258 592062 569494
rect 592298 569258 592382 569494
rect 592618 569258 592650 569494
rect -8726 569174 592650 569258
rect -8726 568938 -8694 569174
rect -8458 568938 -8374 569174
rect -8138 568938 27866 569174
rect 28102 568938 28186 569174
rect 28422 568938 387866 569174
rect 388102 568938 388186 569174
rect 388422 568938 423866 569174
rect 424102 568938 424186 569174
rect 424422 568938 459866 569174
rect 460102 568938 460186 569174
rect 460422 568938 495866 569174
rect 496102 568938 496186 569174
rect 496422 568938 531866 569174
rect 532102 568938 532186 569174
rect 532422 568938 567866 569174
rect 568102 568938 568186 569174
rect 568422 568938 592062 569174
rect 592298 568938 592382 569174
rect 592618 568938 592650 569174
rect -8726 568906 592650 568938
rect -8726 565774 592650 565806
rect -8726 565538 -7734 565774
rect -7498 565538 -7414 565774
rect -7178 565538 384146 565774
rect 384382 565538 384466 565774
rect 384702 565538 420146 565774
rect 420382 565538 420466 565774
rect 420702 565538 456146 565774
rect 456382 565538 456466 565774
rect 456702 565538 492146 565774
rect 492382 565538 492466 565774
rect 492702 565538 528146 565774
rect 528382 565538 528466 565774
rect 528702 565538 564146 565774
rect 564382 565538 564466 565774
rect 564702 565538 591102 565774
rect 591338 565538 591422 565774
rect 591658 565538 592650 565774
rect -8726 565454 592650 565538
rect -8726 565218 -7734 565454
rect -7498 565218 -7414 565454
rect -7178 565218 384146 565454
rect 384382 565218 384466 565454
rect 384702 565218 420146 565454
rect 420382 565218 420466 565454
rect 420702 565218 456146 565454
rect 456382 565218 456466 565454
rect 456702 565218 492146 565454
rect 492382 565218 492466 565454
rect 492702 565218 528146 565454
rect 528382 565218 528466 565454
rect 528702 565218 564146 565454
rect 564382 565218 564466 565454
rect 564702 565218 591102 565454
rect 591338 565218 591422 565454
rect 591658 565218 592650 565454
rect -8726 565186 592650 565218
rect -8726 562054 592650 562086
rect -8726 561818 -6774 562054
rect -6538 561818 -6454 562054
rect -6218 561818 20426 562054
rect 20662 561818 20746 562054
rect 20982 561818 380426 562054
rect 380662 561818 380746 562054
rect 380982 561818 416426 562054
rect 416662 561818 416746 562054
rect 416982 561818 452426 562054
rect 452662 561818 452746 562054
rect 452982 561818 488426 562054
rect 488662 561818 488746 562054
rect 488982 561818 524426 562054
rect 524662 561818 524746 562054
rect 524982 561818 560426 562054
rect 560662 561818 560746 562054
rect 560982 561818 590142 562054
rect 590378 561818 590462 562054
rect 590698 561818 592650 562054
rect -8726 561734 592650 561818
rect -8726 561498 -6774 561734
rect -6538 561498 -6454 561734
rect -6218 561498 20426 561734
rect 20662 561498 20746 561734
rect 20982 561498 380426 561734
rect 380662 561498 380746 561734
rect 380982 561498 416426 561734
rect 416662 561498 416746 561734
rect 416982 561498 452426 561734
rect 452662 561498 452746 561734
rect 452982 561498 488426 561734
rect 488662 561498 488746 561734
rect 488982 561498 524426 561734
rect 524662 561498 524746 561734
rect 524982 561498 560426 561734
rect 560662 561498 560746 561734
rect 560982 561498 590142 561734
rect 590378 561498 590462 561734
rect 590698 561498 592650 561734
rect -8726 561466 592650 561498
rect -8726 558334 592650 558366
rect -8726 558098 -5814 558334
rect -5578 558098 -5494 558334
rect -5258 558098 16706 558334
rect 16942 558098 17026 558334
rect 17262 558098 376706 558334
rect 376942 558098 377026 558334
rect 377262 558098 412706 558334
rect 412942 558098 413026 558334
rect 413262 558098 448706 558334
rect 448942 558098 449026 558334
rect 449262 558098 484706 558334
rect 484942 558098 485026 558334
rect 485262 558098 520706 558334
rect 520942 558098 521026 558334
rect 521262 558098 556706 558334
rect 556942 558098 557026 558334
rect 557262 558098 589182 558334
rect 589418 558098 589502 558334
rect 589738 558098 592650 558334
rect -8726 558014 592650 558098
rect -8726 557778 -5814 558014
rect -5578 557778 -5494 558014
rect -5258 557778 16706 558014
rect 16942 557778 17026 558014
rect 17262 557778 376706 558014
rect 376942 557778 377026 558014
rect 377262 557778 412706 558014
rect 412942 557778 413026 558014
rect 413262 557778 448706 558014
rect 448942 557778 449026 558014
rect 449262 557778 484706 558014
rect 484942 557778 485026 558014
rect 485262 557778 520706 558014
rect 520942 557778 521026 558014
rect 521262 557778 556706 558014
rect 556942 557778 557026 558014
rect 557262 557778 589182 558014
rect 589418 557778 589502 558014
rect 589738 557778 592650 558014
rect -8726 557746 592650 557778
rect -8726 554614 592650 554646
rect -8726 554378 -4854 554614
rect -4618 554378 -4534 554614
rect -4298 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 372986 554614
rect 373222 554378 373306 554614
rect 373542 554378 408986 554614
rect 409222 554378 409306 554614
rect 409542 554378 444986 554614
rect 445222 554378 445306 554614
rect 445542 554378 480986 554614
rect 481222 554378 481306 554614
rect 481542 554378 516986 554614
rect 517222 554378 517306 554614
rect 517542 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 588222 554614
rect 588458 554378 588542 554614
rect 588778 554378 592650 554614
rect -8726 554294 592650 554378
rect -8726 554058 -4854 554294
rect -4618 554058 -4534 554294
rect -4298 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 372986 554294
rect 373222 554058 373306 554294
rect 373542 554058 408986 554294
rect 409222 554058 409306 554294
rect 409542 554058 444986 554294
rect 445222 554058 445306 554294
rect 445542 554058 480986 554294
rect 481222 554058 481306 554294
rect 481542 554058 516986 554294
rect 517222 554058 517306 554294
rect 517542 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 588222 554294
rect 588458 554058 588542 554294
rect 588778 554058 592650 554294
rect -8726 554026 592650 554058
rect -8726 550894 592650 550926
rect -8726 550658 -3894 550894
rect -3658 550658 -3574 550894
rect -3338 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 369266 550894
rect 369502 550658 369586 550894
rect 369822 550658 405266 550894
rect 405502 550658 405586 550894
rect 405822 550658 441266 550894
rect 441502 550658 441586 550894
rect 441822 550658 477266 550894
rect 477502 550658 477586 550894
rect 477822 550658 513266 550894
rect 513502 550658 513586 550894
rect 513822 550658 549266 550894
rect 549502 550658 549586 550894
rect 549822 550658 587262 550894
rect 587498 550658 587582 550894
rect 587818 550658 592650 550894
rect -8726 550574 592650 550658
rect -8726 550338 -3894 550574
rect -3658 550338 -3574 550574
rect -3338 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 369266 550574
rect 369502 550338 369586 550574
rect 369822 550338 405266 550574
rect 405502 550338 405586 550574
rect 405822 550338 441266 550574
rect 441502 550338 441586 550574
rect 441822 550338 477266 550574
rect 477502 550338 477586 550574
rect 477822 550338 513266 550574
rect 513502 550338 513586 550574
rect 513822 550338 549266 550574
rect 549502 550338 549586 550574
rect 549822 550338 587262 550574
rect 587498 550338 587582 550574
rect 587818 550338 592650 550574
rect -8726 550306 592650 550338
rect -8726 547174 592650 547206
rect -8726 546938 -2934 547174
rect -2698 546938 -2614 547174
rect -2378 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 39610 547174
rect 39846 546938 70330 547174
rect 70566 546938 101050 547174
rect 101286 546938 131770 547174
rect 132006 546938 162490 547174
rect 162726 546938 193210 547174
rect 193446 546938 223930 547174
rect 224166 546938 254650 547174
rect 254886 546938 285370 547174
rect 285606 546938 316090 547174
rect 316326 546938 346810 547174
rect 347046 546938 365546 547174
rect 365782 546938 365866 547174
rect 366102 546938 401546 547174
rect 401782 546938 401866 547174
rect 402102 546938 437546 547174
rect 437782 546938 437866 547174
rect 438102 546938 473546 547174
rect 473782 546938 473866 547174
rect 474102 546938 509546 547174
rect 509782 546938 509866 547174
rect 510102 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 586302 547174
rect 586538 546938 586622 547174
rect 586858 546938 592650 547174
rect -8726 546854 592650 546938
rect -8726 546618 -2934 546854
rect -2698 546618 -2614 546854
rect -2378 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 39610 546854
rect 39846 546618 70330 546854
rect 70566 546618 101050 546854
rect 101286 546618 131770 546854
rect 132006 546618 162490 546854
rect 162726 546618 193210 546854
rect 193446 546618 223930 546854
rect 224166 546618 254650 546854
rect 254886 546618 285370 546854
rect 285606 546618 316090 546854
rect 316326 546618 346810 546854
rect 347046 546618 365546 546854
rect 365782 546618 365866 546854
rect 366102 546618 401546 546854
rect 401782 546618 401866 546854
rect 402102 546618 437546 546854
rect 437782 546618 437866 546854
rect 438102 546618 473546 546854
rect 473782 546618 473866 546854
rect 474102 546618 509546 546854
rect 509782 546618 509866 546854
rect 510102 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 586302 546854
rect 586538 546618 586622 546854
rect 586858 546618 592650 546854
rect -8726 546586 592650 546618
rect -8726 543454 592650 543486
rect -8726 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 24250 543454
rect 24486 543218 54970 543454
rect 55206 543218 85690 543454
rect 85926 543218 116410 543454
rect 116646 543218 147130 543454
rect 147366 543218 177850 543454
rect 178086 543218 208570 543454
rect 208806 543218 239290 543454
rect 239526 543218 270010 543454
rect 270246 543218 300730 543454
rect 300966 543218 331450 543454
rect 331686 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 592650 543454
rect -8726 543134 592650 543218
rect -8726 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 24250 543134
rect 24486 542898 54970 543134
rect 55206 542898 85690 543134
rect 85926 542898 116410 543134
rect 116646 542898 147130 543134
rect 147366 542898 177850 543134
rect 178086 542898 208570 543134
rect 208806 542898 239290 543134
rect 239526 542898 270010 543134
rect 270246 542898 300730 543134
rect 300966 542898 331450 543134
rect 331686 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 592650 543134
rect -8726 542866 592650 542898
rect -8726 533494 592650 533526
rect -8726 533258 -8694 533494
rect -8458 533258 -8374 533494
rect -8138 533258 27866 533494
rect 28102 533258 28186 533494
rect 28422 533258 387866 533494
rect 388102 533258 388186 533494
rect 388422 533258 423866 533494
rect 424102 533258 424186 533494
rect 424422 533258 459866 533494
rect 460102 533258 460186 533494
rect 460422 533258 495866 533494
rect 496102 533258 496186 533494
rect 496422 533258 531866 533494
rect 532102 533258 532186 533494
rect 532422 533258 567866 533494
rect 568102 533258 568186 533494
rect 568422 533258 592062 533494
rect 592298 533258 592382 533494
rect 592618 533258 592650 533494
rect -8726 533174 592650 533258
rect -8726 532938 -8694 533174
rect -8458 532938 -8374 533174
rect -8138 532938 27866 533174
rect 28102 532938 28186 533174
rect 28422 532938 387866 533174
rect 388102 532938 388186 533174
rect 388422 532938 423866 533174
rect 424102 532938 424186 533174
rect 424422 532938 459866 533174
rect 460102 532938 460186 533174
rect 460422 532938 495866 533174
rect 496102 532938 496186 533174
rect 496422 532938 531866 533174
rect 532102 532938 532186 533174
rect 532422 532938 567866 533174
rect 568102 532938 568186 533174
rect 568422 532938 592062 533174
rect 592298 532938 592382 533174
rect 592618 532938 592650 533174
rect -8726 532906 592650 532938
rect -8726 529774 592650 529806
rect -8726 529538 -7734 529774
rect -7498 529538 -7414 529774
rect -7178 529538 384146 529774
rect 384382 529538 384466 529774
rect 384702 529538 420146 529774
rect 420382 529538 420466 529774
rect 420702 529538 456146 529774
rect 456382 529538 456466 529774
rect 456702 529538 492146 529774
rect 492382 529538 492466 529774
rect 492702 529538 528146 529774
rect 528382 529538 528466 529774
rect 528702 529538 564146 529774
rect 564382 529538 564466 529774
rect 564702 529538 591102 529774
rect 591338 529538 591422 529774
rect 591658 529538 592650 529774
rect -8726 529454 592650 529538
rect -8726 529218 -7734 529454
rect -7498 529218 -7414 529454
rect -7178 529218 384146 529454
rect 384382 529218 384466 529454
rect 384702 529218 420146 529454
rect 420382 529218 420466 529454
rect 420702 529218 456146 529454
rect 456382 529218 456466 529454
rect 456702 529218 492146 529454
rect 492382 529218 492466 529454
rect 492702 529218 528146 529454
rect 528382 529218 528466 529454
rect 528702 529218 564146 529454
rect 564382 529218 564466 529454
rect 564702 529218 591102 529454
rect 591338 529218 591422 529454
rect 591658 529218 592650 529454
rect -8726 529186 592650 529218
rect -8726 526054 592650 526086
rect -8726 525818 -6774 526054
rect -6538 525818 -6454 526054
rect -6218 525818 20426 526054
rect 20662 525818 20746 526054
rect 20982 525818 380426 526054
rect 380662 525818 380746 526054
rect 380982 525818 416426 526054
rect 416662 525818 416746 526054
rect 416982 525818 452426 526054
rect 452662 525818 452746 526054
rect 452982 525818 488426 526054
rect 488662 525818 488746 526054
rect 488982 525818 524426 526054
rect 524662 525818 524746 526054
rect 524982 525818 560426 526054
rect 560662 525818 560746 526054
rect 560982 525818 590142 526054
rect 590378 525818 590462 526054
rect 590698 525818 592650 526054
rect -8726 525734 592650 525818
rect -8726 525498 -6774 525734
rect -6538 525498 -6454 525734
rect -6218 525498 20426 525734
rect 20662 525498 20746 525734
rect 20982 525498 380426 525734
rect 380662 525498 380746 525734
rect 380982 525498 416426 525734
rect 416662 525498 416746 525734
rect 416982 525498 452426 525734
rect 452662 525498 452746 525734
rect 452982 525498 488426 525734
rect 488662 525498 488746 525734
rect 488982 525498 524426 525734
rect 524662 525498 524746 525734
rect 524982 525498 560426 525734
rect 560662 525498 560746 525734
rect 560982 525498 590142 525734
rect 590378 525498 590462 525734
rect 590698 525498 592650 525734
rect -8726 525466 592650 525498
rect -8726 522334 592650 522366
rect -8726 522098 -5814 522334
rect -5578 522098 -5494 522334
rect -5258 522098 16706 522334
rect 16942 522098 17026 522334
rect 17262 522098 376706 522334
rect 376942 522098 377026 522334
rect 377262 522098 412706 522334
rect 412942 522098 413026 522334
rect 413262 522098 448706 522334
rect 448942 522098 449026 522334
rect 449262 522098 484706 522334
rect 484942 522098 485026 522334
rect 485262 522098 520706 522334
rect 520942 522098 521026 522334
rect 521262 522098 556706 522334
rect 556942 522098 557026 522334
rect 557262 522098 589182 522334
rect 589418 522098 589502 522334
rect 589738 522098 592650 522334
rect -8726 522014 592650 522098
rect -8726 521778 -5814 522014
rect -5578 521778 -5494 522014
rect -5258 521778 16706 522014
rect 16942 521778 17026 522014
rect 17262 521778 376706 522014
rect 376942 521778 377026 522014
rect 377262 521778 412706 522014
rect 412942 521778 413026 522014
rect 413262 521778 448706 522014
rect 448942 521778 449026 522014
rect 449262 521778 484706 522014
rect 484942 521778 485026 522014
rect 485262 521778 520706 522014
rect 520942 521778 521026 522014
rect 521262 521778 556706 522014
rect 556942 521778 557026 522014
rect 557262 521778 589182 522014
rect 589418 521778 589502 522014
rect 589738 521778 592650 522014
rect -8726 521746 592650 521778
rect -8726 518614 592650 518646
rect -8726 518378 -4854 518614
rect -4618 518378 -4534 518614
rect -4298 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 372986 518614
rect 373222 518378 373306 518614
rect 373542 518378 408986 518614
rect 409222 518378 409306 518614
rect 409542 518378 444986 518614
rect 445222 518378 445306 518614
rect 445542 518378 480986 518614
rect 481222 518378 481306 518614
rect 481542 518378 516986 518614
rect 517222 518378 517306 518614
rect 517542 518378 552986 518614
rect 553222 518378 553306 518614
rect 553542 518378 588222 518614
rect 588458 518378 588542 518614
rect 588778 518378 592650 518614
rect -8726 518294 592650 518378
rect -8726 518058 -4854 518294
rect -4618 518058 -4534 518294
rect -4298 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 372986 518294
rect 373222 518058 373306 518294
rect 373542 518058 408986 518294
rect 409222 518058 409306 518294
rect 409542 518058 444986 518294
rect 445222 518058 445306 518294
rect 445542 518058 480986 518294
rect 481222 518058 481306 518294
rect 481542 518058 516986 518294
rect 517222 518058 517306 518294
rect 517542 518058 552986 518294
rect 553222 518058 553306 518294
rect 553542 518058 588222 518294
rect 588458 518058 588542 518294
rect 588778 518058 592650 518294
rect -8726 518026 592650 518058
rect -8726 514894 592650 514926
rect -8726 514658 -3894 514894
rect -3658 514658 -3574 514894
rect -3338 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 369266 514894
rect 369502 514658 369586 514894
rect 369822 514658 405266 514894
rect 405502 514658 405586 514894
rect 405822 514658 441266 514894
rect 441502 514658 441586 514894
rect 441822 514658 477266 514894
rect 477502 514658 477586 514894
rect 477822 514658 513266 514894
rect 513502 514658 513586 514894
rect 513822 514658 549266 514894
rect 549502 514658 549586 514894
rect 549822 514658 587262 514894
rect 587498 514658 587582 514894
rect 587818 514658 592650 514894
rect -8726 514574 592650 514658
rect -8726 514338 -3894 514574
rect -3658 514338 -3574 514574
rect -3338 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 369266 514574
rect 369502 514338 369586 514574
rect 369822 514338 405266 514574
rect 405502 514338 405586 514574
rect 405822 514338 441266 514574
rect 441502 514338 441586 514574
rect 441822 514338 477266 514574
rect 477502 514338 477586 514574
rect 477822 514338 513266 514574
rect 513502 514338 513586 514574
rect 513822 514338 549266 514574
rect 549502 514338 549586 514574
rect 549822 514338 587262 514574
rect 587498 514338 587582 514574
rect 587818 514338 592650 514574
rect -8726 514306 592650 514338
rect -8726 511174 592650 511206
rect -8726 510938 -2934 511174
rect -2698 510938 -2614 511174
rect -2378 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 39610 511174
rect 39846 510938 70330 511174
rect 70566 510938 101050 511174
rect 101286 510938 131770 511174
rect 132006 510938 162490 511174
rect 162726 510938 193210 511174
rect 193446 510938 223930 511174
rect 224166 510938 254650 511174
rect 254886 510938 285370 511174
rect 285606 510938 316090 511174
rect 316326 510938 346810 511174
rect 347046 510938 365546 511174
rect 365782 510938 365866 511174
rect 366102 510938 401546 511174
rect 401782 510938 401866 511174
rect 402102 510938 437546 511174
rect 437782 510938 437866 511174
rect 438102 510938 453424 511174
rect 453660 510938 455862 511174
rect 456098 510938 458300 511174
rect 458536 510938 460738 511174
rect 460974 510938 473546 511174
rect 473782 510938 473866 511174
rect 474102 510938 483424 511174
rect 483660 510938 485862 511174
rect 486098 510938 488300 511174
rect 488536 510938 490738 511174
rect 490974 510938 509546 511174
rect 509782 510938 509866 511174
rect 510102 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 586302 511174
rect 586538 510938 586622 511174
rect 586858 510938 592650 511174
rect -8726 510854 592650 510938
rect -8726 510618 -2934 510854
rect -2698 510618 -2614 510854
rect -2378 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 39610 510854
rect 39846 510618 70330 510854
rect 70566 510618 101050 510854
rect 101286 510618 131770 510854
rect 132006 510618 162490 510854
rect 162726 510618 193210 510854
rect 193446 510618 223930 510854
rect 224166 510618 254650 510854
rect 254886 510618 285370 510854
rect 285606 510618 316090 510854
rect 316326 510618 346810 510854
rect 347046 510618 365546 510854
rect 365782 510618 365866 510854
rect 366102 510618 401546 510854
rect 401782 510618 401866 510854
rect 402102 510618 437546 510854
rect 437782 510618 437866 510854
rect 438102 510618 453424 510854
rect 453660 510618 455862 510854
rect 456098 510618 458300 510854
rect 458536 510618 460738 510854
rect 460974 510618 473546 510854
rect 473782 510618 473866 510854
rect 474102 510618 483424 510854
rect 483660 510618 485862 510854
rect 486098 510618 488300 510854
rect 488536 510618 490738 510854
rect 490974 510618 509546 510854
rect 509782 510618 509866 510854
rect 510102 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 586302 510854
rect 586538 510618 586622 510854
rect 586858 510618 592650 510854
rect -8726 510586 592650 510618
rect -8726 507454 592650 507486
rect -8726 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 24250 507454
rect 24486 507218 54970 507454
rect 55206 507218 85690 507454
rect 85926 507218 116410 507454
rect 116646 507218 147130 507454
rect 147366 507218 177850 507454
rect 178086 507218 208570 507454
rect 208806 507218 239290 507454
rect 239526 507218 270010 507454
rect 270246 507218 300730 507454
rect 300966 507218 331450 507454
rect 331686 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 452205 507454
rect 452441 507218 454643 507454
rect 454879 507218 457081 507454
rect 457317 507218 459519 507454
rect 459755 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 482205 507454
rect 482441 507218 484643 507454
rect 484879 507218 487081 507454
rect 487317 507218 489519 507454
rect 489755 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 592650 507454
rect -8726 507134 592650 507218
rect -8726 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 24250 507134
rect 24486 506898 54970 507134
rect 55206 506898 85690 507134
rect 85926 506898 116410 507134
rect 116646 506898 147130 507134
rect 147366 506898 177850 507134
rect 178086 506898 208570 507134
rect 208806 506898 239290 507134
rect 239526 506898 270010 507134
rect 270246 506898 300730 507134
rect 300966 506898 331450 507134
rect 331686 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 452205 507134
rect 452441 506898 454643 507134
rect 454879 506898 457081 507134
rect 457317 506898 459519 507134
rect 459755 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 482205 507134
rect 482441 506898 484643 507134
rect 484879 506898 487081 507134
rect 487317 506898 489519 507134
rect 489755 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 592650 507134
rect -8726 506866 592650 506898
rect -8726 497494 592650 497526
rect -8726 497258 -8694 497494
rect -8458 497258 -8374 497494
rect -8138 497258 27866 497494
rect 28102 497258 28186 497494
rect 28422 497258 387866 497494
rect 388102 497258 388186 497494
rect 388422 497258 423866 497494
rect 424102 497258 424186 497494
rect 424422 497258 459866 497494
rect 460102 497258 460186 497494
rect 460422 497258 495866 497494
rect 496102 497258 496186 497494
rect 496422 497258 531866 497494
rect 532102 497258 532186 497494
rect 532422 497258 567866 497494
rect 568102 497258 568186 497494
rect 568422 497258 592062 497494
rect 592298 497258 592382 497494
rect 592618 497258 592650 497494
rect -8726 497174 592650 497258
rect -8726 496938 -8694 497174
rect -8458 496938 -8374 497174
rect -8138 496938 27866 497174
rect 28102 496938 28186 497174
rect 28422 496938 387866 497174
rect 388102 496938 388186 497174
rect 388422 496938 423866 497174
rect 424102 496938 424186 497174
rect 424422 496938 459866 497174
rect 460102 496938 460186 497174
rect 460422 496938 495866 497174
rect 496102 496938 496186 497174
rect 496422 496938 531866 497174
rect 532102 496938 532186 497174
rect 532422 496938 567866 497174
rect 568102 496938 568186 497174
rect 568422 496938 592062 497174
rect 592298 496938 592382 497174
rect 592618 496938 592650 497174
rect -8726 496906 592650 496938
rect -8726 493774 592650 493806
rect -8726 493538 -7734 493774
rect -7498 493538 -7414 493774
rect -7178 493538 384146 493774
rect 384382 493538 384466 493774
rect 384702 493538 420146 493774
rect 420382 493538 420466 493774
rect 420702 493538 456146 493774
rect 456382 493538 456466 493774
rect 456702 493538 492146 493774
rect 492382 493538 492466 493774
rect 492702 493538 528146 493774
rect 528382 493538 528466 493774
rect 528702 493538 564146 493774
rect 564382 493538 564466 493774
rect 564702 493538 591102 493774
rect 591338 493538 591422 493774
rect 591658 493538 592650 493774
rect -8726 493454 592650 493538
rect -8726 493218 -7734 493454
rect -7498 493218 -7414 493454
rect -7178 493218 384146 493454
rect 384382 493218 384466 493454
rect 384702 493218 420146 493454
rect 420382 493218 420466 493454
rect 420702 493218 456146 493454
rect 456382 493218 456466 493454
rect 456702 493218 492146 493454
rect 492382 493218 492466 493454
rect 492702 493218 528146 493454
rect 528382 493218 528466 493454
rect 528702 493218 564146 493454
rect 564382 493218 564466 493454
rect 564702 493218 591102 493454
rect 591338 493218 591422 493454
rect 591658 493218 592650 493454
rect -8726 493186 592650 493218
rect -8726 490054 592650 490086
rect -8726 489818 -6774 490054
rect -6538 489818 -6454 490054
rect -6218 489818 20426 490054
rect 20662 489818 20746 490054
rect 20982 489818 380426 490054
rect 380662 489818 380746 490054
rect 380982 489818 416426 490054
rect 416662 489818 416746 490054
rect 416982 489818 452426 490054
rect 452662 489818 452746 490054
rect 452982 489818 488426 490054
rect 488662 489818 488746 490054
rect 488982 489818 524426 490054
rect 524662 489818 524746 490054
rect 524982 489818 560426 490054
rect 560662 489818 560746 490054
rect 560982 489818 590142 490054
rect 590378 489818 590462 490054
rect 590698 489818 592650 490054
rect -8726 489734 592650 489818
rect -8726 489498 -6774 489734
rect -6538 489498 -6454 489734
rect -6218 489498 20426 489734
rect 20662 489498 20746 489734
rect 20982 489498 380426 489734
rect 380662 489498 380746 489734
rect 380982 489498 416426 489734
rect 416662 489498 416746 489734
rect 416982 489498 452426 489734
rect 452662 489498 452746 489734
rect 452982 489498 488426 489734
rect 488662 489498 488746 489734
rect 488982 489498 524426 489734
rect 524662 489498 524746 489734
rect 524982 489498 560426 489734
rect 560662 489498 560746 489734
rect 560982 489498 590142 489734
rect 590378 489498 590462 489734
rect 590698 489498 592650 489734
rect -8726 489466 592650 489498
rect -8726 486334 592650 486366
rect -8726 486098 -5814 486334
rect -5578 486098 -5494 486334
rect -5258 486098 16706 486334
rect 16942 486098 17026 486334
rect 17262 486098 376706 486334
rect 376942 486098 377026 486334
rect 377262 486098 412706 486334
rect 412942 486098 413026 486334
rect 413262 486098 448706 486334
rect 448942 486098 449026 486334
rect 449262 486098 484706 486334
rect 484942 486098 485026 486334
rect 485262 486098 520706 486334
rect 520942 486098 521026 486334
rect 521262 486098 556706 486334
rect 556942 486098 557026 486334
rect 557262 486098 589182 486334
rect 589418 486098 589502 486334
rect 589738 486098 592650 486334
rect -8726 486014 592650 486098
rect -8726 485778 -5814 486014
rect -5578 485778 -5494 486014
rect -5258 485778 16706 486014
rect 16942 485778 17026 486014
rect 17262 485778 376706 486014
rect 376942 485778 377026 486014
rect 377262 485778 412706 486014
rect 412942 485778 413026 486014
rect 413262 485778 448706 486014
rect 448942 485778 449026 486014
rect 449262 485778 484706 486014
rect 484942 485778 485026 486014
rect 485262 485778 520706 486014
rect 520942 485778 521026 486014
rect 521262 485778 556706 486014
rect 556942 485778 557026 486014
rect 557262 485778 589182 486014
rect 589418 485778 589502 486014
rect 589738 485778 592650 486014
rect -8726 485746 592650 485778
rect -8726 482614 592650 482646
rect -8726 482378 -4854 482614
rect -4618 482378 -4534 482614
rect -4298 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 372986 482614
rect 373222 482378 373306 482614
rect 373542 482378 408986 482614
rect 409222 482378 409306 482614
rect 409542 482378 444986 482614
rect 445222 482378 445306 482614
rect 445542 482378 480986 482614
rect 481222 482378 481306 482614
rect 481542 482378 516986 482614
rect 517222 482378 517306 482614
rect 517542 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 588222 482614
rect 588458 482378 588542 482614
rect 588778 482378 592650 482614
rect -8726 482294 592650 482378
rect -8726 482058 -4854 482294
rect -4618 482058 -4534 482294
rect -4298 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 372986 482294
rect 373222 482058 373306 482294
rect 373542 482058 408986 482294
rect 409222 482058 409306 482294
rect 409542 482058 444986 482294
rect 445222 482058 445306 482294
rect 445542 482058 480986 482294
rect 481222 482058 481306 482294
rect 481542 482058 516986 482294
rect 517222 482058 517306 482294
rect 517542 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 588222 482294
rect 588458 482058 588542 482294
rect 588778 482058 592650 482294
rect -8726 482026 592650 482058
rect -8726 478894 592650 478926
rect -8726 478658 -3894 478894
rect -3658 478658 -3574 478894
rect -3338 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 369266 478894
rect 369502 478658 369586 478894
rect 369822 478658 405266 478894
rect 405502 478658 405586 478894
rect 405822 478658 441266 478894
rect 441502 478658 441586 478894
rect 441822 478658 477266 478894
rect 477502 478658 477586 478894
rect 477822 478658 513266 478894
rect 513502 478658 513586 478894
rect 513822 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 587262 478894
rect 587498 478658 587582 478894
rect 587818 478658 592650 478894
rect -8726 478574 592650 478658
rect -8726 478338 -3894 478574
rect -3658 478338 -3574 478574
rect -3338 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 369266 478574
rect 369502 478338 369586 478574
rect 369822 478338 405266 478574
rect 405502 478338 405586 478574
rect 405822 478338 441266 478574
rect 441502 478338 441586 478574
rect 441822 478338 477266 478574
rect 477502 478338 477586 478574
rect 477822 478338 513266 478574
rect 513502 478338 513586 478574
rect 513822 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 587262 478574
rect 587498 478338 587582 478574
rect 587818 478338 592650 478574
rect -8726 478306 592650 478338
rect -8726 475174 592650 475206
rect -8726 474938 -2934 475174
rect -2698 474938 -2614 475174
rect -2378 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 39610 475174
rect 39846 474938 70330 475174
rect 70566 474938 101050 475174
rect 101286 474938 131770 475174
rect 132006 474938 162490 475174
rect 162726 474938 193210 475174
rect 193446 474938 223930 475174
rect 224166 474938 254650 475174
rect 254886 474938 285370 475174
rect 285606 474938 316090 475174
rect 316326 474938 346810 475174
rect 347046 474938 365546 475174
rect 365782 474938 365866 475174
rect 366102 474938 401546 475174
rect 401782 474938 401866 475174
rect 402102 474938 437546 475174
rect 437782 474938 437866 475174
rect 438102 474938 473546 475174
rect 473782 474938 473866 475174
rect 474102 474938 509546 475174
rect 509782 474938 509866 475174
rect 510102 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 586302 475174
rect 586538 474938 586622 475174
rect 586858 474938 592650 475174
rect -8726 474854 592650 474938
rect -8726 474618 -2934 474854
rect -2698 474618 -2614 474854
rect -2378 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 39610 474854
rect 39846 474618 70330 474854
rect 70566 474618 101050 474854
rect 101286 474618 131770 474854
rect 132006 474618 162490 474854
rect 162726 474618 193210 474854
rect 193446 474618 223930 474854
rect 224166 474618 254650 474854
rect 254886 474618 285370 474854
rect 285606 474618 316090 474854
rect 316326 474618 346810 474854
rect 347046 474618 365546 474854
rect 365782 474618 365866 474854
rect 366102 474618 401546 474854
rect 401782 474618 401866 474854
rect 402102 474618 437546 474854
rect 437782 474618 437866 474854
rect 438102 474618 473546 474854
rect 473782 474618 473866 474854
rect 474102 474618 509546 474854
rect 509782 474618 509866 474854
rect 510102 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 586302 474854
rect 586538 474618 586622 474854
rect 586858 474618 592650 474854
rect -8726 474586 592650 474618
rect -8726 471454 592650 471486
rect -8726 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 24250 471454
rect 24486 471218 54970 471454
rect 55206 471218 85690 471454
rect 85926 471218 116410 471454
rect 116646 471218 147130 471454
rect 147366 471218 177850 471454
rect 178086 471218 208570 471454
rect 208806 471218 239290 471454
rect 239526 471218 270010 471454
rect 270246 471218 300730 471454
rect 300966 471218 331450 471454
rect 331686 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 592650 471454
rect -8726 471134 592650 471218
rect -8726 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 24250 471134
rect 24486 470898 54970 471134
rect 55206 470898 85690 471134
rect 85926 470898 116410 471134
rect 116646 470898 147130 471134
rect 147366 470898 177850 471134
rect 178086 470898 208570 471134
rect 208806 470898 239290 471134
rect 239526 470898 270010 471134
rect 270246 470898 300730 471134
rect 300966 470898 331450 471134
rect 331686 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 592650 471134
rect -8726 470866 592650 470898
rect -8726 461494 592650 461526
rect -8726 461258 -8694 461494
rect -8458 461258 -8374 461494
rect -8138 461258 27866 461494
rect 28102 461258 28186 461494
rect 28422 461258 387866 461494
rect 388102 461258 388186 461494
rect 388422 461258 423866 461494
rect 424102 461258 424186 461494
rect 424422 461258 459866 461494
rect 460102 461258 460186 461494
rect 460422 461258 495866 461494
rect 496102 461258 496186 461494
rect 496422 461258 531866 461494
rect 532102 461258 532186 461494
rect 532422 461258 567866 461494
rect 568102 461258 568186 461494
rect 568422 461258 592062 461494
rect 592298 461258 592382 461494
rect 592618 461258 592650 461494
rect -8726 461174 592650 461258
rect -8726 460938 -8694 461174
rect -8458 460938 -8374 461174
rect -8138 460938 27866 461174
rect 28102 460938 28186 461174
rect 28422 460938 387866 461174
rect 388102 460938 388186 461174
rect 388422 460938 423866 461174
rect 424102 460938 424186 461174
rect 424422 460938 459866 461174
rect 460102 460938 460186 461174
rect 460422 460938 495866 461174
rect 496102 460938 496186 461174
rect 496422 460938 531866 461174
rect 532102 460938 532186 461174
rect 532422 460938 567866 461174
rect 568102 460938 568186 461174
rect 568422 460938 592062 461174
rect 592298 460938 592382 461174
rect 592618 460938 592650 461174
rect -8726 460906 592650 460938
rect -8726 457774 592650 457806
rect -8726 457538 -7734 457774
rect -7498 457538 -7414 457774
rect -7178 457538 384146 457774
rect 384382 457538 384466 457774
rect 384702 457538 420146 457774
rect 420382 457538 420466 457774
rect 420702 457538 456146 457774
rect 456382 457538 456466 457774
rect 456702 457538 492146 457774
rect 492382 457538 492466 457774
rect 492702 457538 528146 457774
rect 528382 457538 528466 457774
rect 528702 457538 564146 457774
rect 564382 457538 564466 457774
rect 564702 457538 591102 457774
rect 591338 457538 591422 457774
rect 591658 457538 592650 457774
rect -8726 457454 592650 457538
rect -8726 457218 -7734 457454
rect -7498 457218 -7414 457454
rect -7178 457218 384146 457454
rect 384382 457218 384466 457454
rect 384702 457218 420146 457454
rect 420382 457218 420466 457454
rect 420702 457218 456146 457454
rect 456382 457218 456466 457454
rect 456702 457218 492146 457454
rect 492382 457218 492466 457454
rect 492702 457218 528146 457454
rect 528382 457218 528466 457454
rect 528702 457218 564146 457454
rect 564382 457218 564466 457454
rect 564702 457218 591102 457454
rect 591338 457218 591422 457454
rect 591658 457218 592650 457454
rect -8726 457186 592650 457218
rect -8726 454054 592650 454086
rect -8726 453818 -6774 454054
rect -6538 453818 -6454 454054
rect -6218 453818 20426 454054
rect 20662 453818 20746 454054
rect 20982 453818 380426 454054
rect 380662 453818 380746 454054
rect 380982 453818 416426 454054
rect 416662 453818 416746 454054
rect 416982 453818 452426 454054
rect 452662 453818 452746 454054
rect 452982 454007 524426 454054
rect 452982 453818 488426 454007
rect -8726 453771 488426 453818
rect 488662 453771 488746 454007
rect 488982 453818 524426 454007
rect 524662 453818 524746 454054
rect 524982 453818 560426 454054
rect 560662 453818 560746 454054
rect 560982 453818 590142 454054
rect 590378 453818 590462 454054
rect 590698 453818 592650 454054
rect 488982 453771 592650 453818
rect -8726 453734 592650 453771
rect -8726 453498 -6774 453734
rect -6538 453498 -6454 453734
rect -6218 453498 20426 453734
rect 20662 453498 20746 453734
rect 20982 453498 380426 453734
rect 380662 453498 380746 453734
rect 380982 453498 416426 453734
rect 416662 453498 416746 453734
rect 416982 453498 452426 453734
rect 452662 453498 452746 453734
rect 452982 453498 524426 453734
rect 524662 453498 524746 453734
rect 524982 453498 560426 453734
rect 560662 453498 560746 453734
rect 560982 453498 590142 453734
rect 590378 453498 590462 453734
rect 590698 453498 592650 453734
rect -8726 453466 592650 453498
rect -8726 450334 592650 450366
rect -8726 450098 -5814 450334
rect -5578 450098 -5494 450334
rect -5258 450098 16706 450334
rect 16942 450098 17026 450334
rect 17262 450098 376706 450334
rect 376942 450098 377026 450334
rect 377262 450098 412706 450334
rect 412942 450098 413026 450334
rect 413262 450098 448706 450334
rect 448942 450098 449026 450334
rect 449262 450098 484706 450334
rect 484942 450098 485026 450334
rect 485262 450098 520706 450334
rect 520942 450098 521026 450334
rect 521262 450098 556706 450334
rect 556942 450098 557026 450334
rect 557262 450098 589182 450334
rect 589418 450098 589502 450334
rect 589738 450098 592650 450334
rect -8726 450014 592650 450098
rect -8726 449778 -5814 450014
rect -5578 449778 -5494 450014
rect -5258 449778 16706 450014
rect 16942 449778 17026 450014
rect 17262 449778 376706 450014
rect 376942 449778 377026 450014
rect 377262 449778 412706 450014
rect 412942 449778 413026 450014
rect 413262 449778 448706 450014
rect 448942 449778 449026 450014
rect 449262 449778 484706 450014
rect 484942 449778 485026 450014
rect 485262 449778 520706 450014
rect 520942 449778 521026 450014
rect 521262 449778 556706 450014
rect 556942 449778 557026 450014
rect 557262 449778 589182 450014
rect 589418 449778 589502 450014
rect 589738 449778 592650 450014
rect -8726 449746 592650 449778
rect -8726 446614 592650 446646
rect -8726 446378 -4854 446614
rect -4618 446378 -4534 446614
rect -4298 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 372986 446614
rect 373222 446378 373306 446614
rect 373542 446378 408986 446614
rect 409222 446378 409306 446614
rect 409542 446378 444986 446614
rect 445222 446378 445306 446614
rect 445542 446378 516986 446614
rect 517222 446378 517306 446614
rect 517542 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 588222 446614
rect 588458 446378 588542 446614
rect 588778 446378 592650 446614
rect -8726 446294 592650 446378
rect -8726 446058 -4854 446294
rect -4618 446058 -4534 446294
rect -4298 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 372986 446294
rect 373222 446058 373306 446294
rect 373542 446058 408986 446294
rect 409222 446058 409306 446294
rect 409542 446058 444986 446294
rect 445222 446058 445306 446294
rect 445542 446058 516986 446294
rect 517222 446058 517306 446294
rect 517542 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 588222 446294
rect 588458 446058 588542 446294
rect 588778 446058 592650 446294
rect -8726 446026 592650 446058
rect -8726 442894 592650 442926
rect -8726 442658 -3894 442894
rect -3658 442658 -3574 442894
rect -3338 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 369266 442894
rect 369502 442658 369586 442894
rect 369822 442658 405266 442894
rect 405502 442658 405586 442894
rect 405822 442658 477266 442894
rect 477502 442658 477586 442894
rect 477822 442658 513266 442894
rect 513502 442658 513586 442894
rect 513822 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 587262 442894
rect 587498 442658 587582 442894
rect 587818 442658 592650 442894
rect -8726 442574 592650 442658
rect -8726 442338 -3894 442574
rect -3658 442338 -3574 442574
rect -3338 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 369266 442574
rect 369502 442338 369586 442574
rect 369822 442338 405266 442574
rect 405502 442338 405586 442574
rect 405822 442338 477266 442574
rect 477502 442338 477586 442574
rect 477822 442338 513266 442574
rect 513502 442338 513586 442574
rect 513822 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 587262 442574
rect 587498 442338 587582 442574
rect 587818 442338 592650 442574
rect -8726 442306 592650 442338
rect -8726 439174 592650 439206
rect -8726 438938 -2934 439174
rect -2698 438938 -2614 439174
rect -2378 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 39610 439174
rect 39846 438938 70330 439174
rect 70566 438938 101050 439174
rect 101286 438938 131770 439174
rect 132006 438938 162490 439174
rect 162726 438938 193210 439174
rect 193446 438938 223930 439174
rect 224166 438938 254650 439174
rect 254886 438938 285370 439174
rect 285606 438938 316090 439174
rect 316326 438938 346810 439174
rect 347046 438938 365546 439174
rect 365782 438938 365866 439174
rect 366102 438938 401546 439174
rect 401782 438938 401866 439174
rect 402102 438938 426666 439174
rect 426902 438938 432347 439174
rect 432583 438938 438028 439174
rect 438264 438938 443709 439174
rect 443945 438938 475930 439174
rect 476166 438938 480875 439174
rect 481111 438938 485820 439174
rect 486056 438938 490765 439174
rect 491001 438938 509546 439174
rect 509782 438938 509866 439174
rect 510102 438938 529426 439174
rect 529662 438938 537867 439174
rect 538103 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 546308 439174
rect 546544 438938 554749 439174
rect 554985 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 586302 439174
rect 586538 438938 586622 439174
rect 586858 438938 592650 439174
rect -8726 438854 592650 438938
rect -8726 438618 -2934 438854
rect -2698 438618 -2614 438854
rect -2378 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 39610 438854
rect 39846 438618 70330 438854
rect 70566 438618 101050 438854
rect 101286 438618 131770 438854
rect 132006 438618 162490 438854
rect 162726 438618 193210 438854
rect 193446 438618 223930 438854
rect 224166 438618 254650 438854
rect 254886 438618 285370 438854
rect 285606 438618 316090 438854
rect 316326 438618 346810 438854
rect 347046 438618 365546 438854
rect 365782 438618 365866 438854
rect 366102 438618 401546 438854
rect 401782 438618 401866 438854
rect 402102 438618 426666 438854
rect 426902 438618 432347 438854
rect 432583 438618 438028 438854
rect 438264 438618 443709 438854
rect 443945 438618 475930 438854
rect 476166 438618 480875 438854
rect 481111 438618 485820 438854
rect 486056 438618 490765 438854
rect 491001 438618 509546 438854
rect 509782 438618 509866 438854
rect 510102 438618 529426 438854
rect 529662 438618 537867 438854
rect 538103 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 546308 438854
rect 546544 438618 554749 438854
rect 554985 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 586302 438854
rect 586538 438618 586622 438854
rect 586858 438618 592650 438854
rect -8726 438586 592650 438618
rect -8726 435454 592650 435486
rect -8726 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 24250 435454
rect 24486 435218 54970 435454
rect 55206 435218 85690 435454
rect 85926 435218 116410 435454
rect 116646 435218 147130 435454
rect 147366 435218 177850 435454
rect 178086 435218 208570 435454
rect 208806 435218 239290 435454
rect 239526 435218 270010 435454
rect 270246 435218 300730 435454
rect 300966 435218 331450 435454
rect 331686 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 423826 435454
rect 424062 435218 429507 435454
rect 429743 435218 435188 435454
rect 435424 435218 440869 435454
rect 441105 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 473458 435454
rect 473694 435218 478403 435454
rect 478639 435218 483348 435454
rect 483584 435218 488293 435454
rect 488529 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 525206 435454
rect 525442 435218 533647 435454
rect 533883 435218 542088 435454
rect 542324 435218 550529 435454
rect 550765 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 592650 435454
rect -8726 435134 592650 435218
rect -8726 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 24250 435134
rect 24486 434898 54970 435134
rect 55206 434898 85690 435134
rect 85926 434898 116410 435134
rect 116646 434898 147130 435134
rect 147366 434898 177850 435134
rect 178086 434898 208570 435134
rect 208806 434898 239290 435134
rect 239526 434898 270010 435134
rect 270246 434898 300730 435134
rect 300966 434898 331450 435134
rect 331686 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 423826 435134
rect 424062 434898 429507 435134
rect 429743 434898 435188 435134
rect 435424 434898 440869 435134
rect 441105 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 473458 435134
rect 473694 434898 478403 435134
rect 478639 434898 483348 435134
rect 483584 434898 488293 435134
rect 488529 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 525206 435134
rect 525442 434898 533647 435134
rect 533883 434898 542088 435134
rect 542324 434898 550529 435134
rect 550765 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 592650 435134
rect -8726 434866 592650 434898
rect -8726 425494 592650 425526
rect -8726 425258 -8694 425494
rect -8458 425258 -8374 425494
rect -8138 425258 27866 425494
rect 28102 425258 28186 425494
rect 28422 425258 387866 425494
rect 388102 425258 388186 425494
rect 388422 425258 459866 425494
rect 460102 425258 460186 425494
rect 460422 425258 495866 425494
rect 496102 425258 496186 425494
rect 496422 425258 531866 425494
rect 532102 425258 532186 425494
rect 532422 425258 567866 425494
rect 568102 425258 568186 425494
rect 568422 425258 592062 425494
rect 592298 425258 592382 425494
rect 592618 425258 592650 425494
rect -8726 425174 592650 425258
rect -8726 424938 -8694 425174
rect -8458 424938 -8374 425174
rect -8138 424938 27866 425174
rect 28102 424938 28186 425174
rect 28422 424938 387866 425174
rect 388102 424938 388186 425174
rect 388422 424938 459866 425174
rect 460102 424938 460186 425174
rect 460422 424938 495866 425174
rect 496102 424938 496186 425174
rect 496422 424938 531866 425174
rect 532102 424938 532186 425174
rect 532422 424938 567866 425174
rect 568102 424938 568186 425174
rect 568422 424938 592062 425174
rect 592298 424938 592382 425174
rect 592618 424938 592650 425174
rect -8726 424906 592650 424938
rect -8726 421774 592650 421806
rect -8726 421538 -7734 421774
rect -7498 421538 -7414 421774
rect -7178 421538 384146 421774
rect 384382 421538 384466 421774
rect 384702 421538 420146 421774
rect 420382 421538 420466 421774
rect 420702 421538 456146 421774
rect 456382 421538 456466 421774
rect 456702 421538 492146 421774
rect 492382 421538 492466 421774
rect 492702 421538 528146 421774
rect 528382 421538 528466 421774
rect 528702 421538 564146 421774
rect 564382 421538 564466 421774
rect 564702 421538 591102 421774
rect 591338 421538 591422 421774
rect 591658 421538 592650 421774
rect -8726 421454 592650 421538
rect -8726 421218 -7734 421454
rect -7498 421218 -7414 421454
rect -7178 421218 384146 421454
rect 384382 421218 384466 421454
rect 384702 421218 420146 421454
rect 420382 421218 420466 421454
rect 420702 421218 456146 421454
rect 456382 421218 456466 421454
rect 456702 421218 492146 421454
rect 492382 421218 492466 421454
rect 492702 421218 528146 421454
rect 528382 421218 528466 421454
rect 528702 421218 564146 421454
rect 564382 421218 564466 421454
rect 564702 421218 591102 421454
rect 591338 421218 591422 421454
rect 591658 421218 592650 421454
rect -8726 421186 592650 421218
rect -8726 418054 592650 418086
rect -8726 417818 -6774 418054
rect -6538 417818 -6454 418054
rect -6218 417818 20426 418054
rect 20662 417818 20746 418054
rect 20982 417818 380426 418054
rect 380662 417818 380746 418054
rect 380982 417818 416426 418054
rect 416662 417818 416746 418054
rect 416982 417818 452426 418054
rect 452662 417818 452746 418054
rect 452982 417818 524426 418054
rect 524662 417818 524746 418054
rect 524982 417818 560426 418054
rect 560662 417818 560746 418054
rect 560982 417818 590142 418054
rect 590378 417818 590462 418054
rect 590698 417818 592650 418054
rect -8726 417734 592650 417818
rect -8726 417498 -6774 417734
rect -6538 417498 -6454 417734
rect -6218 417498 20426 417734
rect 20662 417498 20746 417734
rect 20982 417498 380426 417734
rect 380662 417498 380746 417734
rect 380982 417498 416426 417734
rect 416662 417498 416746 417734
rect 416982 417498 452426 417734
rect 452662 417498 452746 417734
rect 452982 417498 524426 417734
rect 524662 417498 524746 417734
rect 524982 417498 560426 417734
rect 560662 417498 560746 417734
rect 560982 417498 590142 417734
rect 590378 417498 590462 417734
rect 590698 417498 592650 417734
rect -8726 417466 592650 417498
rect -8726 414334 592650 414366
rect -8726 414098 -5814 414334
rect -5578 414098 -5494 414334
rect -5258 414098 16706 414334
rect 16942 414098 17026 414334
rect 17262 414098 376706 414334
rect 376942 414098 377026 414334
rect 377262 414098 412706 414334
rect 412942 414098 413026 414334
rect 413262 414098 448706 414334
rect 448942 414098 449026 414334
rect 449262 414098 484706 414334
rect 484942 414098 485026 414334
rect 485262 414098 520706 414334
rect 520942 414098 521026 414334
rect 521262 414098 556706 414334
rect 556942 414098 557026 414334
rect 557262 414098 589182 414334
rect 589418 414098 589502 414334
rect 589738 414098 592650 414334
rect -8726 414014 592650 414098
rect -8726 413778 -5814 414014
rect -5578 413778 -5494 414014
rect -5258 413778 16706 414014
rect 16942 413778 17026 414014
rect 17262 413778 376706 414014
rect 376942 413778 377026 414014
rect 377262 413778 412706 414014
rect 412942 413778 413026 414014
rect 413262 413778 448706 414014
rect 448942 413778 449026 414014
rect 449262 413778 484706 414014
rect 484942 413778 485026 414014
rect 485262 413778 520706 414014
rect 520942 413778 521026 414014
rect 521262 413778 556706 414014
rect 556942 413778 557026 414014
rect 557262 413778 589182 414014
rect 589418 413778 589502 414014
rect 589738 413778 592650 414014
rect -8726 413746 592650 413778
rect -8726 410614 592650 410646
rect -8726 410378 -4854 410614
rect -4618 410378 -4534 410614
rect -4298 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 372986 410614
rect 373222 410378 373306 410614
rect 373542 410378 408986 410614
rect 409222 410378 409306 410614
rect 409542 410378 444986 410614
rect 445222 410378 445306 410614
rect 445542 410378 516986 410614
rect 517222 410378 517306 410614
rect 517542 410378 552986 410614
rect 553222 410378 553306 410614
rect 553542 410378 588222 410614
rect 588458 410378 588542 410614
rect 588778 410378 592650 410614
rect -8726 410294 592650 410378
rect -8726 410058 -4854 410294
rect -4618 410058 -4534 410294
rect -4298 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 372986 410294
rect 373222 410058 373306 410294
rect 373542 410058 408986 410294
rect 409222 410058 409306 410294
rect 409542 410058 444986 410294
rect 445222 410058 445306 410294
rect 445542 410058 516986 410294
rect 517222 410058 517306 410294
rect 517542 410058 552986 410294
rect 553222 410058 553306 410294
rect 553542 410058 588222 410294
rect 588458 410058 588542 410294
rect 588778 410058 592650 410294
rect -8726 410026 592650 410058
rect -8726 406894 592650 406926
rect -8726 406658 -3894 406894
rect -3658 406658 -3574 406894
rect -3338 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 369266 406894
rect 369502 406658 369586 406894
rect 369822 406658 405266 406894
rect 405502 406658 405586 406894
rect 405822 406658 441266 406894
rect 441502 406658 441586 406894
rect 441822 406658 477266 406894
rect 477502 406658 477586 406894
rect 477822 406658 513266 406894
rect 513502 406658 513586 406894
rect 513822 406658 549266 406894
rect 549502 406658 549586 406894
rect 549822 406658 587262 406894
rect 587498 406658 587582 406894
rect 587818 406658 592650 406894
rect -8726 406574 592650 406658
rect -8726 406338 -3894 406574
rect -3658 406338 -3574 406574
rect -3338 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 369266 406574
rect 369502 406338 369586 406574
rect 369822 406338 405266 406574
rect 405502 406338 405586 406574
rect 405822 406338 441266 406574
rect 441502 406338 441586 406574
rect 441822 406338 477266 406574
rect 477502 406338 477586 406574
rect 477822 406338 513266 406574
rect 513502 406338 513586 406574
rect 513822 406338 549266 406574
rect 549502 406338 549586 406574
rect 549822 406338 587262 406574
rect 587498 406338 587582 406574
rect 587818 406338 592650 406574
rect -8726 406306 592650 406338
rect -8726 403174 592650 403206
rect -8726 402938 -2934 403174
rect -2698 402938 -2614 403174
rect -2378 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 39610 403174
rect 39846 402938 70330 403174
rect 70566 402938 101050 403174
rect 101286 402938 131770 403174
rect 132006 402938 162490 403174
rect 162726 402938 193210 403174
rect 193446 402938 223930 403174
rect 224166 402938 254650 403174
rect 254886 402938 285370 403174
rect 285606 402938 316090 403174
rect 316326 402938 346810 403174
rect 347046 402938 365546 403174
rect 365782 402938 365866 403174
rect 366102 402938 401546 403174
rect 401782 402938 401866 403174
rect 402102 402938 437546 403174
rect 437782 402938 437866 403174
rect 438102 402938 509546 403174
rect 509782 402938 509866 403174
rect 510102 402938 545546 403174
rect 545782 402938 545866 403174
rect 546102 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 586302 403174
rect 586538 402938 586622 403174
rect 586858 402938 592650 403174
rect -8726 402854 592650 402938
rect -8726 402618 -2934 402854
rect -2698 402618 -2614 402854
rect -2378 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 39610 402854
rect 39846 402618 70330 402854
rect 70566 402618 101050 402854
rect 101286 402618 131770 402854
rect 132006 402618 162490 402854
rect 162726 402618 193210 402854
rect 193446 402618 223930 402854
rect 224166 402618 254650 402854
rect 254886 402618 285370 402854
rect 285606 402618 316090 402854
rect 316326 402618 346810 402854
rect 347046 402618 365546 402854
rect 365782 402618 365866 402854
rect 366102 402618 401546 402854
rect 401782 402618 401866 402854
rect 402102 402618 437546 402854
rect 437782 402618 437866 402854
rect 438102 402618 509546 402854
rect 509782 402618 509866 402854
rect 510102 402618 545546 402854
rect 545782 402618 545866 402854
rect 546102 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 586302 402854
rect 586538 402618 586622 402854
rect 586858 402618 592650 402854
rect -8726 402586 592650 402618
rect -8726 399454 592650 399486
rect -8726 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 24250 399454
rect 24486 399218 54970 399454
rect 55206 399218 85690 399454
rect 85926 399218 116410 399454
rect 116646 399218 147130 399454
rect 147366 399218 177850 399454
rect 178086 399218 208570 399454
rect 208806 399218 239290 399454
rect 239526 399218 270010 399454
rect 270246 399218 300730 399454
rect 300966 399218 331450 399454
rect 331686 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 592650 399454
rect -8726 399134 592650 399218
rect -8726 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 24250 399134
rect 24486 398898 54970 399134
rect 55206 398898 85690 399134
rect 85926 398898 116410 399134
rect 116646 398898 147130 399134
rect 147366 398898 177850 399134
rect 178086 398898 208570 399134
rect 208806 398898 239290 399134
rect 239526 398898 270010 399134
rect 270246 398898 300730 399134
rect 300966 398898 331450 399134
rect 331686 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 592650 399134
rect -8726 398866 592650 398898
rect -8726 389494 592650 389526
rect -8726 389258 -8694 389494
rect -8458 389258 -8374 389494
rect -8138 389258 27866 389494
rect 28102 389258 28186 389494
rect 28422 389258 387866 389494
rect 388102 389258 388186 389494
rect 388422 389258 423866 389494
rect 424102 389258 424186 389494
rect 424422 389258 459866 389494
rect 460102 389258 460186 389494
rect 460422 389258 495866 389494
rect 496102 389258 496186 389494
rect 496422 389258 531866 389494
rect 532102 389258 532186 389494
rect 532422 389258 567866 389494
rect 568102 389258 568186 389494
rect 568422 389258 592062 389494
rect 592298 389258 592382 389494
rect 592618 389258 592650 389494
rect -8726 389174 592650 389258
rect -8726 388938 -8694 389174
rect -8458 388938 -8374 389174
rect -8138 388938 27866 389174
rect 28102 388938 28186 389174
rect 28422 388938 387866 389174
rect 388102 388938 388186 389174
rect 388422 388938 423866 389174
rect 424102 388938 424186 389174
rect 424422 388938 459866 389174
rect 460102 388938 460186 389174
rect 460422 388938 495866 389174
rect 496102 388938 496186 389174
rect 496422 388938 531866 389174
rect 532102 388938 532186 389174
rect 532422 388938 567866 389174
rect 568102 388938 568186 389174
rect 568422 388938 592062 389174
rect 592298 388938 592382 389174
rect 592618 388938 592650 389174
rect -8726 388906 592650 388938
rect -8726 385774 592650 385806
rect -8726 385538 -7734 385774
rect -7498 385538 -7414 385774
rect -7178 385538 384146 385774
rect 384382 385538 384466 385774
rect 384702 385538 420146 385774
rect 420382 385538 420466 385774
rect 420702 385538 456146 385774
rect 456382 385538 456466 385774
rect 456702 385538 492146 385774
rect 492382 385538 492466 385774
rect 492702 385538 528146 385774
rect 528382 385538 528466 385774
rect 528702 385538 564146 385774
rect 564382 385538 564466 385774
rect 564702 385538 591102 385774
rect 591338 385538 591422 385774
rect 591658 385538 592650 385774
rect -8726 385454 592650 385538
rect -8726 385218 -7734 385454
rect -7498 385218 -7414 385454
rect -7178 385218 384146 385454
rect 384382 385218 384466 385454
rect 384702 385218 420146 385454
rect 420382 385218 420466 385454
rect 420702 385218 456146 385454
rect 456382 385218 456466 385454
rect 456702 385218 492146 385454
rect 492382 385218 492466 385454
rect 492702 385218 528146 385454
rect 528382 385218 528466 385454
rect 528702 385218 564146 385454
rect 564382 385218 564466 385454
rect 564702 385218 591102 385454
rect 591338 385218 591422 385454
rect 591658 385218 592650 385454
rect -8726 385186 592650 385218
rect -8726 382054 592650 382086
rect -8726 381818 -6774 382054
rect -6538 381818 -6454 382054
rect -6218 381818 20426 382054
rect 20662 381818 20746 382054
rect 20982 381818 380426 382054
rect 380662 381818 380746 382054
rect 380982 381818 416426 382054
rect 416662 381818 416746 382054
rect 416982 381818 452426 382054
rect 452662 381818 452746 382054
rect 452982 381818 524426 382054
rect 524662 381818 524746 382054
rect 524982 381818 560426 382054
rect 560662 381818 560746 382054
rect 560982 381818 590142 382054
rect 590378 381818 590462 382054
rect 590698 381818 592650 382054
rect -8726 381734 592650 381818
rect -8726 381498 -6774 381734
rect -6538 381498 -6454 381734
rect -6218 381498 20426 381734
rect 20662 381498 20746 381734
rect 20982 381498 380426 381734
rect 380662 381498 380746 381734
rect 380982 381498 416426 381734
rect 416662 381498 416746 381734
rect 416982 381498 452426 381734
rect 452662 381498 452746 381734
rect 452982 381498 524426 381734
rect 524662 381498 524746 381734
rect 524982 381498 560426 381734
rect 560662 381498 560746 381734
rect 560982 381498 590142 381734
rect 590378 381498 590462 381734
rect 590698 381498 592650 381734
rect -8726 381466 592650 381498
rect -8726 378334 592650 378366
rect -8726 378098 -5814 378334
rect -5578 378098 -5494 378334
rect -5258 378098 16706 378334
rect 16942 378098 17026 378334
rect 17262 378098 376706 378334
rect 376942 378098 377026 378334
rect 377262 378098 412706 378334
rect 412942 378098 413026 378334
rect 413262 378098 448706 378334
rect 448942 378098 449026 378334
rect 449262 378098 520706 378334
rect 520942 378098 521026 378334
rect 521262 378243 589182 378334
rect 521262 378098 556706 378243
rect -8726 378014 556706 378098
rect -8726 377778 -5814 378014
rect -5578 377778 -5494 378014
rect -5258 377778 16706 378014
rect 16942 377778 17026 378014
rect 17262 377778 376706 378014
rect 376942 377778 377026 378014
rect 377262 377778 412706 378014
rect 412942 377778 413026 378014
rect 413262 377778 448706 378014
rect 448942 377778 449026 378014
rect 449262 377778 520706 378014
rect 520942 377778 521026 378014
rect 521262 378007 556706 378014
rect 556942 378007 557026 378243
rect 557262 378098 589182 378243
rect 589418 378098 589502 378334
rect 589738 378098 592650 378334
rect 557262 378014 592650 378098
rect 557262 378007 589182 378014
rect 521262 377778 589182 378007
rect 589418 377778 589502 378014
rect 589738 377778 592650 378014
rect -8726 377746 592650 377778
rect -8726 374614 592650 374646
rect -8726 374378 -4854 374614
rect -4618 374378 -4534 374614
rect -4298 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 372986 374614
rect 373222 374378 373306 374614
rect 373542 374378 408986 374614
rect 409222 374378 409306 374614
rect 409542 374378 444986 374614
rect 445222 374378 445306 374614
rect 445542 374378 516986 374614
rect 517222 374378 517306 374614
rect 517542 374378 588222 374614
rect 588458 374378 588542 374614
rect 588778 374378 592650 374614
rect -8726 374294 592650 374378
rect -8726 374058 -4854 374294
rect -4618 374058 -4534 374294
rect -4298 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 372986 374294
rect 373222 374058 373306 374294
rect 373542 374058 408986 374294
rect 409222 374058 409306 374294
rect 409542 374058 444986 374294
rect 445222 374058 445306 374294
rect 445542 374058 516986 374294
rect 517222 374058 517306 374294
rect 517542 374058 588222 374294
rect 588458 374058 588542 374294
rect 588778 374058 592650 374294
rect -8726 374026 592650 374058
rect -8726 370894 592650 370926
rect -8726 370658 -3894 370894
rect -3658 370658 -3574 370894
rect -3338 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 369266 370894
rect 369502 370658 369586 370894
rect 369822 370658 405266 370894
rect 405502 370658 405586 370894
rect 405822 370658 441266 370894
rect 441502 370658 441586 370894
rect 441822 370658 513266 370894
rect 513502 370658 513586 370894
rect 513822 370658 549266 370894
rect 549502 370658 549586 370894
rect 549822 370658 587262 370894
rect 587498 370658 587582 370894
rect 587818 370658 592650 370894
rect -8726 370574 592650 370658
rect -8726 370338 -3894 370574
rect -3658 370338 -3574 370574
rect -3338 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 369266 370574
rect 369502 370338 369586 370574
rect 369822 370338 405266 370574
rect 405502 370338 405586 370574
rect 405822 370338 441266 370574
rect 441502 370338 441586 370574
rect 441822 370338 513266 370574
rect 513502 370338 513586 370574
rect 513822 370338 549266 370574
rect 549502 370338 549586 370574
rect 549822 370338 587262 370574
rect 587498 370338 587582 370574
rect 587818 370338 592650 370574
rect -8726 370306 592650 370338
rect -8726 367174 592650 367206
rect -8726 366938 -2934 367174
rect -2698 366938 -2614 367174
rect -2378 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 39610 367174
rect 39846 366938 70330 367174
rect 70566 366938 101050 367174
rect 101286 366938 131770 367174
rect 132006 366938 162490 367174
rect 162726 366938 193210 367174
rect 193446 366938 223930 367174
rect 224166 366938 254650 367174
rect 254886 366938 285370 367174
rect 285606 366938 316090 367174
rect 316326 366938 346810 367174
rect 347046 366938 365546 367174
rect 365782 366938 365866 367174
rect 366102 366938 401546 367174
rect 401782 366938 401866 367174
rect 402102 366938 437546 367174
rect 437782 366938 437866 367174
rect 438102 366938 469610 367174
rect 469846 366938 500330 367174
rect 500566 366938 509546 367174
rect 509782 366938 509866 367174
rect 510102 366938 545546 367174
rect 545782 366938 545866 367174
rect 546102 366938 554918 367174
rect 555154 366938 558851 367174
rect 559087 366938 562784 367174
rect 563020 366938 566717 367174
rect 566953 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 586302 367174
rect 586538 366938 586622 367174
rect 586858 366938 592650 367174
rect -8726 366854 592650 366938
rect -8726 366618 -2934 366854
rect -2698 366618 -2614 366854
rect -2378 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 39610 366854
rect 39846 366618 70330 366854
rect 70566 366618 101050 366854
rect 101286 366618 131770 366854
rect 132006 366618 162490 366854
rect 162726 366618 193210 366854
rect 193446 366618 223930 366854
rect 224166 366618 254650 366854
rect 254886 366618 285370 366854
rect 285606 366618 316090 366854
rect 316326 366618 346810 366854
rect 347046 366618 365546 366854
rect 365782 366618 365866 366854
rect 366102 366618 401546 366854
rect 401782 366618 401866 366854
rect 402102 366618 437546 366854
rect 437782 366618 437866 366854
rect 438102 366618 469610 366854
rect 469846 366618 500330 366854
rect 500566 366618 509546 366854
rect 509782 366618 509866 366854
rect 510102 366618 545546 366854
rect 545782 366618 545866 366854
rect 546102 366618 554918 366854
rect 555154 366618 558851 366854
rect 559087 366618 562784 366854
rect 563020 366618 566717 366854
rect 566953 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 586302 366854
rect 586538 366618 586622 366854
rect 586858 366618 592650 366854
rect -8726 366586 592650 366618
rect -8726 363454 592650 363486
rect -8726 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 24250 363454
rect 24486 363218 54970 363454
rect 55206 363218 85690 363454
rect 85926 363218 116410 363454
rect 116646 363218 147130 363454
rect 147366 363218 177850 363454
rect 178086 363218 208570 363454
rect 208806 363218 239290 363454
rect 239526 363218 270010 363454
rect 270246 363218 300730 363454
rect 300966 363218 331450 363454
rect 331686 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 454250 363454
rect 454486 363218 484970 363454
rect 485206 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 552952 363454
rect 553188 363218 556885 363454
rect 557121 363218 560818 363454
rect 561054 363218 564751 363454
rect 564987 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 592650 363454
rect -8726 363134 592650 363218
rect -8726 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 24250 363134
rect 24486 362898 54970 363134
rect 55206 362898 85690 363134
rect 85926 362898 116410 363134
rect 116646 362898 147130 363134
rect 147366 362898 177850 363134
rect 178086 362898 208570 363134
rect 208806 362898 239290 363134
rect 239526 362898 270010 363134
rect 270246 362898 300730 363134
rect 300966 362898 331450 363134
rect 331686 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 454250 363134
rect 454486 362898 484970 363134
rect 485206 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 552952 363134
rect 553188 362898 556885 363134
rect 557121 362898 560818 363134
rect 561054 362898 564751 363134
rect 564987 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 592650 363134
rect -8726 362866 592650 362898
rect -8726 353494 592650 353526
rect -8726 353258 -8694 353494
rect -8458 353258 -8374 353494
rect -8138 353258 27866 353494
rect 28102 353258 28186 353494
rect 28422 353258 387866 353494
rect 388102 353258 388186 353494
rect 388422 353258 423866 353494
rect 424102 353258 424186 353494
rect 424422 353258 459866 353494
rect 460102 353258 460186 353494
rect 460422 353258 531866 353494
rect 532102 353258 532186 353494
rect 532422 353258 567866 353494
rect 568102 353258 568186 353494
rect 568422 353258 592062 353494
rect 592298 353258 592382 353494
rect 592618 353258 592650 353494
rect -8726 353174 592650 353258
rect -8726 352938 -8694 353174
rect -8458 352938 -8374 353174
rect -8138 352938 27866 353174
rect 28102 352938 28186 353174
rect 28422 352938 387866 353174
rect 388102 352938 388186 353174
rect 388422 352938 423866 353174
rect 424102 352938 424186 353174
rect 424422 352938 459866 353174
rect 460102 352938 460186 353174
rect 460422 352938 531866 353174
rect 532102 352938 532186 353174
rect 532422 352938 567866 353174
rect 568102 352938 568186 353174
rect 568422 352938 592062 353174
rect 592298 352938 592382 353174
rect 592618 352938 592650 353174
rect -8726 352906 592650 352938
rect -8726 349774 592650 349806
rect -8726 349538 -7734 349774
rect -7498 349538 -7414 349774
rect -7178 349538 384146 349774
rect 384382 349538 384466 349774
rect 384702 349538 420146 349774
rect 420382 349538 420466 349774
rect 420702 349538 456146 349774
rect 456382 349538 456466 349774
rect 456702 349538 528146 349774
rect 528382 349538 528466 349774
rect 528702 349538 564146 349774
rect 564382 349538 564466 349774
rect 564702 349538 591102 349774
rect 591338 349538 591422 349774
rect 591658 349538 592650 349774
rect -8726 349454 592650 349538
rect -8726 349218 -7734 349454
rect -7498 349218 -7414 349454
rect -7178 349218 384146 349454
rect 384382 349218 384466 349454
rect 384702 349218 420146 349454
rect 420382 349218 420466 349454
rect 420702 349218 456146 349454
rect 456382 349218 456466 349454
rect 456702 349218 528146 349454
rect 528382 349218 528466 349454
rect 528702 349218 564146 349454
rect 564382 349218 564466 349454
rect 564702 349218 591102 349454
rect 591338 349218 591422 349454
rect 591658 349218 592650 349454
rect -8726 349186 592650 349218
rect -8726 346054 592650 346086
rect -8726 345818 -6774 346054
rect -6538 345818 -6454 346054
rect -6218 345818 20426 346054
rect 20662 345818 20746 346054
rect 20982 345818 380426 346054
rect 380662 345818 380746 346054
rect 380982 345818 416426 346054
rect 416662 345818 416746 346054
rect 416982 345818 452426 346054
rect 452662 345818 452746 346054
rect 452982 345818 524426 346054
rect 524662 345818 524746 346054
rect 524982 345818 560426 346054
rect 560662 345818 560746 346054
rect 560982 345818 590142 346054
rect 590378 345818 590462 346054
rect 590698 345818 592650 346054
rect -8726 345734 592650 345818
rect -8726 345498 -6774 345734
rect -6538 345498 -6454 345734
rect -6218 345498 20426 345734
rect 20662 345498 20746 345734
rect 20982 345498 380426 345734
rect 380662 345498 380746 345734
rect 380982 345498 416426 345734
rect 416662 345498 416746 345734
rect 416982 345498 452426 345734
rect 452662 345498 452746 345734
rect 452982 345498 524426 345734
rect 524662 345498 524746 345734
rect 524982 345498 560426 345734
rect 560662 345498 560746 345734
rect 560982 345498 590142 345734
rect 590378 345498 590462 345734
rect 590698 345498 592650 345734
rect -8726 345466 592650 345498
rect -8726 342334 592650 342366
rect -8726 342098 -5814 342334
rect -5578 342098 -5494 342334
rect -5258 342098 16706 342334
rect 16942 342098 17026 342334
rect 17262 342098 376706 342334
rect 376942 342098 377026 342334
rect 377262 342098 412706 342334
rect 412942 342098 413026 342334
rect 413262 342098 448706 342334
rect 448942 342098 449026 342334
rect 449262 342098 520706 342334
rect 520942 342098 521026 342334
rect 521262 342098 556706 342334
rect 556942 342098 557026 342334
rect 557262 342098 589182 342334
rect 589418 342098 589502 342334
rect 589738 342098 592650 342334
rect -8726 342014 592650 342098
rect -8726 341778 -5814 342014
rect -5578 341778 -5494 342014
rect -5258 341778 16706 342014
rect 16942 341778 17026 342014
rect 17262 341778 376706 342014
rect 376942 341778 377026 342014
rect 377262 341778 412706 342014
rect 412942 341778 413026 342014
rect 413262 341778 448706 342014
rect 448942 341778 449026 342014
rect 449262 341778 520706 342014
rect 520942 341778 521026 342014
rect 521262 341778 556706 342014
rect 556942 341778 557026 342014
rect 557262 341778 589182 342014
rect 589418 341778 589502 342014
rect 589738 341778 592650 342014
rect -8726 341746 592650 341778
rect -8726 338614 592650 338646
rect -8726 338378 -4854 338614
rect -4618 338378 -4534 338614
rect -4298 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 372986 338614
rect 373222 338378 373306 338614
rect 373542 338378 408986 338614
rect 409222 338378 409306 338614
rect 409542 338378 444986 338614
rect 445222 338378 445306 338614
rect 445542 338378 516986 338614
rect 517222 338378 517306 338614
rect 517542 338378 552986 338614
rect 553222 338378 553306 338614
rect 553542 338378 588222 338614
rect 588458 338378 588542 338614
rect 588778 338378 592650 338614
rect -8726 338294 592650 338378
rect -8726 338058 -4854 338294
rect -4618 338058 -4534 338294
rect -4298 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 372986 338294
rect 373222 338058 373306 338294
rect 373542 338058 408986 338294
rect 409222 338058 409306 338294
rect 409542 338058 444986 338294
rect 445222 338058 445306 338294
rect 445542 338058 516986 338294
rect 517222 338058 517306 338294
rect 517542 338058 552986 338294
rect 553222 338058 553306 338294
rect 553542 338058 588222 338294
rect 588458 338058 588542 338294
rect 588778 338058 592650 338294
rect -8726 338026 592650 338058
rect -8726 334894 592650 334926
rect -8726 334658 -3894 334894
rect -3658 334658 -3574 334894
rect -3338 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 369266 334894
rect 369502 334658 369586 334894
rect 369822 334658 405266 334894
rect 405502 334658 405586 334894
rect 405822 334658 441266 334894
rect 441502 334658 441586 334894
rect 441822 334658 513266 334894
rect 513502 334658 513586 334894
rect 513822 334658 549266 334894
rect 549502 334658 549586 334894
rect 549822 334658 587262 334894
rect 587498 334658 587582 334894
rect 587818 334658 592650 334894
rect -8726 334574 592650 334658
rect -8726 334338 -3894 334574
rect -3658 334338 -3574 334574
rect -3338 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 369266 334574
rect 369502 334338 369586 334574
rect 369822 334338 405266 334574
rect 405502 334338 405586 334574
rect 405822 334338 441266 334574
rect 441502 334338 441586 334574
rect 441822 334338 513266 334574
rect 513502 334338 513586 334574
rect 513822 334338 549266 334574
rect 549502 334338 549586 334574
rect 549822 334338 587262 334574
rect 587498 334338 587582 334574
rect 587818 334338 592650 334574
rect -8726 334306 592650 334338
rect -8726 331174 592650 331206
rect -8726 330938 -2934 331174
rect -2698 330938 -2614 331174
rect -2378 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 39610 331174
rect 39846 330938 70330 331174
rect 70566 330938 101050 331174
rect 101286 330938 131770 331174
rect 132006 330938 162490 331174
rect 162726 330938 193210 331174
rect 193446 330938 223930 331174
rect 224166 330938 254650 331174
rect 254886 330938 285370 331174
rect 285606 330938 316090 331174
rect 316326 330938 346810 331174
rect 347046 330938 365546 331174
rect 365782 330938 365866 331174
rect 366102 330938 401546 331174
rect 401782 330938 401866 331174
rect 402102 330938 407932 331174
rect 408168 330938 414878 331174
rect 415114 330938 421824 331174
rect 422060 330938 428770 331174
rect 429006 330938 437546 331174
rect 437782 330938 437866 331174
rect 438102 330938 469610 331174
rect 469846 330938 500330 331174
rect 500566 330938 509546 331174
rect 509782 330938 509866 331174
rect 510102 330938 545546 331174
rect 545782 330938 545866 331174
rect 546102 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 586302 331174
rect 586538 330938 586622 331174
rect 586858 330938 592650 331174
rect -8726 330854 592650 330938
rect -8726 330618 -2934 330854
rect -2698 330618 -2614 330854
rect -2378 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 39610 330854
rect 39846 330618 70330 330854
rect 70566 330618 101050 330854
rect 101286 330618 131770 330854
rect 132006 330618 162490 330854
rect 162726 330618 193210 330854
rect 193446 330618 223930 330854
rect 224166 330618 254650 330854
rect 254886 330618 285370 330854
rect 285606 330618 316090 330854
rect 316326 330618 346810 330854
rect 347046 330618 365546 330854
rect 365782 330618 365866 330854
rect 366102 330618 401546 330854
rect 401782 330618 401866 330854
rect 402102 330618 407932 330854
rect 408168 330618 414878 330854
rect 415114 330618 421824 330854
rect 422060 330618 428770 330854
rect 429006 330618 437546 330854
rect 437782 330618 437866 330854
rect 438102 330618 469610 330854
rect 469846 330618 500330 330854
rect 500566 330618 509546 330854
rect 509782 330618 509866 330854
rect 510102 330618 545546 330854
rect 545782 330618 545866 330854
rect 546102 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 586302 330854
rect 586538 330618 586622 330854
rect 586858 330618 592650 330854
rect -8726 330586 592650 330618
rect -8726 327454 592650 327486
rect -8726 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 24250 327454
rect 24486 327218 54970 327454
rect 55206 327218 85690 327454
rect 85926 327218 116410 327454
rect 116646 327218 147130 327454
rect 147366 327218 177850 327454
rect 178086 327218 208570 327454
rect 208806 327218 239290 327454
rect 239526 327218 270010 327454
rect 270246 327218 300730 327454
rect 300966 327218 331450 327454
rect 331686 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 404459 327454
rect 404695 327218 411405 327454
rect 411641 327218 418351 327454
rect 418587 327218 425297 327454
rect 425533 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 454250 327454
rect 454486 327218 484970 327454
rect 485206 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 592650 327454
rect -8726 327134 592650 327218
rect -8726 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 24250 327134
rect 24486 326898 54970 327134
rect 55206 326898 85690 327134
rect 85926 326898 116410 327134
rect 116646 326898 147130 327134
rect 147366 326898 177850 327134
rect 178086 326898 208570 327134
rect 208806 326898 239290 327134
rect 239526 326898 270010 327134
rect 270246 326898 300730 327134
rect 300966 326898 331450 327134
rect 331686 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 404459 327134
rect 404695 326898 411405 327134
rect 411641 326898 418351 327134
rect 418587 326898 425297 327134
rect 425533 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 454250 327134
rect 454486 326898 484970 327134
rect 485206 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 592650 327134
rect -8726 326866 592650 326898
rect -8726 317494 592650 317526
rect -8726 317258 -8694 317494
rect -8458 317258 -8374 317494
rect -8138 317258 27866 317494
rect 28102 317258 28186 317494
rect 28422 317258 387866 317494
rect 388102 317258 388186 317494
rect 388422 317258 423866 317494
rect 424102 317258 424186 317494
rect 424422 317258 459866 317494
rect 460102 317258 460186 317494
rect 460422 317258 495866 317494
rect 496102 317258 496186 317494
rect 496422 317258 531866 317494
rect 532102 317258 532186 317494
rect 532422 317258 567866 317494
rect 568102 317258 568186 317494
rect 568422 317258 592062 317494
rect 592298 317258 592382 317494
rect 592618 317258 592650 317494
rect -8726 317174 592650 317258
rect -8726 316938 -8694 317174
rect -8458 316938 -8374 317174
rect -8138 316938 27866 317174
rect 28102 316938 28186 317174
rect 28422 316938 387866 317174
rect 388102 316938 388186 317174
rect 388422 316938 423866 317174
rect 424102 316938 424186 317174
rect 424422 316938 459866 317174
rect 460102 316938 460186 317174
rect 460422 316938 495866 317174
rect 496102 316938 496186 317174
rect 496422 316938 531866 317174
rect 532102 316938 532186 317174
rect 532422 316938 567866 317174
rect 568102 316938 568186 317174
rect 568422 316938 592062 317174
rect 592298 316938 592382 317174
rect 592618 316938 592650 317174
rect -8726 316906 592650 316938
rect -8726 313774 592650 313806
rect -8726 313538 -7734 313774
rect -7498 313538 -7414 313774
rect -7178 313538 384146 313774
rect 384382 313538 384466 313774
rect 384702 313538 420146 313774
rect 420382 313538 420466 313774
rect 420702 313538 456146 313774
rect 456382 313538 456466 313774
rect 456702 313538 492146 313774
rect 492382 313538 492466 313774
rect 492702 313538 528146 313774
rect 528382 313538 528466 313774
rect 528702 313538 564146 313774
rect 564382 313538 564466 313774
rect 564702 313538 591102 313774
rect 591338 313538 591422 313774
rect 591658 313538 592650 313774
rect -8726 313454 592650 313538
rect -8726 313218 -7734 313454
rect -7498 313218 -7414 313454
rect -7178 313218 384146 313454
rect 384382 313218 384466 313454
rect 384702 313218 420146 313454
rect 420382 313218 420466 313454
rect 420702 313218 456146 313454
rect 456382 313218 456466 313454
rect 456702 313218 492146 313454
rect 492382 313218 492466 313454
rect 492702 313218 528146 313454
rect 528382 313218 528466 313454
rect 528702 313218 564146 313454
rect 564382 313218 564466 313454
rect 564702 313218 591102 313454
rect 591338 313218 591422 313454
rect 591658 313218 592650 313454
rect -8726 313186 592650 313218
rect -8726 310054 592650 310086
rect -8726 309818 -6774 310054
rect -6538 309818 -6454 310054
rect -6218 309818 20426 310054
rect 20662 309818 20746 310054
rect 20982 309818 380426 310054
rect 380662 309818 380746 310054
rect 380982 309818 416426 310054
rect 416662 309818 416746 310054
rect 416982 309818 452426 310054
rect 452662 309818 452746 310054
rect 452982 309818 488426 310054
rect 488662 309818 488746 310054
rect 488982 309818 524426 310054
rect 524662 309818 524746 310054
rect 524982 309818 560426 310054
rect 560662 309818 560746 310054
rect 560982 309818 590142 310054
rect 590378 309818 590462 310054
rect 590698 309818 592650 310054
rect -8726 309734 592650 309818
rect -8726 309498 -6774 309734
rect -6538 309498 -6454 309734
rect -6218 309498 20426 309734
rect 20662 309498 20746 309734
rect 20982 309498 380426 309734
rect 380662 309498 380746 309734
rect 380982 309498 416426 309734
rect 416662 309498 416746 309734
rect 416982 309498 452426 309734
rect 452662 309498 452746 309734
rect 452982 309498 488426 309734
rect 488662 309498 488746 309734
rect 488982 309498 524426 309734
rect 524662 309498 524746 309734
rect 524982 309498 560426 309734
rect 560662 309498 560746 309734
rect 560982 309498 590142 309734
rect 590378 309498 590462 309734
rect 590698 309498 592650 309734
rect -8726 309466 592650 309498
rect -8726 306334 592650 306366
rect -8726 306098 -5814 306334
rect -5578 306098 -5494 306334
rect -5258 306098 16706 306334
rect 16942 306098 17026 306334
rect 17262 306098 376706 306334
rect 376942 306098 377026 306334
rect 377262 306098 412706 306334
rect 412942 306098 413026 306334
rect 413262 306098 448706 306334
rect 448942 306098 449026 306334
rect 449262 306098 484706 306334
rect 484942 306098 485026 306334
rect 485262 306098 520706 306334
rect 520942 306098 521026 306334
rect 521262 306098 556706 306334
rect 556942 306098 557026 306334
rect 557262 306098 589182 306334
rect 589418 306098 589502 306334
rect 589738 306098 592650 306334
rect -8726 306014 592650 306098
rect -8726 305778 -5814 306014
rect -5578 305778 -5494 306014
rect -5258 305778 16706 306014
rect 16942 305778 17026 306014
rect 17262 305778 376706 306014
rect 376942 305778 377026 306014
rect 377262 305778 412706 306014
rect 412942 305778 413026 306014
rect 413262 305778 448706 306014
rect 448942 305778 449026 306014
rect 449262 305778 484706 306014
rect 484942 305778 485026 306014
rect 485262 305778 520706 306014
rect 520942 305778 521026 306014
rect 521262 305778 556706 306014
rect 556942 305778 557026 306014
rect 557262 305778 589182 306014
rect 589418 305778 589502 306014
rect 589738 305778 592650 306014
rect -8726 305746 592650 305778
rect -8726 302614 592650 302646
rect -8726 302378 -4854 302614
rect -4618 302378 -4534 302614
rect -4298 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 372986 302614
rect 373222 302378 373306 302614
rect 373542 302378 408986 302614
rect 409222 302378 409306 302614
rect 409542 302378 444986 302614
rect 445222 302378 445306 302614
rect 445542 302378 480986 302614
rect 481222 302378 481306 302614
rect 481542 302378 516986 302614
rect 517222 302378 517306 302614
rect 517542 302378 552986 302614
rect 553222 302378 553306 302614
rect 553542 302378 588222 302614
rect 588458 302378 588542 302614
rect 588778 302378 592650 302614
rect -8726 302294 592650 302378
rect -8726 302058 -4854 302294
rect -4618 302058 -4534 302294
rect -4298 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 372986 302294
rect 373222 302058 373306 302294
rect 373542 302058 408986 302294
rect 409222 302058 409306 302294
rect 409542 302058 444986 302294
rect 445222 302058 445306 302294
rect 445542 302058 480986 302294
rect 481222 302058 481306 302294
rect 481542 302058 516986 302294
rect 517222 302058 517306 302294
rect 517542 302058 552986 302294
rect 553222 302058 553306 302294
rect 553542 302058 588222 302294
rect 588458 302058 588542 302294
rect 588778 302058 592650 302294
rect -8726 302026 592650 302058
rect -8726 298894 592650 298926
rect -8726 298658 -3894 298894
rect -3658 298658 -3574 298894
rect -3338 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 369266 298894
rect 369502 298658 369586 298894
rect 369822 298658 405266 298894
rect 405502 298658 405586 298894
rect 405822 298658 441266 298894
rect 441502 298658 441586 298894
rect 441822 298658 477266 298894
rect 477502 298658 477586 298894
rect 477822 298658 513266 298894
rect 513502 298658 513586 298894
rect 513822 298658 549266 298894
rect 549502 298658 549586 298894
rect 549822 298658 587262 298894
rect 587498 298658 587582 298894
rect 587818 298658 592650 298894
rect -8726 298574 592650 298658
rect -8726 298338 -3894 298574
rect -3658 298338 -3574 298574
rect -3338 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 369266 298574
rect 369502 298338 369586 298574
rect 369822 298338 405266 298574
rect 405502 298338 405586 298574
rect 405822 298338 441266 298574
rect 441502 298338 441586 298574
rect 441822 298338 477266 298574
rect 477502 298338 477586 298574
rect 477822 298338 513266 298574
rect 513502 298338 513586 298574
rect 513822 298338 549266 298574
rect 549502 298338 549586 298574
rect 549822 298338 587262 298574
rect 587498 298338 587582 298574
rect 587818 298338 592650 298574
rect -8726 298306 592650 298338
rect -8726 295174 592650 295206
rect -8726 294938 -2934 295174
rect -2698 294938 -2614 295174
rect -2378 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 39610 295174
rect 39846 294938 70330 295174
rect 70566 294938 101050 295174
rect 101286 294938 131770 295174
rect 132006 294938 162490 295174
rect 162726 294938 193210 295174
rect 193446 294938 223930 295174
rect 224166 294938 254650 295174
rect 254886 294938 285370 295174
rect 285606 294938 316090 295174
rect 316326 294938 346810 295174
rect 347046 294938 365546 295174
rect 365782 294938 365866 295174
rect 366102 294938 401546 295174
rect 401782 294938 401866 295174
rect 402102 294938 437546 295174
rect 437782 294938 437866 295174
rect 438102 294938 509546 295174
rect 509782 294938 509866 295174
rect 510102 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 586302 295174
rect 586538 294938 586622 295174
rect 586858 294938 592650 295174
rect -8726 294854 592650 294938
rect -8726 294618 -2934 294854
rect -2698 294618 -2614 294854
rect -2378 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 39610 294854
rect 39846 294618 70330 294854
rect 70566 294618 101050 294854
rect 101286 294618 131770 294854
rect 132006 294618 162490 294854
rect 162726 294618 193210 294854
rect 193446 294618 223930 294854
rect 224166 294618 254650 294854
rect 254886 294618 285370 294854
rect 285606 294618 316090 294854
rect 316326 294618 346810 294854
rect 347046 294618 365546 294854
rect 365782 294618 365866 294854
rect 366102 294618 401546 294854
rect 401782 294618 401866 294854
rect 402102 294618 437546 294854
rect 437782 294618 437866 294854
rect 438102 294618 509546 294854
rect 509782 294618 509866 294854
rect 510102 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 586302 294854
rect 586538 294618 586622 294854
rect 586858 294618 592650 294854
rect -8726 294586 592650 294618
rect -8726 291454 592650 291486
rect -8726 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 24250 291454
rect 24486 291218 54970 291454
rect 55206 291218 85690 291454
rect 85926 291218 116410 291454
rect 116646 291218 147130 291454
rect 147366 291218 177850 291454
rect 178086 291218 208570 291454
rect 208806 291218 239290 291454
rect 239526 291218 270010 291454
rect 270246 291218 300730 291454
rect 300966 291218 331450 291454
rect 331686 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 592650 291454
rect -8726 291134 592650 291218
rect -8726 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 24250 291134
rect 24486 290898 54970 291134
rect 55206 290898 85690 291134
rect 85926 290898 116410 291134
rect 116646 290898 147130 291134
rect 147366 290898 177850 291134
rect 178086 290898 208570 291134
rect 208806 290898 239290 291134
rect 239526 290898 270010 291134
rect 270246 290898 300730 291134
rect 300966 290898 331450 291134
rect 331686 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 592650 291134
rect -8726 290866 592650 290898
rect -8726 281494 592650 281526
rect -8726 281258 -8694 281494
rect -8458 281258 -8374 281494
rect -8138 281258 27866 281494
rect 28102 281258 28186 281494
rect 28422 281258 387866 281494
rect 388102 281258 388186 281494
rect 388422 281258 423866 281494
rect 424102 281258 424186 281494
rect 424422 281258 459866 281494
rect 460102 281258 460186 281494
rect 460422 281258 495866 281494
rect 496102 281258 496186 281494
rect 496422 281258 531866 281494
rect 532102 281258 532186 281494
rect 532422 281258 567866 281494
rect 568102 281258 568186 281494
rect 568422 281258 592062 281494
rect 592298 281258 592382 281494
rect 592618 281258 592650 281494
rect -8726 281174 592650 281258
rect -8726 280938 -8694 281174
rect -8458 280938 -8374 281174
rect -8138 280938 27866 281174
rect 28102 280938 28186 281174
rect 28422 280938 387866 281174
rect 388102 280938 388186 281174
rect 388422 280938 423866 281174
rect 424102 280938 424186 281174
rect 424422 280938 459866 281174
rect 460102 280938 460186 281174
rect 460422 280938 495866 281174
rect 496102 280938 496186 281174
rect 496422 280938 531866 281174
rect 532102 280938 532186 281174
rect 532422 280938 567866 281174
rect 568102 280938 568186 281174
rect 568422 280938 592062 281174
rect 592298 280938 592382 281174
rect 592618 280938 592650 281174
rect -8726 280906 592650 280938
rect -8726 277774 592650 277806
rect -8726 277538 -7734 277774
rect -7498 277538 -7414 277774
rect -7178 277538 384146 277774
rect 384382 277538 384466 277774
rect 384702 277538 420146 277774
rect 420382 277538 420466 277774
rect 420702 277538 456146 277774
rect 456382 277538 456466 277774
rect 456702 277538 492146 277774
rect 492382 277538 492466 277774
rect 492702 277538 528146 277774
rect 528382 277538 528466 277774
rect 528702 277538 564146 277774
rect 564382 277538 564466 277774
rect 564702 277538 591102 277774
rect 591338 277538 591422 277774
rect 591658 277538 592650 277774
rect -8726 277454 592650 277538
rect -8726 277218 -7734 277454
rect -7498 277218 -7414 277454
rect -7178 277218 384146 277454
rect 384382 277218 384466 277454
rect 384702 277218 420146 277454
rect 420382 277218 420466 277454
rect 420702 277218 456146 277454
rect 456382 277218 456466 277454
rect 456702 277218 492146 277454
rect 492382 277218 492466 277454
rect 492702 277218 528146 277454
rect 528382 277218 528466 277454
rect 528702 277218 564146 277454
rect 564382 277218 564466 277454
rect 564702 277218 591102 277454
rect 591338 277218 591422 277454
rect 591658 277218 592650 277454
rect -8726 277186 592650 277218
rect -8726 274054 592650 274086
rect -8726 273818 -6774 274054
rect -6538 273818 -6454 274054
rect -6218 273818 20426 274054
rect 20662 273818 20746 274054
rect 20982 273818 380426 274054
rect 380662 273818 380746 274054
rect 380982 273818 416426 274054
rect 416662 273818 416746 274054
rect 416982 273818 452426 274054
rect 452662 273818 452746 274054
rect 452982 273818 488426 274054
rect 488662 273818 488746 274054
rect 488982 273818 524426 274054
rect 524662 273818 524746 274054
rect 524982 273818 560426 274054
rect 560662 273818 560746 274054
rect 560982 273818 590142 274054
rect 590378 273818 590462 274054
rect 590698 273818 592650 274054
rect -8726 273734 592650 273818
rect -8726 273498 -6774 273734
rect -6538 273498 -6454 273734
rect -6218 273498 20426 273734
rect 20662 273498 20746 273734
rect 20982 273498 380426 273734
rect 380662 273498 380746 273734
rect 380982 273498 416426 273734
rect 416662 273498 416746 273734
rect 416982 273498 452426 273734
rect 452662 273498 452746 273734
rect 452982 273498 488426 273734
rect 488662 273498 488746 273734
rect 488982 273498 524426 273734
rect 524662 273498 524746 273734
rect 524982 273498 560426 273734
rect 560662 273498 560746 273734
rect 560982 273498 590142 273734
rect 590378 273498 590462 273734
rect 590698 273498 592650 273734
rect -8726 273466 592650 273498
rect -8726 270334 592650 270366
rect -8726 270098 -5814 270334
rect -5578 270098 -5494 270334
rect -5258 270098 16706 270334
rect 16942 270098 17026 270334
rect 17262 270098 376706 270334
rect 376942 270098 377026 270334
rect 377262 270098 412706 270334
rect 412942 270098 413026 270334
rect 413262 270098 448706 270334
rect 448942 270098 449026 270334
rect 449262 270098 484706 270334
rect 484942 270098 485026 270334
rect 485262 270098 520706 270334
rect 520942 270098 521026 270334
rect 521262 270098 556706 270334
rect 556942 270098 557026 270334
rect 557262 270098 589182 270334
rect 589418 270098 589502 270334
rect 589738 270098 592650 270334
rect -8726 270014 592650 270098
rect -8726 269778 -5814 270014
rect -5578 269778 -5494 270014
rect -5258 269778 16706 270014
rect 16942 269778 17026 270014
rect 17262 269778 376706 270014
rect 376942 269778 377026 270014
rect 377262 269778 412706 270014
rect 412942 269778 413026 270014
rect 413262 269778 448706 270014
rect 448942 269778 449026 270014
rect 449262 269778 484706 270014
rect 484942 269778 485026 270014
rect 485262 269778 520706 270014
rect 520942 269778 521026 270014
rect 521262 269778 556706 270014
rect 556942 269778 557026 270014
rect 557262 269778 589182 270014
rect 589418 269778 589502 270014
rect 589738 269778 592650 270014
rect -8726 269746 592650 269778
rect -8726 266614 592650 266646
rect -8726 266378 -4854 266614
rect -4618 266378 -4534 266614
rect -4298 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 372986 266614
rect 373222 266378 373306 266614
rect 373542 266378 408986 266614
rect 409222 266378 409306 266614
rect 409542 266378 444986 266614
rect 445222 266378 445306 266614
rect 445542 266378 480986 266614
rect 481222 266378 481306 266614
rect 481542 266378 516986 266614
rect 517222 266378 517306 266614
rect 517542 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 588222 266614
rect 588458 266378 588542 266614
rect 588778 266378 592650 266614
rect -8726 266294 592650 266378
rect -8726 266058 -4854 266294
rect -4618 266058 -4534 266294
rect -4298 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 372986 266294
rect 373222 266058 373306 266294
rect 373542 266058 408986 266294
rect 409222 266058 409306 266294
rect 409542 266058 444986 266294
rect 445222 266058 445306 266294
rect 445542 266058 480986 266294
rect 481222 266058 481306 266294
rect 481542 266058 516986 266294
rect 517222 266058 517306 266294
rect 517542 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 588222 266294
rect 588458 266058 588542 266294
rect 588778 266058 592650 266294
rect -8726 266026 592650 266058
rect -8726 262894 592650 262926
rect -8726 262658 -3894 262894
rect -3658 262658 -3574 262894
rect -3338 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 369266 262894
rect 369502 262658 369586 262894
rect 369822 262658 405266 262894
rect 405502 262658 405586 262894
rect 405822 262658 441266 262894
rect 441502 262658 441586 262894
rect 441822 262658 477266 262894
rect 477502 262658 477586 262894
rect 477822 262658 513266 262894
rect 513502 262658 513586 262894
rect 513822 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 587262 262894
rect 587498 262658 587582 262894
rect 587818 262658 592650 262894
rect -8726 262574 592650 262658
rect -8726 262338 -3894 262574
rect -3658 262338 -3574 262574
rect -3338 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 369266 262574
rect 369502 262338 369586 262574
rect 369822 262338 405266 262574
rect 405502 262338 405586 262574
rect 405822 262338 441266 262574
rect 441502 262338 441586 262574
rect 441822 262338 477266 262574
rect 477502 262338 477586 262574
rect 477822 262338 513266 262574
rect 513502 262338 513586 262574
rect 513822 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 587262 262574
rect 587498 262338 587582 262574
rect 587818 262338 592650 262574
rect -8726 262306 592650 262338
rect -8726 259174 592650 259206
rect -8726 258938 -2934 259174
rect -2698 258938 -2614 259174
rect -2378 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 39610 259174
rect 39846 258938 70330 259174
rect 70566 258938 101050 259174
rect 101286 258938 131770 259174
rect 132006 258938 162490 259174
rect 162726 258938 193210 259174
rect 193446 258938 223930 259174
rect 224166 258938 254650 259174
rect 254886 258938 285370 259174
rect 285606 258938 316090 259174
rect 316326 258938 346810 259174
rect 347046 258938 365546 259174
rect 365782 258938 365866 259174
rect 366102 258938 401546 259174
rect 401782 258938 401866 259174
rect 402102 258938 437546 259174
rect 437782 258938 437866 259174
rect 438102 258938 479610 259174
rect 479846 258938 510330 259174
rect 510566 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 586302 259174
rect 586538 258938 586622 259174
rect 586858 258938 592650 259174
rect -8726 258854 592650 258938
rect -8726 258618 -2934 258854
rect -2698 258618 -2614 258854
rect -2378 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 39610 258854
rect 39846 258618 70330 258854
rect 70566 258618 101050 258854
rect 101286 258618 131770 258854
rect 132006 258618 162490 258854
rect 162726 258618 193210 258854
rect 193446 258618 223930 258854
rect 224166 258618 254650 258854
rect 254886 258618 285370 258854
rect 285606 258618 316090 258854
rect 316326 258618 346810 258854
rect 347046 258618 365546 258854
rect 365782 258618 365866 258854
rect 366102 258618 401546 258854
rect 401782 258618 401866 258854
rect 402102 258618 437546 258854
rect 437782 258618 437866 258854
rect 438102 258618 479610 258854
rect 479846 258618 510330 258854
rect 510566 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 586302 258854
rect 586538 258618 586622 258854
rect 586858 258618 592650 258854
rect -8726 258586 592650 258618
rect -8726 255454 592650 255486
rect -8726 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 24250 255454
rect 24486 255218 54970 255454
rect 55206 255218 85690 255454
rect 85926 255218 116410 255454
rect 116646 255218 147130 255454
rect 147366 255218 177850 255454
rect 178086 255218 208570 255454
rect 208806 255218 239290 255454
rect 239526 255218 270010 255454
rect 270246 255218 300730 255454
rect 300966 255218 331450 255454
rect 331686 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 464250 255454
rect 464486 255218 494970 255454
rect 495206 255218 525690 255454
rect 525926 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 592650 255454
rect -8726 255134 592650 255218
rect -8726 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 24250 255134
rect 24486 254898 54970 255134
rect 55206 254898 85690 255134
rect 85926 254898 116410 255134
rect 116646 254898 147130 255134
rect 147366 254898 177850 255134
rect 178086 254898 208570 255134
rect 208806 254898 239290 255134
rect 239526 254898 270010 255134
rect 270246 254898 300730 255134
rect 300966 254898 331450 255134
rect 331686 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 464250 255134
rect 464486 254898 494970 255134
rect 495206 254898 525690 255134
rect 525926 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 592650 255134
rect -8726 254866 592650 254898
rect -8726 245494 592650 245526
rect -8726 245258 -8694 245494
rect -8458 245258 -8374 245494
rect -8138 245258 27866 245494
rect 28102 245258 28186 245494
rect 28422 245258 387866 245494
rect 388102 245258 388186 245494
rect 388422 245258 423866 245494
rect 424102 245258 424186 245494
rect 424422 245258 459866 245494
rect 460102 245258 460186 245494
rect 460422 245258 531866 245494
rect 532102 245258 532186 245494
rect 532422 245258 567866 245494
rect 568102 245258 568186 245494
rect 568422 245258 592062 245494
rect 592298 245258 592382 245494
rect 592618 245258 592650 245494
rect -8726 245174 592650 245258
rect -8726 244938 -8694 245174
rect -8458 244938 -8374 245174
rect -8138 244938 27866 245174
rect 28102 244938 28186 245174
rect 28422 244938 387866 245174
rect 388102 244938 388186 245174
rect 388422 244938 423866 245174
rect 424102 244938 424186 245174
rect 424422 244938 459866 245174
rect 460102 244938 460186 245174
rect 460422 244938 531866 245174
rect 532102 244938 532186 245174
rect 532422 244938 567866 245174
rect 568102 244938 568186 245174
rect 568422 244938 592062 245174
rect 592298 244938 592382 245174
rect 592618 244938 592650 245174
rect -8726 244906 592650 244938
rect -8726 241774 592650 241806
rect -8726 241538 -7734 241774
rect -7498 241538 -7414 241774
rect -7178 241538 384146 241774
rect 384382 241538 384466 241774
rect 384702 241538 420146 241774
rect 420382 241538 420466 241774
rect 420702 241538 456146 241774
rect 456382 241538 456466 241774
rect 456702 241538 564146 241774
rect 564382 241538 564466 241774
rect 564702 241538 591102 241774
rect 591338 241538 591422 241774
rect 591658 241538 592650 241774
rect -8726 241454 592650 241538
rect -8726 241218 -7734 241454
rect -7498 241218 -7414 241454
rect -7178 241218 384146 241454
rect 384382 241218 384466 241454
rect 384702 241218 420146 241454
rect 420382 241218 420466 241454
rect 420702 241218 456146 241454
rect 456382 241218 456466 241454
rect 456702 241218 564146 241454
rect 564382 241218 564466 241454
rect 564702 241218 591102 241454
rect 591338 241218 591422 241454
rect 591658 241218 592650 241454
rect -8726 241186 592650 241218
rect -8726 238054 592650 238086
rect -8726 237818 -6774 238054
rect -6538 237818 -6454 238054
rect -6218 237818 20426 238054
rect 20662 237818 20746 238054
rect 20982 237818 380426 238054
rect 380662 237818 380746 238054
rect 380982 237818 416426 238054
rect 416662 237818 416746 238054
rect 416982 237818 452426 238054
rect 452662 237818 452746 238054
rect 452982 237818 560426 238054
rect 560662 237818 560746 238054
rect 560982 237818 590142 238054
rect 590378 237818 590462 238054
rect 590698 237818 592650 238054
rect -8726 237734 592650 237818
rect -8726 237498 -6774 237734
rect -6538 237498 -6454 237734
rect -6218 237498 20426 237734
rect 20662 237498 20746 237734
rect 20982 237498 380426 237734
rect 380662 237498 380746 237734
rect 380982 237498 416426 237734
rect 416662 237498 416746 237734
rect 416982 237498 452426 237734
rect 452662 237498 452746 237734
rect 452982 237498 560426 237734
rect 560662 237498 560746 237734
rect 560982 237498 590142 237734
rect 590378 237498 590462 237734
rect 590698 237498 592650 237734
rect -8726 237466 592650 237498
rect -8726 234334 592650 234366
rect -8726 234098 -5814 234334
rect -5578 234098 -5494 234334
rect -5258 234098 16706 234334
rect 16942 234098 17026 234334
rect 17262 234098 376706 234334
rect 376942 234098 377026 234334
rect 377262 234098 412706 234334
rect 412942 234098 413026 234334
rect 413262 234098 448706 234334
rect 448942 234098 449026 234334
rect 449262 234098 556706 234334
rect 556942 234098 557026 234334
rect 557262 234098 589182 234334
rect 589418 234098 589502 234334
rect 589738 234098 592650 234334
rect -8726 234014 592650 234098
rect -8726 233778 -5814 234014
rect -5578 233778 -5494 234014
rect -5258 233778 16706 234014
rect 16942 233778 17026 234014
rect 17262 233778 376706 234014
rect 376942 233778 377026 234014
rect 377262 233778 412706 234014
rect 412942 233778 413026 234014
rect 413262 233778 448706 234014
rect 448942 233778 449026 234014
rect 449262 233778 556706 234014
rect 556942 233778 557026 234014
rect 557262 233778 589182 234014
rect 589418 233778 589502 234014
rect 589738 233778 592650 234014
rect -8726 233746 592650 233778
rect -8726 230614 592650 230646
rect -8726 230378 -4854 230614
rect -4618 230378 -4534 230614
rect -4298 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 372986 230614
rect 373222 230378 373306 230614
rect 373542 230378 408986 230614
rect 409222 230378 409306 230614
rect 409542 230378 444986 230614
rect 445222 230378 445306 230614
rect 445542 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 588222 230614
rect 588458 230378 588542 230614
rect 588778 230378 592650 230614
rect -8726 230294 592650 230378
rect -8726 230058 -4854 230294
rect -4618 230058 -4534 230294
rect -4298 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 372986 230294
rect 373222 230058 373306 230294
rect 373542 230058 408986 230294
rect 409222 230058 409306 230294
rect 409542 230058 444986 230294
rect 445222 230058 445306 230294
rect 445542 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 588222 230294
rect 588458 230058 588542 230294
rect 588778 230058 592650 230294
rect -8726 230026 592650 230058
rect -8726 226894 592650 226926
rect -8726 226658 -3894 226894
rect -3658 226658 -3574 226894
rect -3338 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 369266 226894
rect 369502 226658 369586 226894
rect 369822 226658 405266 226894
rect 405502 226658 405586 226894
rect 405822 226658 441266 226894
rect 441502 226658 441586 226894
rect 441822 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 587262 226894
rect 587498 226658 587582 226894
rect 587818 226658 592650 226894
rect -8726 226574 592650 226658
rect -8726 226338 -3894 226574
rect -3658 226338 -3574 226574
rect -3338 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 369266 226574
rect 369502 226338 369586 226574
rect 369822 226338 405266 226574
rect 405502 226338 405586 226574
rect 405822 226338 441266 226574
rect 441502 226338 441586 226574
rect 441822 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 587262 226574
rect 587498 226338 587582 226574
rect 587818 226338 592650 226574
rect -8726 226306 592650 226338
rect -8726 223174 592650 223206
rect -8726 222938 -2934 223174
rect -2698 222938 -2614 223174
rect -2378 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 39610 223174
rect 39846 222938 70330 223174
rect 70566 222938 101050 223174
rect 101286 222938 131770 223174
rect 132006 222938 162490 223174
rect 162726 222938 193210 223174
rect 193446 222938 223930 223174
rect 224166 222938 254650 223174
rect 254886 222938 285370 223174
rect 285606 222938 316090 223174
rect 316326 222938 346810 223174
rect 347046 222938 365546 223174
rect 365782 222938 365866 223174
rect 366102 222938 401546 223174
rect 401782 222938 401866 223174
rect 402102 222938 437546 223174
rect 437782 222938 437866 223174
rect 438102 222938 479610 223174
rect 479846 222938 510330 223174
rect 510566 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 586302 223174
rect 586538 222938 586622 223174
rect 586858 222938 592650 223174
rect -8726 222854 592650 222938
rect -8726 222618 -2934 222854
rect -2698 222618 -2614 222854
rect -2378 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 39610 222854
rect 39846 222618 70330 222854
rect 70566 222618 101050 222854
rect 101286 222618 131770 222854
rect 132006 222618 162490 222854
rect 162726 222618 193210 222854
rect 193446 222618 223930 222854
rect 224166 222618 254650 222854
rect 254886 222618 285370 222854
rect 285606 222618 316090 222854
rect 316326 222618 346810 222854
rect 347046 222618 365546 222854
rect 365782 222618 365866 222854
rect 366102 222618 401546 222854
rect 401782 222618 401866 222854
rect 402102 222618 437546 222854
rect 437782 222618 437866 222854
rect 438102 222618 479610 222854
rect 479846 222618 510330 222854
rect 510566 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 586302 222854
rect 586538 222618 586622 222854
rect 586858 222618 592650 222854
rect -8726 222586 592650 222618
rect -8726 219454 592650 219486
rect -8726 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 24250 219454
rect 24486 219218 54970 219454
rect 55206 219218 85690 219454
rect 85926 219218 116410 219454
rect 116646 219218 147130 219454
rect 147366 219218 177850 219454
rect 178086 219218 208570 219454
rect 208806 219218 239290 219454
rect 239526 219218 270010 219454
rect 270246 219218 300730 219454
rect 300966 219218 331450 219454
rect 331686 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 464250 219454
rect 464486 219218 494970 219454
rect 495206 219218 525690 219454
rect 525926 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 592650 219454
rect -8726 219134 592650 219218
rect -8726 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 24250 219134
rect 24486 218898 54970 219134
rect 55206 218898 85690 219134
rect 85926 218898 116410 219134
rect 116646 218898 147130 219134
rect 147366 218898 177850 219134
rect 178086 218898 208570 219134
rect 208806 218898 239290 219134
rect 239526 218898 270010 219134
rect 270246 218898 300730 219134
rect 300966 218898 331450 219134
rect 331686 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 464250 219134
rect 464486 218898 494970 219134
rect 495206 218898 525690 219134
rect 525926 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 592650 219134
rect -8726 218866 592650 218898
rect -8726 209494 592650 209526
rect -8726 209258 -8694 209494
rect -8458 209258 -8374 209494
rect -8138 209258 27866 209494
rect 28102 209258 28186 209494
rect 28422 209258 387866 209494
rect 388102 209258 388186 209494
rect 388422 209258 423866 209494
rect 424102 209258 424186 209494
rect 424422 209258 459866 209494
rect 460102 209258 460186 209494
rect 460422 209258 531866 209494
rect 532102 209258 532186 209494
rect 532422 209258 567866 209494
rect 568102 209258 568186 209494
rect 568422 209258 592062 209494
rect 592298 209258 592382 209494
rect 592618 209258 592650 209494
rect -8726 209174 592650 209258
rect -8726 208938 -8694 209174
rect -8458 208938 -8374 209174
rect -8138 208938 27866 209174
rect 28102 208938 28186 209174
rect 28422 208938 387866 209174
rect 388102 208938 388186 209174
rect 388422 208938 423866 209174
rect 424102 208938 424186 209174
rect 424422 208938 459866 209174
rect 460102 208938 460186 209174
rect 460422 208938 531866 209174
rect 532102 208938 532186 209174
rect 532422 208938 567866 209174
rect 568102 208938 568186 209174
rect 568422 208938 592062 209174
rect 592298 208938 592382 209174
rect 592618 208938 592650 209174
rect -8726 208906 592650 208938
rect -8726 205774 592650 205806
rect -8726 205538 -7734 205774
rect -7498 205538 -7414 205774
rect -7178 205538 384146 205774
rect 384382 205538 384466 205774
rect 384702 205538 420146 205774
rect 420382 205538 420466 205774
rect 420702 205538 456146 205774
rect 456382 205538 456466 205774
rect 456702 205538 564146 205774
rect 564382 205538 564466 205774
rect 564702 205538 591102 205774
rect 591338 205538 591422 205774
rect 591658 205538 592650 205774
rect -8726 205454 592650 205538
rect -8726 205218 -7734 205454
rect -7498 205218 -7414 205454
rect -7178 205218 384146 205454
rect 384382 205218 384466 205454
rect 384702 205218 420146 205454
rect 420382 205218 420466 205454
rect 420702 205218 456146 205454
rect 456382 205218 456466 205454
rect 456702 205218 564146 205454
rect 564382 205218 564466 205454
rect 564702 205218 591102 205454
rect 591338 205218 591422 205454
rect 591658 205218 592650 205454
rect -8726 205186 592650 205218
rect -8726 202054 592650 202086
rect -8726 201818 -6774 202054
rect -6538 201818 -6454 202054
rect -6218 201818 20426 202054
rect 20662 201818 20746 202054
rect 20982 201818 380426 202054
rect 380662 201818 380746 202054
rect 380982 201818 416426 202054
rect 416662 201818 416746 202054
rect 416982 201818 452426 202054
rect 452662 201818 452746 202054
rect 452982 201818 560426 202054
rect 560662 201818 560746 202054
rect 560982 201818 590142 202054
rect 590378 201818 590462 202054
rect 590698 201818 592650 202054
rect -8726 201734 592650 201818
rect -8726 201498 -6774 201734
rect -6538 201498 -6454 201734
rect -6218 201498 20426 201734
rect 20662 201498 20746 201734
rect 20982 201498 380426 201734
rect 380662 201498 380746 201734
rect 380982 201498 416426 201734
rect 416662 201498 416746 201734
rect 416982 201498 452426 201734
rect 452662 201498 452746 201734
rect 452982 201498 560426 201734
rect 560662 201498 560746 201734
rect 560982 201498 590142 201734
rect 590378 201498 590462 201734
rect 590698 201498 592650 201734
rect -8726 201466 592650 201498
rect -8726 198334 592650 198366
rect -8726 198098 -5814 198334
rect -5578 198098 -5494 198334
rect -5258 198098 16706 198334
rect 16942 198098 17026 198334
rect 17262 198098 376706 198334
rect 376942 198098 377026 198334
rect 377262 198098 412706 198334
rect 412942 198098 413026 198334
rect 413262 198098 448706 198334
rect 448942 198098 449026 198334
rect 449262 198098 484706 198334
rect 484942 198098 485026 198334
rect 485262 198098 520706 198334
rect 520942 198098 521026 198334
rect 521262 198098 556706 198334
rect 556942 198098 557026 198334
rect 557262 198098 589182 198334
rect 589418 198098 589502 198334
rect 589738 198098 592650 198334
rect -8726 198014 592650 198098
rect -8726 197778 -5814 198014
rect -5578 197778 -5494 198014
rect -5258 197778 16706 198014
rect 16942 197778 17026 198014
rect 17262 197778 376706 198014
rect 376942 197778 377026 198014
rect 377262 197778 412706 198014
rect 412942 197778 413026 198014
rect 413262 197778 448706 198014
rect 448942 197778 449026 198014
rect 449262 197778 484706 198014
rect 484942 197778 485026 198014
rect 485262 197778 520706 198014
rect 520942 197778 521026 198014
rect 521262 197778 556706 198014
rect 556942 197778 557026 198014
rect 557262 197778 589182 198014
rect 589418 197778 589502 198014
rect 589738 197778 592650 198014
rect -8726 197746 592650 197778
rect -8726 194614 592650 194646
rect -8726 194378 -4854 194614
rect -4618 194378 -4534 194614
rect -4298 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 372986 194614
rect 373222 194378 373306 194614
rect 373542 194378 408986 194614
rect 409222 194378 409306 194614
rect 409542 194378 444986 194614
rect 445222 194378 445306 194614
rect 445542 194378 480986 194614
rect 481222 194378 481306 194614
rect 481542 194378 516986 194614
rect 517222 194378 517306 194614
rect 517542 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 588222 194614
rect 588458 194378 588542 194614
rect 588778 194378 592650 194614
rect -8726 194294 592650 194378
rect -8726 194058 -4854 194294
rect -4618 194058 -4534 194294
rect -4298 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 372986 194294
rect 373222 194058 373306 194294
rect 373542 194058 408986 194294
rect 409222 194058 409306 194294
rect 409542 194058 444986 194294
rect 445222 194058 445306 194294
rect 445542 194058 480986 194294
rect 481222 194058 481306 194294
rect 481542 194058 516986 194294
rect 517222 194058 517306 194294
rect 517542 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 588222 194294
rect 588458 194058 588542 194294
rect 588778 194058 592650 194294
rect -8726 194026 592650 194058
rect -8726 190894 592650 190926
rect -8726 190658 -3894 190894
rect -3658 190658 -3574 190894
rect -3338 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 369266 190894
rect 369502 190658 369586 190894
rect 369822 190658 405266 190894
rect 405502 190658 405586 190894
rect 405822 190658 441266 190894
rect 441502 190658 441586 190894
rect 441822 190658 477266 190894
rect 477502 190658 477586 190894
rect 477822 190658 513266 190894
rect 513502 190658 513586 190894
rect 513822 190658 549266 190894
rect 549502 190658 549586 190894
rect 549822 190658 587262 190894
rect 587498 190658 587582 190894
rect 587818 190658 592650 190894
rect -8726 190574 592650 190658
rect -8726 190338 -3894 190574
rect -3658 190338 -3574 190574
rect -3338 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 369266 190574
rect 369502 190338 369586 190574
rect 369822 190338 405266 190574
rect 405502 190338 405586 190574
rect 405822 190338 441266 190574
rect 441502 190338 441586 190574
rect 441822 190338 477266 190574
rect 477502 190338 477586 190574
rect 477822 190338 513266 190574
rect 513502 190338 513586 190574
rect 513822 190338 549266 190574
rect 549502 190338 549586 190574
rect 549822 190338 587262 190574
rect 587498 190338 587582 190574
rect 587818 190338 592650 190574
rect -8726 190306 592650 190338
rect -8726 187174 592650 187206
rect -8726 186938 -2934 187174
rect -2698 186938 -2614 187174
rect -2378 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 39610 187174
rect 39846 186938 70330 187174
rect 70566 186938 101050 187174
rect 101286 186938 131770 187174
rect 132006 186938 162490 187174
rect 162726 186938 193210 187174
rect 193446 186938 223930 187174
rect 224166 186938 254650 187174
rect 254886 186938 285370 187174
rect 285606 186938 316090 187174
rect 316326 186938 346810 187174
rect 347046 186938 365546 187174
rect 365782 186938 365866 187174
rect 366102 186938 401546 187174
rect 401782 186938 401866 187174
rect 402102 186938 437546 187174
rect 437782 186938 437866 187174
rect 438102 186938 473546 187174
rect 473782 186938 473866 187174
rect 474102 186938 509546 187174
rect 509782 186938 509866 187174
rect 510102 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 586302 187174
rect 586538 186938 586622 187174
rect 586858 186938 592650 187174
rect -8726 186854 592650 186938
rect -8726 186618 -2934 186854
rect -2698 186618 -2614 186854
rect -2378 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 39610 186854
rect 39846 186618 70330 186854
rect 70566 186618 101050 186854
rect 101286 186618 131770 186854
rect 132006 186618 162490 186854
rect 162726 186618 193210 186854
rect 193446 186618 223930 186854
rect 224166 186618 254650 186854
rect 254886 186618 285370 186854
rect 285606 186618 316090 186854
rect 316326 186618 346810 186854
rect 347046 186618 365546 186854
rect 365782 186618 365866 186854
rect 366102 186618 401546 186854
rect 401782 186618 401866 186854
rect 402102 186618 437546 186854
rect 437782 186618 437866 186854
rect 438102 186618 473546 186854
rect 473782 186618 473866 186854
rect 474102 186618 509546 186854
rect 509782 186618 509866 186854
rect 510102 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 586302 186854
rect 586538 186618 586622 186854
rect 586858 186618 592650 186854
rect -8726 186586 592650 186618
rect -8726 183454 592650 183486
rect -8726 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 24250 183454
rect 24486 183218 54970 183454
rect 55206 183218 85690 183454
rect 85926 183218 116410 183454
rect 116646 183218 147130 183454
rect 147366 183218 177850 183454
rect 178086 183218 208570 183454
rect 208806 183218 239290 183454
rect 239526 183218 270010 183454
rect 270246 183218 300730 183454
rect 300966 183218 331450 183454
rect 331686 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 592650 183454
rect -8726 183134 592650 183218
rect -8726 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 24250 183134
rect 24486 182898 54970 183134
rect 55206 182898 85690 183134
rect 85926 182898 116410 183134
rect 116646 182898 147130 183134
rect 147366 182898 177850 183134
rect 178086 182898 208570 183134
rect 208806 182898 239290 183134
rect 239526 182898 270010 183134
rect 270246 182898 300730 183134
rect 300966 182898 331450 183134
rect 331686 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 592650 183134
rect -8726 182866 592650 182898
rect -8726 173494 592650 173526
rect -8726 173258 -8694 173494
rect -8458 173258 -8374 173494
rect -8138 173258 27866 173494
rect 28102 173258 28186 173494
rect 28422 173258 387866 173494
rect 388102 173258 388186 173494
rect 388422 173258 423866 173494
rect 424102 173258 424186 173494
rect 424422 173258 459866 173494
rect 460102 173258 460186 173494
rect 460422 173258 531866 173494
rect 532102 173258 532186 173494
rect 532422 173258 567866 173494
rect 568102 173258 568186 173494
rect 568422 173258 592062 173494
rect 592298 173258 592382 173494
rect 592618 173258 592650 173494
rect -8726 173174 592650 173258
rect -8726 172938 -8694 173174
rect -8458 172938 -8374 173174
rect -8138 172938 27866 173174
rect 28102 172938 28186 173174
rect 28422 172938 387866 173174
rect 388102 172938 388186 173174
rect 388422 172938 423866 173174
rect 424102 172938 424186 173174
rect 424422 172938 459866 173174
rect 460102 172938 460186 173174
rect 460422 172938 531866 173174
rect 532102 172938 532186 173174
rect 532422 172938 567866 173174
rect 568102 172938 568186 173174
rect 568422 172938 592062 173174
rect 592298 172938 592382 173174
rect 592618 172938 592650 173174
rect -8726 172906 592650 172938
rect -8726 169774 592650 169806
rect -8726 169538 -7734 169774
rect -7498 169538 -7414 169774
rect -7178 169538 384146 169774
rect 384382 169538 384466 169774
rect 384702 169538 420146 169774
rect 420382 169538 420466 169774
rect 420702 169538 456146 169774
rect 456382 169538 456466 169774
rect 456702 169538 564146 169774
rect 564382 169538 564466 169774
rect 564702 169538 591102 169774
rect 591338 169538 591422 169774
rect 591658 169538 592650 169774
rect -8726 169454 592650 169538
rect -8726 169218 -7734 169454
rect -7498 169218 -7414 169454
rect -7178 169218 384146 169454
rect 384382 169218 384466 169454
rect 384702 169218 420146 169454
rect 420382 169218 420466 169454
rect 420702 169218 456146 169454
rect 456382 169218 456466 169454
rect 456702 169218 564146 169454
rect 564382 169218 564466 169454
rect 564702 169218 591102 169454
rect 591338 169218 591422 169454
rect 591658 169218 592650 169454
rect -8726 169186 592650 169218
rect -8726 166054 592650 166086
rect -8726 165818 -6774 166054
rect -6538 165818 -6454 166054
rect -6218 165818 20426 166054
rect 20662 165818 20746 166054
rect 20982 165818 380426 166054
rect 380662 165818 380746 166054
rect 380982 165818 416426 166054
rect 416662 165818 416746 166054
rect 416982 165818 452426 166054
rect 452662 165818 452746 166054
rect 452982 165818 488426 166054
rect 488662 165818 488746 166054
rect 488982 165818 524426 166054
rect 524662 165818 524746 166054
rect 524982 165818 560426 166054
rect 560662 165818 560746 166054
rect 560982 165818 590142 166054
rect 590378 165818 590462 166054
rect 590698 165818 592650 166054
rect -8726 165734 592650 165818
rect -8726 165498 -6774 165734
rect -6538 165498 -6454 165734
rect -6218 165498 20426 165734
rect 20662 165498 20746 165734
rect 20982 165498 380426 165734
rect 380662 165498 380746 165734
rect 380982 165498 416426 165734
rect 416662 165498 416746 165734
rect 416982 165498 452426 165734
rect 452662 165498 452746 165734
rect 452982 165498 488426 165734
rect 488662 165498 488746 165734
rect 488982 165498 524426 165734
rect 524662 165498 524746 165734
rect 524982 165498 560426 165734
rect 560662 165498 560746 165734
rect 560982 165498 590142 165734
rect 590378 165498 590462 165734
rect 590698 165498 592650 165734
rect -8726 165466 592650 165498
rect -8726 162334 592650 162366
rect -8726 162098 -5814 162334
rect -5578 162098 -5494 162334
rect -5258 162098 16706 162334
rect 16942 162098 17026 162334
rect 17262 162098 376706 162334
rect 376942 162098 377026 162334
rect 377262 162098 412706 162334
rect 412942 162098 413026 162334
rect 413262 162098 448706 162334
rect 448942 162098 449026 162334
rect 449262 162098 484706 162334
rect 484942 162098 485026 162334
rect 485262 162098 520706 162334
rect 520942 162098 521026 162334
rect 521262 162098 556706 162334
rect 556942 162098 557026 162334
rect 557262 162098 589182 162334
rect 589418 162098 589502 162334
rect 589738 162098 592650 162334
rect -8726 162014 592650 162098
rect -8726 161778 -5814 162014
rect -5578 161778 -5494 162014
rect -5258 161778 16706 162014
rect 16942 161778 17026 162014
rect 17262 161778 376706 162014
rect 376942 161778 377026 162014
rect 377262 161778 412706 162014
rect 412942 161778 413026 162014
rect 413262 161778 448706 162014
rect 448942 161778 449026 162014
rect 449262 161778 484706 162014
rect 484942 161778 485026 162014
rect 485262 161778 520706 162014
rect 520942 161778 521026 162014
rect 521262 161778 556706 162014
rect 556942 161778 557026 162014
rect 557262 161778 589182 162014
rect 589418 161778 589502 162014
rect 589738 161778 592650 162014
rect -8726 161746 592650 161778
rect -8726 158614 592650 158646
rect -8726 158378 -4854 158614
rect -4618 158378 -4534 158614
rect -4298 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 372986 158614
rect 373222 158378 373306 158614
rect 373542 158378 408986 158614
rect 409222 158378 409306 158614
rect 409542 158378 480986 158614
rect 481222 158378 481306 158614
rect 481542 158378 516986 158614
rect 517222 158378 517306 158614
rect 517542 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 588222 158614
rect 588458 158378 588542 158614
rect 588778 158378 592650 158614
rect -8726 158294 592650 158378
rect -8726 158058 -4854 158294
rect -4618 158058 -4534 158294
rect -4298 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 372986 158294
rect 373222 158058 373306 158294
rect 373542 158058 408986 158294
rect 409222 158058 409306 158294
rect 409542 158058 480986 158294
rect 481222 158058 481306 158294
rect 481542 158058 516986 158294
rect 517222 158058 517306 158294
rect 517542 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 588222 158294
rect 588458 158058 588542 158294
rect 588778 158058 592650 158294
rect -8726 158026 592650 158058
rect -8726 154894 592650 154926
rect -8726 154658 -3894 154894
rect -3658 154658 -3574 154894
rect -3338 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 369266 154894
rect 369502 154658 369586 154894
rect 369822 154658 405266 154894
rect 405502 154658 405586 154894
rect 405822 154658 477266 154894
rect 477502 154658 477586 154894
rect 477822 154658 513266 154894
rect 513502 154658 513586 154894
rect 513822 154658 549266 154894
rect 549502 154658 549586 154894
rect 549822 154658 587262 154894
rect 587498 154658 587582 154894
rect 587818 154658 592650 154894
rect -8726 154574 592650 154658
rect -8726 154338 -3894 154574
rect -3658 154338 -3574 154574
rect -3338 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 369266 154574
rect 369502 154338 369586 154574
rect 369822 154338 405266 154574
rect 405502 154338 405586 154574
rect 405822 154338 477266 154574
rect 477502 154338 477586 154574
rect 477822 154338 513266 154574
rect 513502 154338 513586 154574
rect 513822 154338 549266 154574
rect 549502 154338 549586 154574
rect 549822 154338 587262 154574
rect 587498 154338 587582 154574
rect 587818 154338 592650 154574
rect -8726 154306 592650 154338
rect -8726 151174 592650 151206
rect -8726 150938 -2934 151174
rect -2698 150938 -2614 151174
rect -2378 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 39610 151174
rect 39846 150938 70330 151174
rect 70566 150938 101050 151174
rect 101286 150938 131770 151174
rect 132006 150938 162490 151174
rect 162726 150938 193210 151174
rect 193446 150938 223930 151174
rect 224166 150938 254650 151174
rect 254886 150938 285370 151174
rect 285606 150938 316090 151174
rect 316326 150938 346810 151174
rect 347046 150938 365546 151174
rect 365782 150938 365866 151174
rect 366102 150938 401546 151174
rect 401782 150938 401866 151174
rect 402102 150938 429610 151174
rect 429846 150938 473546 151174
rect 473782 150938 473866 151174
rect 474102 150938 509546 151174
rect 509782 150938 509866 151174
rect 510102 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 586302 151174
rect 586538 150938 586622 151174
rect 586858 150938 592650 151174
rect -8726 150854 592650 150938
rect -8726 150618 -2934 150854
rect -2698 150618 -2614 150854
rect -2378 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 39610 150854
rect 39846 150618 70330 150854
rect 70566 150618 101050 150854
rect 101286 150618 131770 150854
rect 132006 150618 162490 150854
rect 162726 150618 193210 150854
rect 193446 150618 223930 150854
rect 224166 150618 254650 150854
rect 254886 150618 285370 150854
rect 285606 150618 316090 150854
rect 316326 150618 346810 150854
rect 347046 150618 365546 150854
rect 365782 150618 365866 150854
rect 366102 150618 401546 150854
rect 401782 150618 401866 150854
rect 402102 150618 429610 150854
rect 429846 150618 473546 150854
rect 473782 150618 473866 150854
rect 474102 150618 509546 150854
rect 509782 150618 509866 150854
rect 510102 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 586302 150854
rect 586538 150618 586622 150854
rect 586858 150618 592650 150854
rect -8726 150586 592650 150618
rect -8726 147454 592650 147486
rect -8726 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 24250 147454
rect 24486 147218 54970 147454
rect 55206 147218 85690 147454
rect 85926 147218 116410 147454
rect 116646 147218 147130 147454
rect 147366 147218 177850 147454
rect 178086 147218 208570 147454
rect 208806 147218 239290 147454
rect 239526 147218 270010 147454
rect 270246 147218 300730 147454
rect 300966 147218 331450 147454
rect 331686 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 414250 147454
rect 414486 147218 444970 147454
rect 445206 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 592650 147454
rect -8726 147134 592650 147218
rect -8726 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 24250 147134
rect 24486 146898 54970 147134
rect 55206 146898 85690 147134
rect 85926 146898 116410 147134
rect 116646 146898 147130 147134
rect 147366 146898 177850 147134
rect 178086 146898 208570 147134
rect 208806 146898 239290 147134
rect 239526 146898 270010 147134
rect 270246 146898 300730 147134
rect 300966 146898 331450 147134
rect 331686 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 414250 147134
rect 414486 146898 444970 147134
rect 445206 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 592650 147134
rect -8726 146866 592650 146898
rect -8726 137494 592650 137526
rect -8726 137258 -8694 137494
rect -8458 137258 -8374 137494
rect -8138 137258 27866 137494
rect 28102 137258 28186 137494
rect 28422 137258 387866 137494
rect 388102 137258 388186 137494
rect 388422 137258 459866 137494
rect 460102 137258 460186 137494
rect 460422 137258 567866 137494
rect 568102 137258 568186 137494
rect 568422 137258 592062 137494
rect 592298 137258 592382 137494
rect 592618 137258 592650 137494
rect -8726 137174 592650 137258
rect -8726 136938 -8694 137174
rect -8458 136938 -8374 137174
rect -8138 136938 27866 137174
rect 28102 136938 28186 137174
rect 28422 136938 387866 137174
rect 388102 136938 388186 137174
rect 388422 136938 459866 137174
rect 460102 136938 460186 137174
rect 460422 136938 567866 137174
rect 568102 136938 568186 137174
rect 568422 136938 592062 137174
rect 592298 136938 592382 137174
rect 592618 136938 592650 137174
rect -8726 136906 592650 136938
rect -8726 133774 592650 133806
rect -8726 133538 -7734 133774
rect -7498 133538 -7414 133774
rect -7178 133538 384146 133774
rect 384382 133538 384466 133774
rect 384702 133538 456146 133774
rect 456382 133538 456466 133774
rect 456702 133538 564146 133774
rect 564382 133538 564466 133774
rect 564702 133538 591102 133774
rect 591338 133538 591422 133774
rect 591658 133538 592650 133774
rect -8726 133454 592650 133538
rect -8726 133218 -7734 133454
rect -7498 133218 -7414 133454
rect -7178 133218 384146 133454
rect 384382 133218 384466 133454
rect 384702 133218 456146 133454
rect 456382 133218 456466 133454
rect 456702 133218 564146 133454
rect 564382 133218 564466 133454
rect 564702 133218 591102 133454
rect 591338 133218 591422 133454
rect 591658 133218 592650 133454
rect -8726 133186 592650 133218
rect -8726 130054 592650 130086
rect -8726 129818 -6774 130054
rect -6538 129818 -6454 130054
rect -6218 129818 20426 130054
rect 20662 129818 20746 130054
rect 20982 129818 380426 130054
rect 380662 129818 380746 130054
rect 380982 129818 452426 130054
rect 452662 129818 452746 130054
rect 452982 129818 560426 130054
rect 560662 129818 560746 130054
rect 560982 129818 590142 130054
rect 590378 129818 590462 130054
rect 590698 129818 592650 130054
rect -8726 129734 592650 129818
rect -8726 129498 -6774 129734
rect -6538 129498 -6454 129734
rect -6218 129498 20426 129734
rect 20662 129498 20746 129734
rect 20982 129498 380426 129734
rect 380662 129498 380746 129734
rect 380982 129498 452426 129734
rect 452662 129498 452746 129734
rect 452982 129498 560426 129734
rect 560662 129498 560746 129734
rect 560982 129498 590142 129734
rect 590378 129498 590462 129734
rect 590698 129498 592650 129734
rect -8726 129466 592650 129498
rect -8726 126334 592650 126366
rect -8726 126098 -5814 126334
rect -5578 126098 -5494 126334
rect -5258 126098 16706 126334
rect 16942 126098 17026 126334
rect 17262 126098 376706 126334
rect 376942 126098 377026 126334
rect 377262 126098 412706 126334
rect 412942 126098 413026 126334
rect 413262 126098 448706 126334
rect 448942 126098 449026 126334
rect 449262 126098 484706 126334
rect 484942 126098 485026 126334
rect 485262 126098 556706 126334
rect 556942 126098 557026 126334
rect 557262 126098 589182 126334
rect 589418 126098 589502 126334
rect 589738 126098 592650 126334
rect -8726 126014 592650 126098
rect -8726 125778 -5814 126014
rect -5578 125778 -5494 126014
rect -5258 125778 16706 126014
rect 16942 125778 17026 126014
rect 17262 125778 376706 126014
rect 376942 125778 377026 126014
rect 377262 125778 412706 126014
rect 412942 125778 413026 126014
rect 413262 125778 448706 126014
rect 448942 125778 449026 126014
rect 449262 125778 484706 126014
rect 484942 125778 485026 126014
rect 485262 125778 556706 126014
rect 556942 125778 557026 126014
rect 557262 125778 589182 126014
rect 589418 125778 589502 126014
rect 589738 125778 592650 126014
rect -8726 125746 592650 125778
rect -8726 122614 592650 122646
rect -8726 122378 -4854 122614
rect -4618 122378 -4534 122614
rect -4298 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 372986 122614
rect 373222 122378 373306 122614
rect 373542 122378 408986 122614
rect 409222 122378 409306 122614
rect 409542 122378 480986 122614
rect 481222 122378 481306 122614
rect 481542 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 588222 122614
rect 588458 122378 588542 122614
rect 588778 122378 592650 122614
rect -8726 122294 592650 122378
rect -8726 122058 -4854 122294
rect -4618 122058 -4534 122294
rect -4298 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 372986 122294
rect 373222 122058 373306 122294
rect 373542 122058 408986 122294
rect 409222 122058 409306 122294
rect 409542 122058 480986 122294
rect 481222 122058 481306 122294
rect 481542 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 588222 122294
rect 588458 122058 588542 122294
rect 588778 122058 592650 122294
rect -8726 122026 592650 122058
rect -8726 118894 592650 118926
rect -8726 118658 -3894 118894
rect -3658 118658 -3574 118894
rect -3338 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 369266 118894
rect 369502 118658 369586 118894
rect 369822 118658 405266 118894
rect 405502 118658 405586 118894
rect 405822 118658 477266 118894
rect 477502 118658 477586 118894
rect 477822 118658 549266 118894
rect 549502 118658 549586 118894
rect 549822 118658 587262 118894
rect 587498 118658 587582 118894
rect 587818 118658 592650 118894
rect -8726 118574 592650 118658
rect -8726 118338 -3894 118574
rect -3658 118338 -3574 118574
rect -3338 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 369266 118574
rect 369502 118338 369586 118574
rect 369822 118338 405266 118574
rect 405502 118338 405586 118574
rect 405822 118338 477266 118574
rect 477502 118338 477586 118574
rect 477822 118338 549266 118574
rect 549502 118338 549586 118574
rect 549822 118338 587262 118574
rect 587498 118338 587582 118574
rect 587818 118338 592650 118574
rect -8726 118306 592650 118338
rect -8726 115174 592650 115206
rect -8726 114938 -2934 115174
rect -2698 114938 -2614 115174
rect -2378 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 39610 115174
rect 39846 114938 70330 115174
rect 70566 114938 101050 115174
rect 101286 114938 131770 115174
rect 132006 114938 162490 115174
rect 162726 114938 193210 115174
rect 193446 114938 223930 115174
rect 224166 114938 254650 115174
rect 254886 114938 285370 115174
rect 285606 114938 316090 115174
rect 316326 114938 346810 115174
rect 347046 114938 365546 115174
rect 365782 114938 365866 115174
rect 366102 114938 401546 115174
rect 401782 114938 401866 115174
rect 402102 114938 473546 115174
rect 473782 114938 473866 115174
rect 474102 114938 499610 115174
rect 499846 114938 530330 115174
rect 530566 114938 545546 115174
rect 545782 114938 545866 115174
rect 546102 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 586302 115174
rect 586538 114938 586622 115174
rect 586858 114938 592650 115174
rect -8726 114854 592650 114938
rect -8726 114618 -2934 114854
rect -2698 114618 -2614 114854
rect -2378 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 39610 114854
rect 39846 114618 70330 114854
rect 70566 114618 101050 114854
rect 101286 114618 131770 114854
rect 132006 114618 162490 114854
rect 162726 114618 193210 114854
rect 193446 114618 223930 114854
rect 224166 114618 254650 114854
rect 254886 114618 285370 114854
rect 285606 114618 316090 114854
rect 316326 114618 346810 114854
rect 347046 114618 365546 114854
rect 365782 114618 365866 114854
rect 366102 114618 401546 114854
rect 401782 114618 401866 114854
rect 402102 114618 473546 114854
rect 473782 114618 473866 114854
rect 474102 114618 499610 114854
rect 499846 114618 530330 114854
rect 530566 114618 545546 114854
rect 545782 114618 545866 114854
rect 546102 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 586302 114854
rect 586538 114618 586622 114854
rect 586858 114618 592650 114854
rect -8726 114586 592650 114618
rect -8726 111454 592650 111486
rect -8726 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 24250 111454
rect 24486 111218 54970 111454
rect 55206 111218 85690 111454
rect 85926 111218 116410 111454
rect 116646 111218 147130 111454
rect 147366 111218 177850 111454
rect 178086 111218 208570 111454
rect 208806 111218 239290 111454
rect 239526 111218 270010 111454
rect 270246 111218 300730 111454
rect 300966 111218 331450 111454
rect 331686 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 484250 111454
rect 484486 111218 514970 111454
rect 515206 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 592650 111454
rect -8726 111134 592650 111218
rect -8726 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 24250 111134
rect 24486 110898 54970 111134
rect 55206 110898 85690 111134
rect 85926 110898 116410 111134
rect 116646 110898 147130 111134
rect 147366 110898 177850 111134
rect 178086 110898 208570 111134
rect 208806 110898 239290 111134
rect 239526 110898 270010 111134
rect 270246 110898 300730 111134
rect 300966 110898 331450 111134
rect 331686 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 484250 111134
rect 484486 110898 514970 111134
rect 515206 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 592650 111134
rect -8726 110866 592650 110898
rect -8726 101494 592650 101526
rect -8726 101258 -8694 101494
rect -8458 101258 -8374 101494
rect -8138 101258 27866 101494
rect 28102 101258 28186 101494
rect 28422 101258 387866 101494
rect 388102 101258 388186 101494
rect 388422 101258 423866 101494
rect 424102 101258 424186 101494
rect 424422 101258 459866 101494
rect 460102 101258 460186 101494
rect 460422 101258 567866 101494
rect 568102 101258 568186 101494
rect 568422 101258 592062 101494
rect 592298 101258 592382 101494
rect 592618 101258 592650 101494
rect -8726 101174 592650 101258
rect -8726 100938 -8694 101174
rect -8458 100938 -8374 101174
rect -8138 100938 27866 101174
rect 28102 100938 28186 101174
rect 28422 100938 387866 101174
rect 388102 100938 388186 101174
rect 388422 100938 423866 101174
rect 424102 100938 424186 101174
rect 424422 100938 459866 101174
rect 460102 100938 460186 101174
rect 460422 100938 567866 101174
rect 568102 100938 568186 101174
rect 568422 100938 592062 101174
rect 592298 100938 592382 101174
rect 592618 100938 592650 101174
rect -8726 100906 592650 100938
rect -8726 97774 592650 97806
rect -8726 97538 -7734 97774
rect -7498 97538 -7414 97774
rect -7178 97538 384146 97774
rect 384382 97538 384466 97774
rect 384702 97538 420146 97774
rect 420382 97538 420466 97774
rect 420702 97538 456146 97774
rect 456382 97538 456466 97774
rect 456702 97538 564146 97774
rect 564382 97538 564466 97774
rect 564702 97538 591102 97774
rect 591338 97538 591422 97774
rect 591658 97538 592650 97774
rect -8726 97454 592650 97538
rect -8726 97218 -7734 97454
rect -7498 97218 -7414 97454
rect -7178 97218 384146 97454
rect 384382 97218 384466 97454
rect 384702 97218 420146 97454
rect 420382 97218 420466 97454
rect 420702 97218 456146 97454
rect 456382 97218 456466 97454
rect 456702 97218 564146 97454
rect 564382 97218 564466 97454
rect 564702 97218 591102 97454
rect 591338 97218 591422 97454
rect 591658 97218 592650 97454
rect -8726 97186 592650 97218
rect -8726 94054 592650 94086
rect -8726 93818 -6774 94054
rect -6538 93818 -6454 94054
rect -6218 93818 20426 94054
rect 20662 93818 20746 94054
rect 20982 93818 380426 94054
rect 380662 93818 380746 94054
rect 380982 93818 416426 94054
rect 416662 93818 416746 94054
rect 416982 93818 452426 94054
rect 452662 93818 452746 94054
rect 452982 93818 560426 94054
rect 560662 93818 560746 94054
rect 560982 93818 590142 94054
rect 590378 93818 590462 94054
rect 590698 93818 592650 94054
rect -8726 93734 592650 93818
rect -8726 93498 -6774 93734
rect -6538 93498 -6454 93734
rect -6218 93498 20426 93734
rect 20662 93498 20746 93734
rect 20982 93498 380426 93734
rect 380662 93498 380746 93734
rect 380982 93498 416426 93734
rect 416662 93498 416746 93734
rect 416982 93498 452426 93734
rect 452662 93498 452746 93734
rect 452982 93498 560426 93734
rect 560662 93498 560746 93734
rect 560982 93498 590142 93734
rect 590378 93498 590462 93734
rect 590698 93498 592650 93734
rect -8726 93466 592650 93498
rect -8726 90334 592650 90366
rect -8726 90098 -5814 90334
rect -5578 90098 -5494 90334
rect -5258 90098 16706 90334
rect 16942 90098 17026 90334
rect 17262 90098 376706 90334
rect 376942 90098 377026 90334
rect 377262 90098 484706 90334
rect 484942 90098 485026 90334
rect 485262 90098 556706 90334
rect 556942 90098 557026 90334
rect 557262 90098 589182 90334
rect 589418 90098 589502 90334
rect 589738 90098 592650 90334
rect -8726 90014 592650 90098
rect -8726 89778 -5814 90014
rect -5578 89778 -5494 90014
rect -5258 89778 16706 90014
rect 16942 89778 17026 90014
rect 17262 89778 376706 90014
rect 376942 89778 377026 90014
rect 377262 89778 484706 90014
rect 484942 89778 485026 90014
rect 485262 89778 556706 90014
rect 556942 89778 557026 90014
rect 557262 89778 589182 90014
rect 589418 89778 589502 90014
rect 589738 89778 592650 90014
rect -8726 89746 592650 89778
rect -8726 86614 592650 86646
rect -8726 86378 -4854 86614
rect -4618 86378 -4534 86614
rect -4298 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 372986 86614
rect 373222 86378 373306 86614
rect 373542 86378 480986 86614
rect 481222 86378 481306 86614
rect 481542 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 588222 86614
rect 588458 86378 588542 86614
rect 588778 86378 592650 86614
rect -8726 86294 592650 86378
rect -8726 86058 -4854 86294
rect -4618 86058 -4534 86294
rect -4298 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 372986 86294
rect 373222 86058 373306 86294
rect 373542 86058 480986 86294
rect 481222 86058 481306 86294
rect 481542 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 588222 86294
rect 588458 86058 588542 86294
rect 588778 86058 592650 86294
rect -8726 86026 592650 86058
rect -8726 82894 592650 82926
rect -8726 82658 -3894 82894
rect -3658 82658 -3574 82894
rect -3338 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 369266 82894
rect 369502 82658 369586 82894
rect 369822 82658 477266 82894
rect 477502 82658 477586 82894
rect 477822 82658 549266 82894
rect 549502 82658 549586 82894
rect 549822 82658 587262 82894
rect 587498 82658 587582 82894
rect 587818 82658 592650 82894
rect -8726 82574 592650 82658
rect -8726 82338 -3894 82574
rect -3658 82338 -3574 82574
rect -3338 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 369266 82574
rect 369502 82338 369586 82574
rect 369822 82338 477266 82574
rect 477502 82338 477586 82574
rect 477822 82338 549266 82574
rect 549502 82338 549586 82574
rect 549822 82338 587262 82574
rect 587498 82338 587582 82574
rect 587818 82338 592650 82574
rect -8726 82306 592650 82338
rect -8726 79174 592650 79206
rect -8726 78938 -2934 79174
rect -2698 78938 -2614 79174
rect -2378 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 39610 79174
rect 39846 78938 70330 79174
rect 70566 78938 101050 79174
rect 101286 78938 131770 79174
rect 132006 78938 162490 79174
rect 162726 78938 193210 79174
rect 193446 78938 223930 79174
rect 224166 78938 254650 79174
rect 254886 78938 285370 79174
rect 285606 78938 316090 79174
rect 316326 78938 346810 79174
rect 347046 78938 365546 79174
rect 365782 78938 365866 79174
rect 366102 78938 405610 79174
rect 405846 78938 436330 79174
rect 436566 78938 473546 79174
rect 473782 78938 473866 79174
rect 474102 78938 509546 79174
rect 509782 78938 509866 79174
rect 510102 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 586302 79174
rect 586538 78938 586622 79174
rect 586858 78938 592650 79174
rect -8726 78854 592650 78938
rect -8726 78618 -2934 78854
rect -2698 78618 -2614 78854
rect -2378 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 39610 78854
rect 39846 78618 70330 78854
rect 70566 78618 101050 78854
rect 101286 78618 131770 78854
rect 132006 78618 162490 78854
rect 162726 78618 193210 78854
rect 193446 78618 223930 78854
rect 224166 78618 254650 78854
rect 254886 78618 285370 78854
rect 285606 78618 316090 78854
rect 316326 78618 346810 78854
rect 347046 78618 365546 78854
rect 365782 78618 365866 78854
rect 366102 78618 405610 78854
rect 405846 78618 436330 78854
rect 436566 78618 473546 78854
rect 473782 78618 473866 78854
rect 474102 78618 509546 78854
rect 509782 78618 509866 78854
rect 510102 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 586302 78854
rect 586538 78618 586622 78854
rect 586858 78618 592650 78854
rect -8726 78586 592650 78618
rect -8726 75454 592650 75486
rect -8726 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 24250 75454
rect 24486 75218 54970 75454
rect 55206 75218 85690 75454
rect 85926 75218 116410 75454
rect 116646 75218 147130 75454
rect 147366 75218 177850 75454
rect 178086 75218 208570 75454
rect 208806 75218 239290 75454
rect 239526 75218 270010 75454
rect 270246 75218 300730 75454
rect 300966 75218 331450 75454
rect 331686 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 390250 75454
rect 390486 75218 420970 75454
rect 421206 75218 451690 75454
rect 451926 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 592650 75454
rect -8726 75134 592650 75218
rect -8726 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 24250 75134
rect 24486 74898 54970 75134
rect 55206 74898 85690 75134
rect 85926 74898 116410 75134
rect 116646 74898 147130 75134
rect 147366 74898 177850 75134
rect 178086 74898 208570 75134
rect 208806 74898 239290 75134
rect 239526 74898 270010 75134
rect 270246 74898 300730 75134
rect 300966 74898 331450 75134
rect 331686 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 390250 75134
rect 390486 74898 420970 75134
rect 421206 74898 451690 75134
rect 451926 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 592650 75134
rect -8726 74866 592650 74898
rect -8726 65494 592650 65526
rect -8726 65258 -8694 65494
rect -8458 65258 -8374 65494
rect -8138 65258 27866 65494
rect 28102 65258 28186 65494
rect 28422 65258 459866 65494
rect 460102 65258 460186 65494
rect 460422 65258 495866 65494
rect 496102 65258 496186 65494
rect 496422 65258 531866 65494
rect 532102 65258 532186 65494
rect 532422 65258 567866 65494
rect 568102 65258 568186 65494
rect 568422 65258 592062 65494
rect 592298 65258 592382 65494
rect 592618 65258 592650 65494
rect -8726 65174 592650 65258
rect -8726 64938 -8694 65174
rect -8458 64938 -8374 65174
rect -8138 64938 27866 65174
rect 28102 64938 28186 65174
rect 28422 64938 459866 65174
rect 460102 64938 460186 65174
rect 460422 64938 495866 65174
rect 496102 64938 496186 65174
rect 496422 64938 531866 65174
rect 532102 64938 532186 65174
rect 532422 64938 567866 65174
rect 568102 64938 568186 65174
rect 568422 64938 592062 65174
rect 592298 64938 592382 65174
rect 592618 64938 592650 65174
rect -8726 64906 592650 64938
rect -8726 61774 592650 61806
rect -8726 61538 -7734 61774
rect -7498 61538 -7414 61774
rect -7178 61538 384146 61774
rect 384382 61538 384466 61774
rect 384702 61538 492146 61774
rect 492382 61538 492466 61774
rect 492702 61538 528146 61774
rect 528382 61538 528466 61774
rect 528702 61538 564146 61774
rect 564382 61538 564466 61774
rect 564702 61538 591102 61774
rect 591338 61538 591422 61774
rect 591658 61538 592650 61774
rect -8726 61454 592650 61538
rect -8726 61218 -7734 61454
rect -7498 61218 -7414 61454
rect -7178 61218 384146 61454
rect 384382 61218 384466 61454
rect 384702 61218 492146 61454
rect 492382 61218 492466 61454
rect 492702 61218 528146 61454
rect 528382 61218 528466 61454
rect 528702 61218 564146 61454
rect 564382 61218 564466 61454
rect 564702 61218 591102 61454
rect 591338 61218 591422 61454
rect 591658 61218 592650 61454
rect -8726 61186 592650 61218
rect -8726 58054 592650 58086
rect -8726 57818 -6774 58054
rect -6538 57818 -6454 58054
rect -6218 57818 20426 58054
rect 20662 57818 20746 58054
rect 20982 57818 380426 58054
rect 380662 57818 380746 58054
rect 380982 57818 488426 58054
rect 488662 57818 488746 58054
rect 488982 57818 524426 58054
rect 524662 57818 524746 58054
rect 524982 57818 560426 58054
rect 560662 57818 560746 58054
rect 560982 57818 590142 58054
rect 590378 57818 590462 58054
rect 590698 57818 592650 58054
rect -8726 57734 592650 57818
rect -8726 57498 -6774 57734
rect -6538 57498 -6454 57734
rect -6218 57498 20426 57734
rect 20662 57498 20746 57734
rect 20982 57498 380426 57734
rect 380662 57498 380746 57734
rect 380982 57498 488426 57734
rect 488662 57498 488746 57734
rect 488982 57498 524426 57734
rect 524662 57498 524746 57734
rect 524982 57498 560426 57734
rect 560662 57498 560746 57734
rect 560982 57498 590142 57734
rect 590378 57498 590462 57734
rect 590698 57498 592650 57734
rect -8726 57466 592650 57498
rect -8726 54334 592650 54366
rect -8726 54098 -5814 54334
rect -5578 54098 -5494 54334
rect -5258 54098 16706 54334
rect 16942 54098 17026 54334
rect 17262 54098 376706 54334
rect 376942 54098 377026 54334
rect 377262 54098 484706 54334
rect 484942 54098 485026 54334
rect 485262 54098 520706 54334
rect 520942 54098 521026 54334
rect 521262 54098 556706 54334
rect 556942 54098 557026 54334
rect 557262 54098 589182 54334
rect 589418 54098 589502 54334
rect 589738 54098 592650 54334
rect -8726 54014 592650 54098
rect -8726 53778 -5814 54014
rect -5578 53778 -5494 54014
rect -5258 53778 16706 54014
rect 16942 53778 17026 54014
rect 17262 53778 376706 54014
rect 376942 53778 377026 54014
rect 377262 53778 484706 54014
rect 484942 53778 485026 54014
rect 485262 53778 520706 54014
rect 520942 53778 521026 54014
rect 521262 53778 556706 54014
rect 556942 53778 557026 54014
rect 557262 53778 589182 54014
rect 589418 53778 589502 54014
rect 589738 53778 592650 54014
rect -8726 53746 592650 53778
rect -8726 50614 592650 50646
rect -8726 50378 -4854 50614
rect -4618 50378 -4534 50614
rect -4298 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 372986 50614
rect 373222 50378 373306 50614
rect 373542 50378 480986 50614
rect 481222 50378 481306 50614
rect 481542 50378 516986 50614
rect 517222 50378 517306 50614
rect 517542 50378 588222 50614
rect 588458 50378 588542 50614
rect 588778 50378 592650 50614
rect -8726 50294 592650 50378
rect -8726 50058 -4854 50294
rect -4618 50058 -4534 50294
rect -4298 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 372986 50294
rect 373222 50058 373306 50294
rect 373542 50058 480986 50294
rect 481222 50058 481306 50294
rect 481542 50058 516986 50294
rect 517222 50058 517306 50294
rect 517542 50058 588222 50294
rect 588458 50058 588542 50294
rect 588778 50058 592650 50294
rect -8726 50026 592650 50058
rect -8726 46894 592650 46926
rect -8726 46658 -3894 46894
rect -3658 46658 -3574 46894
rect -3338 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 45266 46894
rect 45502 46658 45586 46894
rect 45822 46658 81266 46894
rect 81502 46658 81586 46894
rect 81822 46658 117266 46894
rect 117502 46658 117586 46894
rect 117822 46658 153266 46894
rect 153502 46658 153586 46894
rect 153822 46658 189266 46894
rect 189502 46658 189586 46894
rect 189822 46658 225266 46894
rect 225502 46658 225586 46894
rect 225822 46658 261266 46894
rect 261502 46658 261586 46894
rect 261822 46658 297266 46894
rect 297502 46658 297586 46894
rect 297822 46658 333266 46894
rect 333502 46658 333586 46894
rect 333822 46658 369266 46894
rect 369502 46658 369586 46894
rect 369822 46658 477266 46894
rect 477502 46658 477586 46894
rect 477822 46658 513266 46894
rect 513502 46658 513586 46894
rect 513822 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 587262 46894
rect 587498 46658 587582 46894
rect 587818 46658 592650 46894
rect -8726 46574 592650 46658
rect -8726 46338 -3894 46574
rect -3658 46338 -3574 46574
rect -3338 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 45266 46574
rect 45502 46338 45586 46574
rect 45822 46338 81266 46574
rect 81502 46338 81586 46574
rect 81822 46338 117266 46574
rect 117502 46338 117586 46574
rect 117822 46338 153266 46574
rect 153502 46338 153586 46574
rect 153822 46338 189266 46574
rect 189502 46338 189586 46574
rect 189822 46338 225266 46574
rect 225502 46338 225586 46574
rect 225822 46338 261266 46574
rect 261502 46338 261586 46574
rect 261822 46338 297266 46574
rect 297502 46338 297586 46574
rect 297822 46338 333266 46574
rect 333502 46338 333586 46574
rect 333822 46338 369266 46574
rect 369502 46338 369586 46574
rect 369822 46338 477266 46574
rect 477502 46338 477586 46574
rect 477822 46338 513266 46574
rect 513502 46338 513586 46574
rect 513822 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 587262 46574
rect 587498 46338 587582 46574
rect 587818 46338 592650 46574
rect -8726 46306 592650 46338
rect -8726 43174 592650 43206
rect -8726 42938 -2934 43174
rect -2698 42938 -2614 43174
rect -2378 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 77546 43174
rect 77782 42938 77866 43174
rect 78102 42938 113546 43174
rect 113782 42938 113866 43174
rect 114102 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 221546 43174
rect 221782 42938 221866 43174
rect 222102 42938 257546 43174
rect 257782 42938 257866 43174
rect 258102 42938 293546 43174
rect 293782 42938 293866 43174
rect 294102 42938 329546 43174
rect 329782 42938 329866 43174
rect 330102 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 405610 43174
rect 405846 42938 436330 43174
rect 436566 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 545930 43174
rect 546166 42938 550875 43174
rect 551111 42938 555820 43174
rect 556056 42938 560765 43174
rect 561001 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 586302 43174
rect 586538 42938 586622 43174
rect 586858 42938 592650 43174
rect -8726 42854 592650 42938
rect -8726 42618 -2934 42854
rect -2698 42618 -2614 42854
rect -2378 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 77546 42854
rect 77782 42618 77866 42854
rect 78102 42618 113546 42854
rect 113782 42618 113866 42854
rect 114102 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 221546 42854
rect 221782 42618 221866 42854
rect 222102 42618 257546 42854
rect 257782 42618 257866 42854
rect 258102 42618 293546 42854
rect 293782 42618 293866 42854
rect 294102 42618 329546 42854
rect 329782 42618 329866 42854
rect 330102 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 405610 42854
rect 405846 42618 436330 42854
rect 436566 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 545930 42854
rect 546166 42618 550875 42854
rect 551111 42618 555820 42854
rect 556056 42618 560765 42854
rect 561001 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 586302 42854
rect 586538 42618 586622 42854
rect 586858 42618 592650 42854
rect -8726 42586 592650 42618
rect -8726 39454 592650 39486
rect -8726 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 390250 39454
rect 390486 39218 420970 39454
rect 421206 39218 451690 39454
rect 451926 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 543458 39454
rect 543694 39218 548403 39454
rect 548639 39218 553348 39454
rect 553584 39218 558293 39454
rect 558529 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 592650 39454
rect -8726 39134 592650 39218
rect -8726 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 390250 39134
rect 390486 38898 420970 39134
rect 421206 38898 451690 39134
rect 451926 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 543458 39134
rect 543694 38898 548403 39134
rect 548639 38898 553348 39134
rect 553584 38898 558293 39134
rect 558529 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 592650 39134
rect -8726 38866 592650 38898
rect -8726 29494 592650 29526
rect -8726 29258 -8694 29494
rect -8458 29258 -8374 29494
rect -8138 29258 27866 29494
rect 28102 29258 28186 29494
rect 28422 29258 63866 29494
rect 64102 29258 64186 29494
rect 64422 29258 99866 29494
rect 100102 29258 100186 29494
rect 100422 29258 135866 29494
rect 136102 29258 136186 29494
rect 136422 29258 171866 29494
rect 172102 29258 172186 29494
rect 172422 29258 207866 29494
rect 208102 29258 208186 29494
rect 208422 29258 243866 29494
rect 244102 29258 244186 29494
rect 244422 29258 279866 29494
rect 280102 29258 280186 29494
rect 280422 29258 315866 29494
rect 316102 29258 316186 29494
rect 316422 29258 351866 29494
rect 352102 29258 352186 29494
rect 352422 29258 387866 29494
rect 388102 29258 388186 29494
rect 388422 29258 423866 29494
rect 424102 29258 424186 29494
rect 424422 29258 459866 29494
rect 460102 29258 460186 29494
rect 460422 29258 495866 29494
rect 496102 29258 496186 29494
rect 496422 29258 531866 29494
rect 532102 29258 532186 29494
rect 532422 29258 567866 29494
rect 568102 29258 568186 29494
rect 568422 29258 592062 29494
rect 592298 29258 592382 29494
rect 592618 29258 592650 29494
rect -8726 29174 592650 29258
rect -8726 28938 -8694 29174
rect -8458 28938 -8374 29174
rect -8138 28938 27866 29174
rect 28102 28938 28186 29174
rect 28422 28938 63866 29174
rect 64102 28938 64186 29174
rect 64422 28938 99866 29174
rect 100102 28938 100186 29174
rect 100422 28938 135866 29174
rect 136102 28938 136186 29174
rect 136422 28938 171866 29174
rect 172102 28938 172186 29174
rect 172422 28938 207866 29174
rect 208102 28938 208186 29174
rect 208422 28938 243866 29174
rect 244102 28938 244186 29174
rect 244422 28938 279866 29174
rect 280102 28938 280186 29174
rect 280422 28938 315866 29174
rect 316102 28938 316186 29174
rect 316422 28938 351866 29174
rect 352102 28938 352186 29174
rect 352422 28938 387866 29174
rect 388102 28938 388186 29174
rect 388422 28938 423866 29174
rect 424102 28938 424186 29174
rect 424422 28938 459866 29174
rect 460102 28938 460186 29174
rect 460422 28938 495866 29174
rect 496102 28938 496186 29174
rect 496422 28938 531866 29174
rect 532102 28938 532186 29174
rect 532422 28938 567866 29174
rect 568102 28938 568186 29174
rect 568422 28938 592062 29174
rect 592298 28938 592382 29174
rect 592618 28938 592650 29174
rect -8726 28906 592650 28938
rect -8726 25774 592650 25806
rect -8726 25538 -7734 25774
rect -7498 25538 -7414 25774
rect -7178 25538 24146 25774
rect 24382 25538 24466 25774
rect 24702 25538 60146 25774
rect 60382 25538 60466 25774
rect 60702 25538 96146 25774
rect 96382 25538 96466 25774
rect 96702 25538 132146 25774
rect 132382 25538 132466 25774
rect 132702 25538 168146 25774
rect 168382 25538 168466 25774
rect 168702 25538 204146 25774
rect 204382 25538 204466 25774
rect 204702 25538 240146 25774
rect 240382 25538 240466 25774
rect 240702 25538 276146 25774
rect 276382 25538 276466 25774
rect 276702 25538 312146 25774
rect 312382 25538 312466 25774
rect 312702 25538 348146 25774
rect 348382 25538 348466 25774
rect 348702 25538 384146 25774
rect 384382 25538 384466 25774
rect 384702 25538 420146 25774
rect 420382 25538 420466 25774
rect 420702 25538 456146 25774
rect 456382 25538 456466 25774
rect 456702 25538 492146 25774
rect 492382 25538 492466 25774
rect 492702 25538 528146 25774
rect 528382 25538 528466 25774
rect 528702 25538 564146 25774
rect 564382 25538 564466 25774
rect 564702 25538 591102 25774
rect 591338 25538 591422 25774
rect 591658 25538 592650 25774
rect -8726 25454 592650 25538
rect -8726 25218 -7734 25454
rect -7498 25218 -7414 25454
rect -7178 25218 24146 25454
rect 24382 25218 24466 25454
rect 24702 25218 60146 25454
rect 60382 25218 60466 25454
rect 60702 25218 96146 25454
rect 96382 25218 96466 25454
rect 96702 25218 132146 25454
rect 132382 25218 132466 25454
rect 132702 25218 168146 25454
rect 168382 25218 168466 25454
rect 168702 25218 204146 25454
rect 204382 25218 204466 25454
rect 204702 25218 240146 25454
rect 240382 25218 240466 25454
rect 240702 25218 276146 25454
rect 276382 25218 276466 25454
rect 276702 25218 312146 25454
rect 312382 25218 312466 25454
rect 312702 25218 348146 25454
rect 348382 25218 348466 25454
rect 348702 25218 384146 25454
rect 384382 25218 384466 25454
rect 384702 25218 420146 25454
rect 420382 25218 420466 25454
rect 420702 25218 456146 25454
rect 456382 25218 456466 25454
rect 456702 25218 492146 25454
rect 492382 25218 492466 25454
rect 492702 25218 528146 25454
rect 528382 25218 528466 25454
rect 528702 25218 564146 25454
rect 564382 25218 564466 25454
rect 564702 25218 591102 25454
rect 591338 25218 591422 25454
rect 591658 25218 592650 25454
rect -8726 25186 592650 25218
rect -8726 22054 592650 22086
rect -8726 21818 -6774 22054
rect -6538 21818 -6454 22054
rect -6218 21818 20426 22054
rect 20662 21818 20746 22054
rect 20982 21818 56426 22054
rect 56662 21818 56746 22054
rect 56982 21818 92426 22054
rect 92662 21818 92746 22054
rect 92982 21818 128426 22054
rect 128662 21818 128746 22054
rect 128982 21818 164426 22054
rect 164662 21818 164746 22054
rect 164982 21818 200426 22054
rect 200662 21818 200746 22054
rect 200982 21818 236426 22054
rect 236662 21818 236746 22054
rect 236982 21818 272426 22054
rect 272662 21818 272746 22054
rect 272982 21818 308426 22054
rect 308662 21818 308746 22054
rect 308982 21818 344426 22054
rect 344662 21818 344746 22054
rect 344982 21818 380426 22054
rect 380662 21818 380746 22054
rect 380982 21818 416426 22054
rect 416662 21818 416746 22054
rect 416982 21818 452426 22054
rect 452662 21818 452746 22054
rect 452982 21818 488426 22054
rect 488662 21818 488746 22054
rect 488982 21818 524426 22054
rect 524662 21818 524746 22054
rect 524982 21818 560426 22054
rect 560662 21818 560746 22054
rect 560982 21818 590142 22054
rect 590378 21818 590462 22054
rect 590698 21818 592650 22054
rect -8726 21734 592650 21818
rect -8726 21498 -6774 21734
rect -6538 21498 -6454 21734
rect -6218 21498 20426 21734
rect 20662 21498 20746 21734
rect 20982 21498 56426 21734
rect 56662 21498 56746 21734
rect 56982 21498 92426 21734
rect 92662 21498 92746 21734
rect 92982 21498 128426 21734
rect 128662 21498 128746 21734
rect 128982 21498 164426 21734
rect 164662 21498 164746 21734
rect 164982 21498 200426 21734
rect 200662 21498 200746 21734
rect 200982 21498 236426 21734
rect 236662 21498 236746 21734
rect 236982 21498 272426 21734
rect 272662 21498 272746 21734
rect 272982 21498 308426 21734
rect 308662 21498 308746 21734
rect 308982 21498 344426 21734
rect 344662 21498 344746 21734
rect 344982 21498 380426 21734
rect 380662 21498 380746 21734
rect 380982 21498 416426 21734
rect 416662 21498 416746 21734
rect 416982 21498 452426 21734
rect 452662 21498 452746 21734
rect 452982 21498 488426 21734
rect 488662 21498 488746 21734
rect 488982 21498 524426 21734
rect 524662 21498 524746 21734
rect 524982 21498 560426 21734
rect 560662 21498 560746 21734
rect 560982 21498 590142 21734
rect 590378 21498 590462 21734
rect 590698 21498 592650 21734
rect -8726 21466 592650 21498
rect -8726 18334 592650 18366
rect -8726 18098 -5814 18334
rect -5578 18098 -5494 18334
rect -5258 18098 16706 18334
rect 16942 18098 17026 18334
rect 17262 18098 52706 18334
rect 52942 18098 53026 18334
rect 53262 18098 88706 18334
rect 88942 18098 89026 18334
rect 89262 18098 124706 18334
rect 124942 18098 125026 18334
rect 125262 18098 160706 18334
rect 160942 18098 161026 18334
rect 161262 18098 196706 18334
rect 196942 18098 197026 18334
rect 197262 18098 232706 18334
rect 232942 18098 233026 18334
rect 233262 18098 268706 18334
rect 268942 18098 269026 18334
rect 269262 18098 304706 18334
rect 304942 18098 305026 18334
rect 305262 18098 340706 18334
rect 340942 18098 341026 18334
rect 341262 18098 376706 18334
rect 376942 18098 377026 18334
rect 377262 18098 412706 18334
rect 412942 18098 413026 18334
rect 413262 18098 448706 18334
rect 448942 18098 449026 18334
rect 449262 18098 484706 18334
rect 484942 18098 485026 18334
rect 485262 18098 520706 18334
rect 520942 18098 521026 18334
rect 521262 18098 556706 18334
rect 556942 18098 557026 18334
rect 557262 18098 589182 18334
rect 589418 18098 589502 18334
rect 589738 18098 592650 18334
rect -8726 18014 592650 18098
rect -8726 17778 -5814 18014
rect -5578 17778 -5494 18014
rect -5258 17778 16706 18014
rect 16942 17778 17026 18014
rect 17262 17778 52706 18014
rect 52942 17778 53026 18014
rect 53262 17778 88706 18014
rect 88942 17778 89026 18014
rect 89262 17778 124706 18014
rect 124942 17778 125026 18014
rect 125262 17778 160706 18014
rect 160942 17778 161026 18014
rect 161262 17778 196706 18014
rect 196942 17778 197026 18014
rect 197262 17778 232706 18014
rect 232942 17778 233026 18014
rect 233262 17778 268706 18014
rect 268942 17778 269026 18014
rect 269262 17778 304706 18014
rect 304942 17778 305026 18014
rect 305262 17778 340706 18014
rect 340942 17778 341026 18014
rect 341262 17778 376706 18014
rect 376942 17778 377026 18014
rect 377262 17778 412706 18014
rect 412942 17778 413026 18014
rect 413262 17778 448706 18014
rect 448942 17778 449026 18014
rect 449262 17778 484706 18014
rect 484942 17778 485026 18014
rect 485262 17778 520706 18014
rect 520942 17778 521026 18014
rect 521262 17778 556706 18014
rect 556942 17778 557026 18014
rect 557262 17778 589182 18014
rect 589418 17778 589502 18014
rect 589738 17778 592650 18014
rect -8726 17746 592650 17778
rect -8726 14614 592650 14646
rect -8726 14378 -4854 14614
rect -4618 14378 -4534 14614
rect -4298 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 588222 14614
rect 588458 14378 588542 14614
rect 588778 14378 592650 14614
rect -8726 14294 592650 14378
rect -8726 14058 -4854 14294
rect -4618 14058 -4534 14294
rect -4298 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 588222 14294
rect 588458 14058 588542 14294
rect 588778 14058 592650 14294
rect -8726 14026 592650 14058
rect -8726 10894 592650 10926
rect -8726 10658 -3894 10894
rect -3658 10658 -3574 10894
rect -3338 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 587262 10894
rect 587498 10658 587582 10894
rect 587818 10658 592650 10894
rect -8726 10574 592650 10658
rect -8726 10338 -3894 10574
rect -3658 10338 -3574 10574
rect -3338 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 587262 10574
rect 587498 10338 587582 10574
rect 587818 10338 592650 10574
rect -8726 10306 592650 10338
rect -8726 7174 592650 7206
rect -8726 6938 -2934 7174
rect -2698 6938 -2614 7174
rect -2378 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 586302 7174
rect 586538 6938 586622 7174
rect 586858 6938 592650 7174
rect -8726 6854 592650 6938
rect -8726 6618 -2934 6854
rect -2698 6618 -2614 6854
rect -2378 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 586302 6854
rect 586538 6618 586622 6854
rect 586858 6618 592650 6854
rect -8726 6586 592650 6618
rect -8726 3454 592650 3486
rect -8726 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 592650 3454
rect -8726 3134 592650 3218
rect -8726 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 592650 3134
rect -8726 2866 592650 2898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 5546 -1306
rect 5782 -1542 5866 -1306
rect 6102 -1542 41546 -1306
rect 41782 -1542 41866 -1306
rect 42102 -1542 77546 -1306
rect 77782 -1542 77866 -1306
rect 78102 -1542 113546 -1306
rect 113782 -1542 113866 -1306
rect 114102 -1542 149546 -1306
rect 149782 -1542 149866 -1306
rect 150102 -1542 185546 -1306
rect 185782 -1542 185866 -1306
rect 186102 -1542 221546 -1306
rect 221782 -1542 221866 -1306
rect 222102 -1542 257546 -1306
rect 257782 -1542 257866 -1306
rect 258102 -1542 293546 -1306
rect 293782 -1542 293866 -1306
rect 294102 -1542 329546 -1306
rect 329782 -1542 329866 -1306
rect 330102 -1542 365546 -1306
rect 365782 -1542 365866 -1306
rect 366102 -1542 401546 -1306
rect 401782 -1542 401866 -1306
rect 402102 -1542 437546 -1306
rect 437782 -1542 437866 -1306
rect 438102 -1542 473546 -1306
rect 473782 -1542 473866 -1306
rect 474102 -1542 509546 -1306
rect 509782 -1542 509866 -1306
rect 510102 -1542 545546 -1306
rect 545782 -1542 545866 -1306
rect 546102 -1542 581546 -1306
rect 581782 -1542 581866 -1306
rect 582102 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 5546 -1626
rect 5782 -1862 5866 -1626
rect 6102 -1862 41546 -1626
rect 41782 -1862 41866 -1626
rect 42102 -1862 77546 -1626
rect 77782 -1862 77866 -1626
rect 78102 -1862 113546 -1626
rect 113782 -1862 113866 -1626
rect 114102 -1862 149546 -1626
rect 149782 -1862 149866 -1626
rect 150102 -1862 185546 -1626
rect 185782 -1862 185866 -1626
rect 186102 -1862 221546 -1626
rect 221782 -1862 221866 -1626
rect 222102 -1862 257546 -1626
rect 257782 -1862 257866 -1626
rect 258102 -1862 293546 -1626
rect 293782 -1862 293866 -1626
rect 294102 -1862 329546 -1626
rect 329782 -1862 329866 -1626
rect 330102 -1862 365546 -1626
rect 365782 -1862 365866 -1626
rect 366102 -1862 401546 -1626
rect 401782 -1862 401866 -1626
rect 402102 -1862 437546 -1626
rect 437782 -1862 437866 -1626
rect 438102 -1862 473546 -1626
rect 473782 -1862 473866 -1626
rect 474102 -1862 509546 -1626
rect 509782 -1862 509866 -1626
rect 510102 -1862 545546 -1626
rect 545782 -1862 545866 -1626
rect 546102 -1862 581546 -1626
rect 581782 -1862 581866 -1626
rect 582102 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 9266 -2266
rect 9502 -2502 9586 -2266
rect 9822 -2502 45266 -2266
rect 45502 -2502 45586 -2266
rect 45822 -2502 81266 -2266
rect 81502 -2502 81586 -2266
rect 81822 -2502 117266 -2266
rect 117502 -2502 117586 -2266
rect 117822 -2502 153266 -2266
rect 153502 -2502 153586 -2266
rect 153822 -2502 189266 -2266
rect 189502 -2502 189586 -2266
rect 189822 -2502 225266 -2266
rect 225502 -2502 225586 -2266
rect 225822 -2502 261266 -2266
rect 261502 -2502 261586 -2266
rect 261822 -2502 297266 -2266
rect 297502 -2502 297586 -2266
rect 297822 -2502 333266 -2266
rect 333502 -2502 333586 -2266
rect 333822 -2502 369266 -2266
rect 369502 -2502 369586 -2266
rect 369822 -2502 405266 -2266
rect 405502 -2502 405586 -2266
rect 405822 -2502 441266 -2266
rect 441502 -2502 441586 -2266
rect 441822 -2502 477266 -2266
rect 477502 -2502 477586 -2266
rect 477822 -2502 513266 -2266
rect 513502 -2502 513586 -2266
rect 513822 -2502 549266 -2266
rect 549502 -2502 549586 -2266
rect 549822 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 9266 -2586
rect 9502 -2822 9586 -2586
rect 9822 -2822 45266 -2586
rect 45502 -2822 45586 -2586
rect 45822 -2822 81266 -2586
rect 81502 -2822 81586 -2586
rect 81822 -2822 117266 -2586
rect 117502 -2822 117586 -2586
rect 117822 -2822 153266 -2586
rect 153502 -2822 153586 -2586
rect 153822 -2822 189266 -2586
rect 189502 -2822 189586 -2586
rect 189822 -2822 225266 -2586
rect 225502 -2822 225586 -2586
rect 225822 -2822 261266 -2586
rect 261502 -2822 261586 -2586
rect 261822 -2822 297266 -2586
rect 297502 -2822 297586 -2586
rect 297822 -2822 333266 -2586
rect 333502 -2822 333586 -2586
rect 333822 -2822 369266 -2586
rect 369502 -2822 369586 -2586
rect 369822 -2822 405266 -2586
rect 405502 -2822 405586 -2586
rect 405822 -2822 441266 -2586
rect 441502 -2822 441586 -2586
rect 441822 -2822 477266 -2586
rect 477502 -2822 477586 -2586
rect 477822 -2822 513266 -2586
rect 513502 -2822 513586 -2586
rect 513822 -2822 549266 -2586
rect 549502 -2822 549586 -2586
rect 549822 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 12986 -3226
rect 13222 -3462 13306 -3226
rect 13542 -3462 48986 -3226
rect 49222 -3462 49306 -3226
rect 49542 -3462 84986 -3226
rect 85222 -3462 85306 -3226
rect 85542 -3462 120986 -3226
rect 121222 -3462 121306 -3226
rect 121542 -3462 156986 -3226
rect 157222 -3462 157306 -3226
rect 157542 -3462 192986 -3226
rect 193222 -3462 193306 -3226
rect 193542 -3462 228986 -3226
rect 229222 -3462 229306 -3226
rect 229542 -3462 264986 -3226
rect 265222 -3462 265306 -3226
rect 265542 -3462 300986 -3226
rect 301222 -3462 301306 -3226
rect 301542 -3462 336986 -3226
rect 337222 -3462 337306 -3226
rect 337542 -3462 372986 -3226
rect 373222 -3462 373306 -3226
rect 373542 -3462 408986 -3226
rect 409222 -3462 409306 -3226
rect 409542 -3462 444986 -3226
rect 445222 -3462 445306 -3226
rect 445542 -3462 480986 -3226
rect 481222 -3462 481306 -3226
rect 481542 -3462 516986 -3226
rect 517222 -3462 517306 -3226
rect 517542 -3462 552986 -3226
rect 553222 -3462 553306 -3226
rect 553542 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 12986 -3546
rect 13222 -3782 13306 -3546
rect 13542 -3782 48986 -3546
rect 49222 -3782 49306 -3546
rect 49542 -3782 84986 -3546
rect 85222 -3782 85306 -3546
rect 85542 -3782 120986 -3546
rect 121222 -3782 121306 -3546
rect 121542 -3782 156986 -3546
rect 157222 -3782 157306 -3546
rect 157542 -3782 192986 -3546
rect 193222 -3782 193306 -3546
rect 193542 -3782 228986 -3546
rect 229222 -3782 229306 -3546
rect 229542 -3782 264986 -3546
rect 265222 -3782 265306 -3546
rect 265542 -3782 300986 -3546
rect 301222 -3782 301306 -3546
rect 301542 -3782 336986 -3546
rect 337222 -3782 337306 -3546
rect 337542 -3782 372986 -3546
rect 373222 -3782 373306 -3546
rect 373542 -3782 408986 -3546
rect 409222 -3782 409306 -3546
rect 409542 -3782 444986 -3546
rect 445222 -3782 445306 -3546
rect 445542 -3782 480986 -3546
rect 481222 -3782 481306 -3546
rect 481542 -3782 516986 -3546
rect 517222 -3782 517306 -3546
rect 517542 -3782 552986 -3546
rect 553222 -3782 553306 -3546
rect 553542 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 16706 -4186
rect 16942 -4422 17026 -4186
rect 17262 -4422 52706 -4186
rect 52942 -4422 53026 -4186
rect 53262 -4422 88706 -4186
rect 88942 -4422 89026 -4186
rect 89262 -4422 124706 -4186
rect 124942 -4422 125026 -4186
rect 125262 -4422 160706 -4186
rect 160942 -4422 161026 -4186
rect 161262 -4422 196706 -4186
rect 196942 -4422 197026 -4186
rect 197262 -4422 232706 -4186
rect 232942 -4422 233026 -4186
rect 233262 -4422 268706 -4186
rect 268942 -4422 269026 -4186
rect 269262 -4422 304706 -4186
rect 304942 -4422 305026 -4186
rect 305262 -4422 340706 -4186
rect 340942 -4422 341026 -4186
rect 341262 -4422 376706 -4186
rect 376942 -4422 377026 -4186
rect 377262 -4422 412706 -4186
rect 412942 -4422 413026 -4186
rect 413262 -4422 448706 -4186
rect 448942 -4422 449026 -4186
rect 449262 -4422 484706 -4186
rect 484942 -4422 485026 -4186
rect 485262 -4422 520706 -4186
rect 520942 -4422 521026 -4186
rect 521262 -4422 556706 -4186
rect 556942 -4422 557026 -4186
rect 557262 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 16706 -4506
rect 16942 -4742 17026 -4506
rect 17262 -4742 52706 -4506
rect 52942 -4742 53026 -4506
rect 53262 -4742 88706 -4506
rect 88942 -4742 89026 -4506
rect 89262 -4742 124706 -4506
rect 124942 -4742 125026 -4506
rect 125262 -4742 160706 -4506
rect 160942 -4742 161026 -4506
rect 161262 -4742 196706 -4506
rect 196942 -4742 197026 -4506
rect 197262 -4742 232706 -4506
rect 232942 -4742 233026 -4506
rect 233262 -4742 268706 -4506
rect 268942 -4742 269026 -4506
rect 269262 -4742 304706 -4506
rect 304942 -4742 305026 -4506
rect 305262 -4742 340706 -4506
rect 340942 -4742 341026 -4506
rect 341262 -4742 376706 -4506
rect 376942 -4742 377026 -4506
rect 377262 -4742 412706 -4506
rect 412942 -4742 413026 -4506
rect 413262 -4742 448706 -4506
rect 448942 -4742 449026 -4506
rect 449262 -4742 484706 -4506
rect 484942 -4742 485026 -4506
rect 485262 -4742 520706 -4506
rect 520942 -4742 521026 -4506
rect 521262 -4742 556706 -4506
rect 556942 -4742 557026 -4506
rect 557262 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 20426 -5146
rect 20662 -5382 20746 -5146
rect 20982 -5382 56426 -5146
rect 56662 -5382 56746 -5146
rect 56982 -5382 92426 -5146
rect 92662 -5382 92746 -5146
rect 92982 -5382 128426 -5146
rect 128662 -5382 128746 -5146
rect 128982 -5382 164426 -5146
rect 164662 -5382 164746 -5146
rect 164982 -5382 200426 -5146
rect 200662 -5382 200746 -5146
rect 200982 -5382 236426 -5146
rect 236662 -5382 236746 -5146
rect 236982 -5382 272426 -5146
rect 272662 -5382 272746 -5146
rect 272982 -5382 308426 -5146
rect 308662 -5382 308746 -5146
rect 308982 -5382 344426 -5146
rect 344662 -5382 344746 -5146
rect 344982 -5382 380426 -5146
rect 380662 -5382 380746 -5146
rect 380982 -5382 416426 -5146
rect 416662 -5382 416746 -5146
rect 416982 -5382 452426 -5146
rect 452662 -5382 452746 -5146
rect 452982 -5382 488426 -5146
rect 488662 -5382 488746 -5146
rect 488982 -5382 524426 -5146
rect 524662 -5382 524746 -5146
rect 524982 -5382 560426 -5146
rect 560662 -5382 560746 -5146
rect 560982 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 20426 -5466
rect 20662 -5702 20746 -5466
rect 20982 -5702 56426 -5466
rect 56662 -5702 56746 -5466
rect 56982 -5702 92426 -5466
rect 92662 -5702 92746 -5466
rect 92982 -5702 128426 -5466
rect 128662 -5702 128746 -5466
rect 128982 -5702 164426 -5466
rect 164662 -5702 164746 -5466
rect 164982 -5702 200426 -5466
rect 200662 -5702 200746 -5466
rect 200982 -5702 236426 -5466
rect 236662 -5702 236746 -5466
rect 236982 -5702 272426 -5466
rect 272662 -5702 272746 -5466
rect 272982 -5702 308426 -5466
rect 308662 -5702 308746 -5466
rect 308982 -5702 344426 -5466
rect 344662 -5702 344746 -5466
rect 344982 -5702 380426 -5466
rect 380662 -5702 380746 -5466
rect 380982 -5702 416426 -5466
rect 416662 -5702 416746 -5466
rect 416982 -5702 452426 -5466
rect 452662 -5702 452746 -5466
rect 452982 -5702 488426 -5466
rect 488662 -5702 488746 -5466
rect 488982 -5702 524426 -5466
rect 524662 -5702 524746 -5466
rect 524982 -5702 560426 -5466
rect 560662 -5702 560746 -5466
rect 560982 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 24146 -6106
rect 24382 -6342 24466 -6106
rect 24702 -6342 60146 -6106
rect 60382 -6342 60466 -6106
rect 60702 -6342 96146 -6106
rect 96382 -6342 96466 -6106
rect 96702 -6342 132146 -6106
rect 132382 -6342 132466 -6106
rect 132702 -6342 168146 -6106
rect 168382 -6342 168466 -6106
rect 168702 -6342 204146 -6106
rect 204382 -6342 204466 -6106
rect 204702 -6342 240146 -6106
rect 240382 -6342 240466 -6106
rect 240702 -6342 276146 -6106
rect 276382 -6342 276466 -6106
rect 276702 -6342 312146 -6106
rect 312382 -6342 312466 -6106
rect 312702 -6342 348146 -6106
rect 348382 -6342 348466 -6106
rect 348702 -6342 384146 -6106
rect 384382 -6342 384466 -6106
rect 384702 -6342 420146 -6106
rect 420382 -6342 420466 -6106
rect 420702 -6342 456146 -6106
rect 456382 -6342 456466 -6106
rect 456702 -6342 492146 -6106
rect 492382 -6342 492466 -6106
rect 492702 -6342 528146 -6106
rect 528382 -6342 528466 -6106
rect 528702 -6342 564146 -6106
rect 564382 -6342 564466 -6106
rect 564702 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 24146 -6426
rect 24382 -6662 24466 -6426
rect 24702 -6662 60146 -6426
rect 60382 -6662 60466 -6426
rect 60702 -6662 96146 -6426
rect 96382 -6662 96466 -6426
rect 96702 -6662 132146 -6426
rect 132382 -6662 132466 -6426
rect 132702 -6662 168146 -6426
rect 168382 -6662 168466 -6426
rect 168702 -6662 204146 -6426
rect 204382 -6662 204466 -6426
rect 204702 -6662 240146 -6426
rect 240382 -6662 240466 -6426
rect 240702 -6662 276146 -6426
rect 276382 -6662 276466 -6426
rect 276702 -6662 312146 -6426
rect 312382 -6662 312466 -6426
rect 312702 -6662 348146 -6426
rect 348382 -6662 348466 -6426
rect 348702 -6662 384146 -6426
rect 384382 -6662 384466 -6426
rect 384702 -6662 420146 -6426
rect 420382 -6662 420466 -6426
rect 420702 -6662 456146 -6426
rect 456382 -6662 456466 -6426
rect 456702 -6662 492146 -6426
rect 492382 -6662 492466 -6426
rect 492702 -6662 528146 -6426
rect 528382 -6662 528466 -6426
rect 528702 -6662 564146 -6426
rect 564382 -6662 564466 -6426
rect 564702 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 27866 -7066
rect 28102 -7302 28186 -7066
rect 28422 -7302 63866 -7066
rect 64102 -7302 64186 -7066
rect 64422 -7302 99866 -7066
rect 100102 -7302 100186 -7066
rect 100422 -7302 135866 -7066
rect 136102 -7302 136186 -7066
rect 136422 -7302 171866 -7066
rect 172102 -7302 172186 -7066
rect 172422 -7302 207866 -7066
rect 208102 -7302 208186 -7066
rect 208422 -7302 243866 -7066
rect 244102 -7302 244186 -7066
rect 244422 -7302 279866 -7066
rect 280102 -7302 280186 -7066
rect 280422 -7302 315866 -7066
rect 316102 -7302 316186 -7066
rect 316422 -7302 351866 -7066
rect 352102 -7302 352186 -7066
rect 352422 -7302 387866 -7066
rect 388102 -7302 388186 -7066
rect 388422 -7302 423866 -7066
rect 424102 -7302 424186 -7066
rect 424422 -7302 459866 -7066
rect 460102 -7302 460186 -7066
rect 460422 -7302 495866 -7066
rect 496102 -7302 496186 -7066
rect 496422 -7302 531866 -7066
rect 532102 -7302 532186 -7066
rect 532422 -7302 567866 -7066
rect 568102 -7302 568186 -7066
rect 568422 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 27866 -7386
rect 28102 -7622 28186 -7386
rect 28422 -7622 63866 -7386
rect 64102 -7622 64186 -7386
rect 64422 -7622 99866 -7386
rect 100102 -7622 100186 -7386
rect 100422 -7622 135866 -7386
rect 136102 -7622 136186 -7386
rect 136422 -7622 171866 -7386
rect 172102 -7622 172186 -7386
rect 172422 -7622 207866 -7386
rect 208102 -7622 208186 -7386
rect 208422 -7622 243866 -7386
rect 244102 -7622 244186 -7386
rect 244422 -7622 279866 -7386
rect 280102 -7622 280186 -7386
rect 280422 -7622 315866 -7386
rect 316102 -7622 316186 -7386
rect 316422 -7622 351866 -7386
rect 352102 -7622 352186 -7386
rect 352422 -7622 387866 -7386
rect 388102 -7622 388186 -7386
rect 388422 -7622 423866 -7386
rect 424102 -7622 424186 -7386
rect 424422 -7622 459866 -7386
rect 460102 -7622 460186 -7386
rect 460422 -7622 495866 -7386
rect 496102 -7622 496186 -7386
rect 496422 -7622 531866 -7386
rect 532102 -7622 532186 -7386
rect 532422 -7622 567866 -7386
rect 568102 -7622 568186 -7386
rect 568422 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use posit_unit  posit_unit
timestamp 0
transform 1 0 460000 0 1 200000
box 0 2128 70000 67504
use multiplexer  proj_multiplexer
timestamp 0
transform 1 0 450000 0 1 322000
box 0 0 60000 64000
use tholin_avalonsemi_5401  tholin_avalonsemi_5401
timestamp 0
transform 1 0 520000 0 1 425000
box 1066 0 36000 36000
use tholin_avalonsemi_tbb1143  tholin_avalonsemi_tbb1143
timestamp 0
transform 1 0 400000 0 1 305000
box 1066 2048 30000 30000
use tt2_tholin_diceroll  tt2_tholin_diceroll
timestamp 0
transform 1 0 470000 0 1 432000
box 1066 0 21043 22000
use tt2_tholin_multiplexed_counter  tt2_tholin_multiplexed_counter
timestamp 0
transform 1 0 550000 0 1 360000
box 842 0 17098 18000
use tt2_tholin_multiplier  tt2_tholin_multiplier
timestamp 0
transform 1 0 450000 0 1 500000
box 0 0 11118 16584
use tt2_tholin_namebadge  tt2_tholin_namebadge
timestamp 0
transform 1 0 420000 0 1 420000
box 1066 0 23987 25000
use tune_player  tune_player
timestamp 0
transform 1 0 540000 0 1 30000
box 0 2128 21043 19632
use wrapped_6502  wrapped_6502
timestamp 0
transform 1 0 410000 0 1 120000
box 1066 1504 40000 40000
use wrapped_MC14500  wrapped_MC14500
timestamp 0
transform 1 0 480000 0 1 500000
box 566 0 12000 18000
use wrapped_as1802  wrapped_as1802
timestamp 0
transform 1 0 480000 0 1 80000
box 1066 2128 60000 60000
use wrapped_as2650  wrapped_as2650
timestamp 0
transform 1 0 460000 0 1 600000
box 0 0 68816 67992
use wrapped_as512512512  wrapped_as512512512
timestamp 0
transform 1 0 20000 0 1 45000
box 1066 2128 340000 637616
use wrapped_vgatest  wrapped_vgatest
timestamp 0
transform 1 0 386000 0 1 30000
box 749 2128 75000 75000
<< labels >>
flabel metal3 s 583520 285276 584960 285516 0 FreeSans 960 0 0 0 analog_io[0]
port 0 nsew signal bidirectional
flabel metal2 s 446098 703520 446210 704960 0 FreeSans 448 90 0 0 analog_io[10]
port 1 nsew signal bidirectional
flabel metal2 s 381146 703520 381258 704960 0 FreeSans 448 90 0 0 analog_io[11]
port 2 nsew signal bidirectional
flabel metal2 s 316286 703520 316398 704960 0 FreeSans 448 90 0 0 analog_io[12]
port 3 nsew signal bidirectional
flabel metal2 s 251426 703520 251538 704960 0 FreeSans 448 90 0 0 analog_io[13]
port 4 nsew signal bidirectional
flabel metal2 s 186474 703520 186586 704960 0 FreeSans 448 90 0 0 analog_io[14]
port 5 nsew signal bidirectional
flabel metal2 s 121614 703520 121726 704960 0 FreeSans 448 90 0 0 analog_io[15]
port 6 nsew signal bidirectional
flabel metal2 s 56754 703520 56866 704960 0 FreeSans 448 90 0 0 analog_io[16]
port 7 nsew signal bidirectional
flabel metal3 s -960 697220 480 697460 0 FreeSans 960 0 0 0 analog_io[17]
port 8 nsew signal bidirectional
flabel metal3 s -960 644996 480 645236 0 FreeSans 960 0 0 0 analog_io[18]
port 9 nsew signal bidirectional
flabel metal3 s -960 592908 480 593148 0 FreeSans 960 0 0 0 analog_io[19]
port 10 nsew signal bidirectional
flabel metal3 s 583520 338452 584960 338692 0 FreeSans 960 0 0 0 analog_io[1]
port 11 nsew signal bidirectional
flabel metal3 s -960 540684 480 540924 0 FreeSans 960 0 0 0 analog_io[20]
port 12 nsew signal bidirectional
flabel metal3 s -960 488596 480 488836 0 FreeSans 960 0 0 0 analog_io[21]
port 13 nsew signal bidirectional
flabel metal3 s -960 436508 480 436748 0 FreeSans 960 0 0 0 analog_io[22]
port 14 nsew signal bidirectional
flabel metal3 s -960 384284 480 384524 0 FreeSans 960 0 0 0 analog_io[23]
port 15 nsew signal bidirectional
flabel metal3 s -960 332196 480 332436 0 FreeSans 960 0 0 0 analog_io[24]
port 16 nsew signal bidirectional
flabel metal3 s -960 279972 480 280212 0 FreeSans 960 0 0 0 analog_io[25]
port 17 nsew signal bidirectional
flabel metal3 s -960 227884 480 228124 0 FreeSans 960 0 0 0 analog_io[26]
port 18 nsew signal bidirectional
flabel metal3 s -960 175796 480 176036 0 FreeSans 960 0 0 0 analog_io[27]
port 19 nsew signal bidirectional
flabel metal3 s -960 123572 480 123812 0 FreeSans 960 0 0 0 analog_io[28]
port 20 nsew signal bidirectional
flabel metal3 s 583520 391628 584960 391868 0 FreeSans 960 0 0 0 analog_io[2]
port 21 nsew signal bidirectional
flabel metal3 s 583520 444668 584960 444908 0 FreeSans 960 0 0 0 analog_io[3]
port 22 nsew signal bidirectional
flabel metal3 s 583520 497844 584960 498084 0 FreeSans 960 0 0 0 analog_io[4]
port 23 nsew signal bidirectional
flabel metal3 s 583520 551020 584960 551260 0 FreeSans 960 0 0 0 analog_io[5]
port 24 nsew signal bidirectional
flabel metal3 s 583520 604060 584960 604300 0 FreeSans 960 0 0 0 analog_io[6]
port 25 nsew signal bidirectional
flabel metal3 s 583520 657236 584960 657476 0 FreeSans 960 0 0 0 analog_io[7]
port 26 nsew signal bidirectional
flabel metal2 s 575818 703520 575930 704960 0 FreeSans 448 90 0 0 analog_io[8]
port 27 nsew signal bidirectional
flabel metal2 s 510958 703520 511070 704960 0 FreeSans 448 90 0 0 analog_io[9]
port 28 nsew signal bidirectional
flabel metal3 s 583520 6476 584960 6716 0 FreeSans 960 0 0 0 io_in[0]
port 29 nsew signal input
flabel metal3 s 583520 457996 584960 458236 0 FreeSans 960 0 0 0 io_in[10]
port 30 nsew signal input
flabel metal3 s 583520 511172 584960 511412 0 FreeSans 960 0 0 0 io_in[11]
port 31 nsew signal input
flabel metal3 s 583520 564212 584960 564452 0 FreeSans 960 0 0 0 io_in[12]
port 32 nsew signal input
flabel metal3 s 583520 617388 584960 617628 0 FreeSans 960 0 0 0 io_in[13]
port 33 nsew signal input
flabel metal3 s 583520 670564 584960 670804 0 FreeSans 960 0 0 0 io_in[14]
port 34 nsew signal input
flabel metal2 s 559626 703520 559738 704960 0 FreeSans 448 90 0 0 io_in[15]
port 35 nsew signal input
flabel metal2 s 494766 703520 494878 704960 0 FreeSans 448 90 0 0 io_in[16]
port 36 nsew signal input
flabel metal2 s 429814 703520 429926 704960 0 FreeSans 448 90 0 0 io_in[17]
port 37 nsew signal input
flabel metal2 s 364954 703520 365066 704960 0 FreeSans 448 90 0 0 io_in[18]
port 38 nsew signal input
flabel metal2 s 300094 703520 300206 704960 0 FreeSans 448 90 0 0 io_in[19]
port 39 nsew signal input
flabel metal3 s 583520 46188 584960 46428 0 FreeSans 960 0 0 0 io_in[1]
port 40 nsew signal input
flabel metal2 s 235142 703520 235254 704960 0 FreeSans 448 90 0 0 io_in[20]
port 41 nsew signal input
flabel metal2 s 170282 703520 170394 704960 0 FreeSans 448 90 0 0 io_in[21]
port 42 nsew signal input
flabel metal2 s 105422 703520 105534 704960 0 FreeSans 448 90 0 0 io_in[22]
port 43 nsew signal input
flabel metal2 s 40470 703520 40582 704960 0 FreeSans 448 90 0 0 io_in[23]
port 44 nsew signal input
flabel metal3 s -960 684164 480 684404 0 FreeSans 960 0 0 0 io_in[24]
port 45 nsew signal input
flabel metal3 s -960 631940 480 632180 0 FreeSans 960 0 0 0 io_in[25]
port 46 nsew signal input
flabel metal3 s -960 579852 480 580092 0 FreeSans 960 0 0 0 io_in[26]
port 47 nsew signal input
flabel metal3 s -960 527764 480 528004 0 FreeSans 960 0 0 0 io_in[27]
port 48 nsew signal input
flabel metal3 s -960 475540 480 475780 0 FreeSans 960 0 0 0 io_in[28]
port 49 nsew signal input
flabel metal3 s -960 423452 480 423692 0 FreeSans 960 0 0 0 io_in[29]
port 50 nsew signal input
flabel metal3 s 583520 86036 584960 86276 0 FreeSans 960 0 0 0 io_in[2]
port 51 nsew signal input
flabel metal3 s -960 371228 480 371468 0 FreeSans 960 0 0 0 io_in[30]
port 52 nsew signal input
flabel metal3 s -960 319140 480 319380 0 FreeSans 960 0 0 0 io_in[31]
port 53 nsew signal input
flabel metal3 s -960 267052 480 267292 0 FreeSans 960 0 0 0 io_in[32]
port 54 nsew signal input
flabel metal3 s -960 214828 480 215068 0 FreeSans 960 0 0 0 io_in[33]
port 55 nsew signal input
flabel metal3 s -960 162740 480 162980 0 FreeSans 960 0 0 0 io_in[34]
port 56 nsew signal input
flabel metal3 s -960 110516 480 110756 0 FreeSans 960 0 0 0 io_in[35]
port 57 nsew signal input
flabel metal3 s -960 71484 480 71724 0 FreeSans 960 0 0 0 io_in[36]
port 58 nsew signal input
flabel metal3 s -960 32316 480 32556 0 FreeSans 960 0 0 0 io_in[37]
port 59 nsew signal input
flabel metal3 s 583520 125884 584960 126124 0 FreeSans 960 0 0 0 io_in[3]
port 60 nsew signal input
flabel metal3 s 583520 165732 584960 165972 0 FreeSans 960 0 0 0 io_in[4]
port 61 nsew signal input
flabel metal3 s 583520 205580 584960 205820 0 FreeSans 960 0 0 0 io_in[5]
port 62 nsew signal input
flabel metal3 s 583520 245428 584960 245668 0 FreeSans 960 0 0 0 io_in[6]
port 63 nsew signal input
flabel metal3 s 583520 298604 584960 298844 0 FreeSans 960 0 0 0 io_in[7]
port 64 nsew signal input
flabel metal3 s 583520 351780 584960 352020 0 FreeSans 960 0 0 0 io_in[8]
port 65 nsew signal input
flabel metal3 s 583520 404820 584960 405060 0 FreeSans 960 0 0 0 io_in[9]
port 66 nsew signal input
flabel metal3 s 583520 32996 584960 33236 0 FreeSans 960 0 0 0 io_oeb[0]
port 67 nsew signal tristate
flabel metal3 s 583520 484516 584960 484756 0 FreeSans 960 0 0 0 io_oeb[10]
port 68 nsew signal tristate
flabel metal3 s 583520 537692 584960 537932 0 FreeSans 960 0 0 0 io_oeb[11]
port 69 nsew signal tristate
flabel metal3 s 583520 590868 584960 591108 0 FreeSans 960 0 0 0 io_oeb[12]
port 70 nsew signal tristate
flabel metal3 s 583520 643908 584960 644148 0 FreeSans 960 0 0 0 io_oeb[13]
port 71 nsew signal tristate
flabel metal3 s 583520 697084 584960 697324 0 FreeSans 960 0 0 0 io_oeb[14]
port 72 nsew signal tristate
flabel metal2 s 527150 703520 527262 704960 0 FreeSans 448 90 0 0 io_oeb[15]
port 73 nsew signal tristate
flabel metal2 s 462290 703520 462402 704960 0 FreeSans 448 90 0 0 io_oeb[16]
port 74 nsew signal tristate
flabel metal2 s 397430 703520 397542 704960 0 FreeSans 448 90 0 0 io_oeb[17]
port 75 nsew signal tristate
flabel metal2 s 332478 703520 332590 704960 0 FreeSans 448 90 0 0 io_oeb[18]
port 76 nsew signal tristate
flabel metal2 s 267618 703520 267730 704960 0 FreeSans 448 90 0 0 io_oeb[19]
port 77 nsew signal tristate
flabel metal3 s 583520 72844 584960 73084 0 FreeSans 960 0 0 0 io_oeb[1]
port 78 nsew signal tristate
flabel metal2 s 202758 703520 202870 704960 0 FreeSans 448 90 0 0 io_oeb[20]
port 79 nsew signal tristate
flabel metal2 s 137806 703520 137918 704960 0 FreeSans 448 90 0 0 io_oeb[21]
port 80 nsew signal tristate
flabel metal2 s 72946 703520 73058 704960 0 FreeSans 448 90 0 0 io_oeb[22]
port 81 nsew signal tristate
flabel metal2 s 8086 703520 8198 704960 0 FreeSans 448 90 0 0 io_oeb[23]
port 82 nsew signal tristate
flabel metal3 s -960 658052 480 658292 0 FreeSans 960 0 0 0 io_oeb[24]
port 83 nsew signal tristate
flabel metal3 s -960 605964 480 606204 0 FreeSans 960 0 0 0 io_oeb[25]
port 84 nsew signal tristate
flabel metal3 s -960 553740 480 553980 0 FreeSans 960 0 0 0 io_oeb[26]
port 85 nsew signal tristate
flabel metal3 s -960 501652 480 501892 0 FreeSans 960 0 0 0 io_oeb[27]
port 86 nsew signal tristate
flabel metal3 s -960 449428 480 449668 0 FreeSans 960 0 0 0 io_oeb[28]
port 87 nsew signal tristate
flabel metal3 s -960 397340 480 397580 0 FreeSans 960 0 0 0 io_oeb[29]
port 88 nsew signal tristate
flabel metal3 s 583520 112692 584960 112932 0 FreeSans 960 0 0 0 io_oeb[2]
port 89 nsew signal tristate
flabel metal3 s -960 345252 480 345492 0 FreeSans 960 0 0 0 io_oeb[30]
port 90 nsew signal tristate
flabel metal3 s -960 293028 480 293268 0 FreeSans 960 0 0 0 io_oeb[31]
port 91 nsew signal tristate
flabel metal3 s -960 240940 480 241180 0 FreeSans 960 0 0 0 io_oeb[32]
port 92 nsew signal tristate
flabel metal3 s -960 188716 480 188956 0 FreeSans 960 0 0 0 io_oeb[33]
port 93 nsew signal tristate
flabel metal3 s -960 136628 480 136868 0 FreeSans 960 0 0 0 io_oeb[34]
port 94 nsew signal tristate
flabel metal3 s -960 84540 480 84780 0 FreeSans 960 0 0 0 io_oeb[35]
port 95 nsew signal tristate
flabel metal3 s -960 45372 480 45612 0 FreeSans 960 0 0 0 io_oeb[36]
port 96 nsew signal tristate
flabel metal3 s -960 6340 480 6580 0 FreeSans 960 0 0 0 io_oeb[37]
port 97 nsew signal tristate
flabel metal3 s 583520 152540 584960 152780 0 FreeSans 960 0 0 0 io_oeb[3]
port 98 nsew signal tristate
flabel metal3 s 583520 192388 584960 192628 0 FreeSans 960 0 0 0 io_oeb[4]
port 99 nsew signal tristate
flabel metal3 s 583520 232236 584960 232476 0 FreeSans 960 0 0 0 io_oeb[5]
port 100 nsew signal tristate
flabel metal3 s 583520 272084 584960 272324 0 FreeSans 960 0 0 0 io_oeb[6]
port 101 nsew signal tristate
flabel metal3 s 583520 325124 584960 325364 0 FreeSans 960 0 0 0 io_oeb[7]
port 102 nsew signal tristate
flabel metal3 s 583520 378300 584960 378540 0 FreeSans 960 0 0 0 io_oeb[8]
port 103 nsew signal tristate
flabel metal3 s 583520 431476 584960 431716 0 FreeSans 960 0 0 0 io_oeb[9]
port 104 nsew signal tristate
flabel metal3 s 583520 19668 584960 19908 0 FreeSans 960 0 0 0 io_out[0]
port 105 nsew signal tristate
flabel metal3 s 583520 471324 584960 471564 0 FreeSans 960 0 0 0 io_out[10]
port 106 nsew signal tristate
flabel metal3 s 583520 524364 584960 524604 0 FreeSans 960 0 0 0 io_out[11]
port 107 nsew signal tristate
flabel metal3 s 583520 577540 584960 577780 0 FreeSans 960 0 0 0 io_out[12]
port 108 nsew signal tristate
flabel metal3 s 583520 630716 584960 630956 0 FreeSans 960 0 0 0 io_out[13]
port 109 nsew signal tristate
flabel metal3 s 583520 683756 584960 683996 0 FreeSans 960 0 0 0 io_out[14]
port 110 nsew signal tristate
flabel metal2 s 543434 703520 543546 704960 0 FreeSans 448 90 0 0 io_out[15]
port 111 nsew signal tristate
flabel metal2 s 478482 703520 478594 704960 0 FreeSans 448 90 0 0 io_out[16]
port 112 nsew signal tristate
flabel metal2 s 413622 703520 413734 704960 0 FreeSans 448 90 0 0 io_out[17]
port 113 nsew signal tristate
flabel metal2 s 348762 703520 348874 704960 0 FreeSans 448 90 0 0 io_out[18]
port 114 nsew signal tristate
flabel metal2 s 283810 703520 283922 704960 0 FreeSans 448 90 0 0 io_out[19]
port 115 nsew signal tristate
flabel metal3 s 583520 59516 584960 59756 0 FreeSans 960 0 0 0 io_out[1]
port 116 nsew signal tristate
flabel metal2 s 218950 703520 219062 704960 0 FreeSans 448 90 0 0 io_out[20]
port 117 nsew signal tristate
flabel metal2 s 154090 703520 154202 704960 0 FreeSans 448 90 0 0 io_out[21]
port 118 nsew signal tristate
flabel metal2 s 89138 703520 89250 704960 0 FreeSans 448 90 0 0 io_out[22]
port 119 nsew signal tristate
flabel metal2 s 24278 703520 24390 704960 0 FreeSans 448 90 0 0 io_out[23]
port 120 nsew signal tristate
flabel metal3 s -960 671108 480 671348 0 FreeSans 960 0 0 0 io_out[24]
port 121 nsew signal tristate
flabel metal3 s -960 619020 480 619260 0 FreeSans 960 0 0 0 io_out[25]
port 122 nsew signal tristate
flabel metal3 s -960 566796 480 567036 0 FreeSans 960 0 0 0 io_out[26]
port 123 nsew signal tristate
flabel metal3 s -960 514708 480 514948 0 FreeSans 960 0 0 0 io_out[27]
port 124 nsew signal tristate
flabel metal3 s -960 462484 480 462724 0 FreeSans 960 0 0 0 io_out[28]
port 125 nsew signal tristate
flabel metal3 s -960 410396 480 410636 0 FreeSans 960 0 0 0 io_out[29]
port 126 nsew signal tristate
flabel metal3 s 583520 99364 584960 99604 0 FreeSans 960 0 0 0 io_out[2]
port 127 nsew signal tristate
flabel metal3 s -960 358308 480 358548 0 FreeSans 960 0 0 0 io_out[30]
port 128 nsew signal tristate
flabel metal3 s -960 306084 480 306324 0 FreeSans 960 0 0 0 io_out[31]
port 129 nsew signal tristate
flabel metal3 s -960 253996 480 254236 0 FreeSans 960 0 0 0 io_out[32]
port 130 nsew signal tristate
flabel metal3 s -960 201772 480 202012 0 FreeSans 960 0 0 0 io_out[33]
port 131 nsew signal tristate
flabel metal3 s -960 149684 480 149924 0 FreeSans 960 0 0 0 io_out[34]
port 132 nsew signal tristate
flabel metal3 s -960 97460 480 97700 0 FreeSans 960 0 0 0 io_out[35]
port 133 nsew signal tristate
flabel metal3 s -960 58428 480 58668 0 FreeSans 960 0 0 0 io_out[36]
port 134 nsew signal tristate
flabel metal3 s -960 19260 480 19500 0 FreeSans 960 0 0 0 io_out[37]
port 135 nsew signal tristate
flabel metal3 s 583520 139212 584960 139452 0 FreeSans 960 0 0 0 io_out[3]
port 136 nsew signal tristate
flabel metal3 s 583520 179060 584960 179300 0 FreeSans 960 0 0 0 io_out[4]
port 137 nsew signal tristate
flabel metal3 s 583520 218908 584960 219148 0 FreeSans 960 0 0 0 io_out[5]
port 138 nsew signal tristate
flabel metal3 s 583520 258756 584960 258996 0 FreeSans 960 0 0 0 io_out[6]
port 139 nsew signal tristate
flabel metal3 s 583520 311932 584960 312172 0 FreeSans 960 0 0 0 io_out[7]
port 140 nsew signal tristate
flabel metal3 s 583520 364972 584960 365212 0 FreeSans 960 0 0 0 io_out[8]
port 141 nsew signal tristate
flabel metal3 s 583520 418148 584960 418388 0 FreeSans 960 0 0 0 io_out[9]
port 142 nsew signal tristate
flabel metal2 s 125846 -960 125958 480 0 FreeSans 448 90 0 0 la_data_in[0]
port 143 nsew signal input
flabel metal2 s 480506 -960 480618 480 0 FreeSans 448 90 0 0 la_data_in[100]
port 144 nsew signal input
flabel metal2 s 484002 -960 484114 480 0 FreeSans 448 90 0 0 la_data_in[101]
port 145 nsew signal input
flabel metal2 s 487590 -960 487702 480 0 FreeSans 448 90 0 0 la_data_in[102]
port 146 nsew signal input
flabel metal2 s 491086 -960 491198 480 0 FreeSans 448 90 0 0 la_data_in[103]
port 147 nsew signal input
flabel metal2 s 494674 -960 494786 480 0 FreeSans 448 90 0 0 la_data_in[104]
port 148 nsew signal input
flabel metal2 s 498170 -960 498282 480 0 FreeSans 448 90 0 0 la_data_in[105]
port 149 nsew signal input
flabel metal2 s 501758 -960 501870 480 0 FreeSans 448 90 0 0 la_data_in[106]
port 150 nsew signal input
flabel metal2 s 505346 -960 505458 480 0 FreeSans 448 90 0 0 la_data_in[107]
port 151 nsew signal input
flabel metal2 s 508842 -960 508954 480 0 FreeSans 448 90 0 0 la_data_in[108]
port 152 nsew signal input
flabel metal2 s 512430 -960 512542 480 0 FreeSans 448 90 0 0 la_data_in[109]
port 153 nsew signal input
flabel metal2 s 161266 -960 161378 480 0 FreeSans 448 90 0 0 la_data_in[10]
port 154 nsew signal input
flabel metal2 s 515926 -960 516038 480 0 FreeSans 448 90 0 0 la_data_in[110]
port 155 nsew signal input
flabel metal2 s 519514 -960 519626 480 0 FreeSans 448 90 0 0 la_data_in[111]
port 156 nsew signal input
flabel metal2 s 523010 -960 523122 480 0 FreeSans 448 90 0 0 la_data_in[112]
port 157 nsew signal input
flabel metal2 s 526598 -960 526710 480 0 FreeSans 448 90 0 0 la_data_in[113]
port 158 nsew signal input
flabel metal2 s 530094 -960 530206 480 0 FreeSans 448 90 0 0 la_data_in[114]
port 159 nsew signal input
flabel metal2 s 533682 -960 533794 480 0 FreeSans 448 90 0 0 la_data_in[115]
port 160 nsew signal input
flabel metal2 s 537178 -960 537290 480 0 FreeSans 448 90 0 0 la_data_in[116]
port 161 nsew signal input
flabel metal2 s 540766 -960 540878 480 0 FreeSans 448 90 0 0 la_data_in[117]
port 162 nsew signal input
flabel metal2 s 544354 -960 544466 480 0 FreeSans 448 90 0 0 la_data_in[118]
port 163 nsew signal input
flabel metal2 s 547850 -960 547962 480 0 FreeSans 448 90 0 0 la_data_in[119]
port 164 nsew signal input
flabel metal2 s 164854 -960 164966 480 0 FreeSans 448 90 0 0 la_data_in[11]
port 165 nsew signal input
flabel metal2 s 551438 -960 551550 480 0 FreeSans 448 90 0 0 la_data_in[120]
port 166 nsew signal input
flabel metal2 s 554934 -960 555046 480 0 FreeSans 448 90 0 0 la_data_in[121]
port 167 nsew signal input
flabel metal2 s 558522 -960 558634 480 0 FreeSans 448 90 0 0 la_data_in[122]
port 168 nsew signal input
flabel metal2 s 562018 -960 562130 480 0 FreeSans 448 90 0 0 la_data_in[123]
port 169 nsew signal input
flabel metal2 s 565606 -960 565718 480 0 FreeSans 448 90 0 0 la_data_in[124]
port 170 nsew signal input
flabel metal2 s 569102 -960 569214 480 0 FreeSans 448 90 0 0 la_data_in[125]
port 171 nsew signal input
flabel metal2 s 572690 -960 572802 480 0 FreeSans 448 90 0 0 la_data_in[126]
port 172 nsew signal input
flabel metal2 s 576278 -960 576390 480 0 FreeSans 448 90 0 0 la_data_in[127]
port 173 nsew signal input
flabel metal2 s 168350 -960 168462 480 0 FreeSans 448 90 0 0 la_data_in[12]
port 174 nsew signal input
flabel metal2 s 171938 -960 172050 480 0 FreeSans 448 90 0 0 la_data_in[13]
port 175 nsew signal input
flabel metal2 s 175434 -960 175546 480 0 FreeSans 448 90 0 0 la_data_in[14]
port 176 nsew signal input
flabel metal2 s 179022 -960 179134 480 0 FreeSans 448 90 0 0 la_data_in[15]
port 177 nsew signal input
flabel metal2 s 182518 -960 182630 480 0 FreeSans 448 90 0 0 la_data_in[16]
port 178 nsew signal input
flabel metal2 s 186106 -960 186218 480 0 FreeSans 448 90 0 0 la_data_in[17]
port 179 nsew signal input
flabel metal2 s 189694 -960 189806 480 0 FreeSans 448 90 0 0 la_data_in[18]
port 180 nsew signal input
flabel metal2 s 193190 -960 193302 480 0 FreeSans 448 90 0 0 la_data_in[19]
port 181 nsew signal input
flabel metal2 s 129342 -960 129454 480 0 FreeSans 448 90 0 0 la_data_in[1]
port 182 nsew signal input
flabel metal2 s 196778 -960 196890 480 0 FreeSans 448 90 0 0 la_data_in[20]
port 183 nsew signal input
flabel metal2 s 200274 -960 200386 480 0 FreeSans 448 90 0 0 la_data_in[21]
port 184 nsew signal input
flabel metal2 s 203862 -960 203974 480 0 FreeSans 448 90 0 0 la_data_in[22]
port 185 nsew signal input
flabel metal2 s 207358 -960 207470 480 0 FreeSans 448 90 0 0 la_data_in[23]
port 186 nsew signal input
flabel metal2 s 210946 -960 211058 480 0 FreeSans 448 90 0 0 la_data_in[24]
port 187 nsew signal input
flabel metal2 s 214442 -960 214554 480 0 FreeSans 448 90 0 0 la_data_in[25]
port 188 nsew signal input
flabel metal2 s 218030 -960 218142 480 0 FreeSans 448 90 0 0 la_data_in[26]
port 189 nsew signal input
flabel metal2 s 221526 -960 221638 480 0 FreeSans 448 90 0 0 la_data_in[27]
port 190 nsew signal input
flabel metal2 s 225114 -960 225226 480 0 FreeSans 448 90 0 0 la_data_in[28]
port 191 nsew signal input
flabel metal2 s 228702 -960 228814 480 0 FreeSans 448 90 0 0 la_data_in[29]
port 192 nsew signal input
flabel metal2 s 132930 -960 133042 480 0 FreeSans 448 90 0 0 la_data_in[2]
port 193 nsew signal input
flabel metal2 s 232198 -960 232310 480 0 FreeSans 448 90 0 0 la_data_in[30]
port 194 nsew signal input
flabel metal2 s 235786 -960 235898 480 0 FreeSans 448 90 0 0 la_data_in[31]
port 195 nsew signal input
flabel metal2 s 239282 -960 239394 480 0 FreeSans 448 90 0 0 la_data_in[32]
port 196 nsew signal input
flabel metal2 s 242870 -960 242982 480 0 FreeSans 448 90 0 0 la_data_in[33]
port 197 nsew signal input
flabel metal2 s 246366 -960 246478 480 0 FreeSans 448 90 0 0 la_data_in[34]
port 198 nsew signal input
flabel metal2 s 249954 -960 250066 480 0 FreeSans 448 90 0 0 la_data_in[35]
port 199 nsew signal input
flabel metal2 s 253450 -960 253562 480 0 FreeSans 448 90 0 0 la_data_in[36]
port 200 nsew signal input
flabel metal2 s 257038 -960 257150 480 0 FreeSans 448 90 0 0 la_data_in[37]
port 201 nsew signal input
flabel metal2 s 260626 -960 260738 480 0 FreeSans 448 90 0 0 la_data_in[38]
port 202 nsew signal input
flabel metal2 s 264122 -960 264234 480 0 FreeSans 448 90 0 0 la_data_in[39]
port 203 nsew signal input
flabel metal2 s 136426 -960 136538 480 0 FreeSans 448 90 0 0 la_data_in[3]
port 204 nsew signal input
flabel metal2 s 267710 -960 267822 480 0 FreeSans 448 90 0 0 la_data_in[40]
port 205 nsew signal input
flabel metal2 s 271206 -960 271318 480 0 FreeSans 448 90 0 0 la_data_in[41]
port 206 nsew signal input
flabel metal2 s 274794 -960 274906 480 0 FreeSans 448 90 0 0 la_data_in[42]
port 207 nsew signal input
flabel metal2 s 278290 -960 278402 480 0 FreeSans 448 90 0 0 la_data_in[43]
port 208 nsew signal input
flabel metal2 s 281878 -960 281990 480 0 FreeSans 448 90 0 0 la_data_in[44]
port 209 nsew signal input
flabel metal2 s 285374 -960 285486 480 0 FreeSans 448 90 0 0 la_data_in[45]
port 210 nsew signal input
flabel metal2 s 288962 -960 289074 480 0 FreeSans 448 90 0 0 la_data_in[46]
port 211 nsew signal input
flabel metal2 s 292550 -960 292662 480 0 FreeSans 448 90 0 0 la_data_in[47]
port 212 nsew signal input
flabel metal2 s 296046 -960 296158 480 0 FreeSans 448 90 0 0 la_data_in[48]
port 213 nsew signal input
flabel metal2 s 299634 -960 299746 480 0 FreeSans 448 90 0 0 la_data_in[49]
port 214 nsew signal input
flabel metal2 s 140014 -960 140126 480 0 FreeSans 448 90 0 0 la_data_in[4]
port 215 nsew signal input
flabel metal2 s 303130 -960 303242 480 0 FreeSans 448 90 0 0 la_data_in[50]
port 216 nsew signal input
flabel metal2 s 306718 -960 306830 480 0 FreeSans 448 90 0 0 la_data_in[51]
port 217 nsew signal input
flabel metal2 s 310214 -960 310326 480 0 FreeSans 448 90 0 0 la_data_in[52]
port 218 nsew signal input
flabel metal2 s 313802 -960 313914 480 0 FreeSans 448 90 0 0 la_data_in[53]
port 219 nsew signal input
flabel metal2 s 317298 -960 317410 480 0 FreeSans 448 90 0 0 la_data_in[54]
port 220 nsew signal input
flabel metal2 s 320886 -960 320998 480 0 FreeSans 448 90 0 0 la_data_in[55]
port 221 nsew signal input
flabel metal2 s 324382 -960 324494 480 0 FreeSans 448 90 0 0 la_data_in[56]
port 222 nsew signal input
flabel metal2 s 327970 -960 328082 480 0 FreeSans 448 90 0 0 la_data_in[57]
port 223 nsew signal input
flabel metal2 s 331558 -960 331670 480 0 FreeSans 448 90 0 0 la_data_in[58]
port 224 nsew signal input
flabel metal2 s 335054 -960 335166 480 0 FreeSans 448 90 0 0 la_data_in[59]
port 225 nsew signal input
flabel metal2 s 143510 -960 143622 480 0 FreeSans 448 90 0 0 la_data_in[5]
port 226 nsew signal input
flabel metal2 s 338642 -960 338754 480 0 FreeSans 448 90 0 0 la_data_in[60]
port 227 nsew signal input
flabel metal2 s 342138 -960 342250 480 0 FreeSans 448 90 0 0 la_data_in[61]
port 228 nsew signal input
flabel metal2 s 345726 -960 345838 480 0 FreeSans 448 90 0 0 la_data_in[62]
port 229 nsew signal input
flabel metal2 s 349222 -960 349334 480 0 FreeSans 448 90 0 0 la_data_in[63]
port 230 nsew signal input
flabel metal2 s 352810 -960 352922 480 0 FreeSans 448 90 0 0 la_data_in[64]
port 231 nsew signal input
flabel metal2 s 356306 -960 356418 480 0 FreeSans 448 90 0 0 la_data_in[65]
port 232 nsew signal input
flabel metal2 s 359894 -960 360006 480 0 FreeSans 448 90 0 0 la_data_in[66]
port 233 nsew signal input
flabel metal2 s 363482 -960 363594 480 0 FreeSans 448 90 0 0 la_data_in[67]
port 234 nsew signal input
flabel metal2 s 366978 -960 367090 480 0 FreeSans 448 90 0 0 la_data_in[68]
port 235 nsew signal input
flabel metal2 s 370566 -960 370678 480 0 FreeSans 448 90 0 0 la_data_in[69]
port 236 nsew signal input
flabel metal2 s 147098 -960 147210 480 0 FreeSans 448 90 0 0 la_data_in[6]
port 237 nsew signal input
flabel metal2 s 374062 -960 374174 480 0 FreeSans 448 90 0 0 la_data_in[70]
port 238 nsew signal input
flabel metal2 s 377650 -960 377762 480 0 FreeSans 448 90 0 0 la_data_in[71]
port 239 nsew signal input
flabel metal2 s 381146 -960 381258 480 0 FreeSans 448 90 0 0 la_data_in[72]
port 240 nsew signal input
flabel metal2 s 384734 -960 384846 480 0 FreeSans 448 90 0 0 la_data_in[73]
port 241 nsew signal input
flabel metal2 s 388230 -960 388342 480 0 FreeSans 448 90 0 0 la_data_in[74]
port 242 nsew signal input
flabel metal2 s 391818 -960 391930 480 0 FreeSans 448 90 0 0 la_data_in[75]
port 243 nsew signal input
flabel metal2 s 395314 -960 395426 480 0 FreeSans 448 90 0 0 la_data_in[76]
port 244 nsew signal input
flabel metal2 s 398902 -960 399014 480 0 FreeSans 448 90 0 0 la_data_in[77]
port 245 nsew signal input
flabel metal2 s 402490 -960 402602 480 0 FreeSans 448 90 0 0 la_data_in[78]
port 246 nsew signal input
flabel metal2 s 405986 -960 406098 480 0 FreeSans 448 90 0 0 la_data_in[79]
port 247 nsew signal input
flabel metal2 s 150594 -960 150706 480 0 FreeSans 448 90 0 0 la_data_in[7]
port 248 nsew signal input
flabel metal2 s 409574 -960 409686 480 0 FreeSans 448 90 0 0 la_data_in[80]
port 249 nsew signal input
flabel metal2 s 413070 -960 413182 480 0 FreeSans 448 90 0 0 la_data_in[81]
port 250 nsew signal input
flabel metal2 s 416658 -960 416770 480 0 FreeSans 448 90 0 0 la_data_in[82]
port 251 nsew signal input
flabel metal2 s 420154 -960 420266 480 0 FreeSans 448 90 0 0 la_data_in[83]
port 252 nsew signal input
flabel metal2 s 423742 -960 423854 480 0 FreeSans 448 90 0 0 la_data_in[84]
port 253 nsew signal input
flabel metal2 s 427238 -960 427350 480 0 FreeSans 448 90 0 0 la_data_in[85]
port 254 nsew signal input
flabel metal2 s 430826 -960 430938 480 0 FreeSans 448 90 0 0 la_data_in[86]
port 255 nsew signal input
flabel metal2 s 434414 -960 434526 480 0 FreeSans 448 90 0 0 la_data_in[87]
port 256 nsew signal input
flabel metal2 s 437910 -960 438022 480 0 FreeSans 448 90 0 0 la_data_in[88]
port 257 nsew signal input
flabel metal2 s 441498 -960 441610 480 0 FreeSans 448 90 0 0 la_data_in[89]
port 258 nsew signal input
flabel metal2 s 154182 -960 154294 480 0 FreeSans 448 90 0 0 la_data_in[8]
port 259 nsew signal input
flabel metal2 s 444994 -960 445106 480 0 FreeSans 448 90 0 0 la_data_in[90]
port 260 nsew signal input
flabel metal2 s 448582 -960 448694 480 0 FreeSans 448 90 0 0 la_data_in[91]
port 261 nsew signal input
flabel metal2 s 452078 -960 452190 480 0 FreeSans 448 90 0 0 la_data_in[92]
port 262 nsew signal input
flabel metal2 s 455666 -960 455778 480 0 FreeSans 448 90 0 0 la_data_in[93]
port 263 nsew signal input
flabel metal2 s 459162 -960 459274 480 0 FreeSans 448 90 0 0 la_data_in[94]
port 264 nsew signal input
flabel metal2 s 462750 -960 462862 480 0 FreeSans 448 90 0 0 la_data_in[95]
port 265 nsew signal input
flabel metal2 s 466246 -960 466358 480 0 FreeSans 448 90 0 0 la_data_in[96]
port 266 nsew signal input
flabel metal2 s 469834 -960 469946 480 0 FreeSans 448 90 0 0 la_data_in[97]
port 267 nsew signal input
flabel metal2 s 473422 -960 473534 480 0 FreeSans 448 90 0 0 la_data_in[98]
port 268 nsew signal input
flabel metal2 s 476918 -960 477030 480 0 FreeSans 448 90 0 0 la_data_in[99]
port 269 nsew signal input
flabel metal2 s 157770 -960 157882 480 0 FreeSans 448 90 0 0 la_data_in[9]
port 270 nsew signal input
flabel metal2 s 126950 -960 127062 480 0 FreeSans 448 90 0 0 la_data_out[0]
port 271 nsew signal tristate
flabel metal2 s 481702 -960 481814 480 0 FreeSans 448 90 0 0 la_data_out[100]
port 272 nsew signal tristate
flabel metal2 s 485198 -960 485310 480 0 FreeSans 448 90 0 0 la_data_out[101]
port 273 nsew signal tristate
flabel metal2 s 488786 -960 488898 480 0 FreeSans 448 90 0 0 la_data_out[102]
port 274 nsew signal tristate
flabel metal2 s 492282 -960 492394 480 0 FreeSans 448 90 0 0 la_data_out[103]
port 275 nsew signal tristate
flabel metal2 s 495870 -960 495982 480 0 FreeSans 448 90 0 0 la_data_out[104]
port 276 nsew signal tristate
flabel metal2 s 499366 -960 499478 480 0 FreeSans 448 90 0 0 la_data_out[105]
port 277 nsew signal tristate
flabel metal2 s 502954 -960 503066 480 0 FreeSans 448 90 0 0 la_data_out[106]
port 278 nsew signal tristate
flabel metal2 s 506450 -960 506562 480 0 FreeSans 448 90 0 0 la_data_out[107]
port 279 nsew signal tristate
flabel metal2 s 510038 -960 510150 480 0 FreeSans 448 90 0 0 la_data_out[108]
port 280 nsew signal tristate
flabel metal2 s 513534 -960 513646 480 0 FreeSans 448 90 0 0 la_data_out[109]
port 281 nsew signal tristate
flabel metal2 s 162462 -960 162574 480 0 FreeSans 448 90 0 0 la_data_out[10]
port 282 nsew signal tristate
flabel metal2 s 517122 -960 517234 480 0 FreeSans 448 90 0 0 la_data_out[110]
port 283 nsew signal tristate
flabel metal2 s 520710 -960 520822 480 0 FreeSans 448 90 0 0 la_data_out[111]
port 284 nsew signal tristate
flabel metal2 s 524206 -960 524318 480 0 FreeSans 448 90 0 0 la_data_out[112]
port 285 nsew signal tristate
flabel metal2 s 527794 -960 527906 480 0 FreeSans 448 90 0 0 la_data_out[113]
port 286 nsew signal tristate
flabel metal2 s 531290 -960 531402 480 0 FreeSans 448 90 0 0 la_data_out[114]
port 287 nsew signal tristate
flabel metal2 s 534878 -960 534990 480 0 FreeSans 448 90 0 0 la_data_out[115]
port 288 nsew signal tristate
flabel metal2 s 538374 -960 538486 480 0 FreeSans 448 90 0 0 la_data_out[116]
port 289 nsew signal tristate
flabel metal2 s 541962 -960 542074 480 0 FreeSans 448 90 0 0 la_data_out[117]
port 290 nsew signal tristate
flabel metal2 s 545458 -960 545570 480 0 FreeSans 448 90 0 0 la_data_out[118]
port 291 nsew signal tristate
flabel metal2 s 549046 -960 549158 480 0 FreeSans 448 90 0 0 la_data_out[119]
port 292 nsew signal tristate
flabel metal2 s 166050 -960 166162 480 0 FreeSans 448 90 0 0 la_data_out[11]
port 293 nsew signal tristate
flabel metal2 s 552634 -960 552746 480 0 FreeSans 448 90 0 0 la_data_out[120]
port 294 nsew signal tristate
flabel metal2 s 556130 -960 556242 480 0 FreeSans 448 90 0 0 la_data_out[121]
port 295 nsew signal tristate
flabel metal2 s 559718 -960 559830 480 0 FreeSans 448 90 0 0 la_data_out[122]
port 296 nsew signal tristate
flabel metal2 s 563214 -960 563326 480 0 FreeSans 448 90 0 0 la_data_out[123]
port 297 nsew signal tristate
flabel metal2 s 566802 -960 566914 480 0 FreeSans 448 90 0 0 la_data_out[124]
port 298 nsew signal tristate
flabel metal2 s 570298 -960 570410 480 0 FreeSans 448 90 0 0 la_data_out[125]
port 299 nsew signal tristate
flabel metal2 s 573886 -960 573998 480 0 FreeSans 448 90 0 0 la_data_out[126]
port 300 nsew signal tristate
flabel metal2 s 577382 -960 577494 480 0 FreeSans 448 90 0 0 la_data_out[127]
port 301 nsew signal tristate
flabel metal2 s 169546 -960 169658 480 0 FreeSans 448 90 0 0 la_data_out[12]
port 302 nsew signal tristate
flabel metal2 s 173134 -960 173246 480 0 FreeSans 448 90 0 0 la_data_out[13]
port 303 nsew signal tristate
flabel metal2 s 176630 -960 176742 480 0 FreeSans 448 90 0 0 la_data_out[14]
port 304 nsew signal tristate
flabel metal2 s 180218 -960 180330 480 0 FreeSans 448 90 0 0 la_data_out[15]
port 305 nsew signal tristate
flabel metal2 s 183714 -960 183826 480 0 FreeSans 448 90 0 0 la_data_out[16]
port 306 nsew signal tristate
flabel metal2 s 187302 -960 187414 480 0 FreeSans 448 90 0 0 la_data_out[17]
port 307 nsew signal tristate
flabel metal2 s 190798 -960 190910 480 0 FreeSans 448 90 0 0 la_data_out[18]
port 308 nsew signal tristate
flabel metal2 s 194386 -960 194498 480 0 FreeSans 448 90 0 0 la_data_out[19]
port 309 nsew signal tristate
flabel metal2 s 130538 -960 130650 480 0 FreeSans 448 90 0 0 la_data_out[1]
port 310 nsew signal tristate
flabel metal2 s 197882 -960 197994 480 0 FreeSans 448 90 0 0 la_data_out[20]
port 311 nsew signal tristate
flabel metal2 s 201470 -960 201582 480 0 FreeSans 448 90 0 0 la_data_out[21]
port 312 nsew signal tristate
flabel metal2 s 205058 -960 205170 480 0 FreeSans 448 90 0 0 la_data_out[22]
port 313 nsew signal tristate
flabel metal2 s 208554 -960 208666 480 0 FreeSans 448 90 0 0 la_data_out[23]
port 314 nsew signal tristate
flabel metal2 s 212142 -960 212254 480 0 FreeSans 448 90 0 0 la_data_out[24]
port 315 nsew signal tristate
flabel metal2 s 215638 -960 215750 480 0 FreeSans 448 90 0 0 la_data_out[25]
port 316 nsew signal tristate
flabel metal2 s 219226 -960 219338 480 0 FreeSans 448 90 0 0 la_data_out[26]
port 317 nsew signal tristate
flabel metal2 s 222722 -960 222834 480 0 FreeSans 448 90 0 0 la_data_out[27]
port 318 nsew signal tristate
flabel metal2 s 226310 -960 226422 480 0 FreeSans 448 90 0 0 la_data_out[28]
port 319 nsew signal tristate
flabel metal2 s 229806 -960 229918 480 0 FreeSans 448 90 0 0 la_data_out[29]
port 320 nsew signal tristate
flabel metal2 s 134126 -960 134238 480 0 FreeSans 448 90 0 0 la_data_out[2]
port 321 nsew signal tristate
flabel metal2 s 233394 -960 233506 480 0 FreeSans 448 90 0 0 la_data_out[30]
port 322 nsew signal tristate
flabel metal2 s 236982 -960 237094 480 0 FreeSans 448 90 0 0 la_data_out[31]
port 323 nsew signal tristate
flabel metal2 s 240478 -960 240590 480 0 FreeSans 448 90 0 0 la_data_out[32]
port 324 nsew signal tristate
flabel metal2 s 244066 -960 244178 480 0 FreeSans 448 90 0 0 la_data_out[33]
port 325 nsew signal tristate
flabel metal2 s 247562 -960 247674 480 0 FreeSans 448 90 0 0 la_data_out[34]
port 326 nsew signal tristate
flabel metal2 s 251150 -960 251262 480 0 FreeSans 448 90 0 0 la_data_out[35]
port 327 nsew signal tristate
flabel metal2 s 254646 -960 254758 480 0 FreeSans 448 90 0 0 la_data_out[36]
port 328 nsew signal tristate
flabel metal2 s 258234 -960 258346 480 0 FreeSans 448 90 0 0 la_data_out[37]
port 329 nsew signal tristate
flabel metal2 s 261730 -960 261842 480 0 FreeSans 448 90 0 0 la_data_out[38]
port 330 nsew signal tristate
flabel metal2 s 265318 -960 265430 480 0 FreeSans 448 90 0 0 la_data_out[39]
port 331 nsew signal tristate
flabel metal2 s 137622 -960 137734 480 0 FreeSans 448 90 0 0 la_data_out[3]
port 332 nsew signal tristate
flabel metal2 s 268814 -960 268926 480 0 FreeSans 448 90 0 0 la_data_out[40]
port 333 nsew signal tristate
flabel metal2 s 272402 -960 272514 480 0 FreeSans 448 90 0 0 la_data_out[41]
port 334 nsew signal tristate
flabel metal2 s 275990 -960 276102 480 0 FreeSans 448 90 0 0 la_data_out[42]
port 335 nsew signal tristate
flabel metal2 s 279486 -960 279598 480 0 FreeSans 448 90 0 0 la_data_out[43]
port 336 nsew signal tristate
flabel metal2 s 283074 -960 283186 480 0 FreeSans 448 90 0 0 la_data_out[44]
port 337 nsew signal tristate
flabel metal2 s 286570 -960 286682 480 0 FreeSans 448 90 0 0 la_data_out[45]
port 338 nsew signal tristate
flabel metal2 s 290158 -960 290270 480 0 FreeSans 448 90 0 0 la_data_out[46]
port 339 nsew signal tristate
flabel metal2 s 293654 -960 293766 480 0 FreeSans 448 90 0 0 la_data_out[47]
port 340 nsew signal tristate
flabel metal2 s 297242 -960 297354 480 0 FreeSans 448 90 0 0 la_data_out[48]
port 341 nsew signal tristate
flabel metal2 s 300738 -960 300850 480 0 FreeSans 448 90 0 0 la_data_out[49]
port 342 nsew signal tristate
flabel metal2 s 141210 -960 141322 480 0 FreeSans 448 90 0 0 la_data_out[4]
port 343 nsew signal tristate
flabel metal2 s 304326 -960 304438 480 0 FreeSans 448 90 0 0 la_data_out[50]
port 344 nsew signal tristate
flabel metal2 s 307914 -960 308026 480 0 FreeSans 448 90 0 0 la_data_out[51]
port 345 nsew signal tristate
flabel metal2 s 311410 -960 311522 480 0 FreeSans 448 90 0 0 la_data_out[52]
port 346 nsew signal tristate
flabel metal2 s 314998 -960 315110 480 0 FreeSans 448 90 0 0 la_data_out[53]
port 347 nsew signal tristate
flabel metal2 s 318494 -960 318606 480 0 FreeSans 448 90 0 0 la_data_out[54]
port 348 nsew signal tristate
flabel metal2 s 322082 -960 322194 480 0 FreeSans 448 90 0 0 la_data_out[55]
port 349 nsew signal tristate
flabel metal2 s 325578 -960 325690 480 0 FreeSans 448 90 0 0 la_data_out[56]
port 350 nsew signal tristate
flabel metal2 s 329166 -960 329278 480 0 FreeSans 448 90 0 0 la_data_out[57]
port 351 nsew signal tristate
flabel metal2 s 332662 -960 332774 480 0 FreeSans 448 90 0 0 la_data_out[58]
port 352 nsew signal tristate
flabel metal2 s 336250 -960 336362 480 0 FreeSans 448 90 0 0 la_data_out[59]
port 353 nsew signal tristate
flabel metal2 s 144706 -960 144818 480 0 FreeSans 448 90 0 0 la_data_out[5]
port 354 nsew signal tristate
flabel metal2 s 339838 -960 339950 480 0 FreeSans 448 90 0 0 la_data_out[60]
port 355 nsew signal tristate
flabel metal2 s 343334 -960 343446 480 0 FreeSans 448 90 0 0 la_data_out[61]
port 356 nsew signal tristate
flabel metal2 s 346922 -960 347034 480 0 FreeSans 448 90 0 0 la_data_out[62]
port 357 nsew signal tristate
flabel metal2 s 350418 -960 350530 480 0 FreeSans 448 90 0 0 la_data_out[63]
port 358 nsew signal tristate
flabel metal2 s 354006 -960 354118 480 0 FreeSans 448 90 0 0 la_data_out[64]
port 359 nsew signal tristate
flabel metal2 s 357502 -960 357614 480 0 FreeSans 448 90 0 0 la_data_out[65]
port 360 nsew signal tristate
flabel metal2 s 361090 -960 361202 480 0 FreeSans 448 90 0 0 la_data_out[66]
port 361 nsew signal tristate
flabel metal2 s 364586 -960 364698 480 0 FreeSans 448 90 0 0 la_data_out[67]
port 362 nsew signal tristate
flabel metal2 s 368174 -960 368286 480 0 FreeSans 448 90 0 0 la_data_out[68]
port 363 nsew signal tristate
flabel metal2 s 371670 -960 371782 480 0 FreeSans 448 90 0 0 la_data_out[69]
port 364 nsew signal tristate
flabel metal2 s 148294 -960 148406 480 0 FreeSans 448 90 0 0 la_data_out[6]
port 365 nsew signal tristate
flabel metal2 s 375258 -960 375370 480 0 FreeSans 448 90 0 0 la_data_out[70]
port 366 nsew signal tristate
flabel metal2 s 378846 -960 378958 480 0 FreeSans 448 90 0 0 la_data_out[71]
port 367 nsew signal tristate
flabel metal2 s 382342 -960 382454 480 0 FreeSans 448 90 0 0 la_data_out[72]
port 368 nsew signal tristate
flabel metal2 s 385930 -960 386042 480 0 FreeSans 448 90 0 0 la_data_out[73]
port 369 nsew signal tristate
flabel metal2 s 389426 -960 389538 480 0 FreeSans 448 90 0 0 la_data_out[74]
port 370 nsew signal tristate
flabel metal2 s 393014 -960 393126 480 0 FreeSans 448 90 0 0 la_data_out[75]
port 371 nsew signal tristate
flabel metal2 s 396510 -960 396622 480 0 FreeSans 448 90 0 0 la_data_out[76]
port 372 nsew signal tristate
flabel metal2 s 400098 -960 400210 480 0 FreeSans 448 90 0 0 la_data_out[77]
port 373 nsew signal tristate
flabel metal2 s 403594 -960 403706 480 0 FreeSans 448 90 0 0 la_data_out[78]
port 374 nsew signal tristate
flabel metal2 s 407182 -960 407294 480 0 FreeSans 448 90 0 0 la_data_out[79]
port 375 nsew signal tristate
flabel metal2 s 151790 -960 151902 480 0 FreeSans 448 90 0 0 la_data_out[7]
port 376 nsew signal tristate
flabel metal2 s 410770 -960 410882 480 0 FreeSans 448 90 0 0 la_data_out[80]
port 377 nsew signal tristate
flabel metal2 s 414266 -960 414378 480 0 FreeSans 448 90 0 0 la_data_out[81]
port 378 nsew signal tristate
flabel metal2 s 417854 -960 417966 480 0 FreeSans 448 90 0 0 la_data_out[82]
port 379 nsew signal tristate
flabel metal2 s 421350 -960 421462 480 0 FreeSans 448 90 0 0 la_data_out[83]
port 380 nsew signal tristate
flabel metal2 s 424938 -960 425050 480 0 FreeSans 448 90 0 0 la_data_out[84]
port 381 nsew signal tristate
flabel metal2 s 428434 -960 428546 480 0 FreeSans 448 90 0 0 la_data_out[85]
port 382 nsew signal tristate
flabel metal2 s 432022 -960 432134 480 0 FreeSans 448 90 0 0 la_data_out[86]
port 383 nsew signal tristate
flabel metal2 s 435518 -960 435630 480 0 FreeSans 448 90 0 0 la_data_out[87]
port 384 nsew signal tristate
flabel metal2 s 439106 -960 439218 480 0 FreeSans 448 90 0 0 la_data_out[88]
port 385 nsew signal tristate
flabel metal2 s 442602 -960 442714 480 0 FreeSans 448 90 0 0 la_data_out[89]
port 386 nsew signal tristate
flabel metal2 s 155378 -960 155490 480 0 FreeSans 448 90 0 0 la_data_out[8]
port 387 nsew signal tristate
flabel metal2 s 446190 -960 446302 480 0 FreeSans 448 90 0 0 la_data_out[90]
port 388 nsew signal tristate
flabel metal2 s 449778 -960 449890 480 0 FreeSans 448 90 0 0 la_data_out[91]
port 389 nsew signal tristate
flabel metal2 s 453274 -960 453386 480 0 FreeSans 448 90 0 0 la_data_out[92]
port 390 nsew signal tristate
flabel metal2 s 456862 -960 456974 480 0 FreeSans 448 90 0 0 la_data_out[93]
port 391 nsew signal tristate
flabel metal2 s 460358 -960 460470 480 0 FreeSans 448 90 0 0 la_data_out[94]
port 392 nsew signal tristate
flabel metal2 s 463946 -960 464058 480 0 FreeSans 448 90 0 0 la_data_out[95]
port 393 nsew signal tristate
flabel metal2 s 467442 -960 467554 480 0 FreeSans 448 90 0 0 la_data_out[96]
port 394 nsew signal tristate
flabel metal2 s 471030 -960 471142 480 0 FreeSans 448 90 0 0 la_data_out[97]
port 395 nsew signal tristate
flabel metal2 s 474526 -960 474638 480 0 FreeSans 448 90 0 0 la_data_out[98]
port 396 nsew signal tristate
flabel metal2 s 478114 -960 478226 480 0 FreeSans 448 90 0 0 la_data_out[99]
port 397 nsew signal tristate
flabel metal2 s 158874 -960 158986 480 0 FreeSans 448 90 0 0 la_data_out[9]
port 398 nsew signal tristate
flabel metal2 s 128146 -960 128258 480 0 FreeSans 448 90 0 0 la_oenb[0]
port 399 nsew signal input
flabel metal2 s 482806 -960 482918 480 0 FreeSans 448 90 0 0 la_oenb[100]
port 400 nsew signal input
flabel metal2 s 486394 -960 486506 480 0 FreeSans 448 90 0 0 la_oenb[101]
port 401 nsew signal input
flabel metal2 s 489890 -960 490002 480 0 FreeSans 448 90 0 0 la_oenb[102]
port 402 nsew signal input
flabel metal2 s 493478 -960 493590 480 0 FreeSans 448 90 0 0 la_oenb[103]
port 403 nsew signal input
flabel metal2 s 497066 -960 497178 480 0 FreeSans 448 90 0 0 la_oenb[104]
port 404 nsew signal input
flabel metal2 s 500562 -960 500674 480 0 FreeSans 448 90 0 0 la_oenb[105]
port 405 nsew signal input
flabel metal2 s 504150 -960 504262 480 0 FreeSans 448 90 0 0 la_oenb[106]
port 406 nsew signal input
flabel metal2 s 507646 -960 507758 480 0 FreeSans 448 90 0 0 la_oenb[107]
port 407 nsew signal input
flabel metal2 s 511234 -960 511346 480 0 FreeSans 448 90 0 0 la_oenb[108]
port 408 nsew signal input
flabel metal2 s 514730 -960 514842 480 0 FreeSans 448 90 0 0 la_oenb[109]
port 409 nsew signal input
flabel metal2 s 163658 -960 163770 480 0 FreeSans 448 90 0 0 la_oenb[10]
port 410 nsew signal input
flabel metal2 s 518318 -960 518430 480 0 FreeSans 448 90 0 0 la_oenb[110]
port 411 nsew signal input
flabel metal2 s 521814 -960 521926 480 0 FreeSans 448 90 0 0 la_oenb[111]
port 412 nsew signal input
flabel metal2 s 525402 -960 525514 480 0 FreeSans 448 90 0 0 la_oenb[112]
port 413 nsew signal input
flabel metal2 s 528990 -960 529102 480 0 FreeSans 448 90 0 0 la_oenb[113]
port 414 nsew signal input
flabel metal2 s 532486 -960 532598 480 0 FreeSans 448 90 0 0 la_oenb[114]
port 415 nsew signal input
flabel metal2 s 536074 -960 536186 480 0 FreeSans 448 90 0 0 la_oenb[115]
port 416 nsew signal input
flabel metal2 s 539570 -960 539682 480 0 FreeSans 448 90 0 0 la_oenb[116]
port 417 nsew signal input
flabel metal2 s 543158 -960 543270 480 0 FreeSans 448 90 0 0 la_oenb[117]
port 418 nsew signal input
flabel metal2 s 546654 -960 546766 480 0 FreeSans 448 90 0 0 la_oenb[118]
port 419 nsew signal input
flabel metal2 s 550242 -960 550354 480 0 FreeSans 448 90 0 0 la_oenb[119]
port 420 nsew signal input
flabel metal2 s 167154 -960 167266 480 0 FreeSans 448 90 0 0 la_oenb[11]
port 421 nsew signal input
flabel metal2 s 553738 -960 553850 480 0 FreeSans 448 90 0 0 la_oenb[120]
port 422 nsew signal input
flabel metal2 s 557326 -960 557438 480 0 FreeSans 448 90 0 0 la_oenb[121]
port 423 nsew signal input
flabel metal2 s 560822 -960 560934 480 0 FreeSans 448 90 0 0 la_oenb[122]
port 424 nsew signal input
flabel metal2 s 564410 -960 564522 480 0 FreeSans 448 90 0 0 la_oenb[123]
port 425 nsew signal input
flabel metal2 s 567998 -960 568110 480 0 FreeSans 448 90 0 0 la_oenb[124]
port 426 nsew signal input
flabel metal2 s 571494 -960 571606 480 0 FreeSans 448 90 0 0 la_oenb[125]
port 427 nsew signal input
flabel metal2 s 575082 -960 575194 480 0 FreeSans 448 90 0 0 la_oenb[126]
port 428 nsew signal input
flabel metal2 s 578578 -960 578690 480 0 FreeSans 448 90 0 0 la_oenb[127]
port 429 nsew signal input
flabel metal2 s 170742 -960 170854 480 0 FreeSans 448 90 0 0 la_oenb[12]
port 430 nsew signal input
flabel metal2 s 174238 -960 174350 480 0 FreeSans 448 90 0 0 la_oenb[13]
port 431 nsew signal input
flabel metal2 s 177826 -960 177938 480 0 FreeSans 448 90 0 0 la_oenb[14]
port 432 nsew signal input
flabel metal2 s 181414 -960 181526 480 0 FreeSans 448 90 0 0 la_oenb[15]
port 433 nsew signal input
flabel metal2 s 184910 -960 185022 480 0 FreeSans 448 90 0 0 la_oenb[16]
port 434 nsew signal input
flabel metal2 s 188498 -960 188610 480 0 FreeSans 448 90 0 0 la_oenb[17]
port 435 nsew signal input
flabel metal2 s 191994 -960 192106 480 0 FreeSans 448 90 0 0 la_oenb[18]
port 436 nsew signal input
flabel metal2 s 195582 -960 195694 480 0 FreeSans 448 90 0 0 la_oenb[19]
port 437 nsew signal input
flabel metal2 s 131734 -960 131846 480 0 FreeSans 448 90 0 0 la_oenb[1]
port 438 nsew signal input
flabel metal2 s 199078 -960 199190 480 0 FreeSans 448 90 0 0 la_oenb[20]
port 439 nsew signal input
flabel metal2 s 202666 -960 202778 480 0 FreeSans 448 90 0 0 la_oenb[21]
port 440 nsew signal input
flabel metal2 s 206162 -960 206274 480 0 FreeSans 448 90 0 0 la_oenb[22]
port 441 nsew signal input
flabel metal2 s 209750 -960 209862 480 0 FreeSans 448 90 0 0 la_oenb[23]
port 442 nsew signal input
flabel metal2 s 213338 -960 213450 480 0 FreeSans 448 90 0 0 la_oenb[24]
port 443 nsew signal input
flabel metal2 s 216834 -960 216946 480 0 FreeSans 448 90 0 0 la_oenb[25]
port 444 nsew signal input
flabel metal2 s 220422 -960 220534 480 0 FreeSans 448 90 0 0 la_oenb[26]
port 445 nsew signal input
flabel metal2 s 223918 -960 224030 480 0 FreeSans 448 90 0 0 la_oenb[27]
port 446 nsew signal input
flabel metal2 s 227506 -960 227618 480 0 FreeSans 448 90 0 0 la_oenb[28]
port 447 nsew signal input
flabel metal2 s 231002 -960 231114 480 0 FreeSans 448 90 0 0 la_oenb[29]
port 448 nsew signal input
flabel metal2 s 135230 -960 135342 480 0 FreeSans 448 90 0 0 la_oenb[2]
port 449 nsew signal input
flabel metal2 s 234590 -960 234702 480 0 FreeSans 448 90 0 0 la_oenb[30]
port 450 nsew signal input
flabel metal2 s 238086 -960 238198 480 0 FreeSans 448 90 0 0 la_oenb[31]
port 451 nsew signal input
flabel metal2 s 241674 -960 241786 480 0 FreeSans 448 90 0 0 la_oenb[32]
port 452 nsew signal input
flabel metal2 s 245170 -960 245282 480 0 FreeSans 448 90 0 0 la_oenb[33]
port 453 nsew signal input
flabel metal2 s 248758 -960 248870 480 0 FreeSans 448 90 0 0 la_oenb[34]
port 454 nsew signal input
flabel metal2 s 252346 -960 252458 480 0 FreeSans 448 90 0 0 la_oenb[35]
port 455 nsew signal input
flabel metal2 s 255842 -960 255954 480 0 FreeSans 448 90 0 0 la_oenb[36]
port 456 nsew signal input
flabel metal2 s 259430 -960 259542 480 0 FreeSans 448 90 0 0 la_oenb[37]
port 457 nsew signal input
flabel metal2 s 262926 -960 263038 480 0 FreeSans 448 90 0 0 la_oenb[38]
port 458 nsew signal input
flabel metal2 s 266514 -960 266626 480 0 FreeSans 448 90 0 0 la_oenb[39]
port 459 nsew signal input
flabel metal2 s 138818 -960 138930 480 0 FreeSans 448 90 0 0 la_oenb[3]
port 460 nsew signal input
flabel metal2 s 270010 -960 270122 480 0 FreeSans 448 90 0 0 la_oenb[40]
port 461 nsew signal input
flabel metal2 s 273598 -960 273710 480 0 FreeSans 448 90 0 0 la_oenb[41]
port 462 nsew signal input
flabel metal2 s 277094 -960 277206 480 0 FreeSans 448 90 0 0 la_oenb[42]
port 463 nsew signal input
flabel metal2 s 280682 -960 280794 480 0 FreeSans 448 90 0 0 la_oenb[43]
port 464 nsew signal input
flabel metal2 s 284270 -960 284382 480 0 FreeSans 448 90 0 0 la_oenb[44]
port 465 nsew signal input
flabel metal2 s 287766 -960 287878 480 0 FreeSans 448 90 0 0 la_oenb[45]
port 466 nsew signal input
flabel metal2 s 291354 -960 291466 480 0 FreeSans 448 90 0 0 la_oenb[46]
port 467 nsew signal input
flabel metal2 s 294850 -960 294962 480 0 FreeSans 448 90 0 0 la_oenb[47]
port 468 nsew signal input
flabel metal2 s 298438 -960 298550 480 0 FreeSans 448 90 0 0 la_oenb[48]
port 469 nsew signal input
flabel metal2 s 301934 -960 302046 480 0 FreeSans 448 90 0 0 la_oenb[49]
port 470 nsew signal input
flabel metal2 s 142406 -960 142518 480 0 FreeSans 448 90 0 0 la_oenb[4]
port 471 nsew signal input
flabel metal2 s 305522 -960 305634 480 0 FreeSans 448 90 0 0 la_oenb[50]
port 472 nsew signal input
flabel metal2 s 309018 -960 309130 480 0 FreeSans 448 90 0 0 la_oenb[51]
port 473 nsew signal input
flabel metal2 s 312606 -960 312718 480 0 FreeSans 448 90 0 0 la_oenb[52]
port 474 nsew signal input
flabel metal2 s 316194 -960 316306 480 0 FreeSans 448 90 0 0 la_oenb[53]
port 475 nsew signal input
flabel metal2 s 319690 -960 319802 480 0 FreeSans 448 90 0 0 la_oenb[54]
port 476 nsew signal input
flabel metal2 s 323278 -960 323390 480 0 FreeSans 448 90 0 0 la_oenb[55]
port 477 nsew signal input
flabel metal2 s 326774 -960 326886 480 0 FreeSans 448 90 0 0 la_oenb[56]
port 478 nsew signal input
flabel metal2 s 330362 -960 330474 480 0 FreeSans 448 90 0 0 la_oenb[57]
port 479 nsew signal input
flabel metal2 s 333858 -960 333970 480 0 FreeSans 448 90 0 0 la_oenb[58]
port 480 nsew signal input
flabel metal2 s 337446 -960 337558 480 0 FreeSans 448 90 0 0 la_oenb[59]
port 481 nsew signal input
flabel metal2 s 145902 -960 146014 480 0 FreeSans 448 90 0 0 la_oenb[5]
port 482 nsew signal input
flabel metal2 s 340942 -960 341054 480 0 FreeSans 448 90 0 0 la_oenb[60]
port 483 nsew signal input
flabel metal2 s 344530 -960 344642 480 0 FreeSans 448 90 0 0 la_oenb[61]
port 484 nsew signal input
flabel metal2 s 348026 -960 348138 480 0 FreeSans 448 90 0 0 la_oenb[62]
port 485 nsew signal input
flabel metal2 s 351614 -960 351726 480 0 FreeSans 448 90 0 0 la_oenb[63]
port 486 nsew signal input
flabel metal2 s 355202 -960 355314 480 0 FreeSans 448 90 0 0 la_oenb[64]
port 487 nsew signal input
flabel metal2 s 358698 -960 358810 480 0 FreeSans 448 90 0 0 la_oenb[65]
port 488 nsew signal input
flabel metal2 s 362286 -960 362398 480 0 FreeSans 448 90 0 0 la_oenb[66]
port 489 nsew signal input
flabel metal2 s 365782 -960 365894 480 0 FreeSans 448 90 0 0 la_oenb[67]
port 490 nsew signal input
flabel metal2 s 369370 -960 369482 480 0 FreeSans 448 90 0 0 la_oenb[68]
port 491 nsew signal input
flabel metal2 s 372866 -960 372978 480 0 FreeSans 448 90 0 0 la_oenb[69]
port 492 nsew signal input
flabel metal2 s 149490 -960 149602 480 0 FreeSans 448 90 0 0 la_oenb[6]
port 493 nsew signal input
flabel metal2 s 376454 -960 376566 480 0 FreeSans 448 90 0 0 la_oenb[70]
port 494 nsew signal input
flabel metal2 s 379950 -960 380062 480 0 FreeSans 448 90 0 0 la_oenb[71]
port 495 nsew signal input
flabel metal2 s 383538 -960 383650 480 0 FreeSans 448 90 0 0 la_oenb[72]
port 496 nsew signal input
flabel metal2 s 387126 -960 387238 480 0 FreeSans 448 90 0 0 la_oenb[73]
port 497 nsew signal input
flabel metal2 s 390622 -960 390734 480 0 FreeSans 448 90 0 0 la_oenb[74]
port 498 nsew signal input
flabel metal2 s 394210 -960 394322 480 0 FreeSans 448 90 0 0 la_oenb[75]
port 499 nsew signal input
flabel metal2 s 397706 -960 397818 480 0 FreeSans 448 90 0 0 la_oenb[76]
port 500 nsew signal input
flabel metal2 s 401294 -960 401406 480 0 FreeSans 448 90 0 0 la_oenb[77]
port 501 nsew signal input
flabel metal2 s 404790 -960 404902 480 0 FreeSans 448 90 0 0 la_oenb[78]
port 502 nsew signal input
flabel metal2 s 408378 -960 408490 480 0 FreeSans 448 90 0 0 la_oenb[79]
port 503 nsew signal input
flabel metal2 s 152986 -960 153098 480 0 FreeSans 448 90 0 0 la_oenb[7]
port 504 nsew signal input
flabel metal2 s 411874 -960 411986 480 0 FreeSans 448 90 0 0 la_oenb[80]
port 505 nsew signal input
flabel metal2 s 415462 -960 415574 480 0 FreeSans 448 90 0 0 la_oenb[81]
port 506 nsew signal input
flabel metal2 s 418958 -960 419070 480 0 FreeSans 448 90 0 0 la_oenb[82]
port 507 nsew signal input
flabel metal2 s 422546 -960 422658 480 0 FreeSans 448 90 0 0 la_oenb[83]
port 508 nsew signal input
flabel metal2 s 426134 -960 426246 480 0 FreeSans 448 90 0 0 la_oenb[84]
port 509 nsew signal input
flabel metal2 s 429630 -960 429742 480 0 FreeSans 448 90 0 0 la_oenb[85]
port 510 nsew signal input
flabel metal2 s 433218 -960 433330 480 0 FreeSans 448 90 0 0 la_oenb[86]
port 511 nsew signal input
flabel metal2 s 436714 -960 436826 480 0 FreeSans 448 90 0 0 la_oenb[87]
port 512 nsew signal input
flabel metal2 s 440302 -960 440414 480 0 FreeSans 448 90 0 0 la_oenb[88]
port 513 nsew signal input
flabel metal2 s 443798 -960 443910 480 0 FreeSans 448 90 0 0 la_oenb[89]
port 514 nsew signal input
flabel metal2 s 156574 -960 156686 480 0 FreeSans 448 90 0 0 la_oenb[8]
port 515 nsew signal input
flabel metal2 s 447386 -960 447498 480 0 FreeSans 448 90 0 0 la_oenb[90]
port 516 nsew signal input
flabel metal2 s 450882 -960 450994 480 0 FreeSans 448 90 0 0 la_oenb[91]
port 517 nsew signal input
flabel metal2 s 454470 -960 454582 480 0 FreeSans 448 90 0 0 la_oenb[92]
port 518 nsew signal input
flabel metal2 s 458058 -960 458170 480 0 FreeSans 448 90 0 0 la_oenb[93]
port 519 nsew signal input
flabel metal2 s 461554 -960 461666 480 0 FreeSans 448 90 0 0 la_oenb[94]
port 520 nsew signal input
flabel metal2 s 465142 -960 465254 480 0 FreeSans 448 90 0 0 la_oenb[95]
port 521 nsew signal input
flabel metal2 s 468638 -960 468750 480 0 FreeSans 448 90 0 0 la_oenb[96]
port 522 nsew signal input
flabel metal2 s 472226 -960 472338 480 0 FreeSans 448 90 0 0 la_oenb[97]
port 523 nsew signal input
flabel metal2 s 475722 -960 475834 480 0 FreeSans 448 90 0 0 la_oenb[98]
port 524 nsew signal input
flabel metal2 s 479310 -960 479422 480 0 FreeSans 448 90 0 0 la_oenb[99]
port 525 nsew signal input
flabel metal2 s 160070 -960 160182 480 0 FreeSans 448 90 0 0 la_oenb[9]
port 526 nsew signal input
flabel metal2 s 579774 -960 579886 480 0 FreeSans 448 90 0 0 user_clock2
port 527 nsew signal input
flabel metal2 s 580970 -960 581082 480 0 FreeSans 448 90 0 0 user_irq[0]
port 528 nsew signal tristate
flabel metal2 s 582166 -960 582278 480 0 FreeSans 448 90 0 0 user_irq[1]
port 529 nsew signal tristate
flabel metal2 s 583362 -960 583474 480 0 FreeSans 448 90 0 0 user_irq[2]
port 530 nsew signal tristate
flabel metal4 s -2006 -934 -1386 704870 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2006 -934 585930 -314 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2006 704250 585930 704870 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 585310 -934 585930 704870 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 1794 -7654 2414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 37794 -7654 38414 49367 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 37794 674393 38414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 73794 -7654 74414 49367 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 73794 674393 74414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 109794 -7654 110414 49367 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 109794 674393 110414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 145794 -7654 146414 49367 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 145794 674393 146414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 181794 -7654 182414 49367 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 181794 674393 182414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 217794 -7654 218414 49367 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 217794 674393 218414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 253794 -7654 254414 49367 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 253794 674393 254414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 289794 -7654 290414 49367 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 289794 674393 290414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 325794 -7654 326414 49367 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 325794 674393 326414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 361794 -7654 362414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 397794 -7654 398414 31919 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 397794 92137 398414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 433794 -7654 434414 31919 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 433794 157249 434414 422599 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 433794 442833 434414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 469794 -7654 470414 201919 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 469794 385580 470414 601103 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 469794 669073 470414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 505794 -7654 506414 82599 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 505794 139281 506414 201919 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 505794 259417 506414 601103 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 505794 669073 506414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 541794 -7654 542414 425068 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 541794 460836 542414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 577794 -7654 578414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 2866 592650 3486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 38866 592650 39486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 74866 592650 75486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 110866 592650 111486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 146866 592650 147486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 182866 592650 183486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 218866 592650 219486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 254866 592650 255486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 290866 592650 291486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 326866 592650 327486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 362866 592650 363486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 398866 592650 399486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 434866 592650 435486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 470866 592650 471486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 506866 592650 507486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 542866 592650 543486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 578866 592650 579486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 614866 592650 615486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 650866 592650 651486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 686866 592650 687486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s -3926 -2854 -3306 706790 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -3926 -2854 587850 -2234 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -3926 706170 587850 706790 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 587230 -2854 587850 706790 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 9234 -7654 9854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 45234 -7654 45854 49367 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 45234 674393 45854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 81234 -7654 81854 49367 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 81234 674393 81854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 117234 -7654 117854 49367 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 117234 674393 117854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 153234 -7654 153854 49367 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 153234 674393 153854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 189234 -7654 189854 49367 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 189234 674393 189854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 225234 -7654 225854 49367 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 225234 674393 225854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 261234 -7654 261854 49367 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 261234 674393 261854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 297234 -7654 297854 49367 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 297234 674393 297854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 333234 -7654 333854 49367 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 333234 674393 333854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 369234 -7654 369854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 405234 -7654 405854 30068 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 405234 104460 405854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 441234 -7654 441854 31919 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 441234 157249 441854 422599 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 441234 442833 441854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 477234 -7654 477854 201919 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 477234 259417 477854 322287 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 477234 384817 477854 601103 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 477234 669073 477854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 513234 -7654 513854 82599 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 513234 139281 513854 201919 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 513234 259417 513854 601103 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 513234 669073 513854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 549234 -7654 549854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 10306 592650 10926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 46306 592650 46926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 82306 592650 82926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 118306 592650 118926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 154306 592650 154926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 190306 592650 190926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 226306 592650 226926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 262306 592650 262926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 298306 592650 298926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 334306 592650 334926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 370306 592650 370926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 406306 592650 406926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 442306 592650 442926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 478306 592650 478926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 514306 592650 514926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 550306 592650 550926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 586306 592650 586926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 622306 592650 622926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 658306 592650 658926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 694306 592650 694926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s -5846 -4774 -5226 708710 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -5846 -4774 589770 -4154 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -5846 708090 589770 708710 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 589150 -4774 589770 708710 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 16674 -7654 17294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 52674 -7654 53294 49367 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 88674 -7654 89294 49367 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 124674 -7654 125294 49367 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 160674 -7654 161294 49367 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 196674 -7654 197294 49367 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 232674 -7654 233294 49367 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 268674 -7654 269294 49367 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 304674 -7654 305294 49367 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 340674 -7654 341294 49367 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 376674 -7654 377294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 412674 -7654 413294 31919 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 412674 92137 413294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 448674 -7654 449294 31919 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 448674 92137 449294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 484674 -7654 485294 201919 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 484674 259417 485294 322068 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 484674 385580 485294 500068 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 484674 517884 485294 601103 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 520674 -7654 521294 82599 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 520674 139281 521294 201919 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 520674 259417 521294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 556674 -7654 557294 360068 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 556674 377884 557294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 17746 592650 18366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 53746 592650 54366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 89746 592650 90366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 125746 592650 126366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 161746 592650 162366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 197746 592650 198366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 233746 592650 234366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 269746 592650 270366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 305746 592650 306366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 341746 592650 342366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 377746 592650 378366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 413746 592650 414366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 449746 592650 450366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 485746 592650 486366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 521746 592650 522366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 557746 592650 558366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 593746 592650 594366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 629746 592650 630366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 665746 592650 666366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s -7766 -6694 -7146 710630 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -7766 -6694 591690 -6074 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -7766 710010 591690 710630 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 591070 -6694 591690 710630 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 24114 -7654 24734 45068 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 60114 -7654 60734 49367 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 96114 -7654 96734 49367 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 132114 -7654 132734 49367 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 168114 -7654 168734 49367 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 204114 -7654 204734 49367 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 240114 -7654 240734 49367 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 276114 -7654 276734 49367 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 312114 -7654 312734 49367 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 348114 -7654 348734 49367 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 384114 -7654 384734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 420114 -7654 420734 31919 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 420114 92137 420734 127767 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 420114 157249 420734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 456114 -7654 456734 31919 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 456114 92137 456734 500068 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 456114 517884 456734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 492114 -7654 492734 82599 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 492114 259417 492734 322287 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 492114 384817 492734 601103 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 492114 669073 492734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 528114 -7654 528734 82599 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 528114 259417 528734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 564114 -7654 564734 360068 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 564114 377884 564734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 25186 592650 25806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 61186 592650 61806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 97186 592650 97806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 133186 592650 133806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 169186 592650 169806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 205186 592650 205806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 241186 592650 241806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 277186 592650 277806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 313186 592650 313806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 349186 592650 349806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 385186 592650 385806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 421186 592650 421806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 457186 592650 457806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 493186 592650 493806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 529186 592650 529806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 565186 592650 565806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 601186 592650 601806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 637186 592650 637806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 673186 592650 673806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s -6806 -5734 -6186 709670 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -6806 -5734 590730 -5114 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -6806 709050 590730 709670 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 590110 -5734 590730 709670 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 20394 -7654 21014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 56394 -7654 57014 49367 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 92394 -7654 93014 49367 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 128394 -7654 129014 49367 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 164394 -7654 165014 49367 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 200394 -7654 201014 49367 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 236394 -7654 237014 49367 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 272394 -7654 273014 49367 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 308394 -7654 309014 49367 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 344394 -7654 345014 49367 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 380394 -7654 381014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 416394 -7654 417014 31919 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 416394 92137 417014 127767 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 416394 157249 417014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 452394 -7654 453014 31919 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 452394 92137 453014 500068 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 452394 517884 453014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 488394 -7654 489014 82599 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 488394 139281 489014 201919 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 488394 259417 489014 322287 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 488394 453692 489014 500068 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 488394 517884 489014 601103 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 488394 669073 489014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 524394 -7654 525014 82599 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 524394 139281 525014 201919 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 524394 259417 525014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 560394 -7654 561014 30068 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 560394 51692 561014 360068 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 560394 377884 561014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 21466 592650 22086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 57466 592650 58086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 93466 592650 94086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 129466 592650 130086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 165466 592650 166086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 201466 592650 202086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 237466 592650 238086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 273466 592650 274086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 309466 592650 310086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 345466 592650 346086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 381466 592650 382086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 417466 592650 418086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 453466 592650 454086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 489466 592650 490086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 525466 592650 526086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 561466 592650 562086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 597466 592650 598086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 633466 592650 634086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 669466 592650 670086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s -8726 -7654 -8106 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 -7654 592650 -7034 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 710970 592650 711590 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 592030 -7654 592650 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 27834 -7654 28454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 63834 -7654 64454 49367 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 63834 674393 64454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 99834 -7654 100454 49367 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 99834 674393 100454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 135834 -7654 136454 49367 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 135834 674393 136454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 171834 -7654 172454 49367 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 171834 674393 172454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 207834 -7654 208454 49367 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 207834 674393 208454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 243834 -7654 244454 49367 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 243834 674393 244454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 279834 -7654 280454 49367 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 279834 674393 280454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 315834 -7654 316454 45068 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 351834 -7654 352454 49367 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 351834 674393 352454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 387834 -7654 388454 31919 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 387834 92137 388454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 423834 -7654 424454 31919 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 423834 92137 424454 127767 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 423834 157249 424454 420068 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 423834 444412 424454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 459834 -7654 460454 500068 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 459834 517884 460454 601103 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 459834 669073 460454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 495834 -7654 496454 82599 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 495834 259417 496454 322287 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 495834 384817 496454 601103 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 495834 669073 496454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 531834 -7654 532454 82599 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 531834 139281 532454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 567834 -7654 568454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 28906 592650 29526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 64906 592650 65526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 100906 592650 101526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 136906 592650 137526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 172906 592650 173526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 208906 592650 209526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 244906 592650 245526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 280906 592650 281526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 316906 592650 317526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 352906 592650 353526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 388906 592650 389526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 424906 592650 425526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 460906 592650 461526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 496906 592650 497526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 532906 592650 533526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 568906 592650 569526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 604906 592650 605526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 640906 592650 641526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 676906 592650 677526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s -2966 -1894 -2346 705830 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -2966 -1894 586890 -1274 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -2966 705210 586890 705830 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 586270 -1894 586890 705830 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 5514 -7654 6134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 41514 -7654 42134 49367 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 41514 674393 42134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 77514 -7654 78134 49367 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 77514 674393 78134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 113514 -7654 114134 49367 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 113514 674393 114134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 149514 -7654 150134 49367 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 149514 674393 150134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 185514 -7654 186134 49367 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 185514 674393 186134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 221514 -7654 222134 49367 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 221514 674393 222134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 257514 -7654 258134 49367 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 257514 674393 258134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 293514 -7654 294134 49367 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 293514 674393 294134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 329514 -7654 330134 49367 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 329514 674393 330134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 365514 -7654 366134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 401514 -7654 402134 31919 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 401514 92137 402134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 437514 -7654 438134 31919 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 437514 157249 438134 420068 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 437514 444412 438134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 473514 -7654 474134 201919 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 473514 453692 474134 601103 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 473514 669073 474134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 509514 -7654 510134 82599 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 509514 139281 510134 201919 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 509514 259417 510134 601103 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 509514 669073 510134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 545514 -7654 546134 30068 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 545514 51692 546134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 581514 -7654 582134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 6586 592650 7206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 42586 592650 43206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 78586 592650 79206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 114586 592650 115206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 150586 592650 151206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 186586 592650 187206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 222586 592650 223206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 258586 592650 259206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 294586 592650 295206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 330586 592650 331206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 366586 592650 367206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 402586 592650 403206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 438586 592650 439206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 474586 592650 475206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 510586 592650 511206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 546586 592650 547206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 582586 592650 583206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 618586 592650 619206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 654586 592650 655206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 690586 592650 691206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s -4886 -3814 -4266 707750 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -4886 -3814 588810 -3194 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -4886 707130 588810 707750 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 588190 -3814 588810 707750 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 12954 -7654 13574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 48954 -7654 49574 49367 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 48954 674393 49574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 84954 -7654 85574 49367 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 84954 674393 85574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 120954 -7654 121574 49367 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 120954 674393 121574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 156954 -7654 157574 49367 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 156954 674393 157574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 192954 -7654 193574 45068 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 192954 684676 193574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 228954 -7654 229574 49367 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 228954 674393 229574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 264954 -7654 265574 49367 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 264954 674393 265574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 300954 -7654 301574 45068 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 300954 684676 301574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 336954 -7654 337574 49367 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 336954 674393 337574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 372954 -7654 373574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 408954 -7654 409574 31919 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 408954 92137 409574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 444954 -7654 445574 31919 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 444954 159644 445574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 480954 -7654 481574 201919 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 480954 259417 481574 322287 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 480954 453692 481574 601103 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 480954 669073 481574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 516954 -7654 517574 82599 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 516954 139281 517574 201919 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 516954 259417 517574 601103 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 516954 669073 517574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 552954 -7654 553574 30068 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 552954 51692 553574 360068 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 552954 377884 553574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 14026 592650 14646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 50026 592650 50646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 86026 592650 86646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 122026 592650 122646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 158026 592650 158646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 194026 592650 194646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 230026 592650 230646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 266026 592650 266646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 302026 592650 302646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 338026 592650 338646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 374026 592650 374646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 410026 592650 410646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 446026 592650 446646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 482026 592650 482646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 518026 592650 518646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 554026 592650 554646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 590026 592650 590646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 626026 592650 626646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 662026 592650 662646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 698026 592650 698646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal2 s 542 -960 654 480 0 FreeSans 448 90 0 0 wb_clk_i
port 539 nsew signal input
flabel metal2 s 1646 -960 1758 480 0 FreeSans 448 90 0 0 wb_rst_i
port 540 nsew signal input
flabel metal2 s 2842 -960 2954 480 0 FreeSans 448 90 0 0 wbs_ack_o
port 541 nsew signal tristate
flabel metal2 s 7626 -960 7738 480 0 FreeSans 448 90 0 0 wbs_adr_i[0]
port 542 nsew signal input
flabel metal2 s 47830 -960 47942 480 0 FreeSans 448 90 0 0 wbs_adr_i[10]
port 543 nsew signal input
flabel metal2 s 51326 -960 51438 480 0 FreeSans 448 90 0 0 wbs_adr_i[11]
port 544 nsew signal input
flabel metal2 s 54914 -960 55026 480 0 FreeSans 448 90 0 0 wbs_adr_i[12]
port 545 nsew signal input
flabel metal2 s 58410 -960 58522 480 0 FreeSans 448 90 0 0 wbs_adr_i[13]
port 546 nsew signal input
flabel metal2 s 61998 -960 62110 480 0 FreeSans 448 90 0 0 wbs_adr_i[14]
port 547 nsew signal input
flabel metal2 s 65494 -960 65606 480 0 FreeSans 448 90 0 0 wbs_adr_i[15]
port 548 nsew signal input
flabel metal2 s 69082 -960 69194 480 0 FreeSans 448 90 0 0 wbs_adr_i[16]
port 549 nsew signal input
flabel metal2 s 72578 -960 72690 480 0 FreeSans 448 90 0 0 wbs_adr_i[17]
port 550 nsew signal input
flabel metal2 s 76166 -960 76278 480 0 FreeSans 448 90 0 0 wbs_adr_i[18]
port 551 nsew signal input
flabel metal2 s 79662 -960 79774 480 0 FreeSans 448 90 0 0 wbs_adr_i[19]
port 552 nsew signal input
flabel metal2 s 12318 -960 12430 480 0 FreeSans 448 90 0 0 wbs_adr_i[1]
port 553 nsew signal input
flabel metal2 s 83250 -960 83362 480 0 FreeSans 448 90 0 0 wbs_adr_i[20]
port 554 nsew signal input
flabel metal2 s 86838 -960 86950 480 0 FreeSans 448 90 0 0 wbs_adr_i[21]
port 555 nsew signal input
flabel metal2 s 90334 -960 90446 480 0 FreeSans 448 90 0 0 wbs_adr_i[22]
port 556 nsew signal input
flabel metal2 s 93922 -960 94034 480 0 FreeSans 448 90 0 0 wbs_adr_i[23]
port 557 nsew signal input
flabel metal2 s 97418 -960 97530 480 0 FreeSans 448 90 0 0 wbs_adr_i[24]
port 558 nsew signal input
flabel metal2 s 101006 -960 101118 480 0 FreeSans 448 90 0 0 wbs_adr_i[25]
port 559 nsew signal input
flabel metal2 s 104502 -960 104614 480 0 FreeSans 448 90 0 0 wbs_adr_i[26]
port 560 nsew signal input
flabel metal2 s 108090 -960 108202 480 0 FreeSans 448 90 0 0 wbs_adr_i[27]
port 561 nsew signal input
flabel metal2 s 111586 -960 111698 480 0 FreeSans 448 90 0 0 wbs_adr_i[28]
port 562 nsew signal input
flabel metal2 s 115174 -960 115286 480 0 FreeSans 448 90 0 0 wbs_adr_i[29]
port 563 nsew signal input
flabel metal2 s 17010 -960 17122 480 0 FreeSans 448 90 0 0 wbs_adr_i[2]
port 564 nsew signal input
flabel metal2 s 118762 -960 118874 480 0 FreeSans 448 90 0 0 wbs_adr_i[30]
port 565 nsew signal input
flabel metal2 s 122258 -960 122370 480 0 FreeSans 448 90 0 0 wbs_adr_i[31]
port 566 nsew signal input
flabel metal2 s 21794 -960 21906 480 0 FreeSans 448 90 0 0 wbs_adr_i[3]
port 567 nsew signal input
flabel metal2 s 26486 -960 26598 480 0 FreeSans 448 90 0 0 wbs_adr_i[4]
port 568 nsew signal input
flabel metal2 s 30074 -960 30186 480 0 FreeSans 448 90 0 0 wbs_adr_i[5]
port 569 nsew signal input
flabel metal2 s 33570 -960 33682 480 0 FreeSans 448 90 0 0 wbs_adr_i[6]
port 570 nsew signal input
flabel metal2 s 37158 -960 37270 480 0 FreeSans 448 90 0 0 wbs_adr_i[7]
port 571 nsew signal input
flabel metal2 s 40654 -960 40766 480 0 FreeSans 448 90 0 0 wbs_adr_i[8]
port 572 nsew signal input
flabel metal2 s 44242 -960 44354 480 0 FreeSans 448 90 0 0 wbs_adr_i[9]
port 573 nsew signal input
flabel metal2 s 4038 -960 4150 480 0 FreeSans 448 90 0 0 wbs_cyc_i
port 574 nsew signal input
flabel metal2 s 8730 -960 8842 480 0 FreeSans 448 90 0 0 wbs_dat_i[0]
port 575 nsew signal input
flabel metal2 s 48934 -960 49046 480 0 FreeSans 448 90 0 0 wbs_dat_i[10]
port 576 nsew signal input
flabel metal2 s 52522 -960 52634 480 0 FreeSans 448 90 0 0 wbs_dat_i[11]
port 577 nsew signal input
flabel metal2 s 56018 -960 56130 480 0 FreeSans 448 90 0 0 wbs_dat_i[12]
port 578 nsew signal input
flabel metal2 s 59606 -960 59718 480 0 FreeSans 448 90 0 0 wbs_dat_i[13]
port 579 nsew signal input
flabel metal2 s 63194 -960 63306 480 0 FreeSans 448 90 0 0 wbs_dat_i[14]
port 580 nsew signal input
flabel metal2 s 66690 -960 66802 480 0 FreeSans 448 90 0 0 wbs_dat_i[15]
port 581 nsew signal input
flabel metal2 s 70278 -960 70390 480 0 FreeSans 448 90 0 0 wbs_dat_i[16]
port 582 nsew signal input
flabel metal2 s 73774 -960 73886 480 0 FreeSans 448 90 0 0 wbs_dat_i[17]
port 583 nsew signal input
flabel metal2 s 77362 -960 77474 480 0 FreeSans 448 90 0 0 wbs_dat_i[18]
port 584 nsew signal input
flabel metal2 s 80858 -960 80970 480 0 FreeSans 448 90 0 0 wbs_dat_i[19]
port 585 nsew signal input
flabel metal2 s 13514 -960 13626 480 0 FreeSans 448 90 0 0 wbs_dat_i[1]
port 586 nsew signal input
flabel metal2 s 84446 -960 84558 480 0 FreeSans 448 90 0 0 wbs_dat_i[20]
port 587 nsew signal input
flabel metal2 s 87942 -960 88054 480 0 FreeSans 448 90 0 0 wbs_dat_i[21]
port 588 nsew signal input
flabel metal2 s 91530 -960 91642 480 0 FreeSans 448 90 0 0 wbs_dat_i[22]
port 589 nsew signal input
flabel metal2 s 95118 -960 95230 480 0 FreeSans 448 90 0 0 wbs_dat_i[23]
port 590 nsew signal input
flabel metal2 s 98614 -960 98726 480 0 FreeSans 448 90 0 0 wbs_dat_i[24]
port 591 nsew signal input
flabel metal2 s 102202 -960 102314 480 0 FreeSans 448 90 0 0 wbs_dat_i[25]
port 592 nsew signal input
flabel metal2 s 105698 -960 105810 480 0 FreeSans 448 90 0 0 wbs_dat_i[26]
port 593 nsew signal input
flabel metal2 s 109286 -960 109398 480 0 FreeSans 448 90 0 0 wbs_dat_i[27]
port 594 nsew signal input
flabel metal2 s 112782 -960 112894 480 0 FreeSans 448 90 0 0 wbs_dat_i[28]
port 595 nsew signal input
flabel metal2 s 116370 -960 116482 480 0 FreeSans 448 90 0 0 wbs_dat_i[29]
port 596 nsew signal input
flabel metal2 s 18206 -960 18318 480 0 FreeSans 448 90 0 0 wbs_dat_i[2]
port 597 nsew signal input
flabel metal2 s 119866 -960 119978 480 0 FreeSans 448 90 0 0 wbs_dat_i[30]
port 598 nsew signal input
flabel metal2 s 123454 -960 123566 480 0 FreeSans 448 90 0 0 wbs_dat_i[31]
port 599 nsew signal input
flabel metal2 s 22990 -960 23102 480 0 FreeSans 448 90 0 0 wbs_dat_i[3]
port 600 nsew signal input
flabel metal2 s 27682 -960 27794 480 0 FreeSans 448 90 0 0 wbs_dat_i[4]
port 601 nsew signal input
flabel metal2 s 31270 -960 31382 480 0 FreeSans 448 90 0 0 wbs_dat_i[5]
port 602 nsew signal input
flabel metal2 s 34766 -960 34878 480 0 FreeSans 448 90 0 0 wbs_dat_i[6]
port 603 nsew signal input
flabel metal2 s 38354 -960 38466 480 0 FreeSans 448 90 0 0 wbs_dat_i[7]
port 604 nsew signal input
flabel metal2 s 41850 -960 41962 480 0 FreeSans 448 90 0 0 wbs_dat_i[8]
port 605 nsew signal input
flabel metal2 s 45438 -960 45550 480 0 FreeSans 448 90 0 0 wbs_dat_i[9]
port 606 nsew signal input
flabel metal2 s 9926 -960 10038 480 0 FreeSans 448 90 0 0 wbs_dat_o[0]
port 607 nsew signal tristate
flabel metal2 s 50130 -960 50242 480 0 FreeSans 448 90 0 0 wbs_dat_o[10]
port 608 nsew signal tristate
flabel metal2 s 53718 -960 53830 480 0 FreeSans 448 90 0 0 wbs_dat_o[11]
port 609 nsew signal tristate
flabel metal2 s 57214 -960 57326 480 0 FreeSans 448 90 0 0 wbs_dat_o[12]
port 610 nsew signal tristate
flabel metal2 s 60802 -960 60914 480 0 FreeSans 448 90 0 0 wbs_dat_o[13]
port 611 nsew signal tristate
flabel metal2 s 64298 -960 64410 480 0 FreeSans 448 90 0 0 wbs_dat_o[14]
port 612 nsew signal tristate
flabel metal2 s 67886 -960 67998 480 0 FreeSans 448 90 0 0 wbs_dat_o[15]
port 613 nsew signal tristate
flabel metal2 s 71474 -960 71586 480 0 FreeSans 448 90 0 0 wbs_dat_o[16]
port 614 nsew signal tristate
flabel metal2 s 74970 -960 75082 480 0 FreeSans 448 90 0 0 wbs_dat_o[17]
port 615 nsew signal tristate
flabel metal2 s 78558 -960 78670 480 0 FreeSans 448 90 0 0 wbs_dat_o[18]
port 616 nsew signal tristate
flabel metal2 s 82054 -960 82166 480 0 FreeSans 448 90 0 0 wbs_dat_o[19]
port 617 nsew signal tristate
flabel metal2 s 14710 -960 14822 480 0 FreeSans 448 90 0 0 wbs_dat_o[1]
port 618 nsew signal tristate
flabel metal2 s 85642 -960 85754 480 0 FreeSans 448 90 0 0 wbs_dat_o[20]
port 619 nsew signal tristate
flabel metal2 s 89138 -960 89250 480 0 FreeSans 448 90 0 0 wbs_dat_o[21]
port 620 nsew signal tristate
flabel metal2 s 92726 -960 92838 480 0 FreeSans 448 90 0 0 wbs_dat_o[22]
port 621 nsew signal tristate
flabel metal2 s 96222 -960 96334 480 0 FreeSans 448 90 0 0 wbs_dat_o[23]
port 622 nsew signal tristate
flabel metal2 s 99810 -960 99922 480 0 FreeSans 448 90 0 0 wbs_dat_o[24]
port 623 nsew signal tristate
flabel metal2 s 103306 -960 103418 480 0 FreeSans 448 90 0 0 wbs_dat_o[25]
port 624 nsew signal tristate
flabel metal2 s 106894 -960 107006 480 0 FreeSans 448 90 0 0 wbs_dat_o[26]
port 625 nsew signal tristate
flabel metal2 s 110482 -960 110594 480 0 FreeSans 448 90 0 0 wbs_dat_o[27]
port 626 nsew signal tristate
flabel metal2 s 113978 -960 114090 480 0 FreeSans 448 90 0 0 wbs_dat_o[28]
port 627 nsew signal tristate
flabel metal2 s 117566 -960 117678 480 0 FreeSans 448 90 0 0 wbs_dat_o[29]
port 628 nsew signal tristate
flabel metal2 s 19402 -960 19514 480 0 FreeSans 448 90 0 0 wbs_dat_o[2]
port 629 nsew signal tristate
flabel metal2 s 121062 -960 121174 480 0 FreeSans 448 90 0 0 wbs_dat_o[30]
port 630 nsew signal tristate
flabel metal2 s 124650 -960 124762 480 0 FreeSans 448 90 0 0 wbs_dat_o[31]
port 631 nsew signal tristate
flabel metal2 s 24186 -960 24298 480 0 FreeSans 448 90 0 0 wbs_dat_o[3]
port 632 nsew signal tristate
flabel metal2 s 28878 -960 28990 480 0 FreeSans 448 90 0 0 wbs_dat_o[4]
port 633 nsew signal tristate
flabel metal2 s 32374 -960 32486 480 0 FreeSans 448 90 0 0 wbs_dat_o[5]
port 634 nsew signal tristate
flabel metal2 s 35962 -960 36074 480 0 FreeSans 448 90 0 0 wbs_dat_o[6]
port 635 nsew signal tristate
flabel metal2 s 39550 -960 39662 480 0 FreeSans 448 90 0 0 wbs_dat_o[7]
port 636 nsew signal tristate
flabel metal2 s 43046 -960 43158 480 0 FreeSans 448 90 0 0 wbs_dat_o[8]
port 637 nsew signal tristate
flabel metal2 s 46634 -960 46746 480 0 FreeSans 448 90 0 0 wbs_dat_o[9]
port 638 nsew signal tristate
flabel metal2 s 11122 -960 11234 480 0 FreeSans 448 90 0 0 wbs_sel_i[0]
port 639 nsew signal input
flabel metal2 s 15906 -960 16018 480 0 FreeSans 448 90 0 0 wbs_sel_i[1]
port 640 nsew signal input
flabel metal2 s 20598 -960 20710 480 0 FreeSans 448 90 0 0 wbs_sel_i[2]
port 641 nsew signal input
flabel metal2 s 25290 -960 25402 480 0 FreeSans 448 90 0 0 wbs_sel_i[3]
port 642 nsew signal input
flabel metal2 s 5234 -960 5346 480 0 FreeSans 448 90 0 0 wbs_stb_i
port 643 nsew signal input
flabel metal2 s 6430 -960 6542 480 0 FreeSans 448 90 0 0 wbs_we_i
port 644 nsew signal input
rlabel via4 451808 75336 451808 75336 0 vccd1
rlabel via4 333704 46776 333704 46776 0 vccd2
rlabel via4 521144 666216 521144 666216 0 vdda1
rlabel via4 456584 97656 456584 97656 0 vdda2
rlabel via4 452864 93936 452864 93936 0 vssa1
rlabel via4 460304 101376 460304 101376 0 vssa2
rlabel via4 436448 79056 436448 79056 0 vssd1
rlabel via4 481424 122496 481424 122496 0 vssd2
rlabel metal2 422510 446138 422510 446138 0 design_clk
rlabel metal2 411960 159868 411960 159868 0 dsi_all\[0\]
rlabel metal2 448362 161058 448362 161058 0 dsi_all\[10\]
rlabel metal2 447166 172142 447166 172142 0 dsi_all\[11\]
rlabel metal3 449152 332180 449152 332180 0 dsi_all\[12\]
rlabel metal2 447166 332741 447166 332741 0 dsi_all\[13\]
rlabel metal2 447258 333115 447258 333115 0 dsi_all\[14\]
rlabel metal2 447166 334101 447166 334101 0 dsi_all\[15\]
rlabel metal1 445464 334050 445464 334050 0 dsi_all\[16\]
rlabel metal2 447166 335461 447166 335461 0 dsi_all\[17\]
rlabel metal1 445464 335682 445464 335682 0 dsi_all\[18\]
rlabel metal2 447258 336515 447258 336515 0 dsi_all\[19\]
rlabel metal3 449980 503472 449980 503472 0 dsi_all\[1\]
rlabel metal2 447166 337059 447166 337059 0 dsi_all\[20\]
rlabel metal2 447166 338249 447166 338249 0 dsi_all\[21\]
rlabel metal2 447258 338555 447258 338555 0 dsi_all\[22\]
rlabel metal2 447166 339609 447166 339609 0 dsi_all\[23\]
rlabel metal2 447258 339915 447258 339915 0 dsi_all\[24\]
rlabel via2 447166 341003 447166 341003 0 dsi_all\[25\]
rlabel metal2 447258 341309 447258 341309 0 dsi_all\[26\]
rlabel metal3 449796 342380 449796 342380 0 dsi_all\[27\]
rlabel metal3 450156 505531 450156 505531 0 dsi_all\[2\]
rlabel metal3 450087 326196 450087 326196 0 dsi_all\[3\]
rlabel metal2 425208 159868 425208 159868 0 dsi_all\[4\]
rlabel metal2 428184 159732 428184 159732 0 dsi_all\[5\]
rlabel metal2 431496 159460 431496 159460 0 dsi_all\[6\]
rlabel metal3 450156 328629 450156 328629 0 dsi_all\[7\]
rlabel metal3 448646 329460 448646 329460 0 dsi_all\[8\]
rlabel metal3 448646 330140 448646 330140 0 dsi_all\[9\]
rlabel metal2 487370 298054 487370 298054 0 dso_6502\[0\]
rlabel via2 452042 135133 452042 135133 0 dso_6502\[10\]
rlabel via2 451582 136493 451582 136493 0 dso_6502\[11\]
rlabel via2 452594 137853 452594 137853 0 dso_6502\[12\]
rlabel via2 451582 139213 451582 139213 0 dso_6502\[13\]
rlabel metal2 452594 140641 452594 140641 0 dso_6502\[14\]
rlabel via2 452594 141933 452594 141933 0 dso_6502\[15\]
rlabel metal2 452594 143361 452594 143361 0 dso_6502\[16\]
rlabel metal1 474260 276726 474260 276726 0 dso_6502\[17\]
rlabel metal2 451858 146115 451858 146115 0 dso_6502\[18\]
rlabel via2 452594 147373 452594 147373 0 dso_6502\[19\]
rlabel metal2 487646 297340 487646 297340 0 dso_6502\[1\]
rlabel metal3 450930 148716 450930 148716 0 dso_6502\[20\]
rlabel metal3 451114 150076 451114 150076 0 dso_6502\[21\]
rlabel via2 452594 151453 452594 151453 0 dso_6502\[22\]
rlabel metal2 452502 152881 452502 152881 0 dso_6502\[23\]
rlabel metal2 452502 154309 452502 154309 0 dso_6502\[24\]
rlabel metal3 451022 155516 451022 155516 0 dso_6502\[25\]
rlabel metal2 451766 157097 451766 157097 0 dso_6502\[26\]
rlabel metal2 487922 304378 487922 304378 0 dso_6502\[2\]
rlabel metal2 488198 298734 488198 298734 0 dso_6502\[3\]
rlabel metal2 488474 315972 488474 315972 0 dso_6502\[4\]
rlabel metal2 488750 315292 488750 315292 0 dso_6502\[5\]
rlabel metal2 489026 319474 489026 319474 0 dso_6502\[6\]
rlabel metal2 489302 295266 489302 295266 0 dso_6502\[7\]
rlabel metal2 489578 318726 489578 318726 0 dso_6502\[8\]
rlabel metal2 489854 296660 489854 296660 0 dso_6502\[9\]
rlabel metal2 503785 385900 503785 385900 0 dso_LCD\[0\]
rlabel metal2 504337 385900 504337 385900 0 dso_LCD\[1\]
rlabel metal2 505310 387862 505310 387862 0 dso_LCD\[2\]
rlabel metal2 506046 388576 506046 388576 0 dso_LCD\[3\]
rlabel metal2 506683 385900 506683 385900 0 dso_LCD\[4\]
rlabel metal2 507327 385900 507327 385900 0 dso_LCD\[5\]
rlabel metal2 508063 385900 508063 385900 0 dso_LCD\[6\]
rlabel metal2 508753 385900 508753 385900 0 dso_LCD\[7\]
rlabel metal3 540492 82348 540492 82348 0 dso_as1802\[0\]
rlabel metal3 540584 102748 540584 102748 0 dso_as1802\[10\]
rlabel metal3 540630 104788 540630 104788 0 dso_as1802\[11\]
rlabel metal3 540676 106828 540676 106828 0 dso_as1802\[12\]
rlabel metal3 539948 108785 539948 108785 0 dso_as1802\[13\]
rlabel metal3 540538 110908 540538 110908 0 dso_as1802\[14\]
rlabel metal3 539948 112865 539948 112865 0 dso_as1802\[15\]
rlabel metal3 540722 114988 540722 114988 0 dso_as1802\[16\]
rlabel via2 539925 117300 539925 117300 0 dso_as1802\[17\]
rlabel metal3 541550 119068 541550 119068 0 dso_as1802\[18\]
rlabel metal3 541320 121108 541320 121108 0 dso_as1802\[19\]
rlabel metal3 541412 84388 541412 84388 0 dso_as1802\[1\]
rlabel metal2 500342 318080 500342 318080 0 dso_as1802\[20\]
rlabel metal2 500526 295693 500526 295693 0 dso_as1802\[21\]
rlabel metal2 500894 301488 500894 301488 0 dso_as1802\[22\]
rlabel metal3 538959 137836 538959 137836 0 dso_as1802\[23\]
rlabel metal2 501446 302882 501446 302882 0 dso_as1802\[24\]
rlabel metal4 538844 137700 538844 137700 0 dso_as1802\[25\]
rlabel metal2 538936 137836 538936 137836 0 dso_as1802\[26\]
rlabel metal3 541458 86428 541458 86428 0 dso_as1802\[2\]
rlabel metal3 541596 88468 541596 88468 0 dso_as1802\[3\]
rlabel metal3 541228 90508 541228 90508 0 dso_as1802\[4\]
rlabel metal3 541504 92548 541504 92548 0 dso_as1802\[5\]
rlabel via2 539603 95132 539603 95132 0 dso_as1802\[6\]
rlabel via2 539741 97172 539741 97172 0 dso_as1802\[7\]
rlabel via2 539787 99212 539787 99212 0 dso_as1802\[8\]
rlabel metal3 541274 100708 541274 100708 0 dso_as1802\[9\]
rlabel metal2 463121 385900 463121 385900 0 dso_as2650\[0\]
rlabel metal2 470665 385900 470665 385900 0 dso_as2650\[10\]
rlabel metal2 471217 385900 471217 385900 0 dso_as2650\[11\]
rlabel metal2 472190 387471 472190 387471 0 dso_as2650\[12\]
rlabel metal2 472926 387403 472926 387403 0 dso_as2650\[13\]
rlabel metal2 469982 453628 469982 453628 0 dso_as2650\[14\]
rlabel metal3 459655 637908 459655 637908 0 dso_as2650\[15\]
rlabel metal3 459701 640356 459701 640356 0 dso_as2650\[16\]
rlabel metal2 469890 494258 469890 494258 0 dso_as2650\[17\]
rlabel metal2 468510 493544 468510 493544 0 dso_as2650\[18\]
rlabel metal2 477342 387471 477342 387471 0 dso_as2650\[19\]
rlabel metal2 463949 385900 463949 385900 0 dso_as2650\[1\]
rlabel metal2 461610 494564 461610 494564 0 dso_as2650\[20\]
rlabel metal2 461702 494428 461702 494428 0 dso_as2650\[21\]
rlabel metal3 459801 655656 459801 655656 0 dso_as2650\[22\]
rlabel metal2 480286 387352 480286 387352 0 dso_as2650\[23\]
rlabel metal1 467636 388926 467636 388926 0 dso_as2650\[24\]
rlabel metal1 468234 388722 468234 388722 0 dso_as2650\[25\]
rlabel metal2 482494 387182 482494 387182 0 dso_as2650\[26\]
rlabel metal2 464639 385900 464639 385900 0 dso_as2650\[2\]
rlabel metal2 465329 385900 465329 385900 0 dso_as2650\[3\]
rlabel metal2 466065 385900 466065 385900 0 dso_as2650\[4\]
rlabel metal2 466801 385900 466801 385900 0 dso_as2650\[5\]
rlabel metal2 467583 385900 467583 385900 0 dso_as2650\[6\]
rlabel metal2 468273 385900 468273 385900 0 dso_as2650\[7\]
rlabel metal2 469246 387284 469246 387284 0 dso_as2650\[8\]
rlabel metal2 469982 387148 469982 387148 0 dso_as2650\[9\]
rlabel metal2 409906 367778 409906 367778 0 dso_as512512512\[0\]
rlabel metal2 447258 372045 447258 372045 0 dso_as512512512\[10\]
rlabel metal2 447166 372419 447166 372419 0 dso_as512512512\[11\]
rlabel metal2 447258 373439 447258 373439 0 dso_as512512512\[12\]
rlabel metal2 447166 373813 447166 373813 0 dso_as512512512\[13\]
rlabel metal2 447258 374799 447258 374799 0 dso_as512512512\[14\]
rlabel metal2 447166 375173 447166 375173 0 dso_as512512512\[15\]
rlabel metal2 367770 461584 367770 461584 0 dso_as512512512\[16\]
rlabel metal2 370530 467092 370530 467092 0 dso_as512512512\[17\]
rlabel metal2 447258 377587 447258 377587 0 dso_as512512512\[18\]
rlabel metal2 371910 478856 371910 478856 0 dso_as512512512\[19\]
rlabel metal1 445556 365602 445556 365602 0 dso_as512512512\[1\]
rlabel metal2 407790 485044 407790 485044 0 dso_as512512512\[20\]
rlabel metal2 447166 379287 447166 379287 0 dso_as512512512\[21\]
rlabel metal2 406410 496774 406410 496774 0 dso_as512512512\[22\]
rlabel metal2 447166 380647 447166 380647 0 dso_as512512512\[23\]
rlabel metal2 403650 508470 403650 508470 0 dso_as512512512\[24\]
rlabel metal2 447166 382007 447166 382007 0 dso_as512512512\[25\]
rlabel metal2 447258 383061 447258 383061 0 dso_as512512512\[26\]
rlabel metal2 447166 383367 447166 383367 0 dso_as512512512\[27\]
rlabel metal1 445510 366962 445510 366962 0 dso_as512512512\[2\]
rlabel metal2 447166 366945 447166 366945 0 dso_as512512512\[3\]
rlabel metal1 445418 368458 445418 368458 0 dso_as512512512\[4\]
rlabel metal1 444774 368390 444774 368390 0 dso_as512512512\[5\]
rlabel metal2 447258 369359 447258 369359 0 dso_as512512512\[6\]
rlabel metal2 447166 369665 447166 369665 0 dso_as512512512\[7\]
rlabel metal2 447258 370719 447258 370719 0 dso_as512512512\[8\]
rlabel metal2 447166 371025 447166 371025 0 dso_as512512512\[9\]
rlabel metal2 483421 385900 483421 385900 0 dso_as5401\[0\]
rlabel metal2 490590 389256 490590 389256 0 dso_as5401\[10\]
rlabel metal2 491517 385900 491517 385900 0 dso_as5401\[11\]
rlabel metal2 492062 387896 492062 387896 0 dso_as5401\[12\]
rlabel metal2 492989 385900 492989 385900 0 dso_as5401\[13\]
rlabel metal2 539067 425068 539067 425068 0 dso_as5401\[14\]
rlabel metal2 540355 425068 540355 425068 0 dso_as5401\[15\]
rlabel metal2 541834 422630 541834 422630 0 dso_as5401\[16\]
rlabel metal2 542931 425068 542931 425068 0 dso_as5401\[17\]
rlabel metal2 544219 425068 544219 425068 0 dso_as5401\[18\]
rlabel metal2 545698 424092 545698 424092 0 dso_as5401\[19\]
rlabel metal2 484157 385900 484157 385900 0 dso_as5401\[1\]
rlabel metal2 546795 425068 546795 425068 0 dso_as5401\[20\]
rlabel metal2 498877 385900 498877 385900 0 dso_as5401\[21\]
rlabel metal2 522330 406062 522330 406062 0 dso_as5401\[22\]
rlabel metal2 500349 385900 500349 385900 0 dso_as5401\[23\]
rlabel metal2 500894 387318 500894 387318 0 dso_as5401\[24\]
rlabel metal2 501821 385900 501821 385900 0 dso_as5401\[25\]
rlabel metal2 502366 387420 502366 387420 0 dso_as5401\[26\]
rlabel metal2 484702 387352 484702 387352 0 dso_as5401\[2\]
rlabel metal2 485438 387250 485438 387250 0 dso_as5401\[3\]
rlabel metal2 486319 385900 486319 385900 0 dso_as5401\[4\]
rlabel metal2 486910 389607 486910 389607 0 dso_as5401\[5\]
rlabel metal2 487837 385900 487837 385900 0 dso_as5401\[6\]
rlabel metal2 488382 387182 488382 387182 0 dso_as5401\[7\]
rlabel metal2 489309 385900 489309 385900 0 dso_as5401\[8\]
rlabel metal2 489854 387216 489854 387216 0 dso_as5401\[9\]
rlabel metal2 522330 369002 522330 369002 0 dso_counter\[0\]
rlabel metal2 565294 360009 565294 360009 0 dso_counter\[10\]
rlabel via1 566766 360077 566766 360077 0 dso_counter\[11\]
rlabel metal2 547262 369172 547262 369172 0 dso_counter\[1\]
rlabel metal3 511282 379780 511282 379780 0 dso_counter\[2\]
rlabel metal3 511650 380324 511650 380324 0 dso_counter\[3\]
rlabel metal3 511604 380868 511604 380868 0 dso_counter\[4\]
rlabel metal2 547170 370396 547170 370396 0 dso_counter\[5\]
rlabel metal2 544410 367268 544410 367268 0 dso_counter\[6\]
rlabel metal2 561154 359254 561154 359254 0 dso_counter\[7\]
rlabel metal2 562626 359356 562626 359356 0 dso_counter\[8\]
rlabel metal2 519754 370804 519754 370804 0 dso_counter\[9\]
rlabel metal2 456734 387522 456734 387522 0 dso_diceroll\[0\]
rlabel metal2 457661 385900 457661 385900 0 dso_diceroll\[1\]
rlabel metal2 458206 389324 458206 389324 0 dso_diceroll\[2\]
rlabel metal2 459133 385900 459133 385900 0 dso_diceroll\[3\]
rlabel metal2 462806 389028 462806 389028 0 dso_diceroll\[4\]
rlabel metal2 462622 391544 462622 391544 0 dso_diceroll\[5\]
rlabel metal2 461150 389256 461150 389256 0 dso_diceroll\[6\]
rlabel metal2 462077 385900 462077 385900 0 dso_diceroll\[7\]
rlabel metal3 449152 352580 449152 352580 0 dso_mc14500\[0\]
rlabel metal3 449014 353260 449014 353260 0 dso_mc14500\[1\]
rlabel metal3 448876 353940 448876 353940 0 dso_mc14500\[2\]
rlabel metal3 448922 354620 448922 354620 0 dso_mc14500\[3\]
rlabel metal2 485224 500140 485224 500140 0 dso_mc14500\[4\]
rlabel metal2 486420 500140 486420 500140 0 dso_mc14500\[5\]
rlabel metal2 487478 500140 487478 500140 0 dso_mc14500\[6\]
rlabel metal2 489102 500140 489102 500140 0 dso_mc14500\[7\]
rlabel metal3 449842 358020 449842 358020 0 dso_mc14500\[8\]
rlabel metal2 450701 500140 450701 500140 0 dso_multiplier\[0\]
rlabel metal2 451773 385900 451773 385900 0 dso_multiplier\[1\]
rlabel metal2 452463 385900 452463 385900 0 dso_multiplier\[2\]
rlabel metal2 453054 387522 453054 387522 0 dso_multiplier\[3\]
rlabel metal2 453889 385900 453889 385900 0 dso_multiplier\[4\]
rlabel metal2 454717 385900 454717 385900 0 dso_multiplier\[5\]
rlabel metal2 455262 389607 455262 389607 0 dso_multiplier\[6\]
rlabel metal2 461058 498552 461058 498552 0 dso_multiplier\[7\]
rlabel metal2 485990 319508 485990 319508 0 dso_posit\[0\]
rlabel metal2 486266 313286 486266 313286 0 dso_posit\[1\]
rlabel metal2 486542 304344 486542 304344 0 dso_posit\[2\]
rlabel metal2 486910 292259 486910 292259 0 dso_posit\[3\]
rlabel metal1 445556 358870 445556 358870 0 dso_tbb1143\[0\]
rlabel metal2 447166 359431 447166 359431 0 dso_tbb1143\[1\]
rlabel metal2 447166 360485 447166 360485 0 dso_tbb1143\[2\]
rlabel metal1 444774 360298 444774 360298 0 dso_tbb1143\[3\]
rlabel metal1 445602 361658 445602 361658 0 dso_tbb1143\[4\]
rlabel metal2 447166 362185 447166 362185 0 dso_tbb1143\[5\]
rlabel metal2 447166 363239 447166 363239 0 dso_tbb1143\[6\]
rlabel metal2 447258 363545 447258 363545 0 dso_tbb1143\[7\]
rlabel metal2 502550 320766 502550 320766 0 dso_tune
rlabel metal2 403650 203218 403650 203218 0 dso_vgatest\[0\]
rlabel metal2 408234 104924 408234 104924 0 dso_vgatest\[1\]
rlabel metal2 503378 319440 503378 319440 0 dso_vgatest\[2\]
rlabel metal2 450662 211174 450662 211174 0 dso_vgatest\[3\]
rlabel metal2 426680 104924 426680 104924 0 dso_vgatest\[4\]
rlabel metal2 450570 211956 450570 211956 0 dso_vgatest\[5\]
rlabel metal2 450846 209236 450846 209236 0 dso_vgatest\[6\]
rlabel metal2 445172 104924 445172 104924 0 dso_vgatest\[7\]
rlabel metal2 451198 104924 451198 104924 0 dso_vgatest\[8\]
rlabel metal2 457546 104924 457546 104924 0 dso_vgatest\[9\]
rlabel metal2 580198 6715 580198 6715 0 io_in[0]
rlabel metal2 580198 457453 580198 457453 0 io_in[10]
rlabel metal3 582046 511292 582046 511292 0 io_in[11]
rlabel metal3 581908 564332 581908 564332 0 io_in[12]
rlabel metal2 580198 617185 580198 617185 0 io_in[13]
rlabel via2 580198 670701 580198 670701 0 io_in[14]
rlabel metal3 558923 699788 558923 699788 0 io_in[15]
rlabel metal1 446108 422994 446108 422994 0 io_in[16]
rlabel metal2 429870 702093 429870 702093 0 io_in[17]
rlabel metal2 365010 702178 365010 702178 0 io_in[18]
rlabel metal4 444268 504560 444268 504560 0 io_in[19]
rlabel metal2 580198 46597 580198 46597 0 io_in[1]
rlabel metal2 235198 702076 235198 702076 0 io_in[20]
rlabel metal2 446430 510918 446430 510918 0 io_in[21]
rlabel metal3 444153 421940 444153 421940 0 io_in[22]
rlabel metal2 40526 701957 40526 701957 0 io_in[23]
rlabel metal3 1786 684284 1786 684284 0 io_in[24]
rlabel metal3 2016 632060 2016 632060 0 io_in[25]
rlabel metal3 1786 579972 1786 579972 0 io_in[26]
rlabel metal3 2154 527884 2154 527884 0 io_in[27]
rlabel metal3 1970 475660 1970 475660 0 io_in[28]
rlabel metal3 2016 423572 2016 423572 0 io_in[29]
rlabel metal2 580198 86547 580198 86547 0 io_in[2]
rlabel metal3 2108 371348 2108 371348 0 io_in[30]
rlabel metal1 4554 253946 4554 253946 0 io_in[31]
rlabel metal3 1878 267172 1878 267172 0 io_in[32]
rlabel metal3 2108 214948 2108 214948 0 io_in[33]
rlabel metal3 1832 162860 1832 162860 0 io_in[34]
rlabel metal3 1855 110636 1855 110636 0 io_in[35]
rlabel metal3 1970 71604 1970 71604 0 io_in[36]
rlabel metal3 1602 32436 1602 32436 0 io_in[37]
rlabel metal2 580198 126463 580198 126463 0 io_in[3]
rlabel metal2 580198 166413 580198 166413 0 io_in[4]
rlabel metal2 579830 206329 579830 206329 0 io_in[5]
rlabel via2 580198 245565 580198 245565 0 io_in[6]
rlabel metal2 580198 299081 580198 299081 0 io_in[7]
rlabel metal2 580198 351985 580198 351985 0 io_in[8]
rlabel metal2 580198 404651 580198 404651 0 io_in[9]
rlabel metal2 562350 169490 562350 169490 0 io_oeb[0]
rlabel metal2 580198 484517 580198 484517 0 io_oeb[10]
rlabel metal2 580198 537319 580198 537319 0 io_oeb[11]
rlabel metal2 519570 455226 519570 455226 0 io_oeb[12]
rlabel metal3 581908 644028 581908 644028 0 io_oeb[13]
rlabel metal2 580198 697085 580198 697085 0 io_oeb[14]
rlabel metal3 523457 502316 523457 502316 0 io_oeb[15]
rlabel metal2 447810 528530 447810 528530 0 io_oeb[16]
rlabel metal2 444130 510952 444130 510952 0 io_oeb[17]
rlabel metal2 332534 702144 332534 702144 0 io_oeb[18]
rlabel metal2 449282 511224 449282 511224 0 io_oeb[19]
rlabel metal2 544410 192134 544410 192134 0 io_oeb[1]
rlabel metal4 449604 510748 449604 510748 0 io_oeb[20]
rlabel metal2 137862 694426 137862 694426 0 io_oeb[21]
rlabel metal2 442474 328219 442474 328219 0 io_oeb[22]
rlabel metal2 442750 328729 442750 328729 0 io_oeb[23]
rlabel metal3 1740 658172 1740 658172 0 io_oeb[24]
rlabel metal3 1855 606084 1855 606084 0 io_oeb[25]
rlabel metal2 4140 683060 4140 683060 0 io_oeb[26]
rlabel metal3 2062 501772 2062 501772 0 io_oeb[27]
rlabel metal3 1878 449548 1878 449548 0 io_oeb[28]
rlabel metal2 462254 272102 462254 272102 0 io_oeb[29]
rlabel metal2 579830 112965 579830 112965 0 io_oeb[2]
rlabel metal1 4186 292570 4186 292570 0 io_oeb[30]
rlabel metal3 2016 293148 2016 293148 0 io_oeb[31]
rlabel metal3 2062 241060 2062 241060 0 io_oeb[32]
rlabel metal3 2200 188836 2200 188836 0 io_oeb[33]
rlabel metal3 2967 98668 2967 98668 0 io_oeb[34]
rlabel metal3 2016 84660 2016 84660 0 io_oeb[35]
rlabel metal3 1878 45492 1878 45492 0 io_oeb[36]
rlabel metal3 1878 6460 1878 6460 0 io_oeb[37]
rlabel metal2 580198 152915 580198 152915 0 io_oeb[3]
rlabel metal2 580198 192831 580198 192831 0 io_oeb[4]
rlabel metal2 580198 232781 580198 232781 0 io_oeb[5]
rlabel metal3 581908 272204 581908 272204 0 io_oeb[6]
rlabel metal2 580198 323561 580198 323561 0 io_oeb[7]
rlabel metal3 582138 378420 582138 378420 0 io_oeb[8]
rlabel metal2 580198 431103 580198 431103 0 io_oeb[9]
rlabel metal2 580014 20213 580014 20213 0 io_out[0]
rlabel metal2 467774 321038 467774 321038 0 io_out[10]
rlabel metal3 582000 524484 582000 524484 0 io_out[11]
rlabel metal2 580198 577269 580198 577269 0 io_out[12]
rlabel metal2 468602 321072 468602 321072 0 io_out[13]
rlabel metal2 468878 321752 468878 321752 0 io_out[14]
rlabel metal2 469154 321701 469154 321701 0 io_out[15]
rlabel metal2 445694 509388 445694 509388 0 io_out[16]
rlabel metal2 449466 327794 449466 327794 0 io_out[17]
rlabel metal2 348818 695038 348818 695038 0 io_out[18]
rlabel metal2 446706 503846 446706 503846 0 io_out[19]
rlabel metal2 580198 60163 580198 60163 0 io_out[1]
rlabel metal2 219006 697826 219006 697826 0 io_out[20]
rlabel metal2 154146 702008 154146 702008 0 io_out[21]
rlabel metal2 89194 694392 89194 694392 0 io_out[22]
rlabel metal2 24334 695021 24334 695021 0 io_out[23]
rlabel metal3 2039 671228 2039 671228 0 io_out[24]
rlabel metal3 1947 619140 1947 619140 0 io_out[25]
rlabel metal3 1832 566916 1832 566916 0 io_out[26]
rlabel metal3 2108 514828 2108 514828 0 io_out[27]
rlabel metal3 1924 462604 1924 462604 0 io_out[28]
rlabel metal3 2154 410516 2154 410516 0 io_out[29]
rlabel metal2 580198 100079 580198 100079 0 io_out[2]
rlabel metal1 5336 59330 5336 59330 0 io_out[30]
rlabel metal3 1970 306204 1970 306204 0 io_out[31]
rlabel metal3 1924 254116 1924 254116 0 io_out[32]
rlabel metal3 2154 201892 2154 201892 0 io_out[33]
rlabel metal3 1786 149804 1786 149804 0 io_out[34]
rlabel metal3 1947 97580 1947 97580 0 io_out[35]
rlabel metal3 1970 58548 1970 58548 0 io_out[36]
rlabel metal3 1878 19380 1878 19380 0 io_out[37]
rlabel via2 580198 139349 580198 139349 0 io_out[3]
rlabel metal2 580198 179265 580198 179265 0 io_out[4]
rlabel metal3 581908 219028 581908 219028 0 io_out[5]
rlabel metal2 466670 296626 466670 296626 0 io_out[6]
rlabel metal2 580198 312647 580198 312647 0 io_out[7]
rlabel metal2 580198 364735 580198 364735 0 io_out[8]
rlabel metal2 467498 321004 467498 321004 0 io_out[9]
rlabel metal1 486496 319090 486496 319090 0 oeb_6502
rlabel metal3 539281 137972 539281 137972 0 oeb_as1802
rlabel metal2 462477 385900 462477 385900 0 oeb_as2650
rlabel metal2 447166 384421 447166 384421 0 oeb_as512512512
rlabel metal2 503293 385900 503293 385900 0 oeb_as5401
rlabel metal3 449566 358700 449566 358700 0 oeb_mc14500
rlabel metal2 448346 159868 448346 159868 0 rst_6502
rlabel via1 427754 444397 427754 444397 0 rst_LCD
rlabel metal3 449980 345100 449980 345100 0 rst_as1802
rlabel metal3 449980 345780 449980 345780 0 rst_as2650
rlabel metal2 447166 347429 447166 347429 0 rst_as512512512
rlabel metal3 449934 346460 449934 346460 0 rst_as5401
rlabel metal3 449750 347820 449750 347820 0 rst_counter
rlabel metal3 449244 348500 449244 348500 0 rst_diceroll
rlabel metal3 449221 349180 449221 349180 0 rst_mc14500
rlabel metal3 448876 349860 448876 349860 0 rst_posit
rlabel metal2 405957 334900 405957 334900 0 rst_tbb1143
rlabel metal3 449198 351220 449198 351220 0 rst_tune
rlabel via2 447166 351917 447166 351917 0 rst_vgatest
rlabel metal2 598 1843 598 1843 0 wb_clk_i
rlabel metal2 1702 1911 1702 1911 0 wb_rst_i
rlabel metal2 2898 1979 2898 1979 0 wbs_ack_o
rlabel metal1 194580 44846 194580 44846 0 wbs_adr_i[0]
rlabel metal1 213624 44914 213624 44914 0 wbs_adr_i[10]
rlabel metal1 215050 44982 215050 44982 0 wbs_adr_i[11]
rlabel metal1 217212 45050 217212 45050 0 wbs_adr_i[12]
rlabel metal2 58466 22736 58466 22736 0 wbs_adr_i[13]
rlabel metal2 62054 22770 62054 22770 0 wbs_adr_i[14]
rlabel metal1 220938 45254 220938 45254 0 wbs_adr_i[15]
rlabel metal1 222824 44778 222824 44778 0 wbs_adr_i[16]
rlabel metal1 224618 44710 224618 44710 0 wbs_adr_i[17]
rlabel metal2 76222 22498 76222 22498 0 wbs_adr_i[18]
rlabel metal2 79718 21240 79718 21240 0 wbs_adr_i[19]
rlabel metal2 373566 171020 373566 171020 0 wbs_adr_i[1]
rlabel metal2 83306 21274 83306 21274 0 wbs_adr_i[20]
rlabel metal2 370806 171496 370806 171496 0 wbs_adr_i[21]
rlabel metal2 370898 171428 370898 171428 0 wbs_adr_i[22]
rlabel metal2 93978 21376 93978 21376 0 wbs_adr_i[23]
rlabel metal2 97474 21410 97474 21410 0 wbs_adr_i[24]
rlabel metal2 101062 21444 101062 21444 0 wbs_adr_i[25]
rlabel metal2 368046 171462 368046 171462 0 wbs_adr_i[26]
rlabel metal2 367954 171632 367954 171632 0 wbs_adr_i[27]
rlabel metal2 365286 171428 365286 171428 0 wbs_adr_i[28]
rlabel metal2 115230 21172 115230 21172 0 wbs_adr_i[29]
rlabel metal2 17066 1775 17066 1775 0 wbs_adr_i[2]
rlabel metal2 118818 20186 118818 20186 0 wbs_adr_i[30]
rlabel metal2 122314 19812 122314 19812 0 wbs_adr_i[31]
rlabel metal2 21850 1962 21850 1962 0 wbs_adr_i[3]
rlabel metal2 365194 168521 365194 168521 0 wbs_adr_i[4]
rlabel metal2 30130 2030 30130 2030 0 wbs_adr_i[5]
rlabel metal1 198030 39474 198030 39474 0 wbs_adr_i[6]
rlabel metal2 37214 19948 37214 19948 0 wbs_adr_i[7]
rlabel metal2 40710 19982 40710 19982 0 wbs_adr_i[8]
rlabel metal2 44298 1996 44298 1996 0 wbs_adr_i[9]
rlabel metal2 4094 19846 4094 19846 0 wbs_cyc_i
rlabel metal2 8786 2183 8786 2183 0 wbs_dat_i[0]
rlabel metal2 366574 168674 366574 168674 0 wbs_dat_i[10]
rlabel metal2 369242 168810 369242 168810 0 wbs_dat_i[11]
rlabel metal2 56074 20084 56074 20084 0 wbs_dat_i[12]
rlabel metal2 59662 20118 59662 20118 0 wbs_dat_i[13]
rlabel metal2 63250 20152 63250 20152 0 wbs_dat_i[14]
rlabel metal2 371910 165614 371910 165614 0 wbs_dat_i[15]
rlabel metal2 372002 165852 372002 165852 0 wbs_dat_i[16]
rlabel metal2 373382 165750 373382 165750 0 wbs_dat_i[17]
rlabel metal2 77418 18554 77418 18554 0 wbs_dat_i[18]
rlabel metal2 80914 18588 80914 18588 0 wbs_dat_i[19]
rlabel metal2 13570 2115 13570 2115 0 wbs_dat_i[1]
rlabel metal1 230368 36890 230368 36890 0 wbs_dat_i[20]
rlabel metal1 231518 36958 231518 36958 0 wbs_dat_i[21]
rlabel metal1 233358 37026 233358 37026 0 wbs_dat_i[22]
rlabel metal2 95174 18724 95174 18724 0 wbs_dat_i[23]
rlabel metal2 98670 18758 98670 18758 0 wbs_dat_i[24]
rlabel metal2 102258 18792 102258 18792 0 wbs_dat_i[25]
rlabel metal2 520490 330344 520490 330344 0 wbs_dat_i[26]
rlabel metal1 449190 292298 449190 292298 0 wbs_dat_i[27]
rlabel metal1 447626 292366 447626 292366 0 wbs_dat_i[28]
rlabel metal2 116426 17364 116426 17364 0 wbs_dat_i[29]
rlabel metal2 18262 17058 18262 17058 0 wbs_dat_i[2]
rlabel metal2 119922 17398 119922 17398 0 wbs_dat_i[30]
rlabel metal2 385710 210120 385710 210120 0 wbs_dat_i[31]
rlabel metal2 23046 17092 23046 17092 0 wbs_dat_i[3]
rlabel metal2 385894 147628 385894 147628 0 wbs_dat_i[4]
rlabel metal2 519478 313276 519478 313276 0 wbs_dat_i[5]
rlabel metal2 520766 314534 520766 314534 0 wbs_dat_i[6]
rlabel metal2 38410 2064 38410 2064 0 wbs_dat_i[7]
rlabel metal2 41906 17228 41906 17228 0 wbs_dat_i[8]
rlabel metal2 45494 17262 45494 17262 0 wbs_dat_i[9]
rlabel metal2 9982 2047 9982 2047 0 wbs_dat_o[0]
rlabel metal2 519110 316880 519110 316880 0 wbs_dat_o[10]
rlabel metal2 365010 153442 365010 153442 0 wbs_dat_o[11]
rlabel metal2 57270 15732 57270 15732 0 wbs_dat_o[12]
rlabel metal2 60858 15766 60858 15766 0 wbs_dat_o[13]
rlabel metal2 64354 15800 64354 15800 0 wbs_dat_o[14]
rlabel metal2 523342 320654 523342 320654 0 wbs_dat_o[15]
rlabel metal1 450524 289714 450524 289714 0 wbs_dat_o[16]
rlabel metal2 75026 2200 75026 2200 0 wbs_dat_o[17]
rlabel metal2 78614 15902 78614 15902 0 wbs_dat_o[18]
rlabel metal2 82110 2234 82110 2234 0 wbs_dat_o[19]
rlabel metal2 384698 160004 384698 160004 0 wbs_dat_o[1]
rlabel metal2 518926 324870 518926 324870 0 wbs_dat_o[20]
rlabel metal2 89194 1860 89194 1860 0 wbs_dat_o[21]
rlabel metal2 523250 326094 523250 326094 0 wbs_dat_o[22]
rlabel metal2 96278 16004 96278 16004 0 wbs_dat_o[23]
rlabel metal2 99866 16038 99866 16038 0 wbs_dat_o[24]
rlabel metal2 103362 1826 103362 1826 0 wbs_dat_o[25]
rlabel metal2 369334 158678 369334 158678 0 wbs_dat_o[26]
rlabel metal2 110538 1792 110538 1792 0 wbs_dat_o[27]
rlabel metal2 114034 14542 114034 14542 0 wbs_dat_o[28]
rlabel metal2 117622 14610 117622 14610 0 wbs_dat_o[29]
rlabel metal2 19458 14440 19458 14440 0 wbs_dat_o[2]
rlabel metal2 121118 14576 121118 14576 0 wbs_dat_o[30]
rlabel metal1 446246 386478 446246 386478 0 wbs_dat_o[31]
rlabel metal2 24242 1894 24242 1894 0 wbs_dat_o[3]
rlabel metal2 520950 320824 520950 320824 0 wbs_dat_o[4]
rlabel metal2 462438 114716 462438 114716 0 wbs_dat_o[5]
rlabel metal2 36018 14372 36018 14372 0 wbs_dat_o[6]
rlabel metal2 39606 2098 39606 2098 0 wbs_dat_o[7]
rlabel metal2 43102 14406 43102 14406 0 wbs_dat_o[8]
rlabel metal2 46690 2132 46690 2132 0 wbs_dat_o[9]
rlabel metal2 5290 14304 5290 14304 0 wbs_stb_i
rlabel metal2 6486 1792 6486 1792 0 wbs_we_i
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
